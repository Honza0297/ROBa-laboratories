PK   -�OV]� �  �    cirkitFile.json�]]o�F��+ͫ٨�*�mfg�ld�}�n�H��uK^YN'��nK��\�=e��ql�=:�uxY�>��\����m�����v���m�\�,>���S}�Wv���l�î�u_�X���/ܷ�r���r��T�u#�Z5�j-e��]K��B��U��1]��-n߾�������dTV	2*�$��U�́��*M�@E`�!s�"�ʒ9PX����*��]��J2D���'�����n�nU�k��[��B-�-J�4W�e+.�u%Ղx�8����Q�˱;(�z�xY����r�X��,ZǄ��-[�7��!��c<�c�/�x����}��K��ww�~s��ض�R�JepC�� �}�-�ٴ�;�������=��~�@�#����_~d�ntL��!:�D�ѱ �
����'d���UB��X�2Dǂ�2�!:���ѱ��d��=v�_)���6ͺ����U(֬�reV[1��M���Ǝ$&~�D�1��ή{q"�]�!|eǱ��;1d7�	`�'�co��7F�ĺ]b%eǱ�X���SX�A�q,;Vi��4�wPvˎU�;���ǲc����b}eǱ�X尾sX�A�q,;V�XߕX�A�q,;�W��,?��Wp��C'&����ppn¡cx��������,ˏ����3������\���/�%��g+����W88a���`~~��?p҂������U���3������Ã���pp������:8xf��`�q0?���8����`~~����ˏ���]`���,?���{���~��8��ߩ�x�ˏ���=6`���,?��w��N_��8�����8����`~~G���>��$i�2u�{k<rk�xon��v��p��D��nש�i�����uA�Q>�G���Љ��m�͇�1'�7RN� U�D���U���j?��<՞(��p�T{���CScQ�����D������l��jO�_��}�=Q�F�/A��$Q��'�O*�Z��z%Q��P�}K�xK�x��#��"><���(�ã�C`b�VD�+b�V�ୈ�SD�i��4Q��?Mԟ��`D�i��4Q��?Mԟ!���g��3D���Q��?Cԟ!���g���D�Y��,Q��?Kԟ���g���D�9��Q��?Gԟ#�ύ�/��&q5e
5�5��`��r�r�.V�1Y��5+�kV�J���kS�I��L2d�������d~E�)���0�|<&����$��H�&�숺�2��fOTޕi�4�+o�*O�y36�V|���r��s����jw���ˏ.������@�#�0��I1�@@}�R#P_���1�0�%M1�@@}�S#P_���?�0K��B$.j��m�ږ�	�yoW­�5�,r�>�6˥���	�9,x����I=��dN������˲�%�,��S�u�rE��Ἇ��}�,�sXG!�z���8.`�oұ�'�,���t,
���6G!��8�⸀�QH�"� N�8.`q|�^`4��Epk��Qa\�
�pT�_spˊb<0<#
G��u8z���5ƕ���Q8*P�9��5E1�)�����kXo��YS8*Я9���H1�A�����kX����T8*Я9��5L1�Y�����kX���T8*Я9���OA#�IL�*h�'���6R��m��+O��&��"}�'���6RV��m��+�H�U<,ҷyR�,l#�X��٘,l#EVANȓ�%MANȓ�ea�Ê�E�6O:��m�F+fA!�e
rB��,�HV<,ҷyҲ,l#�Y�@�fa��
rB��,��
rB��,�HQW<,ҷ�����eAAU<,ҷy�,l#�`�H���˲�����"}�'/��6RD��m��,�H�Y<,ҷy�,l#�g�H���˲�����"w%��ˢl���+�PF�rO�C@�/=�*- e����� .#�~�W���쭝Qs�Q��!��h0����Q����ر�%kQ���43��"`0*;h2��-��3*�"`0*�K��%h(�Q�<�xx�yF�[�^���%k=�����g7�Q�¨XaT�0*V�1&+��&+L,V+��5F��b�Q�ƨX�;��5F��b�Q�ƨ�`Tl0*6��F��b�Q����`Tl0*�[��-F��b�Q�Ũ؂��0*�[��F��b�Q�è�aT�Uqj)��3Ωexc�
���}�+�P��Lj]] ʳ�I��@y6����<�R+�"T/F�ϯ-$W�E�`����X�7Vumz�ݯu��J�>�C(��m���߼� �c	]#б�.��XB�t,�a:�Ѕ0K�B���%t!�@@��F �c	]#Щ�.&D�6.l��6�nҩ�.�,vsX�F!�J�b8��7�pҩ�.�,�sXG!�J�b8�⸀�qҩ�.�n����⸀�qҩ�.�,�XG!�J�b8�⸀�qҩ�.�,�XC��E���P#%tѨ0���hT�_sp��Ѕx 8��F�5�H	]���hT�_sp��Ѕx 8{�F�5�H	]��s�hT�_sp��Ѕx 8s�F�5�H	]���hT�_sp��Ѕx 8k�F�5�H	]��s�hT�_sp���Ō��$\aQZ�>Oʕ�m��.��LiW��+,J�E�6Oꕅm��.��<�W���pX�o�`Y��J��a��͓�ea+��E�6O*��m��.��<�X���pX�o�dY��J��a��͓�ea+��E�,��˲���Ѕ�"}�'/��6VB��m�%�<yYX���m��,�X	]8,ҷy�,lc%t�H���˲���Ѕ�"}�'/��6VB��m��,�X	]8,ҷy�,lc%t�H���˒��(�KG��=��.ed���t��=�3J��QF���(�KG�[;��. �ޱC`sJ�`0;5��. ��cCsJ��F�c�i���`T<v�dN	] F�c'0���`T,1*�K�P�b�Q�ĨXbT,1*�K��F�
�b�Q���1*V+��F�
�b�Q�ƨXcT�1*�kPb�Q�ƨXcT�1*���F��b�Q���؀�'0*6��F��b�Q�Ũ�bTl1*�[�4F��b�Q�è�aT�0*v;��ݳ*N.�KGy���K��Q0\��Lr	]:ʳ�I.�KGy6�%�Х�<�K�T/F�ϯ-����`����ZB��r�O�o����P�vw�}�i~_�ru���ٷ��]�j�j��v���/n߾%,��׃�r�.;�\td��֮UM�ؼ^Y��²*�o�3�/�Dha�Z�RJ8Y�\��ڶ�mZe�i��(��T�W.���h��n/�& A����ā�:M���7���k�VFw�γ�^,�6�Y�0k�u����)mi36Yd��њ��l��J3i�+l��U7�{;!i�,׌)9���I����>:O_'}�+�5���yR�y.
ǥ$R����W���{E&@����Ur�1���q5��3�\�kr�@��,�<�<6��yd��۬��T:n4�U|�YJ��}����YU�)3�O�q�T䏧$]��{��O����_fv����omS��&6��#�5���J�}��'~~;��Px��$�W�	�3BOF}k����x,|4�9�!���S�3�N�^e�*3�tF�V����ރ�#c2#���y�_dV�΀:aJg@�7�3�N��+�e>�ڳ�2]@f@�!��Q|&���	�A�x�"�(t�x@b _U8^��i����)��}���T�Z�}���Et����7dF�����5�53u�\6߀���(K�<s�5�\���׌/�������l>Y_�s������-kV�2y2��Y��$t�F\�e�o�5���F�	������v�`X�7�\5��>����n�!A�u�aA�|�aAރ��Xt���C}h�_߭�G�갫7���O
Y^��(��!XތȂ��S�Dd֟�%� C��T.����z�,��?LdA�`��b"2�O%Y�!X��Ȃ�����a=}�c��,� ��Ǵ�� ��Ǿ�� �r@ĥc��9�{8� �5s�$� (�5x�J"-@��k�h	"-@�怸M�`�"�ԑ p������e��< �Y ƾtv,�L���0��c�c�g*@��10��MSy � ����$�z��E$�<����X����������.��!���o o�R��!]��_�Ã�ˏ���*�*?�X~̏U����� ����`~�
������cU�{8<����8�������A������X|}�?,?�����itBf���ڇ�������K8v���9��_�A����r4C�҄�!:#3�h���K(`t��tj��	�a��y
G'*`���r�2Ƈ�d̐��[M�/���1.E'0`�~�-Ktf���#DP@��9��_oG��ŀr4C�W �Ctf���>��Y�!G3�{4�>Dg1`����/A���f������i�!G3��z�>D�-`����IB����r4��JY� �$�^�h�<B�p�a�`��D�`k�D�`K���xD�`����3�3�N�sr�}��q�}�Sq���z�
2<�2�*����T�`?�T ��S�B� LLT%����P�
@Ub��}* U��^� T%������J�T%J�[��D���,�?U�2r؍RDG>wJm*U��*[E����VQe�ȣKj UT�*j U� ��JTT%j�5U���DMU�&':T%j�5U���DMU��*�P�h�J4T%�U���DCU��*�P�h�J�T%Z�-U���DKU�%��P�h�J�T%:�U���DGU��*�]Qbb	��g&'P�~���\���˂��vpkS��fwͪ^��r~u�:���B��$���>���#���:R쯄�$�+Q*��J�J�����C U�צ�� ��6-�p�m�V��z}�Ʌ5#E�>�,�`6�����?��)�xq�v���
�7�z~>��5!_���Y�i"?����r�E1�"��7�5���:��po!��豽���[o!����[o!������-����Bz�-����By�-��P�x�-��P�By�-����B{�-t��B{�-�����x�-��0��x���[oa����[Xoa����[Xoa{�z�-��p��y�-��p�����^��Ş:�$H����h����u�}<�u��X��b��o��oi�)
9�76���W�����`�T�
*C�׷����~�ot_F��Zu: d���������
>\�!2�V�~z���]�l��a�ӏ���=��wpE�.��>]��%~���K�tI����/��%^��K6��N�\x�<]*� �����zg�]請���w_ҷEٽ���l���kׇ��:Y���R��U��7�<��L�������5��I_�������2��i��o��Mۏ�?�o�/�Λ��f�������_�Y�V�=���������#�������ӏ��p�����.>��_6��]��o��7��Y�:�]w}����zuxܷ�kΛ�19f0�to��a����\�9���7�so����)~��-JU����FvO��]��u�j�KW�e7r�YtYơޮ�6I���b��tV�,�]���f��kO����ھ�7�`�\K����E^�7�O��E?O�v���W�%*?�����E6�#�.��9�փk�7������R�>�/��ܙx9~M^�3g�v��vO��K���|�X��W�Ը�>��m�+.�A���n�]�N�vQg�͢��{ ����h�.޻��f� Ǽ�x���ai6|�F��ɑf.-x��M�P�H,�!�2퓵JRo˱+N�])]$�:��ˆc�D�]	�xWB�������O���	��_刅pcf�BmN���V��zE���t�ّ+���v�ƌڨQ9j�Gmؘ�3���S7��W���@؝�v�ލ�;;�.��x����"ʈ7�%�0��hØ��#��7��,�0��xÈ�#��7�4�0��h��|�v����o?���v�p��7���H�r9d��+�3.?bڛ.��.���u>vW�6Kݬ��r?��T����r����.��ݓ���c���`�n�S賆�x��Y.�����(�?�������Y�w�]�:�w�����	;T�M��s9a����{���®库��z�J��S�����TNJq�o}��ؕȃi&��>��Vڦ�R��&��� ��o�w���G�/���;z$~)pI�Y��x��)�v�W"���O�vt�[S�����_��6�ަ����0Z+st��2i����O�u1ճld��mS��{�]Ө�tm]�V���f��lL�����×�Ƌ� ��d�^��+�l�T_d�_yN~�q��mz]v�����O���������/���o�6�ჇP���Er�C�ǰۅSOֿM��������C�����O��p��M�鿺�z���4|�ۿ[ܾ[��1o�nq�O�?���~���f�t�`�@Q>{�}��g$�����m����Ç��w��-�4�������������o?n��|T�"��n"�.�_[ig��*T��23Zi6 �����N�����:P�����m�9Z��S5h�����^��LD��e��V�����`R+9|�����-`�`93N����Ux�+?�n9'}�b~7�݈~Z�Z��od���-�9�J�b�xyN�O|���e��}���c��Di���%ͣ�?h�{�ٳ��7�H����#���Ť�h��9/"^��,��o�����Z��<�ݳ�N�]�Ի���H|����J��_��_��%�����sX���U!������I͒Guk[�Z��G�wf�˳��<�S�"��"z�꠰ϴ��`%ܪ\�e �20e �20�d�S^�V�[@Fe����-�,P6�,Zv��@%��/[]n��A��(?�����q�C}h����B������߶���>�w�}���~|�T�^|�PK   ]�'V�cŌ ~ �� /   images/40a6b5df-e714-4004-b865-d48720df955d.png�eP]��.
�����-�-�������݂��w�.��!�%�����{������=�V1�{�7z|�Cz-��dD�ap`@@@��ń@@@{�|� >z<�F�A@p;ݕ��]l�m��,��l��\͌A@\W�������k�u���S�+\��.�=�Xn���" C�lBC���{�Z��*v��KY(�?~J����>z�1i��9xx~U�:Q|rz؅�!ß=����~������tww7��?�=���!��M%6���wz�O����=v=���K:~���������wv��I���y��r0A��E��"����+��������E��bOj������Ъ�4�����]��ד�E��"]�o�/g't��b|���k>#�ի�������]�ޛ,�ĪE���s��&���0��\�*^�6�Hg�X|�U:��c��*5H������<U��Cx1sT�-����&vƯ���Ik��#w�Y�/��K�.M�]���5ݪo�1�m�-�rP=_Z����e���С,�ҷ.�u�K��`0~�H���$_ғ�UO�!b��a�Y�|�ܙ�	�\�!F:��INV���3�S�X�c�O�j<�/ާ�m�Dq[��4!�W1�����Ȁ}��/'MQ07+Ĥ�/J�(ml�R��m<�0kl\Ho�V��]ѼX�]c
=C�R��V`?��A�e�d����Դ\���4;IUݩq>��vW�mɩy��̮77I�wonV��y�p�ڞm��ĪY�mWt�s�wqv�|�r�#U!b�W����NDd!ra�|���iҜ�|�}�a�2���l��I��MT"�o�k�.��0�Е��*[$��i�'9P�oV�e�ܷ�Y�L��?��%���E.��jh��:vu^�~}O@LԤ�.�8Q�T18-G?��jF�>�����b;]�о9׀$ݞ]<�q�P,�>�j�&E��<*���=����Ӹ.������n?�vYJ���F �
u[s�e#�pR�}�z�I��O#����њ>=B����%��8 ~R�p+�-��Q��^������[��m�l?��w$銜�<���.͝��a����U��݄fxG�ި��|�F�A�������b n��Nt��S[��&񍣉5y1�Hk�w�U�V��]��j9�g �-[|Ԃ~��n�<}��C��a���u��jz��r�3x�ЗA?z\�~Sc��%@�������E�=��R�������@�ѹ8_#Y��W�ʁ&���U��f-ƗXJ���bv;�bi� 8��"�����(�$��a�Ndk�,��q�Nv�7[���L_�%����75?��l���wq��D�(2�;t��d+�#�|��^x�6��q9k��(�;3h�Y���82_¡�c��c��t���0��3a�ih�y��w�����"�v�Wݚ�9�.@����{L���OHgp��E�o;k8�2�Ԩ�y;�΅����S���r�i�4˃.0��mՂ����g�Z�I��rU�C2�n'n����:�_Pkk�-����H0�t�猾���KpS�� ���S�\؆s���E1���L��� ��Ær[�����&#�j�GS	K�l��}��fV�§��F��T�,2^�[�,�����������_x�h�น��N,��rm������!�H���98Q��~��&913j ]*�*NG���2V 1����?5���
���(�M"QX��?D�2�zXkS!H��%�-zl1-\��D�(M��*��i#Df[q��qK˪TRD��JA�1鏗�H��ll�!�Q�R�؁�*okC�p��-�A�98C�CQ��>	ί�0��}-k��x��Ϝ$�Yѹ��Ð<���̓�-d���+`���(��P9�o�[b���+�P��%���1F	�cEZ.��g3G9��v�Ce+����3tx��y!/`c/�;_3��B���`w
>5�%0��zj���"���9�o����Z��m4�2���/��� 0�7�R��u������I�x8�!��4K�f4D�1����<�j(s�%���05�%`IŢ
�]��%ǁ�+t�P��:������S>t�pUȼĘ&i� ��o�X����W���[	���uS��F�e�i�K��kCB��^�jZ�6�|_vl^��v�QU-�f����Dp���F���4�5(�\��POc^Ƒ0�4�����o>d��Ӡ	�C�����̩Ϛ_���&�f��|�����@�E{�*��1�N�'�#8�}&�mf�ݛ�()��0·������#��¼ U�X��$�kK��~�L�����&�h0 ��D�\ ���� �̨";/����Ӑ��bj9�-����T�}b�3%�&��~b����8G��F�P��W2ҭ�T�6B�C,Ra=�/H�8��3�t�C�����V�c�T����p�>��ف��K'<��)��#P�"hzg��ψеvO&��	9c���D��OpI��\���^>D#�oYߧ�q��_��4f.�{^�N8����
ϸH;A���z�@F�n�� G�y��� �w��!*��rU��zpgic�Kn���ᗏ>�E���x������,t��Mey�U]���B�i	N#K���K�Ks;Sc�x��1�Cy�ÖR�߳4~:'6ts
d6e��HL��5��P!�Gs�2���JгtsP��A/2�C��'�k��`��]�ځ�9[�6�\�[:t.A�$�:ظ�$�fQ.��V ��B�2�)z��L�
�:���mx� ,�]��`�'	���q)�g�qZ�2�������c����XW��/=C>foo�t�o��C�#�Z}�
r��q=�_y\l������5���po��4��8h ���4@����]�6s���T����R��>�V�K<v}ފmI�,f=�3L��1��ب@��h���]�������}\jM0��T"�)p�cuIw-y �m0��n�f�=�6�6J�C���HeQp����&[T� �.H�}5Xe��EW��9���,���>B+ș����%_�7�E�)�+/�@�� w�(1�fs��Lߎo=:#"4�=�����tv^f�M�>J��T�4��ەya�����h�0(��ӡv�8 � �.wi1H���0#=q�d66O��BȎ�Dl����W�Fo6}�!�w"��3��23�oJ}ˢ*�:<��Em�'����t��q}^(�ٹ�P~�����f"�N����q�ݘT?e]S� �e���6	�>�\H�_[&M�"r����$z�y|C��
��VA��ۿ*|�<BcGr]�R�SQD�A�E���.-����Y��!wf�}K�L�ҽE�Td�܈���(a��!��������������W��mT�$���\a�v>�PY���ˢ}p_�mv	��m�߰#!�SX�=jǣ/F��!�
Wb��g��@��D!�UNn�2�2�@�`��T3گ�)�Q��
���fn3.����}t���vcS�*א���q^9��"�#�2��J���q_fd�Jg����COz�*t��Z��T�O ��K:��ǻ�~��&D�Ƅ�ߝ��B7`)�u�"[��R�`7O�Q�~}FN0Z��S��
V�K�p��D&��+'FŠ�?��L?�7?UQ�{�[h#n"z�i�ᗞ9'�_��j����~�XTph��0|̋2��	�]ƈ��y��
;�E�#�����_Y
RJ" 3[�2��h�� 5�(u��=1���JD^�Q��!��[мQ+LLC�_�U��SY��s�,��#Bww�M�״e����<~r�0�a7�ўѥ���n�k=r_u��-+��؍oG\����+˔#2����@����M����Q7��d��0���r�O�n�tV�w�9ݠ=~堂6瘲���(o�!���V�Û�s�/�Ԉ��MG����h�8�������$yw��Q�����D�������yBU�+���
���Mh0w�1�PĿ��V��Q��at�ңp�����c��#D�axݪ�!�<r �{\�y�G}us|w�5M�k�H��(��v,�_�ʾ�R�%�̆Ɗ�Gl��
ZXhD��	 %����\/�W�P���O��HLN&Ks�R���@��̍H�������Z�S�+�Y��'�� a!l��s�CzR��'zt	o?E�FE ��iH*���s��=�RY$a+U�38-�짌>@}�8[�P�4��v�Qy����2�1yeMkT��[yױ2t�D����ρ1�`�_��|銣( pv��I�?ӆ�'T6*"��6�#�@Сq~B���V����9G��e<�:=�^��?�]����!??�|�Q�����堓n:�+k����6<�<�
hG�a�m���ՂC�&- n�q�����ɉ5�@FR�T�K�#�`���j�{�D&^?�iz����b�r�]�!� e���bY�sU���A�B�b��?194
��&�Џ�q���}eIp��H\ڗ{��!C�NK�֩j'���	a�����U�g����ΒH#/#��%�lj��H��Q�-}��$.9#绉��m3�AX�F�ݒ���S
R8P�sᯎ/e�])�/"�~�c8��5��A7���YvGz=���S"���~V*�����A�G��Zz6��fb1;{����a�J/��� ����'ɑ��J
/ٮ�0O)4*vuu��N��U���&�=���!-C�ϼ��B�+��$��������Z�_A�vZ�7�7�H����USkK���*�(�ۢ��.x糑�P�p#�*�xN���9aTu6����X2'���j�1�e��ƒ-Qx��s65�i��W�C�5(�5�/g�WW8�x��4��K��u��B�CP\�_d�`%6ֽ�M{�W�y���$��_���ʮ��)�C؛�t������]L��ۢh�Y�Qv!��W�z����A`ꡦE ���#g�48Ƶ�W��s��^O����DK��I��Q����ԟ�l'a�%A	������*Fx�����������8�G�QCm�&aQ��0���٣�����|/��sFKK�P^����XY�^��}��g�D��/d̂'	�%�Q��ZP�1�Jiu3(� !d��m�YZ�o�����xK �����,����ɭ�maE���l�q�H��3z�v'��&�t-��:Js`}bx�t	2a�G����q�L��|ھ�:ό��
ħ"u6���cw�=H��mW���Y��C�H���5��A%���%�bV�;��:�>ꁤZz٪Q�$�}�K�(|�G1{�UD����rK��L����c�����JF�a�`4�&U� `����Z5��C�у2��H,f�zQq�9�N�k��1�``�H\Asb�!L,����T�m�~U.E��|��5m'�)�R�1�w�{�:��տ0H'���gXQH��2��`j���}���]g��F-!�`@���!ވ��9g�u�O�.����{T3h=����5�7��Ie<ԿBZiu��cC��DF�2Y�54Q����h��Q?T���L$��KPG��J)�������9j_Z{��T�L�5>��^e��`��$)���ņ��[%25�:l��?Dk���$�D�f�\dT��$�hOEmB��}>��h�tn'����J8Ka"���gL|"��p�^�'�"x;b/�0~�&�7(W�[Ìh
*�aj1�U�OMܽ��?t�"t����|,����s����~��KM�Ɓ�,)�-��Y��N�q�P�B������[`�s��ؙ���DT,�;u�
�1�cx�R��N�#;�.��|�R��a@��Ť���n�NN�z�1'�cv=�o��Pv�ع��߭��('!��ǈaW�oJLU�
���8�#��(�#Qī���bo�k�bpf|,�L�%��+4W��!�R�������R>��.�ା��LƜ�A���?n�."�JmE+e�ȍ2��x�N �����
D����q�~�$ŶӠ�v^�X[/��3�Z�vKYPZ�7��
������e���*����IN�̓���	�RjM�H�?�`u{�ZE�A.6n6�,����;;��!A��-�m�h�������!�&���;� !�t�
I�Ps��3-88��y�T�=iթ)�~%�����̌������_o�������]eRw�-?��0|п�\�$uu�3j���j�K��g�琧�:�x������*�x��b%� �}�㢑[��u�`k�M"�]H�u���E�|V7h͈[E�JН/_��fe��ѥG�)ś���{��E[-ҝ4�s�һ��1��8�Q�BOY�֙-Z_�"����ɛ��?y)���a?�X/���:s"-��?�|8_i��#_�3J����[��`p4��	H�"�jޥtLv5h��m53�]պ�#�8��")>�kY�bF�C%����"H����cj�����.'�*���mD��0褵p7
�p��'�(x�֒R�y�ć]$@���:~�i9���zl}���&t��ߢ�����Ɣ8r�q	"c�(Ĳ,�j�l: --Bԁ��=�@� �a"������'�*�E�*�g��w��[J�����>���2G����A4ɡ��*ޙ!Hբܶbq��=���C@�~���Q�@9ɗ�	T���;zS�J�{�7��e�YH�/��,���؞��� ��� �}gcW@0+(+>e�Q(ge��9	ؓ�V��ψ���K�1�x�	��4F�O�i�Flݠ*���V
�16��y[�~��P?�A�I��j�� $��W��D��:Z�*C_l�Q����	Y�~ ����(
��Ŕ����k4���K�J��s�����U�S쩙BdL_ۘ���[8M���]�p�Q:���:��Z3ru�P�YFg��7�D;"���Q��b
�{�m�(�P�� ��V�C�J�+�|��:l����`�{������msJء.���=�3|2S������f��,Ӈw�;�%?$=��7�7>���};�@�o��Ŀ}��_�@@\3��x���Ђd���B�Kd0���HÅk�V`*9S�oӘI(��-zz��"���	?���n��i��n_�N�\o��N�0�<Na^gU��W������!���n�</M?�4yzxU�2�0��'���� MZ�@x�@Q�P]q\��c�x�jݹ�=���0���@ժ����̅���z�Ԏ�Eԫ��.�<���y��tʂ�Q������:]�`@(|�tG>R['�Y)W��u��K����HF��!b�3,W;G�%�8d��c�%a�\�w�p�����=ऩx�;�E�p$Vz9ɿ!Pԕ/�f4���"-E���?�N�����΃������}��3(V�}�^��'xg3%5G5i)N����������-ȟ����Vha�H``dbf�Ct��ED`f�C��"� m����L���H�]F	�n�0$���v�� �2r�'p���v�t�!����������ை�����7{#f:f:ZaW3gF"^n{CcN!�B|�x�Lm9��]\\�\��l�M���􌌴�n֎����� ��!d� �7�u4��&���7�qr�!"�'���Y�JK�7���?Y����Uߖ@�@oeE��3����3��l���l��F��F֎��
a����N���1�YY}�:|` �M����ܿQ`bfe�w����M�������?#�����l�_�q
� ��,O\���~NC��!��Wc��>�!�!;�-3�-�#- �����J���Q�h�꣇��ǀ���d�J��Чefef��ggf���g 0�22������ǩԷ��U��2��b34b�`bg�56be�e2��| 32q�0�L�����"6�V��if�obDokm�w��r�<D�t��#g��h�1��̬m\�gH���H�Q�� V6& ������������T��>��T �ߑ?�ǜ#�����N�o�F��6�J66�<D ����a��2�w��w4� e`d�d p2�)889YX��4�E�������K���p��f13��n���S�Fv�h��ii���_�����}g#C���[�}���7�� �33-�1#;-3;-�>+-;����>�ǿ�8�;���	�|����ǩ���?�����]L���A-��H`'������j-7�����K������>"!��������%�Q�%�Q�%�Q�%�W)���˔��G��qU���5�q͂0��{�y������VL����4����Q\Z� �3�U�� D\H@�u�ã�D������paw�����|�44�U"?X����Y7(�5D��494!by*3�S��(+zj��[bj�B�MM��A�0X�@i��$+��65�=3�cȩ��O6V�i{nS�Q��Q՗yo�xx� ��������DB����������K%����(0u���B+D�(��T�(H�(�3=�T)W~[���q}#OR���u)��-�O�������^�.==������S����뚻x�كЈA.UѸg�Ӯ�X�>��T�徊j�DSs�ܦ8T_�����p��eռ�8Y�Z��}������M��W�ŧ����+"LzC���F�|�ݫ��`qc�	.�H����J��o�V>�I/e%�ſ�	�ݲd׫P*}�8�T�'oJ_��*�%b��*P���Wm�54�8E�N�6t�9�%)k��ީ�}$�>S�aFW�d�m�����³;ܷ{�=1Y��8͐.,,,���J��$�u%)�>�A�H�܄��A�W�߈Յ��TO�7��n�rc�B�'b_�e��]�~/��S��l�������i��HDV�W (�'"��>�(><�b%��D��;�I��_�����x]�� @�A=��O���+�HbfuyY�[����"ʵ���i~��C���8����^ռ��$�(S��D�@��3�*����*�_K�a�o�$!B@��7 e����U�2hZ��^�ۀ�43��p��Z+��Q���H����p�zu�H*�F'���8��rZ(�������
������z�D:�M
Uw�� ]�0v�I&u�m���[�u7�AdET\���#4װ�z%ZVRޯ�|#����>�H�nur1)�U3M$�>[ �ȴr�&�{r�.�{2��!�*v�D&���q<��`k/L��${im�m������������A<ސL� �pǂ�R��v�ް�ੴgw�0�R�4�QB�@�Zti�d�0&��r\�����Y�pA�{HM�Ji
^�iX��&箼�c���D�֐�_���R�vG�z��z6�~�,����ﾓt�(�z�lVU����455=��|���^�����CHsp���,�ϗ!s��{$#�{>@���� �$����z8S��Oe����i�����>P� ˂:�7JHY�M1�����M'^/���ʍ�.;�}V�8�'-ù|�51/���%5����V���n@�y &}U]�s,&ݕf� " Y�Q�$��gI�#xĔm4ը�Ք���o�%SX;d��F�Mݱ��97B�ݚ4��x�C��x��^���.�b-��R���wa^�g�&�D��a�J��)��:\~͘ϠP��])��\����a�uvN��������]��rqq��7�W����0^���Ea���=/�!�>7�@�Vw<��Ѥ��2�����o��ڦ�t9D�u�ՠ�~�v����jG��������+��祡�΄Q�����m�i�/�#&v@�oצܴ���o�&ѠU����q_��Πf^l����g�6�(���~R~&-�Q�B�@��í�����....b�K��5��=o��x�tC��n�+��c��Q��(?hb�	~T��V4��hd�	��g�mlo�G7�,�Ud!X��Ő�� �8�&��rLZ|�~�uO�2����h�O��D���o���E���"�扃꼅=�gCL��EGJm�>Rf����.?���O�_7���<@.7mr	ѡ�>K�N������(9x*��L���z�ֻT9��e�]�������zm��A����#Kh�����9�����I*S]Eh׿�9�1;<V�.�����<�$���3��ۢs������c�M�]�DX���]��~���kR7B��!�����x��=}��)�� y2�}�`���]��VV�r�"�Y�'��VG_Ҙӑ��A�ՙtP��I��ZN��QVw�(JW��*I��Qn��,h!��n����4���;ƹ<��/,��(��.��l���A���L �}�)�9������I(ؘ]-ᾠQ����m�;��$��;�����77j٠F���t�zn6�Z.��P��a͟�*4��0��*�x�Kr|q1�x���6C�����6`g�PV�����d���@��N��E�Hy'����εo��Qj�6Iu��\�����;��%�������5�-� M�ȕ�`�wf9�x���L�T����Q)�@�~�i�����s��Q��3�)w^�k�88�ڽb-��j��0�Y�-�u8���HH�I�O��}��ӦEs�UY3D�
�a���IH��Ҏϔ]�Ϗ^���X�TӏA⳩E�:�+ŪgL���e>N;��\c���^��?�r{f���K/���(�ŋ�����奥nϯOâ���(c����l�����E�U���c�̔-ZQ��;���?�gܬ@����ʐRa��W1��3S!�H;8�X:鞯f#p�"wٱ�>� z�ۇ� X��#�:���������9s|�OF�n�e-�=G�B���0)+c�h�s7�T���HZ�U5
q�&������R̳�-M�;U����_�Lk����Xt�K�3�	����@&y|F�x<�?��,���n��A,����T�������v�P6�����j��Tx?	e_�g�D@z?�ڃ����C�׭F�<D��M�Z
C��cQ�Cǥ�G�ti
U��7y�"���Ib�@?�OU��fv�lޟ��&���{)>O)���F����g�k2��/V��NF�ej^>,&�1��FXd�Z�t�<Cc+hU�n:7]E�����W6�☄e7�Z�UI9���ݽ=�f*�7s1= (��;�`�[VTV~�t؇��{���_���~��
�KC̡��B��,E���of�����e�X�aȝ�����>ym�:]d�>���1��4���z��&�ψuZ	ߗ�R�]��^�t	ӂ*�=���1a;R����>R�k��������IS��=8]���E	�Ɂ�!	Ӆ��V����s��tA0v-B�S�:��rRx`��l�e�����m޾ڱ��\/�Q=u��9o|o� P�䘬���HO��du����%��O�����#�����}մu�U?���Ər������o�vؕ�>xr�ɶ�ze�9�R�=1��-4-�Y�VП!P�Ѽ��Y�c� ��v�����U�+�o����ޅWHۑ�	:A��Q�Q�V�-C���Ion�������r\j�_H�X䪘8)�ٸ�@�[�T���;�Ϝg0aYL90>6�[k啇6p��u���"W	��-�~��RM*^�����t^ܞ���#��#n$����������N�h�w]o���!F����(�b͍��-O���;o���9�����"X`�p0A��bB�υI{���`�H*�'P5(P{�l��M(��`*i<��:F�OEGn^�Nӿ��+�_ۺ�w%ȆS e�������V��<���X��=��a�)�e�wv��I6��o��&\�o�b�3��ż��C|��=/�ݬLUY�v׸�,��z�ɏ�������siF�i�JD�<����� a�F9hX��i	��2/��Zs&!�	)-��<&�dy��MB��ԑ�zE��ڽ31�
�
J�i�����2���%�P�6���׻��[�z5��;'w������%2|�����bZ��ܣ��R�Jw��4��@%���xI��zO��4���O0��B,�'׾�a���A�������G�����;�|C)F��`!��Ե<�hd�(dA���5�h�@~�+��'䢒A4� ZA9�U�hX�5��ޙh�#nbK�.*����D[�X�X
�^��r� ��&�� ��MJpH�6�g<��KeZZ��,����b(������L��+��0�%~T~%Є���E���1�d��Cf�;�QY�]�f�Z�ˎ�ӎy��/��̻FA�yS$CaM	�Я��kgyݫ;;;/--m=�\ b�%�T��SM�>��@�B�8�V�&!n�Iǵ/�d�*�B��@�fz:g�������p~P�d�Ί��,bh̆kP(��QG�.W��W�����d���x6��K��a}�o�Ih�;_-����rަc��f�ҡ"3�ʑ�-�0>�nk���M~]��J�vf�@�R�Q8��|@9J�{�r�ډ�f;@��hR�y�P�L�x8�|F���?���NG��7��������������6D��V;���} RQC��(��/�3#����tY$ֵH�B��,���J{��5��cq��yq��Dj�u�������o�L+��%1cO\��Ĕ[WhV�����,��(C7�Z1�0Z���M�r?�2Y�;��B�E�)�WSSU�9�R���Ԉ�V���=�ak�;M�l��7皘�h�П|�������ks����R��]y�G�M">��+��?&�X��.�
���ǥҰ2��&��k�3�Zۿ�zz�������s�q�����}�8��K�f]�h<XnF�NFT�¸��iZ�oSC�,��Z����L�<����2ѝ7"̺X�����I]�@���)�Lѵ�<w�$@�������L�Mf3�����#���ﹺ�>"J;�����3f�;� &����3q���vB{>Q�6�H`�$?2c��[�̤�Ծ�癒!*�[���ެ��b�6tC�4fB�Qi�D��8͗v�̇HE���k�?w1WنMR�9C7�4�=� �۾i7�U�]\
�R"�ʬ��;H(�؎�(Fl���Qθ۵d-<~;��{�vT��t��g�:&Lt5�,vm�/@���ml~K�E�`�z���������� M��
��61{���_\��߷�*�����fљ@Q�5�EQ��/�I�Ҍ�k����x5?o�����o}}�d1:�i�@uzm7	^�Q���r�p�|aY=������`s6F���P�q��g]��/�l3��3���F�k�b>��D����M�Ƿ!n���/�Hw�9]����5Ry���^�9��V�Qdժ��8N$��=ߝ|�؋w���A��ߦ��[���_�)���(�)�ЦMHb5�z�g=�r�q3��3
w��׻O�eW,�����Y���V�:� ���.�����_=���4	L+�����$���M����z�� }�5p�df���U�lZ�Fٜ�� m�Qz5�?%��X���GWnM�p��];<�":
���Z��^;�F05�o�e���A�ey�ғ骗r�
ٲ���e��w��L�r{��<�\ABp�oK�ic+c	�1��ܣduғ���7:����ל�ő"����IHF��k�̦��2��GR��[Peu�g�]��-��<	����hP?NO0�N�q���NMR+�J�
ɏa���u6�賨���h�\�~0ϯ�φ�g)�^<����P�����1����?C��zSڄ�*i.���[2������I�	̺���Z�4���3#j�[��]N0lOYD��,p������۲��Ĝ�#I�H�	�\�nV�)Y�a3�g��%�D��݂gh0!��H�!���Md�
]U��٣�+1�4hg����a�"��d4����cO��j��l�L+�2 K���q��в�Xe"�*3F�+N����Վ��_E6��]L�K��*И�I}��d [��_��Ebv�H�QY��(W�>��fH� y���Ջ���4|��V=f:GLhx�[M�@�HѮK���k���*�4o�J���Ob��\eb'�^	�V��S/V`����p���e�It�%J���L-=�QE� �Jײ�����^Å��нI\f,���ز���l��A4K���1Cb��T""U�?s�(����2�õ�t#�{�Ȃ`c`����*�5X�5+� 5`��X�����D�HGXՈ��k��6�*�k�j�\z��B��T�
�Jyf���	_���t�8�Y�������D۴�3o����;��b8!,��LAN��m��N���,����9ʖ%F�
7���ܶ���lE�~��X�j�x
�\�04B��U�IR9FA��;J��Qd��$r5m\(� �yb8���L)�vf&�+�n�Z��:�B!5,<�0�$*�M��c�4 �V��S����a�U�얽�fZ����#��ǻ6?�(�(O��}q8�Læڕ{���v�����ݥ�`4�v�1|��^I	���x|����#gf^j���3��qX�b�t�AY��	i��3ʉF3��K�&$�D�L�mޚ��"��@"L��+\J��Ue��0z�i�NG�T�9�@�m����y���ET�*���$�+NI_Q�������/�(bᇠ���Mr��1?��>ke��W�m�셸"9d��Y{ �)��$X�*����Eʰ\	��+�p�M|���A�@��B^�Aj%Ҋ��ѯR��_���ú˳��o���ERB	����+Y�%p��U�&[A���F�e�$�IV���E�J3@1Qv�A#b�G���u�sA�yU���Cͽ�������o0]/s<� #ǥ�W�T�t��rNK�|q+/*Q����$7#�)���m�2�&�v�e�r��0{&��-�'S"�s\� )n6���� T�)�
J~0|�T�yu ճH��g�*"Mgy.�b�W_�Ms�z��,B���F�%ع�`�G"P���E�M�^���|i�Gjgc�q%b?}��QҍS�T�h���pj��0|�����^T�&�Ð�ٌ,���'6c�"oh@U�~{��Sr��Qa�Mڕ�w Q���(�ZHiEr�%k�����dhu��SL�.�&?n�i�T�k�-%�z��2cuR����]���_�	i -���n�0���:.L�R�_dүß!�=�;ѫ�~�3�8�c=m^15oKoܧcd������_B^�p ��V4������1~����p�&�tX9c�G�ml�^�_�N1��]�khP��=?��ێ�)��߶NWu2��~���EЩ�\z\�Ќ���c�,�;ĭ5�n-PdWS��nY_a�ll��G~K�&�cЫ��V۽	z�s<o����xӐ�g�m�L����-��}"/e��+���3����Uϐ�Wꯤ��F�f�Fr����%G�(���:��Re�����,-����}�ÇfS�lĎ?E��"|�9��p���1hɁ���]ͫ�&H��&�Ky*8�]��BU�E9�$��M3���7w������Q�C�eNl�ӵK��~�(%��M�H�}(w�/f������K��kO�P��_*F�g��H($UFt��]��"��o�_|?2`��ynsi���z�<��\8������O<I���EL���3ŉ�b��[o�7bŠ��fʄX��r���������`x,��������0�����Un�{4��˙�R�r��Ap7����ps�4۴aG�ּq����}v/�9���߂��m04�J����N�C>\>0R�.��|����wu�!6�<�9?XD׼��
�+�G�һ�M���j��\�2�ǚ����y�JAN��07����m�.һK�f��~ل��\K�^�[�9��U�s[  �GO�=�-����Ц)��6udǛ��d��R�;/�R�h�0Mc��J�P)Q��	*� ��_���\��r{��Z6z�{�M�D\=���
v��,M������[@�K#L���+N *b�I�+]�`�ަ#v�e���AԞ��[����M�g��)
g���t���]�� ��.2mb��8���`�Q,��3G�o7n�F'9%e�Ie?�1,�'~oψ��T������N����swsKS�{9<�QC�b��f���|a��ʼ�NGK!oV-qP�`1�_,Ku\�L��viY��2��(w���vjJ�kg��)@l�̅���kP у<*�#fٷ�]�g��N]�����)����0,�țۤ�?�w��D$C�^Ǝ�z�<f�7>���������y�0	 ��\>/h�st�,������������qu��O�$���h��l0acO�ƶ�hb۶�4��ƞ��;������9��g�uc��Q��5�Kw��=���p<�j�W����5�\�&x�^QQ�}ve������p�]���A���M�c	��w���Ў�,!/�.��+��p�&LTJ�K�E-���<`��3�@F���ڿ�`�a5�*��#o��h���v�H
.�\�hMS?&*ϒ}��B�hX�T�<����^�}�� �.�E5�J.����q���ə�X�@�/�2$�nXF��#a�Z~$[:���Ю#_Ǵ����@�l����T;'���/珜��ʣ��8L�U�wS����O?�x��,;uE��=���DK�W
�JĬ�DBBB���;ħb~/�b��i��p4wK^�K������Fnn-:M/� ����Ƒ*r�x�ɰ����h�O;�r��`RY@z�M<�.�	������g�R?��N�E����a��K�?���8�UmR����*u�a�~�����%�xP!w}��t�\E�E�g"�6�dp���{����75!;d��T��mL6�N���ճ�D
��x�hb�!��[�i���b-�y�&�cl��딧��d
�{�h�ܟ�J��R�|և��K�n�z��&T�&3��-�4��w��	�fB����-I�����+*D�Z[��LeC/l�VVv������hx���df/�#f�����:k��e��-���~O6�6�It�Q2ohlTTD��^�4���1 I&߃�Y�l��!��c�'ss�lx�q�ݛ���˳D9%:�������Vl\bĵ[�5җ7�),M_�����TrC$�͔٢�r�A�8aO4���t(A99)�̵�j8*
%�����%Te���M8�3�V��7��𛳴P�^�Y�܆��[�N�ǻ�cW��A wO��8���Ѽ�e�޿Ƨ��^C^�����+�	b���~4�	���_��>�����?ϥ��ؖ�J�7�����vjֶ��ܱ1h��5�~:-s���F���Yg�ϻ�>^o2y�~AF�����gt rz}t���5����v��~�I#��:�UZ���S�ΪU+ރO~��R|����ƚ(��h��<*�Pmc� ���
�3a�-ؙGSD#����]���w�&�`m���=���1��,��.�����V���c����h;N��?;����-R�������Ţ �D���yuu��y>�/��b�H���=o�o��U���#��Wj�������Ii���P�y�Uv�!�1r���	���Ǒ�����r}}}��������������$�Ͱ���������t�夝o�X(�U�[g��S���b�/�����?����kk{��b��Ḡn�nҗ�?�n�b��ݺo�:���G%9	9�To�9 �A	?��o>�w�����1��+��!����	�4�B�����nW{�W2�d����u}����D[:>�,��'�^�x��c��8���c�ᑦm�������n��}�I3�i����&�OI�Z�V�e�k��O�U멉� ��@�]�5���� B�qa�Ә7.�`��K�{Qtm���66W�	;\t=@�;�>����w�]��<�QR��Ѥ��-'�7E!�<�T�ZC��?���n����9����a�����8�F�y�gc�xѲ��A�eU�J�eu����3@���\������뤚ZHqo��~K��/��]ڶ�C�B�l�B$�[PC�l\ ���uG�K��H�+����{[����B�&�}� ��d��Cm�Y�v�0�nׅ�̫�Fs^��%��]o<t���LC�8�mZ����f K��q7���+ƭ�%TI�
���49���%�'�p�;4���o����l�9o�����l��9�V|���'Ҿy�7� $��*1[��ȅ���������W���ϳt�(Ix��ֆ�lQ���9Y5��`]�_hO׸�p�!�����bkV��4@R��|��6F�7�q�I�TO~ש�k������%Sfxg �|z���6Offf������K*v=m>�n�������RD&����<;/|.��{��-���m[ƽ��!)�o�Ї�p�.�66/��帓�w!���E��P�o;�O�7߄�Gh�*z���YUˆL<��%)]��$��D���%�&H�?�����伷��wf%I�!�!��(�v3���v�A�E|���������~9߅��mÃ�m�޳�(L���TQS��C�s�3��J7��G�玮ܵd�NMb����Q����h��@&�FA��HV�+"/�2��|���ĥ�2������l�&�b|@*%��E&������|l��z�䤜�m{��ypb�-�O]�t�bx�����n������6ZJv.�Uw�ߍ�;���ɿ ^���/��vݩ��%-�C�
$A�Y��s���a/�r���7�o(����뛝�HF&&�M��Yۖ�p7�*i�}}����|��X��Jr��W�,S)yܘ���O���B��G�e��fIއ?�U���o��v��q*�txܲ3��2�Ѯ��I?�6��U^�(s�(59�k�3c���ٳ���<�?9][^���v��vF4���O�9��w��wK��ЗOܺ��F���?| �6S��9A�-(j�n�wI�5�|���p�{
�?ޒ�J����"Z╎�OT�������p��]�㐴+��Ь���B	;���WG���?�3|lj�돣<��>��lx]�k+(y�xd�T}"��FKNOOU6nX>����`��\c}Ҟ秙R�{Msw�n)��� r�6�)�Ъ8!�Tb�������ق$*��5<??���'�-��Ǹ�k$sq=>/�L�S��H��)��~9���t��d,��m4�T�\x��ᣆ�&<O(�.(8�уY�r��KH_��&�3~W��y�������>��a���g���X�{��%��!0����U:9P����cP�&w]w�s����A������C6oxmq�vF�o..�1u�k��p�h��u^M���V���1�++i#���z]� ��"aإ�=\,e����x��v^S��W	��m�&T��-=�5oϒ�_.�,�B�f,���������]f��N~�7٤�ͫv4���DZ�b�ƽV��p��N�${n�>o'�9)h���'I�}�M��_�dB-�@ځ=�?�o4ؚ�+k����Gؿ)|�SߊRQ�7��U�����5�@�n6f�����M�-������O��[f����/�rY��K��]B1]�|6�^�vH�~��8(����gx��Z:G�:������7n
.z��Ȓ��;�a���nP�� �S���㒰�T�� �'pN��	y��kReU�ͤ�Od(�/>��t���[��ϱJ�}S�~օ7͙�"��m"W��m; =���Z%q�)�/JC0'�0���C3�T�zi:��h�E�m�j,uE6F?.�ٲ}%� �M(���ꍹm��f�qĻ�+jhū����B��@� �q���Mt���o�~�n�4/)=I�ta�YCd�� 5�����)\�d{_ۍ#*oޞg70�܄�=J��t����[��_�8k��K���g���vZ%nq:����~�&������I�]--4����	#}0V�����Q�*}H-��d��m��tД��1�E��0�X�����*��:,����5���<<�������mѫ��{�2z����|��o-|_Z�2�%ޠ��UN��_\�;Gd}vn�4I+Ǫ55�;�����d!B��0PX����Y�9�7&y�F>�bVH�;�5xf����	,���9�?~�`���֑��g� OO�!����-*Y�1���f|��kq)t2�!i�jN�zIJ�2� FR~G�׍�8<�jL@�
ۯV?��4�2�xE@ȸ睧N����ܺ.�)[̩l�k7ѕ�:�2��W��ysl�(~�Pn0U�*��R`z��my:MՆ�d��ȵc��o�K�Ƽq:�o���G4��JY$d�DY9���=���ܖ74�؅�H��l��u�j!nhj�_�e��c�-vz��`�k�*����ֲ�������a%bH-k y'�ф��k��*5�rJ�G���.@)�#��ɻ��e�ʶ��3���4B���#��!�ʿ6��6J��T_2��JW N��=�F�{�7�J���@�Rf*�΄J��������D���K��df��Փ6yNC�J_�_�D�c�tA$���aȠym_�G�1�4�
/\�q���Q�q���+jP�o��u
��>޻TגKͤC�&�_��Jؼ5�3%�T�}���q���ݿK��b�����kf�bO��BxZ9�D8dc��,`	Ef�\�vD8"�	o�a{��ܿ�Bܱ���`�;�F��[q^����խ�ԢZZ�h�XrF�b9_���'1�7_0g ���<������~�T��f�0lڈ���X)�a��.��ɰ�ӕxqj���h�'Z������Z{_d_������lCvW`1��b�2_�4�`\��)�O�~��`�����7��#��'�M�aMII	WS�sg�S5	�W���vk �O"����U� D*>��I"�5���z�K���r�ku�P�d�=�~r?���<[�;�<�HḾ��k#]��>�D�C>�EA-�n��g��*���б������#؟�a�E4���DT݃WLhDW���ӣ�����9�*�qm�+GÍ�kV�R��Eḋ���F�ek�
Vm�F���5�U���^>�*�w�����Ge�	����N(�����2�6e����l[dmkƾ�#+�`@L�K�na���z��W�mv��g�ު+>+If���x�:���޶��f*_����g�9�!ꭠU�<����~0u�T#��s�_{�D��4�# �	������XE!��y(�J� a���j�躇9PŎ�ܘ�UЊ�S���i��Y�S�))�ϜQ�ϺO�ȆS"�=� \Q�|��6k E�?�N��G��H������ cXr{�[�ò�-Ċ�/1QR��\�Es��rcs�Z�|)��{=����-v�v`����g�ĕ����Rk����r*U��q���ex��g: �_-�$-a�g=�h	���ȥ��T�[�(5��15��"��M���ؗ�7�(0�Z7�+�hŵ�yG�prB��z\H
NB����ԩZ5���u-l��)�6�.���c���l�ߨ�m��Z$��+�T����Ň�bb�h�ʖ�����P�0�u?U"�Frڊ&�fe$����B�h�n�N�%��N)-	y �8eZX>��R�s��`�36��C6sB@k+T�P+U��d'�݃�m�Z$�N�"��`��!�(T1�$'�]�* �I@M��$f�Nm��[��&��|�Ă��n_���7/R

_����c����	8Ӻ����P0н�G��̼���񬿡�8YNr*R!Ɯw��Г=j�$�� ��x @����&�Y�/Bվ��������I���>b4���7��D�%���m���+�"O���L6j�X����7Ԫ����t�^!�2�$�ǎoa[�I����'L�L%o��M�X�rX���}��`Q�A�"'��u���+`:��Y%vrρ����Xr�+�2f��iG`tE��aUNG��|�U%�Ac�z+����h{�"YN�z����'y�Q�V�1���)�NU�_����ZDࠑ��;���e�j���s�a���Q �`@&NQ!㸹[���
�X%�Z����Q5� X�T��a�!�d��o���*�͚"3��#����76���WTP�����G��d�W4�7���Ц���2������6..�Y_�����j���=wf��.�5mf��)84�b��}��"������l�B�G�*��yv��͂��zo�wBv� .[GQ��QY���͵�䦽#��0#�Ot���	�ߕN��ftN�z�r�~�ID��}u\mJ�����r�}�6��2,9�a���|�e��V�l�'C�Q6�;r2=4�#���y���Tx*wUm��ٕ���\FFD�f$�tt�����0f�x>�w�0-������V�+�rw_��n��n�8e�BCc�
����o^ۻ���c�G�!Y(
��)���F9��nQ�?�3W��VǓE	K��v��H�=���$"�,P��iMBUO�o�o�qMB����Aq���2w �%N�` �tFg��b�����1�s�� ��<j�t�][�7������:��6��P�,f��ö���%�~j)�57Rh$R!�k���MY���Ed����g���
ӎ�䩠��5�3�ly��kB��Q���m������Č�d}_��O�p��]�s�7%r��&�"Ȉ�3��0����p�h�I����z6��� �p����.�6'cXU�2��e�1G�Db�Y�	UE�}e��Yd�����$�,;WV{�� %� Ǎ!�=�0�'4%�sl�2L��Ʀ�P��}���o���{�^�U6��-���g�Ѱ��.{�0&oR�R�4�8f�j�h6����d�5H�׶��B̺��6H��9�?"�*=߲e�2�.p���";�b�U�����g���#���x: �Ɔ��*���^˨��Rs�e ��ԭ�t�Y+�2��j�B�Ƃ��n�٤篹���Ks�bG ��YCJ���A��@��ˏ�ӓ�� !J�-J/MEŎK�@[�(ΐֽ�U=�����B�^o�C��~���h<�Q�#�:��h�vTg�u�M�}lDÑ�Y{��;_���K3���#�3=ޝ	�'n2���q	���N�4��`6V��CnkL�@�ɌQ��k߾��]��X�Q�
�q�Y�  �	�� 9	J  �+O=�:{�&oܒ�ڳ�SD�5�g2Y�ޙo9��^�>�ok�]z��Z������*�� �\6qQCD�y|7"�9DP�ޠoc����zD[ޮ{�_}[�)J<2���ݴ��-���2�%`�zƶ�;;I̺���h�0���܀�+ ���{�つc�O�w=����V3P>���'K�G�2��NyF���11)	Ƕm?9�us��Z�v�*�]��e��ٝ?W+����w��FA�\����u�TQ��YX�"��G��Qw�o�ńz���(19����	>K@����W�O|ƥM"�A�1�5LCDv�-��,0ԓ(�5ñ��D�cE�6�0m�B�C�4���B��[���S����匑�֧��t˘|ǵ�}��#���\��36Ә7�l&��s[���id��]Gʘ;����4X���h������SӍ���(��q�mn���^s0����jjn-�=29{���/x�T�.]8��e�/�|^���zX���\�2 �:G�n���ח~_���_�4a���G��o3+g��'�gC�?�y�Ki������'��c�3pL*�6�E�	�/>-8b�����4��֫;T��j���nPHg�^����I���D��e1Ѭ���\m��.K�d ����ŲS�P�&B�[�]�:��L�>�0�4�
�Ho�փz愘Di�?����w��|�%�}��OaHSz%|�g��R~�w���jLu��� *��y0���o�`s����c����*�H��D���P��Gw�Ƞ�u[��In��+��͹*=��P�<�$�4�HQ��+�ݸ��h��@��C�-����k�z�\�9牮��������Md86��'dRU)���z��������}37mt���~����ꦵ��S�э����F��*u�����ֲ*DrJ_�;�	�@�H�t�N�6f_�J�C'߇��� ���SP|��^��d�y�$>�TK5و�455��9e�a����<$J:F̭���,u�8��s���7Í$
`�a���J$��[���f�"մ�.���55r�M`����߷D�i>�?���w��-h��l��ځR�_s��
#���)A�{��1��R��Zqn��;e�j��屃�DM�8u\
�Ҵl�#sw�C���o�9wUr;<?9��Ifы��g��U;�z?�Ę`�S�̦I l#$�U����L|��|�:W���ۢ���4�*��+{bޮ=%�(�B�pq�ੵ4���.n�>���=��i�16RK߃J|3��FeK#$� _>���X{��C����F��)\���v ��H�Q�@�Hb�X�r2-�t�h�Ec����S�-���>,KD�?������1��]�3�=�p*�t��躆�1G�4qQa�O�xP�q|�q%�sC*A�$��!Q���"��A��+W��/	��{�_Y���a��3�{i���~���C�y(�A�d6�&I%��u��ԱŊ�)o�§M��傴���i�Q���`��X���J�8R�:��Ƴ9|�X��i%�i��[�2	�?ܦ�Z���&�޾����J�zO�l����6D2��Fw���H�Q���9zئ8EA2tf%1�C>ؓ"�]YҺ���8|�b���Ҫ���L�]E�mn�S3C�E���#��Z+�b�-�SiT
�IB�ۥà�,���`�Q����Â�s�L�j�0Q;�O�#�M�{����+���Y�M�[���Cf��y��dQ`�U%H�@��}~����1��O2j��ڱ���p�ɘjH��5��+�u�����_(��u1�M�,^��y�;�(���
!�V\�=,�<.��Q������<�B4I	C4��ӒͶ����^�rFJ��Ey_�� 5kڍ���x/��~Cox��oϽ�A�S		���9̶e���$���G��� *ܧ�%�U��N��5������M���+O˦/��T<U}j[��������Z||%I?�T�.�!�L����Z��S�I�CO�$�.ya�ԗ��v����RMG���S ���p�6��\�W\k�Arە��ޗ �B��SunΒ�����Y��#��R��R*pﻸR��!w��F��y]ck�,�l[�H��R�yE�EQ�|��T�O�}֎�tq���s4^��F ���2�Zd�B� 1��V�|�]nn]v���{p:�B��u4��6���C �y9U5�@ �Oh�Yo^�k퓚ͺ3Ĩ��6���?+�e|�Ev��]W>�b�vs�q�.j	�J*���#���Ƶ55<<�Uړ��y� �SVޜ&�"��-�6���a����KJ'[��?Tv�q�N|�r�,���apQ#}|,ۄ��x�?Ih7�W��u� G&�$7)�x�d�PC�u�n�@s��(3�F����|Pxƕ�!��P�1���]4ȏo�c��#ƾ���B�s���Mwf*9��ҺJA@���_G�[��s`�c]���H�y�ں����;@̍�h>�����*��|�����l�����t�㣺�l��*�U'8��[t�}�	�7�	X1�.�%K�K�i�ӕ��\�ur�S�8P�'iA��l�G�N9����tGd�;AJ�����{nK���J)��f��/٠?�0�|�q�plQYF]]}̾��&��T����j1�����V`�6'*
�כ�s���1��ЋKYxA���+)\g�yJ�G�V�П0�j�F;��~U�p"r[s}K�E3�`ZL��B�� �s+�khƍ�5��A����4L�m�NY$�1���)��`��c鹥��Y~�ŵ524�aƸ�8qvs��꼿�3s���\mW�)�~�9XG9�x�,9Eڞ$&c\��5���2x|��_8>���t., ��>��6�Qۜ1T,u���%g%��������n��T m��1K���bAd,G3����x���Z��ܻ�b]���R�eӠ3��Ed�O�2_��� ���M�<\����2܂_$�P.��_p���$R�2���b����M�0������~���U&ˇ'�>s-�dL��,L�X�V�<�#���K�{��"<��L�D��q��H(�_��`J�\f��E)�X��Q0��R?���~�I�3;�Ș�w�YI�LP��(�hX����>A继��0�FB#��9L�q�om7�=~����*y��`Qog��F5k��c!�y:�}�Ԛ�������U�`���q����}z�6��^��yx�M����h��D�w���E�9{���
�.�|���5�U:�e�|� �R�Wx����B�	��n��-�
�ay'�#O*�U�[�:{����85����ig]-���s�m�4�4��e�()���ꑑ�׫�+���,�F��CK~ez���u��3�َT:@�X���F�2j"(1�A���|�mr��lq����x5��I��(�y�΋j���@����D`�b�w'\�jM��<��sN�tGww��b]�$Q�)�Ά��/�����+�1�+���\e#��;J����f+ڽ��q�[~��"�����o�A<��_E�������F�A�C?ѲI��[As�m��� &������Q���
>�Ns�/���'M44�N������࿐i���T�ZY�/�Ǳ�}컽��Hz~w.äbm Q,j������K�gѵ�Q�����ݻ����?���/Mu�|�,ݡ�_��)����ڠ��g�T欔KPBD�~2��G��̙S�QRͥ�����\
���������,������`�`b9�]��=��|�y�9���mO]�L�{��`�����]��s�vmYL�A�z�0p6`Gx_�� �!~�/��o���p�e�}>����O
�%J������0�U٪MU�V�{@����͵�߹%�.����|8�K�����q���,3C���`��C0��'"3-��/���"����Ԍc�&���hRx�T������w��,�L��(G�����BT (e�Nϯ��'�#e�G�lLq��wR\�Fԛ����g*.�SI�Z�/6w�g�,�����C��g��X��S���z�<�WI�v84n�h/χ��㈠P���n�v�[V�����3g���nr]~ˇ��I���B2�k�úqls	2� �V/!Pɩ��������^W�g,d�nۇ���o�1� �x&�SY��rY_�8��� kH�T��w�¶ӱk�za|��3�>͓��w\�.s\`ܛ}x�(�,�=v:��������ՎR��jIg�HiSPk��U[O�K�܏�D쐝N���]�z��0$�w�]��Ԍ�&�NeNy�-�-�|�����`�.��0�S���Z;70��+��}��^xp��[7&�#��Z!\�,���V$^<Z )��f)B��wf\���L�����@n���Xi�U�y��ێ�`�0�z� Bj�s1(�ǡ`��V�.��(�/V�Q�s���(�����4�e-�6;����v7�hF��')�\�	��Ϛ�e0���FU[�3���x�$�t����ꪣV�e��B=ޞ�lT
��֠���V�u�o���*loW�Ĳ�N��5(�tҜ��/m�˚��|�D9�����t�����^��R��"#�5��������>�_�*	ѷ,�_]��Ɖ��1�q	'�@s�����,�Tԃ�5Mh�P0�i$���	-D0=r�@�u�"˜sſ���g�n	Y�"ou���Z�pl0�V��ʼ�:���>V����O�����0԰Z�X�B+�R�J��	�͜M6��U��*AKr��Yn����
�2�-�*�,	XH�9����Ĥɗ�A<��D����i����Z�bOy�D�BQ��.��Z\��U�o���Smٸ�N�ȥ��������Y&t�ᢡN�2OJ%3�5ʶ�_���QK<�%��u�(q�����#��1� )R�W����o�c����ɬ4aL�<�*6����@���+�v���A��M ۯz�I��pL�f��d��e��Q����8lB�gЮ�g8�ľl4o�<򲸈�"�����1�<���ji	�X7T�)b2��:��Xz����]!
9ݬ�<=V|��ǝH�?�]ps�[�J&k�_�L��*�e���D��d��4�N��7/�ȡd���M>(��`��;:����G���~�OV|t ���.����$X-l�TD�q.�$-�wL�3I��_P?e����@I�sz�@�)8��dY�F����:B�U���I�Ʉ���}O7iE���3M'9.�w�\>�W�QQ��	W�c�����P -G��\��~�nޟ�2Ƿ0���;���'e�����ː%QM�I��Lڭ��y��������N5����N�p��ے&�Ś���P0H��|��l�~|z=����O�k���Pn#�i\p	Gs���c��iB�O��%�^6g�P����w�rx�����B��|'l_/�Y�kA��p��ƃ�?"��ǡ�DIA�U�5�dp�a��_&��%����qۈH�6�!Kɜ ,��	}g�����%&H��}�lI!I71k]G^rƠ�f�#\t�&r9�������|Ʋ���.�V̪-Ǿ�͙H*��\��R���W�ל�ѐt���egBG��1���q�\�Y��y������%����!$�Ԕd�ĈQq�
L�|;�������zFdѽ��� ��ܮB���oi��j^@'�L���+0D�2��3'��{^z-� 6p;�јhX� ���e���;H�ZQp��C}�V�߫����
%��6rZZcs�0��5(2�4��V��\Y~z�A��M�?~:�UnE��}��ڈd��"��۶D�x7#T�Zwu�?�Ed�
��L�}�F�Vg�U�52ʒ{�罸R��2������zo�9��R����G�A����)�ȁ�m>���kԍ��/�*���E����I$�E��v�Ϫ�������oGͶY+�6�kQ� k�${>���M��M>O����Ң�*CES<aJ�<�r!b0�
e!TmE +am���	���GP,��4��&��#n�#s�tv!�/�*ܳ��~�o'���+e�(b�ۄ���睩�<����GC<Y���yT�!��o�k�����AdDa�p��o���MǋT�NW<]�G�������e�V�.����U�<NMR���X��k�ݑ\�o�<��*.r�m�,���BLJ��j�vb�Q\�������^K�o����Y��|��A��q�MS-�;�X��aP�w�j-����Úײ�n�p-��񽇍8{�'�1|l����roq�s����P�hE��dZ@�@��h�pG��
���B}��԰I|*����	b�Z��&�H�g���ĮՏ���$$�+��*�����2ۊ�G��LJ��(*�U	7r
o
���S+5V*�p��L�w�P�����d�UT�ڶ�bb0�c.��R�Ғ�H}]�/�#�E̓X`Bp^rn���%�{������Y��n~<�=m3��ݙm��S�&ۧ/>5qz_�5����挈~�_�����g]�gv���D�Փ��M4���=r��=N���8��/�����������ꗝ�ŧ�9�ҧ��ʿ�B�ڗrM>cΦ=��t�Rҁ΂��Op'�-��o�mSQ��'�95�%�Y��y�$�QI�Ͳ\��'����](�8����?2GD=r��K ���Fv�a�In����Q�X�DB�Ŋ�a>�\�ȒȢ��E���?�S6X���Vqf[��rHm�F��FU�e~]9)������YQ}֩�K�@� ˣFP�����Y��j��;1�D���;$pm��������b*)��N�ie;7>ƶQ�PY-4Xx x$!!���+���kXT��&��_�O"� �t�1d\�d�%�.�˧���������u�[>fƧ[;˲��H������C��(�B�9�h�d��6뼹����{:�|8_IP��{�Pâ�޷ݼq���DMs��������ǲL���J�LTz�d㒋�P�N�x�[��!/-�w2F5���r��]I��'�;�(��*���ɑ�אm�,�,���릐d��Y>��W���3қP_��oTg�g��m7sr�g}�켿�w��zH���P={��%�t�8ьɓBG`�=�̰�=~�z��]<�)R4��`�=��uZ�N)��ن'$ɰ](D��Ȼ#�D�0�aN���RM�Z2�'� <~d�H���=�=�Hi�[&��;�gQ��@��P�ƕ;�~"بw�y��*�	TZs��h� ��JL��T���'��\G�T���DF����^�tv�3������	u��"o��Zgݰ����s�R�t�;;��VSMτ��������a��s<>c�_F��������d���:�\u�d��+��׼�&�(spŁ��f�("(���y���ݺ�ݘ+�e]�_|�i�x��	��t�t���8m�eŊ�f;j-ܗ�n�
��9~����g�<�2�AC7N�W�dyςܗvߖ����n(����6u5����]��=�E�,OP�����.q������Ă*@�v�m�\� �^<!�s�Ã��>XD؈--�иY:��^y��WK>{Fc�$l𵹪�w��
�����Ǜ�y��Z%�d��)naW��̟��R	uUa��[d7d��9&��0��"@]W���;u5uߝ	�K�����b�)ѭ's�E�.^��U�f�z�z�������ѫY�H4�����C�}y���=C�ӎ���&�����l�_:��h,}�������t���(2��|39�Xp��)��~!o/���K+�Y�sr��=�ދ��~���5ˤ絻����C�`7:�9�,)X�V��{oǌ2&"�R"�]z�|:���D�M����;�c�'(�o֕��_��������Љp��t,Ӫ�r��B��(�����ZQ�(]���J]j�=De�ލ��(nvp���v�ƿ7�X�����R�{��D۲�ZMF!�Z��G�L�9���I6���1��&4��G�$�csu%=�rO�D���>�$\&�7)�dZ�LP#��ciyC/�ތ�
�w�J�^MX_-���->N$ G��W*��pk��;*a��~��V��&@;�a�:�«�hxM-PY��M�	�#�<�p�v�j��2͛=��/��Nd���~�D��hL�؆�����.>JY�����j�{��%G�o��yꉛ�a�U�W�ܯ&B+���xu����{�����[AV��d�i��/�����[ Gm���Q�m~�����/�jҧ��;�wK+;<�m�_[�>�ي����7fu�d����]zs�<�����U�����n�V������.�i��s4���D��V�����W�p>m*FJ��Ƙ�Z[q��D�tC�୙� N8�OR��'�qg��ej&�M��݋D�{.���SU�J.�I��x�(�]e�d�swN�MK��^]tM�O�Șox������������	�?�Rx��_ߦ}%�GF���/��.��AGw0�Q�L1��E����q.��z��jI
�~�XQ�\"�:�W{N�u��Bl���t+�rn�v*���/E�;�u�ZR��F�����).Z�j�WWl��n�������t��AI���6�6~~���\�ᬷ����E��4"n`��B��*K�چ��5�h�y#N�F�f�G��(p���Z4�tb���@����(�}j�]4��%�ee�	�X0"���&\�8���',����^�
�����u5�x9�0��"Jl�i��'�Ւ�Ҟ����.�S��S�hO n��^����T���(���I����!--�_��[b���v[Zx(��7U&Z���ߖФ ��p���G��JW�e�"��2�n:Yen5}
�� կΑ���<m�%(�j0E�x�
���o/l�5��F��a�'� �\(aO������3lY0əh���%9���BKN�(��9�.aPI�;�(��^7��>o�·�������#��pt >
�D��ׂH'��懕���[�~ʼ*�N�Y7�-��#�4���AK>���Q\OK}YD��{��%��ߧ�i����MmVU�T�pvq'U�e6c1��$IDqw�F*�{��N^�
�%�9��Lj���F������V�G/9��ɬ .ek�hp��O1������;�[�)�sV��\�<�.�����a[��a������W_���:�U�J�C��l��ο�I�N�*��9�r]��y���b��O�-	�.*�I�t�a^nL���P���3=A�\�E��?vSs�$�K�,�lAoW����p�ț�Ef?���G�6Q���/U��L�r���5�p�hy� ~��;��r>m!�@e#-\^�8�~�fR�����'o����mԄ��;�
�����j���0N��.���J���!�k)�R������
ww(w�/<���e֚�L��}���9s��S�Y^X���y��K�%��A���Mye��42�P+�F�9�x�_y�Ys�<����w�rt�@bXq^�#����I��AI.X {�9��셊��?Ǡ��r�b�('�ζ��U�N��x{w땱VV�屳��'9��z`ۅ]�n���$�h��^�ܼ�K<+�p��r塼i��n��t�-0/���ѵ�>`�}Sy"D*�o�i�r:/�Eͼm��0.���������g�v/���b�a�`�D���w��^�_�ŕ�	V���Ӽ1���.�U��^���S_��j�8W9eL���@/Y 2C@-�����u�c%�^z����0��4��$3�$�B
M�ܹ��XxM@�ӪP����T䔢�x�O��^�"c&���"��Z������2+no��v�}�n��hLӪ=OI�uQ&|Ji�k��HNlz������g~�s=�sj�w�lp��t���#��r�g�B���J��i�_0�+tG4����vj�Z�@�A<��R�T�ϨH�_Jٔ����Z'7��J�=�%��<��j�p����?�r���_>����v���A�}~�����*�<��#p�y�0���A%�����2����t�Ϧ�)�����?6@�d���bI��,��y�g����w�ۯI���������EKm8����+o��C�Pu+���C�HK�ྲྀ�>��T��8V��_�F��)�^��������
��P�5Yp
��Kxt����]��v~Fp"q�d)`7��^�5����ʒ�_3��r���-),�M��o��%��va�[t����4��A`�րѤ��9�	�-a|���5�.R:
������!�9��1���#���mpND�:A��t�_b{E������!����v�ͨ��V8�0a��S�#]�����*��]Obj-���!�{h�:PY[�t��H�Md%���[�f��堮��y�߉,Ք��b�Vb���\�6��`�]5�.��-��@*u�Cd��l0�j�w*�L���0��U/
�+��R�Y����×ฏ�S�1�h�m�8��,���f4���*R��n8Ӂ��s��L�z���jGMP03��f!�[	��������u{@>'�Y�Ι�-ڄ�ȧG�	�v�[2�=�5���E���)�l$!mb�[��.��->��tn�h��43U�i0�Ed�|K�/�U� ��F��7��ЙO��z�V��Sr�r1M�Xu�"dv]�ܱ��h<�\�l���R[!�ܚS�ψ>#]�&����[t���G�
��D�q��đSm��p���C�e��@=�������I	17�*�)4b����{�����\�$V�]�L���9��U�~�p.��7ĿT�2p>�I������'w��K��1=[�&e(s����D�gv��8����LP��}�H���������9{�$�V,����ݡ=�]�����.�r���y��m.�����t?��_�u������{{�p�ؖm�\h��X��D6&�� �`C����l�Wd�n�WV�)�S b��mn��]�2�y�
��#9@�9"��^?1�)���a"���S�ȥ(�綂+��@�Ƅ��vC���g|j�	���̓t�&�c��P>Y��Rk�+������+#5��B�cMnT�yI�i]��5�C��/z��Uq��XT�R;*��8��-�-9E߈��_�-3��DOG�������:�+����%X�_���D�A�R�\�G2Q5i�����p�о=5�4�_� ��61��ة�%�%�����-�r%y�h阍�O�ݫA�fޚ�˒���k���8,�77�u�\�)G�/�d��k8��<�_$1��Q�Y���żC*�8�H�#s�Pa�6�Zf���ġ���K��$\�?ϷW� 6WmK�k�d�yR��A�g��o�w�C�/�s�a��*��Elh��95?~�gw�1��$J�5��l������d$�(��a��U�~[-��Ec���c�Tp�~$눯:�(�O⿐~@�8��gr��D8$��pMe ,�
�,=���R�l{f%&g�����4�8�&�E��.WyRZ���D�̲������a�2N�����t��ȯ%�����z�ݸކ�T<�h-ˢ�-������f�����h������غ��吂VZ�]"��"�������N..��(����T�#
��_/w�@��f�O�*+�[A���E�|��_��<���B gA�!P�v����I-E�@��x�7%���؅S'�b��ܫ����gk�O|���F�D��k">A�;��?xo�f	'�'#�Ef� ,B��'���GaZ�o�E7�>�g�+L�sӃ�e�7�I��r"	.WQ9!����PH5�%]�P��r2C��y��ޏ�q��
T,�$s�;�*\3I�p���F\�b��H�qO���|=m�q	�z�僝e�`n^�Nc�$j��n�
��ڮ0r��T��9mo�&�V�j�$x�}���x	t�1�g>}kq�TvdpVRQ�m-ޮ�:��������y�K�GvP-`��HC2J�
���h�L�SW��Zb�Cv<
r߁���:6s�����ǧha����RGg!�!���W�/�>��;���A>������i褣һ�g�m{�����zk��2�#��k|v5�ol�J0o�L�:�J	�ŀ��d$M�N(�O+��t��4vRm����+������qim$�}�iFs�t*��qI�t�>��LUc�}wX6�m�p�0z�Q3��I�1��`f�D����a�Q��@?�}���_lk���CY/6���<�����B��Y���'� z�Yp�;�l|�E����v"���:��J�X
إB�}$mqX�=����C*�:�~
��.Dv� $+q�bح�������=�RHw|u	�'�"%26�s�+Q������j-�<�NSE�XS۳���H�Gng���ݷ�'��ˊ���X��zB�
"o�+���(�Ja�i	�)�z�Z<=G���餑�(Znݠ����YU�Y/|%���(��Ħ^ᒩ<b ��S��G�]1	�i�����B.@�8+5
����wY���A�B.�q�5���#�s��3A���[�
������?��_��M�m�u��+?�l����O�V��0���Tuw��np������NI�7�+� =Ã�b�3|�ݖ�ǐ�H�$�!8��FN�3%SVm,0?jp<5(��̙K��>@s��j������h�ܰ.�����ӅB�7<��PDT��<r���OY�{�1�i������q�[�㮯ۃ"�a��2���*�W"���\$w��%�[����M s���6n �F�J�q�z�R�ʷ� <�����,�IO��cJ�@#9w�N�6����|�|��0��KHk]��
kw�yw�X&�jN�R��~�.g}�A�������?������hp���4��Z�\�:]�r�Pm�E�a��)��l�a��$<\ƠG��m����#���|�B����)�.]Y��26�a����ϱ�g���o	:L�zڄ�拻0�<��Z� �"�aFڐ�X���6�!r{ɨ�,E-3�
�˶-RN�o���9��A�
LI&0D�i��]h��u�#�+8��j&��2�N������c���P�*l�m���e-ն111AkG�`ˆ1�:#v�����|��߳FS�y�j9}�+�3��M��&��o�ͲOx��/]Xv�g�,^Rb�3}�{`)�_r!��:xu����u���$��i���MA��e�	��4��+
t���?��k>��SU��n�=ھ��u�O i�Ჳ��AJU䥿�a�[O%,5��A����i��1��T�,������m��綟���&JѴ�we��h)/L������=4B,{TAQ�O�kFCdVd��K���]�[���9ڑ㣵Z���?����h3�3N��+E�\x��8�n%I�M�?���Dl44��1��B�����]݃���\� ��������+�MQ�81����AP�,%8'~�x����wM��V}W>�	lP�"�
�	ώ[���MPx�>��� ����U�����HkK`�aP�ނq���t�)��0���������y�0pQN@_9��l�(�( �c����a٫VYN�Ȟ��C�������̇ҋU;��2
�j���m�ȸf���Ɏ��i�D�ز@P����6?�L�qE���T�q�w6c���*?�s��^}��a[4��=,�$B���C��WJ�Zvʋ4g�F�,uozZYL��31+�<n{>�q�/���|�ebI�]E���h�@��J2t�M7�s�I��-�9���aƴ Ç��t�ﳩ3Ժ&�<΄�>�at@_@=`�#�.����G_�>������MM��!�wG3۬�9����2�+��?�r�^vZ6@���a�F5|J%l�g����J1E��3SZ��oƈ�U�弝��#Q��|�L,?Q4�d�tBQ$���j+��p��n��:��H�F)�ϭ��l"_yҭf[bL�AӘ�O�or��7Px�S�<*55���&����C�.��S�]�ԴM�K�<l³��^X'Ҕ�`�d�I��a-�l�ޏ/��a��l�%U?y�$aN�vx֒���ϳU0/��&qHv�n�j��^���5�>����F+X�S�&~��K�����)
F0��إ�
�5Y�~v?�jo��	��LZ6":���e2�O�i�Gl�r��NHѕ����7�4A͞��̛��2�]�
rw�+�dl
;���>Q�A(�[���i��5��i5����E?>�ꢉ�~9��D-WW������`ܝm�ݻ�>���C{��݌�y�+��W������F�_�@/I���"�����EZ0�B�d�X����Mш������K���i��쓖�L��h��i��f�3��U�ؕԞ��s9r</�� q}�Y[��5�\%	<�;�v�'V�T�����̽v��:D�b���tFe�c�Eh?�����8�����(\�7ؠSPsS����:j�/�c"
j����B|�@i�v?�M�P�]������n��Z�W2���j�wt���I�YZZ2f'�@�7몐Q5X��\5�҂�B&��{j
3r)���t6��^Z�/T^�:��cZ�l�G�!gy�W����[[7J4�'�S��A��������Z�\j	�3e��hx���cVz�G��R�����'�+�&��(ء��]Bۻ��^疇���(��crl��7Zۅ��_�8#bE��k:�bEHH;'*�6��8��Oڥ(P�L��8�C9RT�BJD ��&��-nT}e��Q/���g�vt�0I{= ,���pdo��7!�eG	�;5���{˿��9��s�	�f�-?#����t��r�̩��{���'I(QTj܅����߶����f۫�Z<�W������#��g�މ�����������H��%5m�ó�9�s�9��T�.����50��a,ޥ/"�ۥjl����9�@���5ZfE5Pb��q���0��3�߳��eGr����WC�����[�.lI�ee?�����0�y�ݰ�LW��8��q&�cB�~F����k5;������l����p��g��ɱc����:�2)�Lr�N�Ғ�����]�����,���O��a�W�KL���b�Cэ�8e���)�1;	')�6Uky�1΀MUӥ��\����(\�������bعS^�e��
�y�ߡVr��YƲ���q�2Y�m��3��I0a�A��:g�X�����~s?��S�W�_�����︓@�����2b!p��V��"���)47^��"Y �
}OY�f>�Q��Q�,���A�c1�c��
'��^�J�.,z �w�ާ�x3�z-丘����]�t�./;�/��.j��Xn�ё���s	/�W��:{���wH�Ѕ����mwH]����͘P��ϕ"~�-���Ow�����<�Og�W�o��X�4ѽ!��*�!e��ĳ�^?P�M|�N��������Nmy䋎�Y{J�7�9TIzXz(V���P�șф���U���'�$k��l,����*}�[���g"Ĭ���j��/9�{�#��tم�~��,�^�����wr�{��������o�7�	���1�wb%����B\��v�2
�0^��E��Q{�&���5*	����j/UR�� 3A�dPB�/z��u�h��%��9��!�2ס�
��GVW � Y��N�J��4K�w�Y���/Ep�f�W��;?���ȿ��`s|/��G�W]Hr����ѝ'���Ar�'mzh��}zJ������.���F)B��sD��ء�v�I�dU�ݪ��C�����|V"����깿�3V��f��o��h���/��SV��͹��^��}� �s��X��=Uh�Q��=V���F�6Vp����jr�-���0E�⺒��"��^ �>�d:wq>��������.Z�[ς;[-EǠ�o=�9��~P[E)s�}4�v�T�A~xL�](3U�q�oQ�9�鶏���x�0�2r��=�!'OK����B|��Q��ȵYO瑯�gΔ�-�^$ðnT�j����Ya�=9|/��d��_�K����������`Ff&uTf�iU2����'0zd�2h-+c�lM�wC��:�%�����KkT������>
�6��)+8��3w$�/�2?��U���eIP.m��}�,����7])$�8n!o�<�rK�XW��1*�"p�����A���QmV��������!�_�V$(NDaXAK��r�=Mqt]*�gb1d�3~�pU$���F�S.�"���XųO]xbH&E��[�� ���$���py���"ܫ�%tl�Z�1����?q|��#�2��E����x=��(iΝCfb� S)~w�lu��MV���s�>�B�����|���O|��<�)E_�*�M��+���L�kCS|�Z-�':/x
���nۛwG:h?�t�ZLΛ��r�(�1����֌7ӝ�N�(Y��y{��̫�c��©��[��뫰8�a�C!����?�%��B��q��P��۶��M{wM����˨N��n��7�L>.�6�:�
8�c��F����>E�kX8$�ŭ���/��i�o���'JL���#%�ri�����y
�����ihuϘڠٵ�,�UVD���=��Y�E�8�j����ֹ�_�s�q&SDu�-���&�z�(������T�A�ncbm��CuU��d⳧���>��I8��9cͬ�₂H0�8 ��K���b��Q�����Yq�f�k��$�D}r��B�l�i~[�=�Dי�JF��WUmw��߱<�3n�mG5��6A�tʤK>�g#��7yzQ
J�e��M)��8�Y�#�~z���@�<� 6��CU1w��7
�$^���"��5�ٜ3�|���G���q�
*Nz�N�"LD	^yn�	1�Vv��έďث���l1�j�p��aќ�>�o�
�\�صѕ�Y��f��u;��면��{]�q���lYR��1C?�j���Ӹ�=�c�Q�V4랛v,�-�}8�d�<eK�X�4�n<Q�-$�Y�Qh���������7+V��sn���m ��MQH�O���F[~4hK�{�t�C��n?~��m��1^ļ�1I��1��sW�A�/� ��1x%t{{�*އ�ݡ���V����Q�G�P�X�ђ�b<1n���J1���&���-1��?~s���{���O�cf(�+u$����l'v������*��U)��ާ*�G
���G��3�]2���O̥���{��Q`w4n��k�k����E*9T�[��к��R������%gz�9a���W
H�������|����t�]�|(`����5j� ���(�V.�b��B�D�X����W��XiK��<!t&�N����kk�m���eW��)b_v�iMM|�H;��Yc�k���cSS8�k�Aʣ�����M��B�S-ox�!\��C5ZޑpAf���ٵ�����As��k+�.�'��+)��"�Ս���-�4�U0d�4y��L?	��i��xY%��s��bPFV��x���s�1ypo��h+2@8o���D�y�?��R�?�h�z���yr(�K��<���t�@���(f�\,��#�c2�������`̯J�o��[�����>��Ixwn׸��
�;Eu����ƽ(�X�I&�L-S����X�bנp���{��F9��|�6sۉ�Ơ��
�ګ������)d<��m�P����V�����*҇�܋h����.q��3�s�Cv{�b�`���R_Vq�A�'v�1]b%�m�vd�)������ݫꕒ�y=oұ�h�����%�_���W!I���a���J��9\��3�Q�k�W��s2�K%�ȡ_U��JĄ���W�OO�#MJ��Z�TЄ��\3˘���e���Nq���_�<���������(n�Ȧ Q��B�
��亶�����Z�;�6��
x�����|+�&i<4���@���݋�1�~F1�C������#�
�)��HHL���ihR��I1��R"�k�(o���$�I��ڢ�̙!���ۚ�8�9�z�i��*��GI%���h�q�1�4���z�^jj&����=QLa
���,��!%�P�>"�ջᒓn���8��=Mg,Ͳ�I$jg�k�#iCZ��?�~�]Y�.�/��yG��}�I�G����>���l�=a�hJ�+G��Y"i)�l�V�������3���ʢ^6n���m)E�5���fse+^|[�?���&y&`n����x�����zC�VI�IE�x�҇�����2^�l������/}ǔ���_�e�o��E%��b�Y�
���TO΄蠈f�	NH�\9y��܇$�J��;w5+oM�z�|ȓ6�>y*����	8�ĉJ/t����^FO_O��+6ΰ�)��o440C��g��\ND�pWb� T6�:MU�6�^b�{��5�������3�F"`� 	"D$�$����G~��	��<%�P���n9��oE�9��������p��Z"l��1��#�8>��f�qAcK����U�`�b�b�I1�v�T� ��ו�o:��k���o�P�&zէ��T��uG�	�%>��%e�覘��7��^*b���?u�X��:Tb-ӊc�+��g�(M0� ��^��Q̲��!��$����˥�~�������p���&�6CZܓ$�i�'S";�ְ2���İK�7Ǖ�um��Q�w�|~��!�^@/�j���P'Z<Q�ߟP�R3�6[)�;�:�yt��ws�dމ�̲ S�w�%|g���[��Q�ٿ9<JK���sWpK�{�.��^��|��&��T+W*��\냾qG�5`Q`Q���I@0O��i�s;@.�OxK*�O�'�86�z�>�a�it���Ƌk\#��%���?�Ab��M��U<���?X�N��HB2:ZI��5�Bg�0'���A�c����v��]���O��T�
�gƴ#BG��m�5��]a��I�-:�.GO���ö'�Q����1n��͙:����9����]e���Hֺ���vT���f��FGʆ�3;H�9*���-c7���y���N�A�ka�9՚�3x�����D�oV���jE�K�&b��NY�s��=���OUMc��K�!��}��r2��BT&͇��Q\����v��'ܴ�����|�Aú�k���C�vvv:)�F��%k��n�|�Ai�!�J[�A Jrڴ�B#@!��C�@/�T3�R��HB���p]�{�������kବOar#tedj�K�{��M�������xL��YY��}b�ȵ�ܼc*>�r�������� �i����(n���zHf��kVF�
`3�|��x3�?D�W�g�./e�9��z���3�h�O��F>�+|��Sݪ��M[����5�3���]̀��v��a%�r�\��E͂���Y�(�g��i�B�0���.��4l}�h� я�����xz
d���rT�m�(�>�����M#U�ѱ��i���\�X�RF,��t֑������f���׳mܾ��w�9aff����7�0�ٹ&�TY�w,���8���--�3�N�4��JR)d�X�F������f���)��j���0�g�|$yk��e��U�mѪ��@H�>b�Ie�W��R~�R@OQ �4u6��#�W����=M��8�I���sr%���[OM�����0m�w�:�����g��u5W�\�J�����:�å{z��0���_�p�k�T[�	G�p�녷���Ɔ-+V�*Ga�o��]2{�e��1��2�ܔN��}suu���q�zu][i�*�)��+�g]��X�_vܣ���o�0�b෶���3}�9sA��Yi��?��T��>wO5�j���� ;�Y���}�[���	p�}y�E�ȵ�Օ��> ���Q)SJ�+�۔�ⴤ����R �`�|�o=0�%����9�,E��.�߰?�d��)��(���Grt7�QG��8�����R��o�����E=��emD���M�{���L-ط����Z,��l�� <RkZ��Ɉ��]Cܶ���p�'�\ۡY��y�9���q|�ڤq���[���\��RDu:��u��2Y�y���
�:�H��H�3��HR�ͤR!�W��2�Ψ�D͕f�d
�7���^����I����d�K%�UI��R�񈕕Ih4�"F}Zi�%�/��=2ӑ"���h��C6���R-��/�V����X���t� Pm����#|yQ0���C-Y~.U��!,�f���q��r��˪�(�v*h��R��J�`��,�hp�h�X���f&�_u��կЊ��eE�P�|@�ui(7��`g4;-���b�����uA{^`���J��pc�ܡ�8!e�(]F�.��J�hi�/��@����	��֋""mdi�����|s�����")�"\�[����]41&�[pb"�L��'N�rѽ�r>Vm1���W@P��s(D�8ED�*�`t����k�*���H��ElwT�Ŀ�߄:c�R�8��2��GP:T;�������b������ %�� �@��e&�+6�6.R攐�-�JG��@�ܴȥ�pO���+�����NR�c�0��S�,Z;;�m���q�3��
��e t��|�����-]�:9A��z�������_We��֯�����R�^;mD�@o�n�t8Wy-��� �l/I�)��Q��.����7zZ�u�'�/uy�'޲d�l��η��ZVې�K����5��2|��y�u�"�9�q�	�>�l4��]H�"�Z���C�ʫ8�x����o'3������V����B�%�A�2Ú��RĦ~m�Y��N���5�����I>MmۏTp0Y[�9���爊 �a(�5�Ղ_������4�����ʕ���šHGT����"��I�X�>\�z:�v���đU�Y�%�_3~!2Kr�@w=A������i�V������X.uqi��XT�k��0:1�V��1��"g��LFbqpu�G�����?l�,����\ʏ��-s����NJ�ʹ�����t.���a|��S���.�����\����ެw��u���^k����4ѳX��P��g3�ESt9)�����f4).I ����$�K"+��K]"��W�%��Ve�Sڣ3���fn�ԛ�[VuEN���`�s�������3�øs{:������!��H����ju�M�[��8}@%��	���C~��3`����i���Z:y����>��l����r�,m�,9��+*�?}fR�	4:���o��Pm����`go/P+�ZO]��u�#ӣ�v���^�%�m�`I,��u#K���������f+�Y�C�e��5��[d�*H�ZY���b�v�ȧI��6��:K�<+RP�#l�'�ro�L��_�s�ޅ�������V�y��s�e[��G٥]l.	��F��� �YV�l��*�HL��ԁp8>�b�sm�S�y�� qUMM��Hj�����*�9{n"_��gw0��8����/;� ���I��m�Vp�X��Ń�|T|�Y
�������-���OI�����~ooS���H�qDP���!����Ե����MZK�R���133�%�@�>bqm��&�I􍙭��	|�$� m-��`��U����-ˀIW]m"����\���f���Nd�a�msc��k��7J^�2�S�������F9�$Z��%�Q�@�����7���6��*��1ɺdʱ��y�*�b���������Ԋ:��Tc��>���L��E�'n�H߶��{e��~��Ltd@�3�n����{��t����@E��>c�
!���y���G���Ҩ�����_�v��|1X����)J5�����[�����ˉ��d�䐀�����G�?ߺIv��`�a�y]��:���+�\9<P�s�4�b�\4Wa�pڞhֺVSjґ)��1��츨�ƕ//Zъ���� 2��M��3��J��4����>`4WL(��!��Q�#��?��@A�VKK���;���ZM�a#j�D����d������5�7��~ߺ]��U��c�L���&�8g.������ѲT��)��ɽE�r.�-��{�N�Ã'/��S��7D�}ϼ�Ѕ��e�s>� �������:�<��	�{&4����e͍����������1��S��]䑑�����U����w[э�Sw�wFbǎ���щ���?;��gۧ�g{Ct��ޝ����ޣ�nͷ�[W�I�ݢ�5�s<�S�����4��Vk�<_7R�@��qOA�cL�K���N	�2]-� �E9)���cP7��o������ub����v���(��0��	���M��pQڠȅ+��;l��v�bY����U�uD��l�*��ug�S�ϣ=f�80ㆿ�+�1�����Rh���W+fwc��] e�UO^�3F��D�Q3j�HW=澩?|�-���I����W�KL?ȇ��\����wkKHz�;`�Fm_�puMv�~Z�y{�@���>�r|�s��L@z��v8�U�������)�g]�_I=�W��[[[{��tA��a�χ���<�O�I���3�v�Ž��k����G�����8���u�Y�h�����{�����!<rzK�0��r�q5���wg�r3�����������ӎ'�[77�-��L=/ �˹������S��j}W�U����:��{`����/��x��@-�LI�l�T�&ٔb�L��SԾ8ex�4qƊ�5���Xƍs���Ȱ��޳���)n-_�+M�`�Z�⨹���{��N��y��y�j�K����W�`+�:2 �C�4eį��OP��^�����/�)j[~��̣�B�~,�K���V��́��2c��MB�q��}Q�W8n"���5��U�ۺ؋w����!��_��o���?N�ݯ��oW�\�.es6�h�]2�mYR�-��H�qb?�j��\����u?(8��4`߼;2�i�l��ޭ���t\��r��*��w6��i���	_ �z_�%u�?_	=�Kz��y�f��z�E�;���/�o�o�s5���}ӗ�LLL��W>g�;/g�"�"���lf1﹁o�S�o��	�w��!t���q=-�slJ�c�vcX�Y��������(!SYY	9P��KKO�����o� ���������e��>����Xq����s뻟����i���0 zzG�	_�|V�&���6m����~<N��x���&2��.o�rg�[�hs;!�}���m�]� 8�~-�2�q���k�xa��H�F�t>�|mHSx%�<�*�ࠋ<�w��u�#C������ݪ6~�������*s�_��c)Jm���C�z�n);m�����=�0�-�g����,��~ݽ�K���.�aQgC�mMG�Ү9�㺙�u�f��@4q�ۋH��e����;/��d�_]�R��;M�[��|��S ���W������O���힬����y�x�>��4����=��i6�����o��;���}5��_I�꾊�?�Z>�������'�	ݓ��p��[��>k���|lY7��������=|ErD��n$�K�ԑ�Ә��QH2�ɟ���Y��	j7D<��N�Bǻ���7��#��$L��O��~IYu�?hs�@+?�I4��4���$*	A��k���t��L/��P G�ɉ��~�k1_��軣(�9C�bo�2W�A��U��2RF3J"���s�}�1K粆�s���߻k]m��	��R��j`���'�~]�T�J	ǧ���ˉ*`�T��.$.���l�0�^��2�|N�^����^�����	��.����B��Umg�B����G�����g!%��5�T��������Y5��|t_ ̈́�3H����3ܻ�=������� 8����}�T���ԹQ8sP[_����n*������v�*���!G*i:=:�a��Ќ��\� nO4�����:��\�
���,Ξw�Z�.Tt0�7�{Z�=��G��u��;�c�����O�B4�o� 4�^�a๋��e���y���un;�ZZ5�hc�s�9{����=��I>�v���ܝ�1b��CcG�ؑԚ���h��$��{���H��х��}�r�t�����:����=�&����T֋��c;G��m&�F��?l����Mt�]�hl��v�M���pg(t�V>�nܣ�v�����hS�u]s�H�^�}�6<��v���{��t�?	6y%J�7�D��>:���7CÇ��w�`cusg۟�\���F5kź����5o�*8���k�3d>i�]��c
�Ն�S�����wK��׉�!G�Sg�v�h��D�1ND�5��Ll��h�����g�=�?7�8o�P�����l`밐����s�HE�÷w�w�	�e�sK��hU�(�����Q�`��3u�fݲ��I9�i�~���d؃��[;��!�ÿ5��o81e$|���_ ]���H�6�;Ʒ�n���w���� 
�kcc$�ڻ ��6�#<Sꤜ��M'�s|7�xO^Ƿ[W�L��4*.-��E>�6�Vl_1�?A {؟0�٭L���d[-Ísd۽X�40�N�41j�r���7�O4�vS�>�-.���S�~[����4m��n\���s��G�}���u$[��&���~�@z��Q�7��r�o�;��.�[5Y ;A�>�����ng�@��st9���LQ(�||����)c,�>k����8��F�U�E�F�����Q���K�AU&ӭ{;0�ctl���]o?�7Sa��d� C�I���ۻ=���FG�/�:OӢ��3�����_|�R���ZFҹ,��t^>�&P��1F-�);�O��X%NgY_\�l}b�'�ǚ�p���:M��n����}��'{[x�Ҥ"��_оP<_�R��p�eh��S�jZ�Oc=�9�.�b��՝9Kg��f���h�R�w���{��O<���)S�� :�J�B#O���f4��?9�Wd�K�X�����^:�xQI��r��֦��y��=�e��e �7ƨ8�"�)�m,�d��/iQ/5���n
1p?dD���>����O-�}�B�J�:9���)�Et]"����� Z��$�d��1��.���ܪiř#��@���L)���� ���#��d���!X\_7���U�#�Dq���ײ������5Z��1я�ɵ��3���mm���X���_9 @���}n��3�~?+T#��p�md�>���� u2�OA�m��5;��+хO�<��E��⮽�"*40C�x��2!-x0��Y�}[#t�{�Vi��� �Iu�ݽ�<Ê,�t������EB�x��{`����%dH��\*�>���YU��[j��pm��=�N���,�W�4;��Lv]�?]�wSA��igqQ�2�t�I_OP����W�(!�%�����+�i�Z��#e�0���%�p4.��!��%�"�����]��:���X�f�=\�̛��h���{�M��W��sל�D
`�����Cbׯ�gЌ�W4%� 0	�MQ�qnr(sk�[}<N[z�v,�f\�������Jf�*"�׉���ޔA} �!\��^��9_7�K5=M��-��\�w���B��a��!11��>-G����@������M>HI�5�3*�� ~o��B�H(pa^���q9�íb��TVT����hJH�?��2(����n�Kp��%��www�����Np������W�?��t��K�W�)V�����yq��&Q7��b� Cm��A쫹v��2�Rs�kU�c��W+و�~n����A
�	���.�k�o���j���*�`a�e fw�A��q�hhP��0N�m�?jo=��L�ݑx]�IE�1�)U���ڐ,6��I�r���S�i`��4���柞B�DL��ؿ�JZƗ;v}}=S�S3UP+��W�M:�=����DJ|�PJ��4�K�M�qr��Tu��;��$l<��$�oPb��i�����|��S��u6.	��H���XK�M�$�~8���(Rq�ڠ;�{����9K -�b/�V<
HMMGW7�a�e�yu��J���5�a�G55��!�6�2T8�ճ�
2i�mv���?�ۚ��i�u�aw�
���B�c�l�}74+����[�b_�lEnQ�������<K�a�Z
	n-� �Z�Ml�h���{v��x=� :�sW�%�&wb���F�����LU4�_�+Ϊ����r��N��o�'?3����#��W�c\�Bݞ�P����x;��v%�M/~[���$Q
`����cMA��r"jˁe1@'B�8�l��,����2_HorƱqB=��iV�zN�6��ˇ	���d�������Ȝ��T�X��Ԧ�)��̉�&2��A���cT��_8R��� ���I�'�UU��E��c�(��{b��B?Å����yz�����vvlU�C�Х�ۋP"���#,�0���DB
H@K��>x:�T!��ǤK٫o�����{#?�߇_>�`�J*��pe���G�
��p0bzX@d}@��Z(�%g��	��d��3�A�{��T(��J���_�.�K_U~�r���y�	�qv�xЕ�֍�/��"�Vo8��>.o^cQ��,�ni_��T!��Fú�A�찑ҁF�}��cF��y%A*�q��2������(d���3҈R��H�c���x��z��ch
U՘��>�:��_0��,#���x����tR�3}��`�J����ΊEwS���\X� ��h97�<�u��V�!���Ab��Cu��T��a5�����+x�{!���Ԫd P�����Ϊ���E�A�6�ER��a�H���Z���r�"��?�}�j�>���6�Y�i��).�1J�5����e_D��$R)(L�&X�mo'�	�)zL��O��i3����
��r�� |�C�Q"H��>p�nDgc*3��3�g/���,�9�r h��6?e��ڈ~'Q$=��^�L�C�Z0��@�#��=�u��C�Ze�)@#E���9��뀈�Ė>J�L���U��� �\�)� �n�a%�d���*�~6��MX)z����-�!���a��U�io��>(��^$0�i�����^�o+��v���4ݼ�6��	O
�<�Όr�B$��KG1]�i�u�]K�R�V���d��P�$�_D�����]�@ƆGŖ�K���ff��t���r�O30�][���0�_n����i�>rR>?�P ��rk�º�"��Q�n��N���K���H�p�a/�eh%���)!���#�4�ap%H0�{�ctp-2B�����l9��r��L�Gb];�!����eY�n?;������,�A��W̩�@U��kJ� �LWCy�*kS.8i�ng�1d�g28GE�S�������2�&�O�k���7��':�\y�Q�z�H�_!u�[�т�g����g*����c��q������@vøRW��w|��[^�3���8&�,,��K�i�&�7������E=�LZ<�?z�H��%>V��9�S9��S�|�pW���خE6����JNvu䓳̻5(����o�(\4�Č��H4�8"����<R0�jc�=�����t,���z�����)��9���iC��fվA�xi�ML265�K��G7�>��i�f�'�������7�|�BN��PE�����ʊ�1��L��+�Lm�K�i����]��|̓��l�nM����Ru�fNH�/pd��Hsߌz��1Ĉ��d�%o5��A��4�ˊn)�K�(/�����K�b�>N�7sR#Ir���o��\l�V�N��}4�ph���?ɑu����y�V��a�jzq�Z��S�HxP�ȡ���kQ�\)i@�+I�·8��}�=���>�5F�^�9j��˕˞�N	>:��x��Z�boY�~��C$dT`h�#�t׺��"r��o}��Ӎg����<�(7�����{�a�,�5�N��2us;:��enǴLsy�G����|w�T���Hq�M���5[�-|�k	<2��G��U�Y���k���w��AƣZ�<D�nA�u����c�rRk5���K̓�F��
�zu]��6�|��2|t��<�1&h�TH � ���� =�9�L^4���-|!F����4w<1�{����Bp���!'&`J����gӼޓ�/㦏���K�� �.9�@��*���9��q}�vٍ�����ł�׽z�Ͷ�7��cz��.�H,r<Õ-�7j�-Ny��;�b�v���n��J��nh�PM��pJ����OUd� ��ɽ/���L�n����r�n3���+�W��P�s+�V�J���L�"~SR|X������L&*�9���c��C8AZ?�.B��ԭ���z�NWn+~�l~~��c��8�*�Q�Hڒ��2��zIqrJ�Q�zC����z��2�PY��ٵagP4�|Oz����"!�?%n���/z�ۂx;sF�6ѐ���\l6r<H���"�����%�_
TƸ�y�%�Ӡ�K�!K�����Cy�ʨ�b��2�ˡ[tT��k\���E���~�?[�grU"LrM���A��J
��U罾��]G�c,�\��T�}�I�'�V�0"��gFp~�'
ݦ����vK�ֳ���Ͼ������Φ�P�}I{쥀��v?f��|�uH��b}�&��#$�>����`].�Do壩)�K�R� �Ӏ�y�{C��6i��� ��0���{O���Z�aM���L�)��@��f�]����TM���C�c�b<(ž$��!y���&�EO����NL$d(ؠ.�86�EG��T Fʂ_�gI֭3:/#��z����i��0�ב�b�k�.}��p�����zg������E���OOW�VW��c������&x��u+ˀ�����}_���#��]ߔBzN<�U�u��Hi���#X]�٤�h�<�绺Z�8	~ػ�V�Ⱦ:`�<�Q��#��n a��卩p�wi sX��ټ�K����a���o�%c�/srS��#`�[�o��r���Eҋ==sv>���1J��Ds��#>���m������a���e.{'A��i�&u���ff7�A�x�w�ܾnZ������d=,�^[և_�e����ipAw�'v��ټ��ד�)a��i�xqV\�EJ���P���H�I��#7k-�CT����9�o�4xq��_V��C��]}�C��G�` ��hX��&# %�r<oʓ�P�4�����B�b��=����	�l��//�h�ULI"�x�gs�W~k�0��=5�-R���uN����wUk��^t�u,��BҏfǷ~�A�/�KDM���Mj}��r���*i�B�ͺ�Aq�4s�D�6R����-��Bz���N�6�u�V4�4���)�I�J�B>���3�B���0U���S�MA�9vs_	�]����2��"0��k����%e�?.�S)�E'z��.�H�;5멞^4�@9�v��OQO+��$��aS7���E=���^�`�):��F���}��L"`V}��O� �7�٭���뀺(��2]���~7w�b���i4�����ͪ�����;d��G<�p��O��iǎ�O�ݵ���|���giU8�����<zڭ3�ύ�=|�M�]��<
1�	�Dy�WML��Z3O�夨��/����w�:�-j�6�&l�j�d�+�����7�
)
X��C^2{h���x�D�ܔ����3�#���p��e�g�S�R�S�A0�K7Tӟ��]���ۢ "�0ctKp��q��exͮ��z1��L2�z�ݐu�aF!��]����ګ���eMR��d%��n�����B����~Ӎ���B��N�.��Dc+
�	���'��6H9�\�&�/�@�C.m�%^N;k�>dQ��~���U��srr2a�?=;�I��D�寞Cin��QD*�%�5a[`�/SA`�Q�ͦ��7���lB`�AԱJ��B�����oQ�G�@e�{8��?@L�s��3p[_���#��#�˅��lj!��M'�$�(oX���.����f������)xZ�@���WaJ�c�g���|'��P��j���#�+L3:q����U�V�B�B(y.�������B�/��bu��rE}G4v� �������q�R�GS'��sfj�@������G��誮;h/�K�h����$����O�@�2�(䡝s{���fe�w�����k�hpR��=�S���y4"R�X
� m�i���4��TQh��R�9R�G�������9�E��0uE�r��ͱ%s��,*�|�u|}��c+x��[�W�� 3��t���>���[����v������0�E5|��������}�sAKS�-b"�W����Y�_P����?pqyY��=-2���Ӥa���ٻ�{�)�jI<o}�eu6ge�.�?��>#lI��N��ɸ�o���a�fHB��_�P��vww���B��=gv+6.	_ ��-�A��G�����S{�y�\��`G�Uϖ���4;%0�$ns|�v��m����3��X��=���y��ƍ���~�b�8��(1_�q^��J�`e='���#��²���ŷ:(�`��'�r��Q�Jq �
���2Q��G�<��#.61��}H�:��$zDd
?q6L�p�ݦ��y&��t�3���fgA���x.F���+��]��h�Z;_[S����ɵ��Δ9�n��n��F��)��C�&���@O���yh��������4��ӞnQ�Nܚyx�5���+(Dppp����7���U���#�{z������wN� u�̧l���-�����oJD:�U�K
��GUd]�9���4�f��(n%k.���!�{��y����,-e�ώ�q��+�7W(�����_pW�5e/h�㈃K�G�t�7�S1�Z�^yWVVꛚ �-"�����p��"�*P����h��?z�����'j�8eC�;b����Q ��J��|����̜}����U�>���YY�eݡ=7Wvzz�����,V����d�$]6�q����[��J��Y i��z������G@�#���I�hrg�=^QG���
B-��zJ��kjq.uI6�W�.Ob��� t���(*�SbѪ��v�����ʪu0�l�(niii��w��������~[��'�>宎�%��S�}^kU?=[�o@�l�X������h��O\��n`F(�glJI�T�H����{Y�~;�|
��o�Q���uҝ�<�<���g^��ӊAq�� ��.��6� MC��J�Z�p�4���&猌���V�X�Ҁ�d��ĉ��Ή�e����IFL����ڸ���/���Op^U��11�����˨�[�H}���A�W 閮���};A���V���m��}?�2[�H\ �_�뛟���ȉ��C���#�O������8xM��Μ£f����j���q��hz�q��%i1��1�|f�QM���r"����R1�x�
������*�V����]����_d������KaK�ZZ�2��?ݞXTX�W-4�V�����r�*F�`K�dUc����u#�v\7mL�^��i�����ed�{N}�nl�)r<9E�td6� ��#�Ȃ�`�Qy}��A�ݻ}�yVVV����Xc��m;�de�+)��66֐>P�mR��:�����W�hnN\�W��(�߮E��b��@/�Ѷ�.h�N�!��f�����i(I�[��V���=��-���Ĵ�8(7��4���k|�6�K~�k�P�7�7�$����j����j@�������ڲd1:>UK���j%���{��7v���|�����+�C��&�.����"s�M���z�����hΤ����Ҿ��p��w~9�z�ŝ�8�#yc����������D�|�m�����@䦚v� ��R�XqryxK��|UKy%}[WC�ls�DC5��C�ʿ�׾s΀��gw�8�V���H>��'�S�z�����m�{a�6���M��8�h�t���mA�`�&�H]'	l>;����0z1U�V�����D0���%	����G����ok��!Љ;���OO���pT�´FFF�`C��0߲/�]�c��w��z��;O?N�~ȦdR���$���m~0�)��_�Rgn��o�D�f�V��_�TӅ����#c���	�9xK��L�qZ���?��	<#��������B$
�$JJN/��lY��3�*U�fO��V��D���|ʐ9H�� 欽�4P��a�wW�y�c�4a�9>���~�C)�T��ג�N���Ykkͼ�������g\T��f8����i���2h�t��oφ�ρ.m�Y[��Cr��DF�3�4����������j�G����h�����{�2��@���ނƀ��;b�U�����l2��&��p��g��R�����?l�ӻup����Q5��9�2���즥|�'��c��p�T2��l^�@O�¤���#�	��C�"��t�:�c]uu��4ҭ[�Y��O�ϳϔ߿&�6��=p�J�� �*0;%�rY
����8ԑ����FU�8����5M��#d�b9�h�<V6y��)��������N��U��޽�$��K�^�		���ʰk�4f�"11�ɔ1?�B��)/����q!䫖ն�G����s����׍��D�B��M�+�u ����!�Vy♳ �R����Jb�0�����&%����Ώ.r�&��$��֭o,;fz\3��L{���2
ď��L	����b��)'�'?�\2u`��ЦU�mU����]=�,����G*>�A��������Q�!�JK���69�9����������`#U����AA��b��^���W}�y�U(����,����%���&86A�c��ƪj����\�B��iŪQ�m �a)@'�@٠�]58�F��y#�	�P,b�+�qm�Y���F��>�oҲ����@�Yvm�f(�Dg��,��e-w�|��VJ�Z��텪z�$�����3��k,X����B���ؔ��%�!;��lY��W���1���� ==��f*�!��)�g���8����H.�C�^�S�A��S��sC�L0h��f�Y�4�C7��*�]�@|8�'��a:.f�������j��5͐E郧t�6�j2�%����H��ϰ�Z�:����H|p��hz$H���xl�����wq�W���JR�삃�?r��c�!�;?� P�@H��qZ���z8&��z�ᱺ�X�/����aln��u��^N0�^����y�|��5���6i�������މ;�΃o��Z�}1VM��o�C���&n7��ΏBnM+kV�Do\�r���&��]�1���ڈ�������R��m_f`g��UKz�K��|����y]�}����e��3k+Z���:'�#�4ҫn�R_�}�4ӭsf�	��4���Ϛ6��ަv.{&��Ih������G���:�EM5^����M�	�����z��W�o��|؉�9�/�yU��ֱ����l ���e�&>M᭯w+���ۃy�6ʖS�Wh�?�KN4Mz�C�<����~�#�ʃ�3��U��ʿ}3;�!��|/M��]�����iu��)Nt����=�ץ�����E�%t�>���z�0:N������'��o���p��ү���W��8������:2u?�`��m��?�:�"�p�[*�~�\BGW�:6��S���e2�q�����/(���� �.G��r� ��
���L:�s���ن��+^\��_5Dw>._5̸Q�DU�ٱ[�Bd�����n�������w֊Gx$PPX�/��o����r�|��~-�Hʧ���������>#n��L��`���`	�*���e�<�M4>.;��P�)jڹsf
%�k֒��C�����h���.�Q�#�%ԣZڣqM9���#T�ǵa .b0�r�/Z�e%HCc�x��������{�
[0ӎ�V��n.�~�U�2H)vlӲZU�9w?L��lK�q����7�p�9�+�g	b3��)`��Z����Ǖ�uC}}�#+�XJں�q亸��o���S�XV��=	�A�;�|$d��F�{��^���~g�X���2�3+����bH�����q{��z�	�P10����9�p�"=�[�.�|�_2��FmKヺ����]jb��5�a���u��F����Ť��� LY*���n��Z5�qN�s
>��7[���q6��Q0�N�ĸ<���f��|ΐ�nh���@�L��ѡ�健����J�UK!N#�]�������rf�b٤е�H{na�PŇ�z֡ոД��Q�ߒ�10 � J�^+�M��"��3�/��vN�vE�e�YX����� ��J��7^�$�3�I�OEC�����Ҹ�9#�2]��r&<�B��YJ4;=�j�hS~�鸺�&^g�4(���D+z}��xG�>a���.���,R��>;�0Ce�A��r�r�j��1X.Lts��7٣���hI��I��/z��su�����:�BHث���wh�'�>�酡OWj��&��w/������p@�u�����=s:��1��pCY��0ut#��i�/p�5o�W�f[�¥�Ӊ�C�Mwbcn��/̟�
%�W��~���zE��[^���K��l�ֿ�5� ��58�b�4�ڪ9p�� ����`�
P~��GA��� �!���(��+���F � C���P�Y@���FbO�lw��0����m����3?~���+��mG�2����n�h��;O�Hl]��O*"Ӌ�	H���##x���	�Ygg�Ɵ�C��3s���R�/>���2��#c�"ɐ��������VD,��o�O+�/*wP��Wӧ;� ��L[�����r�C���d����,D��F �mn��*�[��㣢���e��Y�D�YAL=�0��b�;�eܲ�[��zAl_����[[7��\�ł'�"���Ơ;�y��5�Y�1KK .Z�g�ā�J���P ��ÑUp78O�M�W�����.�$��R"���gg��M��`��q1	u���i\-n�t�/['�A+B� 'ggx3c�f���q���ꕏ�yk�H}��m~&G�g߫��|�U�cv|T���-�Om�5N4|�y��+�"{Rw���ʊ��Mq������P��B��l���I4��Ý�X�u���K��އ���2�o��|6��2�L�ih�[YE�����N&�~�����\gsrqI�;�u��рi�:-�ooaˬ�:�º�s�s�E*|ߕ{r1�\r������9� &�	�!,N�N�5J�e�C����}������8 s�F�`��|{d�kiq5m�PWח�8��n�o�SJ*�A�W��"G=���4 :��g���� C!��B�hu,B�1�"��YXay�����+g�\��06a�c����4���u�w�o�---�C���0f��]U�"���d��/����A>�Ѩw�y�������x�l��zE��Rл�GV�UZ�����Tp��< �&�X�����/��Y�+'X�*l��ک�<�։��U��)����X5��˥���$&%�"***r����*``���*��c��f�> ��;��j#B/�qΑU$�_���1�����֯�\�q<�9
&9�|L��g��3�r=:�-�'K�J��㔄���?ُ���0-i�F[b�esp�����3r��n��3�\H%�Cd��uP�(��N)`��kL�ē��S�J��vt��W�7� ��3U�љd`�@E�Ka��S�4�|�)�������&���9SN�C
�@�9f
�V��b.��	�W#�)�r{EB�5�X��q�oY1P�"�I��n@�s[��߽-����v��^#W=��ex�u���A��b�9U"�en~��z·B� ��e �k7��5���q����^��݁�]6_mL�[c�����Ѐ|�ԣ;�Ó<m�nc�v������*z��R���YK��c՟?�.XG�T&�y>n$͙%}�	|߰��$�Iٗ�L�\c���[��f���_a�1)�;;�R����)C��r�t[�g6�"��������_�NbI�G6��f����,P̙9b�Q*�Y�T�ߣ���v�9�ѥ����]���D�lL-����\=�F��_�`àK�Y<26:g;�u�����`���5��H��
GmP�P�P�Ymעe3>-C��a�}փy�p�;@��i*+����јUӉ#¡oyEEMc�~��녔_�Lĥ�9?�On�$\����^U�Z?$���T<�<��q%1�(��n�CZ1^Q9�Rq�ݘ��S�o�l /�]v	�.�+bY��j�̾���sδ�-��z����<Ҕ�?|�9r�H���'�ݜp����3/�3�����R^v��cyE��W�����y�H�@]>0�^�h���c>֐vΌ;Z��J�^u�0��%y��&�/�e�/Z�U�����T�`xt~��Z�̕��n�W�۶�qyH8�ǅi�]]��0��~����%_9sB��� �Z�*���S�f�1j�����˹L��o�: _��
z��83��}�Fн�A\�
��%c�aht~�t� ��+�R�%[l'gE	��Z�z(N���BuhjҀ�<�"0����)@Z�u$f�B����X�B� �h);�%-�ƺ0��a��v��]�r�"-/�#/ 	u�%�� �ݕ�H�X�ї���jOS�n�f782Ji%���#񳢕
�����c��;e�.�IH.�ӻ�Ÿ�h%}��D�u�N���w#�R��rrqLl�i,3�lT��FD?
?a�)��>*A+�F���F�QN|f]��pU�xurڰ~�5���`�F���}��F8�����>$""�k��B����N�.����I�,V��wjۉ�:�nn���~����}��,�ଇ�,]5.��_/�����5;�`u1r�Z�02��\�}����O�l>Ŕ���?m�=&�U:��J��tP��`�X�C�Ĭ�dxY2>w���Kf��������U�ژ�9�۪��5	ز)��O#.mb�/@��>�q}��'�q'K�h���a �E�����Qx�+x�h�)�j�eL�QǑ�=��eײ�2���-��X�EǢZ��؎���`+�(^8qk�*�='~�#��0�#����nj
����z�$�����>����F6�ߢ�錨�{��F!���!U	�Zq�8=\��#ɓ]���b)|�O@,��f������k~��6���աY{s�Y�v�An<��欜�ɪp(��&���a(e���l� ��S��'���J#a:zƚ.�A�O5R�o�U��7�R��u-FT�tc�E�XR ���"�a�D�g��<�J�Ǝ������	R�q1Z.��b�BcqmM; �WmIp0�5x��5��β��z��v��8w=ky�
����O��M��V������#�)%��h���ORW�����J���
��O)�cFB+�qKm>찀��I�هEWMsAt�P"qO|�N�`Y���5���Z�*U�`�����i �S��P� ��[�Ǐ���өZ#���w6㔜o��G�+�j�U��6e"m(����+��F���Jq�I̯tjKC}~|]~�ܺ���&띁���4.kr E�@�f�˧�{�/[�}.~BuĨ�=��}}r|y���q��ɾ�����fag(�෈��,^�i��'s̔���ܭ���H�����T(�mbb"3!�����f���G
�� E������߆%Y����ϮRmɰA�4����Q0�sb2����~������z�z~˧�c�iI��a�9���{���Yq�+�_*;:��dҁhr�p��g��.{	?7�Ѧ��篈q�RNut|���f��>��>�؅����%3�!K�)H��Ϭ�tt�J+37�cn~�d��ʩ��J��V�LI��$"���!�G{�odT� -&�y���|�4���.���EW�D��AazM ��cRH���%:�%+C��ȼ�#��ճ��o4���J<�N����VI�x�ܙ�[�se	�ΖZz�f�zN/�>��8����r�O��G�{LPZC4h�=���@��/\V"�#�g��U�r�գ}��c"���?�xg���h"xI�t���ލ|�%	�A�C��k���{p3�r��a]e��1`mVˀ�K[U�~���W��+��&�$ZQ��ؕ�Љ�(B⋲�d�`�|�<+$j�fk-�ҙ es��Jৈ��H���1�!��A\���������Q5uu�$o��GEY�<j��5$�%E��WǼ��q���3��+«+��_��"���%}�8�_�Bw�U4�?��]�E��	�����sN��~��oai���M��Ƿ	�2K5ad�^��[2�Q,���#1pV{��Oke�c��,Bмv��<WD�2�3Q�:_m��-8�����CcX�P	;�&�+�ǚI
8�Ê��HTcR�E�<0�a��b,G����? �_X�\�x����?;��O��:����[����h(��rx�������0����jZZOǩ�WF���X��hV-���]m�4a6g��JY����O�Ǒ8�=���do�ڃM���OJY��w�j���)аVU�r�8��.��׫�֍(R�J@i�>뷳�����t]�պ��e_�)n�#��������b������O�O��!����"[�<w��u���E�M���'<"�M�p i�B�w�>�+5,Z��\@`�UUPu�Õ��ˬ-w�l�]�E@������Ac!Λ9"Em�/�tC?���E׻@.i�Z[��ύ74�>b!
�&������� \�S�V@���㑕p�/����~T�O���P��&���)���(��G@2�"L�P��rfQ�(�2�ǆ0��h)�~�?��SG1��`��nn������q�o�U;�7�<=��#��QPQV��3:#�����ߧ��{�#�4���$��`|���K��A�!Ń����f�-�� ÐX�%�}���\U��-ǋ�������Ut����\�����U�,�����3�E�f��h�.��V����	e?zk(��^�SQ���
�"���]�DnۣiJ���ˌ�'�K����xWΌ
�}%l��s�{3�+��˥��ㄸ)�?im���4����,zja	)�]67e�� -��Y>C2��Y�X;� ���j{����� ������˩��'�>P(�~~Xhd�1$��?��(��e��uu�e%�`�t �qx��E�ᓵt���� (�K��Zʧ䳋��@\
a者�f�(᫑ʓVn�7�R���!(���*��*�����S&��l>Ex�,-<�[���i<��{�D{�����*m�M�&s�y��"��`��4*'֍�<`�Jӥ���L�jPS�~�sH��:&|n���$���v-�;�vw�����*��j�k#�:�2e���@1(�0�(Ʈ��>�9�º=��L�>����p�+Pjc��C�#9�R��Wp(�t�!��θ�Ȗ�r�#�<�C(���i��V����ĭ�G@3O�ų�����1�ԣ���f�#��8�ޕ��M�nM�G�L�# E�����%4ǣ$2�	��Dӻ]�'H����d��x�\*���J��ib�_����d���|!�	��35J�{?:p�������i������ΤW���G�tQ�G�'l�0\�"6��'݂����b�����������"�I�S���i"�x0ƓL�r�X�hvx�3��ㆪc��0n�V�q2S�),1�FL��c%�q�ǻ��:Hon���o�����	���sk<7_�K���z��ݙ:�
���6��#X���yE�l����X�K�$�����zE���ɢ�"��w[mtF�9��0����O��X��z��rЋRA@ŏ�Be�4�9�_�V p���sI��b��dP��T�F��S@�=Bo��<�RS-�h>�]��qo��P*�Z|��	ų�gt(<���yVo\�.� z��u_��2P����;
�� .+������m���q�1�/���d%��1�m�3Ӌ�OB>eg�����Pn����@C0S�jb1+�*�<1���Z�r�?K���aF1�����l����'`Q�6=[�eH��Eχ��ؑ��m���{�j��q�KD����F!��(K���2������W���M �O[�ݝ ,���H�� r��'�m�Xȶ�o�ZH�?"f���$��n�Ϳ���"E��ф@��D
�l�+���f���-��k��,�j
os�Y�1������x�93�(l�O����T�}2Xy[�BɅ��Ц�=�Z`�X��#��ی�)N'P�-���ܓ���v�� ���Ϲb��YT��/�(C�2!=�ԠOd0pd��G��^~mmw�,�X1���=�/�Y�oN"l�emP���63R1����R>���EXi,�N%<��m\|4z���(E?����@�o^�հ5�>N�5<���u���I����ι����B��$���E~��Dtw;��\�mkp�|m!;�m�DC]GG���}B��:���ֲ�.�4R�`��*QE�o��M1D\~yi�g}�X��x�q`��I�J�#4���D1�q��w;��/�a��k�ƈ(F2�ɺj���fX�%�������k}LE��)������{��vY�����,�h=-�4��.5�Ū�⇷n���"]+	a���|LLf�)�����5���'���Hh�rR?_�H�5cjj*%'S��.U>䖛�]�MH�7���h�%�|'S���K����d׃�S���m���E������-!�ȶ{ӭ���jzDV["g��Ȱ�yn,,}.nz��}|7r��+�d�
;��wul��;м�JXt��Y�
U��q�+ӥҖJ���X[��M�C�e�k��Ț����>I�L~:y^d�G㌏�8���f#�X����^<gVm��3a���;��h�F�. D8�ޒ��z]�mMn����\LNF 
�4���V���<�;I���������i׀��� X{*��8�k`@�K����T,��'6��W����7 T��aGE5�6C���\+c�He��Ke̲�Ir���zB���
`(�bÏ�yW���=]��|�i�����ŕ��J���������t�!3�^Sl�ӕ%0�vkƦ7�Ȫ��rE�Fu<��v��>�h-�"�޼��P��x�d�*��%�=>JY9�&[er�?��dn�,--?��c�谢��B���eUD�������1���}�%<T!4 m�$wY�b
iGa*z�+� �8R�뇑�^4��{��n�_Hm�\k��������=>̜�\ٜ�ij�x�yѺ}�j��s����u�)�pG�{��b�1b��\��D!�J�D	t��	�(��0jzzzx&N��;X�nƯ_�Y�6�k�[�F1`��{����姆-�ڋ��t'CJ2�!B
}��%X���jT��U�)�%���O��	�YC���?h��m�q�R-�q2�㭬�P�?�`>���:���a���ub����M�.�c������ ��� ��l����� �$\&ٯQ���ҖM��tK�GGv��Q��}�8D�k����tt	a�_��/��GUn�H�ܒu��~}��!�QֳXm������'O�x���yDT?�:��Z�� ��sr0��,p�'f��a���D/p7�����#C`�9_�qɤ~�~nv� >��U����CuKK(�I���|E�������4�5�o�5��FX��F��q�7g��]����l�lYߔ�&)���d�i|#��R<�j�6���Fklj���B�HEU�Z����-����I؎��*/����,��vm�=A�!�f3i{�?e�������aP��➛Aa�;D�TA."b��5S&h|l��7� ���u�t/w�[n����7�DK�2�~H6b�f�������0u��+E+}��eV?�Gcy����X�A�궶p����RB��eG�j����jq�����Q�⮭�M'"g��� ��h�ʰ(��kb��Ap�!��A@�A:��Ni����F�[@�A��ޙ��y��e�k���}�Zk��ظ���a�a��ӫ�Gt������h���?�;�?d�?���j|�{{ ��}g� �L�����>J�Y�;���RSGgng�J����F���_M��a�yl6��l���������?~-�Li<�L�{����-���8<��Y���h>�*G��Ij�H*6|"�|a����\��y��Q���A�D���U����/�����_\]{��fg�-/V�ܶ��~&����۵`�5|�s�`�������n̿~�ᠣ����J��h��B����̅�V���t=}����+��^�Xq���;B~�=�y�Swr�#5�sd�kAUL.y����~��B,�Ŋ�UT�� �K5�y�����U�Q��/$Ϥo�F@�P�nVs���
�EDD�7O޿`��Jh��aJQ$srF|��w������ׯ[k�=({���p%��]�!ja�����Ua�z"�b�qi�xzdL�"&!1�"�+`�%���=���搛5_
��UQ��"�_~����M��~���3�q�B���O�l8W��GG��sSz�;�x����̒��`&���������0-�SG:�Ҡϧ?���5�A[���l�@��O�o>z��ڕ�L��D1j;���c���m8CS��U����W��M�[:��h����ǝ܍
�)q�h������J�ھKqe�br'M�S�/[to��(p�[6iGcap��^Y��P_+����w��9��j�j�h�vF_�V���������*22�-�w����am�#��*v, �0xP',�~\�[<=K�:@x� F��:�P s�v���xrRì|/($��F,~�̴s�@��Wa��$/�����p�ˮrIH.a`1�:�}���E��/����������� )C�r�[�����F�M�Yߝh�ÿ*����>5t�����9�eN��j��Wy��DD@��-1X��j�r��RLD�Ӳ�O��-�5CS[[�h�h��Q$��%���������P�@&���e*�[1��e�dɅ����(��#�*� ���6�2�T�?�a��E��A_\�u��W/���XaSvt)�'e!�c��;�������ϙ�tʝ���>k�"ng��\��nY���U̊�[C� .B��'��璊��Bk⧝�2%Fp�������ݧQ��G�-���Y*%}P)@��4��gTġ��C&�nֻJ@릊��yG6ԚCc^��y��]+�
�%��=*d31�� �N�������}���E�t�*���]���t�45qW��~��T�l�sc���������BjԦ��o�=i%�x���\1�3��?8��̱�T��3|Ok���Z0��Z��Gnbb⺆ځ��SX@^��_�NN6H����Xf3�}u�
��B$�&�eQ�DZ��	=S�P#M$zQ� �j��!�Hn�p�\�V����(<7�Beq���i��0��/������7�U=�X"�-����{86L	v��^�]�3����n�'*�~�w�˯�����ј�,���|ԕ�J��ܑ��4��|wa������oKw4��y$?���Z3g�r�����o�пB���'}A����~%<%�j���}m�6�S�W�&뛻8�u�e����~O�i��og�>(�EI�mj�P�4D�R�>�'e��sRSr �(ӌ�7�duH�le}�" �� ?��׷/��S�����S��L��ZF�x�Rj�J���Lh>p����$RPN+�2�uUUi�eɓ	?�3�n���ꢥCJ��6�jAU�W��j�!��d42�"q���;�A���w���5œ#���E�
��
k;"�zs��s�Tr��A�~b�0QUF�����ϵ��Ͻ>W&���K
 ����M��vo��ޥ�v^�{�C�����/S'�k)�F9��P�8����l��\@h���<�O[_����£� I�b�ލІ�鴺�X�b�L�yI"��	$P��ֶO��L��#>o��j ߤ�J��Đ��-���Z?�4��I;N"/a䪤�t������h�pUZCo��b�<ʛ����@�yc����2�� �"�B|͆g��� ��=^	�����c��1�y�Wwΐ�$,�mR��o٩3�W{ЋO�+£�J��NNU���̈̆��w�������T�A���I��}/�M=�W�%[{�}w��{�q{d!�=uGC`������q홮�<�~�g�3�H���@RJ�Ĥ�1�b_m��/�|j�� Z>W�7�I���G�^�J7q(f�d�L�v��v�`|9�= ��+&
	���<�:�M�P=�S6�-�YewP�'�.�ˇ0��Y�Gcy�Z���|S��*ϩd���g��P��F��"�$d#2j�K��<6�M��PŲȒ�r���C�վ�S�ٟ�v��F$>C,wM�bG�Hw��>5��~sd�S�k��0����ť�[�6t�A�D�Fp�lmqso��!�����#x�o�x�"�D���amw���;Z��X8�I�6�M�ɢ(q��:p��?�B]SS�'.\�Xr�i�h�'�&��D>�x?��{ �p�俯gm�Wq8ҟ��6<�X��"m[Ic�N��5G�"�nX�!1G���u�vMpί�]Z����?�J�S���5s��rCv��MGH?B������j�Me+`(�Vٝ�!��:�Ok�8�^h�DJ��	�e�;ѫ\��e6��*��"L*��ϝdl�DZ%'?��vNW �ݶpᏎq��
�ψ"���]}�^�Q4X.HSН���f�B�Լop{��%1�R6@f�19xI�N����}��bl�[p��NKՑn{�_ή�Qn�٘Un����F����jO-���	����3oJ����L���Re@y��-�,Sm��>��n8�ZeX�)�k&�Ҩy���|�@��j��G��m�ܾ!۟���"K.2�ƧU�	�#�g�N_������%�[�
����*߲8Q�h�s�K#�F�;@�k���8�i�s�%��e�.�ǌ�h��g����b��+cI"�g�}4Q��"㶱?-h�{MGV�8ϒ�)��hM��W"綾|e���cD2�{�Q8��241A5x����U5,�p��p<�.6��a�@�vX݂H�a������ق�����Xs�mLf�G� �ʣg�ش��	MV�5	���{�2p�
�T��I ��&���-�f�&4�����c���A!&���L�ݵ8�F�ni�� �C�
|SW�p�\�6;^[�]]{�a�����lӯBL�	����C(�fl�D�,����:����#���>fKi�$�����K�1��!���1&��7u]]1mO��r��u/�6Yv��4#�@��>��n�9l�
8� �w�K/��]�����V�c2���քe�� M�[��N��P�3���"�G�Q�Z�튕Me�G*��H�R����+t!�6��g�qP���9BL�����D0����[ ���'�yk��!�����Z.�l�&y�&;D� Y���G�g:���+�� ��*�]T�����?�㝅A��QV��f�4jϯ�⚹�vDS*zP	[c�������|�����J�ì��I�$[�B��PIX$<��1|	���M�JC�1&U55��9���;��?��|Oo�>v���5�����#O�>�Q̩G���u��8d�����۪y ���>:��wW��j=�������]t�Yjpd��<N	#����t�sI�^/�[=��qi-�S�o�H�d� �	�r������D`P�y�K�[��H<���.>�,i��98��%�" l�}���[��hT" �'�����K�ð�q?!��U$6r\�^q���OM\r�.zAFa�ٯ�*>o�z_�m �濑����9	vL�������zA� ��t��B\�P���hʴ�
�=K
�x��X�`P&��Pi����з�˕��L[�ͽZ?��-l<���㶉	g������j�$��>�v�]h�E�J5���^�eu��w^&��U���E���{��88p���po���:})������"�m/����nsNh�#�t��&�����w�(FZ�k�7��4Ƒ�+�
?(C� 9{�	 e�|��D���O��Mث�VT�%�}�_3\��'}�c"iΌ�Q�X���o��/�
A)��fys��m��U�5�A>��bX�}�Z�S�����C�R�W%���(�o���=n��"w����#���t��K��P��m�Xe�a� �r���a�YѼ�19��]�u�ba5�{�f[[[yBS�9�,Ӽ�4���?Sc���EVI�0�7!�5EVX�iVt���%UH_����q�V7�/����5_��p���k�[fV�Oq���)��?F�$��J�K���_�{g4c Y��}]�fi�����>lF�����U*���7A^�D,PJp��.Q��S�`tm�U���.�"����O��Bu��v����?WV��.�L���f�u+�D_Ȧ�f[�$�}�-��h�DKϨ��~1�,r�:�q�.1+Ǯ��gHg���[�>�_on���d����]!�h_�q��.,.#�m�9>��׼�f�� )#�����O�X��WNo6�u��mW�N�3��+���;U�_P&�	�֡ ��<�*;���ս��g����Q'F?}ɱU�7����`�z얕�pM��a�b@�,��)���.�C�Ȕ��(��Gu��<�LMP��	Hր��vq_x�d_���b���"vz�vfI4��t5����Sq�;�Di=cJѼw�c��e����E�%����G
T�'�8�d�6Y(��
-d)`��N~����)�j�?~i�HAV�X �vnB<�[��
˲҇eͮ�J�z���!�����9���Ff�ҹ^�6��g[�SK�9�]��][ԧ���< i�\�/���o8�1��:E�Z�Φv���sP3/�J�����şU~�c!���N���F����3�e�����X��\��XC�w�n�!������`��@��n�-�,㳗[��|2�ZD����	��Q��Fm� ���
]��.m��a��v-"��5[�\d}�A�\�N�r���p� fi�3�-�=�ttt�.�-f�Z�އZ����l��/�\�Сisc��i��� ��4_��E Qb�W�Nk�I�C?7$4��&lZ:�8��,�DK��]���]�a�#��^?���FX���%��(���Pl�]zn�ؒ�<�(�)��;C49�,�!�"[v�hl,�wφ�o&q��A�1���� �=}��ɂg���Ƒ8�|-Dz#5KČ� ��w9O�W��]F��ؙJ��*OF5z{v�������%C���$)��;�*�&�|uabIU�Λ�[e��%�|9���8%�]���Ϧq�LSڏ��>l�=�����B�6\�M4��U�R�l�S�=4RȎ<�R�) �N��\pVQd����{e��B׮��/�e
Cq�*�]{�mՈ�����ܙ=��>��t��@,0(T/m�� �$��{�����I$f�D]nN���w��A�}�R �(m
9NQ�C62\�J��j���� Q�#��7�V�S-�~�-;���p�(t�i��p��^[z���ǆ��C���ѱ1�o�äI͏9W����o�����P�$žɗ-����n����t���7��a��Gc�u��S:yOo{�¥C��F�������}�G�g�뽓�['���jFjh�g�<e��RsD5�T@�l���YV�%uu��a8m�5��J�k�7�
�p����\E��G&�Ȍ���n�k�:f鑈��R�������+K�=����k���m9��X�aɟ�Ã.F�Wx�n��+5�geY��C<��/5��-�P�0S��5Ny�q�r�@$���^p0Z���7h"��z��bix�����{~Y�@���^�(X�NG˶|�ܮ�r�c̖T(��̣ٵ�km�����uT��$���v�������7=�T���S��V	���_p��;S��cT��������Q�S�>���9�D�|r"��h�	���l3*��G���l�����Ut(�x��L����W�|�O�f��M6O�AFr{��|�����fIĞ��Z�eq�ж���	��o��\DH�����YX�¶:�F��z��EO���;d8���)rA g��[c[@��:yb	�����b��+�0���zr��e��B�r�y#f"�
�0���H7B�՗7�lAWV����X�"��^��sY�}䓞-��3k:p��N��ϩG��_���"mD�M'��_�ӣ名D�2�����O�C#>��n,B�o�H@dR(�R�P遀�8�p�f\��&bJ��?ifL#jT��!?��sh����l�{3�C=j��X'$,m�+���;���!L���[tg���!c�"y�7��e��g��'��C��lG����!���D��I�l]�L���
��-Ġd �כ��0.za(N����Լ9��7���(�$q�Y��S���C�C�="q��3�6�<[��bq��4�����%��sv���s��{��^W3�̶jN�P�T��s�� ڡ����@��1�M,���Z�z�C40�g�'>0��S��~���%�c�3顖�(���.����S�_���c쵼�*P?����\���R'z�j}�9��h��p�4�k���;��e\�]݇/�ri�������\����W�̻��e����:0�a�JD���R`ځaN
ۿ����L�>�/�O�RA���MCͥ8�pB�s���?w�֏�G�HH����[ɩ#	��}��'�{"��6�.m�=�U��R*�*T��77N0*�3gi]�4�)���p��~�5I��Yƌ��?�f)�U��^�R��$#������?������G5�����Q�R���zMoTi%0ee��?���{pp�?T'Q�>�mkJ�$��"?�,X��ȶFJk
�k��V��>��8"CQ)�,�3i�%oD��c(ItK�*ȵR�.8(���*Jj�-��x���s}+}Ye2F�z�l %=~U���	~Z�A�ce1������2J~���u����-��k�15��0��#[u�/�l*>��q鮽��Ѥ3{G�%�Kz�=��'S�-'t,�u����>�T("�E�f��H��B�1��g���/�k|R���؞��py9�p3�B%�rL��Z-�����^VB�Bk�u���J��1I?���� ��i���{ޚ�hl���=r����Q�Y��|�8A�i%�"�����3�&ҍ�ih�+�v�ݭ����������֫�D�0�6��BcW�ԥR�:��S�
.:�D��͖��{N�P }��27��OV`�*f��҄����ǘ���I.x7����{�z�a!�� x������B���uR�3V�Ea�0릊�X����Λߞ`MK�?d���"�}8�Gd�;;�}�c���Y�z�]oy��ɥ��[�(�A�v�D�f�T͍�`�J���c!�ɉ�^�x��1�^��g�i`)&�����d�2�6<к�;���Z��4P�ŏfT�^�e��x�� �-/H��m��ݮ�>pCk'���zZʳva�a]evM�F\�S��QٙP��x���+�F�\����^Ȉk"�X���������?�*˥�y ��]^8�K���W4�J���/�����5�I|���+B��[m�<����H	��BjH����A�<򆫎\7B��A��h�*�s���MBfmE�Tq~9+�_xP�Z����������vȤ"���/V�I�3C���KۿnL�%��5�=A DNrp}�^����|�t���}X�џ!���>���{�n�n�X�����t�Jx]w?��^<_r�%kք*o�Q��ya��{9�UE0���DMե�"M��Kb�B�"�1[\f�ũ���K�p�
W�->a:-v��ݑpD�a@7��v����H/9�uw�jW����q�a�h����(_�C����mUAQB�G�
�ٰL��g�Xc~˪���0�׺�}g��E�r�D.A Y�h��u������"�4��kX��wh�6���g��w�t��?&���Щ��^)�
`�g2
�w!�P� 	�^��d���R��������~�c}@���ScF��l��lC�9a� ��)�t�SU������֐�����+�4>�6ˡ���'M=}�W�J���`�H�~��D���J�!���r�W��?��8�=e}X�������-�Z������T 6��T��3�

��B7EH ���$:2�����!O��x2W�5=�E�r]�N�AՑ�<�Y��w�ֿ��M�Ʊ��|���~6d�4�d��u,d�W��q�m<�c�e��7�ec���[��w>�ϷB� UPOPT����^�V�JlIt9v�9.4NgJ�^\-�Q^�2��ITM�Q�&�:��V)�����d�:�v�i/�0L�=��u�`!�8�R��"ݞ:�j��m��H��H*Y�#W~` R�i�́O�?�f������&VZ)>���Jϊ	8�`�?:��Fc�-rL�*��U�����%W�i�-���'� H_D:@�Y��i��a޲%T���	(ʃ�R�q��Z�S��_,�=O?�I�a�-@j�d˧i��7�%"���CFg�M�ଊ�/�h����t!�_=v�FH�[ʿ�L�
������s�|]�efeUL���'
nl�Yc������H$<���^�A����֚���+��_�3������X�E=ޏͲSg�Bc��j?�͞,gS+��7���2&ER�(,0���0�l^ŲZ�5�k�w�|�ѯ�յ����f�L��e$������R&������OL74�j�j��Ot�6gJ��	:�0*4Z�s�E��h���߾�z�����G���
T�,M�_LO��Y��y�zް���5Nm:��C�:�t�1A�B�v�su�Cŗw��=���^�:�J��Q�Wz�AI�_��=���c4�xh�~`�G�G==�i;���9xa�z\3���`�>����'_ K�U󾛲� ��3&t�3���X��>7$Pb�5x���a��`�tl7$�������xH[YV����������d�$� %�\�Io��������r�@��I[|L?$��ʨ��\��JLL�T�z��HB*���κ����1A��g~�~�7b����lllz�pt[�ّt	�خ�׵ t����V	���j=1��F�c�MUm�X�R��Z)J:KI����I���O��b&_y��ӓ ϻw��x�Hؑ�e�+�àl�ε�m�p�ҷ�9E�q1)�Ԩ�sJ p���� ���sI��"���A�*n&(�P��`�k�����ڋ1��P9���3��v;B�N~!"�9��7��LLu���D������>��sU�9$O�D�v%��6�,�9�*U+2�I��Md�M�x2�e�aR�O��1P�p����y����$ʠ���Mw��--";�{�X^�5����긅f�N��#Z� n�9FR&�0mK9�NF� Ȳ��NV�� Շ�����d0�J@��� tKn�:�@RBIh����9h�|��m�qn��d9��d}KK��.���RWH$�d��l�c��$�8�!A�2�P�< I�p�1��g������MK�mܟeF��#£N5�[.��:O��o���c�" �����R�Hv��N�P�N#� P[
	cVdT٠�V�!T$�_���ݚ��$n��k�Ӈ����n}B��v6vX0�b��uА�'�$�K�PK0�F< w��M�6,�����8[3`O���Z(k���/�o��/���Q��IFU�� ;����蓘(.��o��R��=��y0.A<�dX�>����D��Bz;��KG]�k�ر��:��ꍝ~8C��ŗ\���0'��vX��<��*����#1�A����<��T�B��:^�2F����Ğ墭Jݹ���Q��+TE"	{F%r>5e�eaF���i�wD��r�另4ܤ�1�eH.�H����`�R� ���|�c��̛�p��N+����+�}V�J�=��:��%�7�bi��������h��ذSYu%�Ѐ�����|/{?&0�7�5>���~�럋�� ��)�rPW�D����o۲� ��*�@�P_�u��v������
'Oq�X|���i����ŹN��A��f{�U��v�z��L�Q�k#ŵ}�G<c�겂(q���8�U۱o/.Ȓ{�F슬2@H�}h?ݟ����p$7b��~�T劥��%+����4ƧU�J7�^�l�4@*W�!�8�ǅ��]������	��R�3?��?�WGg9�W�G��@l��~��5R��sɵ�D�;��vF-�Mp���>/˝�%��r�)r���C�Y������љs]��|y1d�bdhff&��2����}�(z���n3�%|J7:Fr<;�~:�]ν���2/Q� �0�S�/�ׁ\��0��\�=�� &J���,��@9�����ӌH��Niג��_�p0�\�D1���B�ɜ�`���IW��x�;c݄ha �|�s,�!���J% �%�,R!�7��s�6}�;;*YӬCҏf��
�H$"�]�c�<�릐y%y*͘�C`���@X҂��� ��`�H�dpc�GFOǔ-��6sr��h@d�l�waOD����B�E�� �ˇ�м�;�W�
V��a(lӢ�'�.9��ڃ�F�&2����v\wܦ��B����E���! ��[�����M�P����h���z�`r�RiҽjZ_�F�F
��/
t{�(�;��O�x3�B3��H����_�ގg��#��/�}y�`�9�p$�G��N�(i�S����Z�t��t�������+�~0�����D����7y�˫8�8�"�	�A�m�E� (�,(�l�&=�y�Ɍ�<�\�cR,N`�4��5:��mȆ�_�5�|��G)�N	��ɝ�^���_�B�k�����9�0�L8Yb���sD-j��@R�� Su_�|�V�r^&^l��G[���F>F�˧�pr��Xq�:B>�Az`>0"Ic��*!V�S9v��>�����,�n0�g�_��$�ˉT����BbS~4%$Rڽk@*�j�n`\ɼ\<E���y���ś��Zr#^e�)F~O+��D6�4��.��xI�M9s��u�.T�D�"�`5��7��8Wj��������F�\Q��Ѓ�y4;ʤ�H�ֶ��{�{��z�p����h�<�5��l��ևS
��W47*T8"���/j��m��A��,{{|���g��Ɲ2��"�?����#�Dh6C����	��=���ZTF9�X�xGȊ�Ñ���l@z3$K�Ĥ�B(�j�m2N�L�����#+��jH��	胆X�*S=,[���}!�"
�����R4H�l�[�,r����,��$
�=��di>�72�������t^� ��Γ��.M�G~YBA殠�E��i�H��6:�� �6H�{yQEr�>&Ф�����(����H����֛6�b�-�K�������7�/T?t1�!�ư����ͦѡ�����,��]O-)�5�JA[m����\�O�	�E�S�'η�kwپm_(���26욅����e��Ĺ�9�����AQ�Q�r�/�O��ER��(L����$���20����Xc��и���N���pP�a3��3t�S��Gw���SwtSd�������paP0ŁiV�VIuEm��!G#!���Q-+�<�)��7�p%l`����T�|��,��!l4������T�bQiH��5�25�`ҁ�{jKZ�f�z���s�L�O� ��5�����!�����Ͽ|}�}�F�T\s��m��0S��w�������k�ш�b`�Ե�ŹdV�Z`�6���`���dܥ�A@QJ������L��7H��\�#�X�Q;de��£_l��%b�麿�0�P��a0˛����a�����!f��ؘU�p�Hg�z>C΢�e8������Ȓj�SC����dp���*�>���NّE�L�+SaLaq�x6Vp����xU�n�������gx�i����~�QF��_|�����<���sN�K�|���E�h{;7jZ��y�'9���t����D2V6	0e�U�a6tg�aJ�,��!�J�{��P�KE�4�=U��wC6�D�2�
��R�p���o8QȢJ��U�O�l�r��PYΞ8�H�J��� $B���<")�$�x�+��;:����QF���E<� -�����u��Y��4� �����=-0q������3���+���m��/[T�����(����F�M�ا�6a�������i?���D\��p���v��HJ�;D84���>�!%ped�y�Xu~mz��-��[6SCo4�a  r��#�s����n�Q����/��愵	���1�Ž�?��HX��|[	c��^�-Xb)�(_��}2�^���Sv��~������L�^�a`��2 a���+Ӵ���$fS�^�b>�i�.�WPs�3c�^��w�`�n�J��B�	{C��D�E��±�FKP^���<K�*�����$?2z��D��Ð�cR�%���Wҥr�_ p�˙�
K��^v'v\a�z���M�=%@xwJ
���/��'��Q�%��i���D��nc�楧�*�><u~�3]�ۻ��k�<�٠W�v���Ʊ�6,��5�a��_�@7�5i���,�1�	�E-�%E�7^�ɾu��N��8-��\�r��|:�y�a��Df�9<��[�-}ϳK�����#���Aր�ě�#父�����|���Ur���w�ǻ�)g?�}�Cϩ��"$DA�Vq�No�>-�:9>��rZL��|���;XR�jJ��~&՝�a:m���70�ñ˿��w�0��Jn�pnk�=�k����Q/��.�q�3�;kcG�čq�ASt[��L!3�Zߤ��d��σ�8��;[�_a����05��HieG9Q��P���2zoE��w�2�l�"$�w����7`� k�w4��s뎿c��^����'�?�,�֤A۴�IrU���G�B��M���t���V��l�m�3-�w��J���&x�˾�o����$��" А��7-mmc.���2����w'���L���>c �
l�I����;C��l8��J
>�}��t�j�E/ECcZ�e\��Dn#_�����SIzѡBDD4HG��s�!��Y�D�-q�݇������*"��7Lv������GU+�AZ����%���%đ'�?0��zfV=�&��(k���F%iU׹/�K�/����X�u�t���(afe%1rԩ]bx����S�Ūe�c��vC�gG��c[	-@MU��<�"	�5���:��
Ax�4�������f�� �V?��A7��K���绀���t4�oa�s�i9~��Ey��%_��ϡ%l��Zs�ؒxN��t�z.ݷJ	w��:7�j�f���;�屁����~Ֆ*���}F<'���0�c�mDX�$�|V�b��w/�i�,r�K��SV�}��5�C��g�[V�g,AC�[�i�:��Vj�dB}�=DU��%:�L�q	��Sr�J=5��� 5�㽖+������S�ے!�;m�ۂg)��P�v��Okv�o�������ݿe���X��,�Q��.�����GF���(�߯�1��s�nC��-�.�!��I1��V+��@v��Έ�;���_r,a!Q�j�fز�Т;�`��$�m%�}����=�\����f3�͔���cy9��\o�Z/�S��K�O����Q��P!�5{�bbh�^�qJ,`D%qV&�*�;�2o� ��x����S���#5�Pb��[��`��j��߲��Ś�m�~@���nT�%�}5�����N��(b��7ƺJ����wC"��g��}=o��2H�%�Ӓ��$�I]՛�ī ��N�ɤ%��>9��Y��$��91qLi��Q�f�Vڊ��*����5��a�&��G��yfN���tW�P��c�p�B�Y��a�իWg��l�w�Ok��"���i}�U���+���ׯ̲��Ro��[kt�0��;l3Jc6�Dҥ/��+8M�^0Ѝ�j�_$k��U�"V��/�)	˪�9�k�5��4���L	8i�t�X[���y�'����\��|/}4����h_\�\��4���}b�@���"��Z@Z�R&��F�a�Y����"YŕK�/�Ě7e��P�Zs��u���2tq�t�Aq.�I���b[�g��O�Sl�	��^Y��|u�a��GV��~�z��5�I��!���2����tk	p��n�0 i�e~��Pj��E@w�7�%����P�"*�U���y*}*o�p�����I�z�0jX�G�ߘ��5LjL�)3�DU��/���i�Iy�ы�OgBZ���Z4�{V4���F��K���K�b;Ҳ�&�})0�8�&����\b�S��L;`�,�	˳ȋ0i��I�`�Ֆ����u��5�+�������D����2u]01��Y�f��7d Ҝ��?I^���87MWxɨ#������i�4w���W([c��,�l�%��^	� �#k�E�j����
 )T��f��=��5
����z�'���Zwl[Ύ'��=���	yr���m���L��VgR�Cr����YQ�
W�o���VZ]�4S��d�l3��ڴ4M&2ט�ᾬ��!)��t�s�U��s��4�=-	WO����T���dXJ���f>���3�4������kA	Pf�b���y��Y͗���ɟ����9 ɜ�+�kV��/�K�hD�D>���j�s���ǧG�Sj�Z↫C!���F����Q���� 3�p�vQ���bۚ�ko�N�Ǵ��Z=R����~�r�z����ޯ/��ʗ�fҌ�k(,�t���8d#�����~�ɖ�y^_��tJ���{?W�g�V\�/
+���Տ�^Ta*Ǵ�1��T�4�%O�ײ3�`����5���fABй�e0�n�48qY=�-�.S�e�#s�1�\,��u���ڞE=lgٲ�V�
�Me9�X{�xx�z����?\�������p+?����g[s�|O�l����u$�&�4Q"�����|M,l���\�_�4�P��Bb�X*K~S�z%�$uH?%��җ5�wK�����u�)�3F��Ke�3��)݁b�GEC����MHݣ�tR�q�56�v���7ɗrK`�q�?��K͆qE�#	� �4�ʨoa��z��$�v�ٲonc�~h��NA5�U�l��A���
�L=M���U���32B��Ȳ�ۗ�	�'�/�K%&<⢬݈��M�דa�ZԒ]��6�=.3�*�ҧ;����2��=y$E�n��bd�������0fޡX�
G�׎a1aפ�f�f���$����|�֒�"2T���NxolAɱ�}���>5�2TAeS��'�K
&&�7�ԏ<m��N<��7����H� �F�ԏ�����{����I1�Ѝ��~�1F��%ܴ��Q�8�R&�Ǩ~Ȉ@b��ǐ>`�o*1��X:�i��\�����%��	L���7d�8H�hY5���wG�&+)�3�s�eY}�׾X-��3�#�� sVn�^2=��`\��h�a��d�A�8�ӮN�_e�,[����i�)�=�~W�t�b�&����N�GA��ϖ�sFf.�^q�n�-��笂�_g�Z
~��n�%]�q��/&K��s��(��u�FYB�m�ی�-4a�̲�w+��erϟ�·�<:}.�Ov�&��%V`п-rV:���
�^�O�Hg&���,�A�:8��U�W�55��6��`6]�����Z�φ\y��]H��4��&�a[��+WR��
r��\������'�-akC�(��9`�/�����o�W�����?o��l����垃�G����� DE��u��@	CF�����\޷32\���B���\{���a�A�OŪ̷��tQ��[���U+���@J�l��V>K�QMg�N�h��tI��H͆8����p#^���_�ֽ��E��5Dl��MD�,$(�)�wy\3�*do.�>.�=�������'\��c����hMO+�.bŻ�؇H��|z�I��y��o��'<fa��9$�:D�������Ly����C�%_c�4��^r���C��ɕ3I�����$�K����~����������fξ��+T*��
��I�'3���2r��>1��H��JtC,J��(��3���~�_ D�����S�}��n���L!�_�ޞ��Ͻ������t��$��z+���:�~U�4ޣK��np�Yt�p�~����4��Ճ�&�}��p����k
��o'���⋐@�1�ec������Qm�K��R�b�)N�R�
hq).�Hqww/^�ݡ���5���]_������ˏd嬬�s����{����T��3��t�2y.�Yi��Usz�)�(�uas�?BlU�Z v�ِ��볁2�α��Ǩˏ�M���� �U��D� �_����t�S:7��|l�6�/�M�~�cFy{�  �SF�d���'�l{ 1��f=3�7'?����	YQ��״��T��S�D�ZՋ�{��闔����N��¯����AR��HZt�Wl�]/�@$�=�^�~PI�UX]�xi�+��)�	Z�U�Fn�����=Ϋc�ȇ�\�3�j�x�hy,�2w4��uE-�$J������3m��5c&��Gx�6��&�ჶ^{:79��9G+��e[�����ݘǿ��eU+ᨀC!�����:E��`n��${�_J9VO�Ncg��"glY{.�}h.���r�(����������e�z�l���*�B��k��.b�4F|0O�������sе��:p�О:r$����_��RCx@u^/���@�A��&oO�i��Pۄ��h��k���R�쉨i�(�W�I������m�ṡ�������RVL��";~��!=a�V���M|�T�]����h����v���X}�]R&A��F�:�L�Z�q#�d�좂�����_�ydҖ�,�*����357��$�54�Ե��͑y��;9�U�S�b�౺���_w�mS��Q��%��0>�I��d��/���X:Nd4Q;T<�TLBd��L!��I��c�@bys-Y�e�6��ɗs�����ޫ�m�٘�ɢcRc���jV�'�Y�7�#f	�[ք�y)T�Ʉ�
GEz�Nw8�.�=�;���!��䪛R7�P)� U�Z����1�-nOq�H���mb2�.ծP�"Spro��~�7w;��ps^$*նT8�;�i2���IWT��������W���ձv�i��΍۩��r"ï_;��̐���8-���fAdSvtآ���y��Jx�[��_��,8m�ǆ�ɥ�r9G�#`��^��i�S�(��j�����{T~��ό!#N�7�lԥ#���������|���/7����)|�47U ���V�k���£�Vh����r��2�+TE�yS�����)W���6�x~"��X���\��.{`��L�Wb)��ڴ�JhT���|�<^���Xn�!+s�G���F������p�P�����9����q���rv���p�2/����rZKF+eH�D)��$2�ٞ��#Rr]ZA��{?\�r��^���-usa�������!����=%�q'{���z���}�� ��K��1y+��@�`���e3����9Ww��*�Ԟ�6��o0�<�����P�ޅیP����!��2*�5���i��,�j��F$���"���"�$�F�u�};��\�p��9�m��2�8���˜�r�u�	��m�ttJ������2}����`��Li����]T�jъ^��&��|���Y�e,n�֫�!4����Y���hN�� ����ԛ��ESk���D�E��_���Tשa
��%\T�@���������P�?�Y���"���3��\�g��A=�b��	p2y���w)��h)o ��ϖ(�{!����?��c2E�?p~�⤥����aM.�`F�ם�ķK�+��W���H��+��"9A��s&W�nY����w�斢gX��,l�t�H�Hğ�){��<���u�:�`z�1�2fTo�yd-5�Ť;:��]�/�c�}������rJ
�� ��v9�����+u��Zt�vu�.�~�[��9&7��Mrlr� �R2#�����t�T�,��ī������aJ1��U-�0�r�?�L��(p�����~Im��B��g>#xK
P�9��5����|���2�
�'N�3�hk������軼D}��]G��?]V�M%��y����d/��l�%�FH�_�Eo�(@W}<��3(W��
�5�E7�;g�c�sf�'�}�7>aT��38���Nc�7`hH>�'��i���KOM�O��jԟJ�{AXWғɦ�Y�Ȇ��ؙ��U���`��kyr ���A���٘ыQ��.�<)7�%АW��7����R��C\y$]:�d<b��!ʔE+7Ih��ޒ�����<{cp�1�Dq�,��s��5��t�E��_H&�6*�]1�U ?!P��.O��3Mh�KX�bD.�ݷ	�loQ;ny����i�O8����z�����$�DSnͮaS��7;oj	.�y�����D��.���!nSM>B�NacO�T����T�I?�| '��p�U`/E
�G��Sn����݉��n@��O�б��"�$���(w�*sm0IA�l��&���鴭#e�ۅ�Y��F�Ut�M�D5��1�T�`d�3C�C0#������3G��u�*�BE8��e�뷣12@H�4mv��5�Dو�o,r�����Aeb�����D�v2y~%�.��kс�{�G��p6�7����:�;<��yy�$�R*�ǂ� �[���^�zEm��t�8#���uLz�������(�n焸��<���f��U�9�D�./v]����9:	��
O�"R;�����b���y=�cm�4R����R?[����cۙ����Q�>�t/�G�c�ow��]��������9�z�Ü����4�ޢ�V��j���t��9�ϓXS&{��T� ����Y�������֡��4�ܰ���M"K`n��^��P�_�\V���R��5i�i�v��aF����_�]��ݿ�L�1�:d]����E�0�2X�Z9�@X�D�h��&Ǐ��� ���z&�A|*�_�3���C����I?���S̱��%tV�V���3+�ZΔi�=��=\���#�Q��U/��slջ������L=�9L�vn�ȓq�(3	ۀ�.,��B�_R�K<ޏ=e(q7���O�]pT76(����9,��{�<\Tz���)Z���WpA��'bm�x�8�n�3�Β7���:�����.vxn1�I<�Ā�����;�L�rD�F�*t�aƍME���{�p�qT�+0��5�����	����"�fV'G���{b�O�ﻥ�Up˚9�t�햰HF�Y6aIĕ���/�����2-����F��t�{�g�^��l@Z.�+���mX!@HΌ'0x����ws(e��n�}����# ��� �N(����z�t5��$&_�o5����i.���,�I��^(��Yr���� �:pY�:ZM��Kc:��ٺI1p��9�j����{vBf褭�k�wy���}.�-�@��+%:��W�(�y�R�(6�H��|4,�[%\P�� �z��{���{s�'Ɯ}���p�x��.5�7�+.6इ��"��-���઻������:����.=���E��y��)��������'��(�D��M~��2�P�����yt�FvMq�iC�af�	t�mm�#c�)?���6VWWo>�گ�;��r:l�S@�Pl��_�v$��Gt�<�h;{����	��TY�Y��#�!���X�eݳW-�{���C�s cw�O�����I�nd9��m��E��kwd;�:��t�7]٫����Dgɵ�Q�
Ĉ��O�SS�3ڪ��3�2��ŷtYE2�t��p��U�fP�t��#������-���=�`,�4Y-�T�g�/ϸ3�	����C]<�>.[�7��f9�Ϣs�b��{��3c,�)[�Q/�O�6�40�#��Cv�������%��i5��֞!o�^CJ�����1��L����W�
k���e�w�K�u�[�	��Bh����4l9��dv�l��&vn��(eH�{޻U��5G��.�70{K�Ns%Bnp�B����yG��&�G���{#�kQ�/F��G�����:[���
3D}��;N�~�E�nl=&R��:jy�p~��3��/�ܶ�*���T��}1�X6�f�+�H�y�ߕ������*���;�mz@����K�SˏM��5_�����X�\�
|�š~��:��u�pD�Ԅ��|CYs�ЎZ����$F�+O�J��w�ϣV�
� �ܚ6o�p��^��w�^$� 2{G�̯kyh��B��{������w�kg7c�ц�]9�2��Ug_\RN�z߷GdE[�T���u����Mļ�l�5�{IG���/ �����q#�����^�M���������ݑ����̓�K��2�|`,h]:#=�xO�j�Y�R��y;���s�;ʱs�� ��]�E���)W�zD{�H�~�|<ݹ�Hrr�YyEuA��7YW��¡A��s��8
z��TCRثkjT�����7���5�It<{N=&�*`>ΔJ���A��"�����AfN�S�����=�z*�����Ʌ­��f�n��;?�p�W�L�'��>�7��}K
�2)u��E�C�In~{��)
z���P�%��|��$z�&گ�ط�B�\���xM�y������a��Q6��l�,�t���7�*O��m���&Trj��Xr�a�$�T�0�D��jdí��?�z���GE�Ӿ�O����T	���|�i�b�?$��A��A}82�(<���J�m����
mmm$Ƴ�榦AN|P؎S۾���0�zm6:r�unڠe�55P	'��+�A@�F%<����SG5�6{�y��"�BB�?6߱�4g���sϩT"ݽP��&|ul<�5d^fԺ��l�����K2uOa�=;w�Ŧ���h� sv�3ϑs`�vt�of�oP]mgBxĮ��f@צ|��T��y��ٵ���Y�Hw��_���~	�KXI�gHK�(�23 -�bz�gR<�2@��>2�G�?����ux�i�+�ND[�N�zȕ��!S�B��)++������B\�� J��lX�"������1kv���i�I���L{�-D�u$wvv���s�b�4�y"o_�5�A�g�^m7PS�0���$F�ĞT�U� �v���VQ�v� �y�(�;��P��bW�\E���~���}6|*X^�5K^�N���Z��ɵ�A�I=z-m���8C;�ު��@r��9�����ag�;�5hWX����r`!�^/�e]�r�����,�ٯ�r-�n��`ka����>E-�E�b�5b��x�r��oS5ft8R0D*�M�l:�nT"�o�+�`{P��������|���}#?�����Km	�E(�.�`���F)�B�߿��[�����g��ʵA�
e����B}H>�޸^	�S�*z���/�����.�&���2!�T+f���_������%�����`�"e���a�\�g�ů��U�����	���燑⋓ ˬ��`z���	&h�{۽�b�i�;/�k��sJNI���2PP�'�Fl�9�G)}�)�ב�\|��g;��L���ݖ���F��/e����R{|V���GVHA}.�\���n�Z���4��i.����������q��92����Uk�0 �,(ms�H�R_����*����e�T�+�ʕ%_�����(����Efm[[�z8`�f�"��s��#a�1*	-F���e+�ꪼ�Uc��a<�4�O�`��K�}O�h��:��,4,��FP�Uy��%6_�Xq�����x�s(�����L*x3i��Cb���D�𑮢���Q�g��Kؑ����j�T��ݤ82T���WPP�m�twԙ}�q��Q�lJ�����9���o�\Й
gShMPͲC�k�-�	R�~t��20^�\��VU���������C��X�L%RL��|�9 �@܉&�3��D_�Z�m�'�=��)������\�o���e�m������`M��<���Ƚ��^���+�X	�s�n?ا��3UQc�f)�i1�K�NSЃ���s�^#��.�X�S����� -��<�6�FQ�?�{�0��wk��D ���V����g�_�2c�X��UAQ��I��M��f�Cc����y67�b���a,����b�G�ߩ���P��ll�@-m����3ϡ&O�·�N��#�ۍ���#|5�k�u|���d|�d��"j
�`���"fo-��xx�A%#��`���a��es��R���2�y�Q.c�������8��;�B-�rP��u��2���� �pc��&�� ��U�2����x�Rk9�sEH�b�i7I����J/Ў$J:2Xb�8�]�u8�FnM4:o~��B̀5\��zy��9�Wb]��\~{�1H�@��:ʇ2�ʈﴅ�:g�@��"��*"��FM�c�eH2E��K� q �ԕ�7���� E#�U���B�8A�!U��[�4�-k�KL�ЗS��i�L�'�V̅��Y�_��K�}D���\�oWDmO&�Օd0dh�F?�ɱ!"$��k:M���~���Gpg4�v Ty�R&���v��C�A ��ȹqY�.��'D���?ƛʾ'�Z�z�q����y�q��R���މk_ʒ����"T]�jf\�0
]BgHm�y��G�����msv~>wΚ�,*�k�Ry�Bg��Ik�ܨ�Β�9�o�Dor9����=.����@o_O�H��R��[�bY�0���FZ6�+2�T�8��ጎ��#�T	���.�sF	Si�[qAc���[��!Ž�"3�(>_�f���E��2j�����s��{��o s���_O�f��:uyh�xaE~l�e�$sB}�,�e#`�,�/�N$11�:%5]��1ᾂ!b��=]v�1�����=R�I�c'�r�6��C~r�w�I�A{�=�12�X�`!���=�;2\tn$P>�T$l�;��~���n��ֿ_'�K̅U�\�7���D��jFI�c��0U�(d����~�=��C��������Iw�|�(h7_w��P�%>�c�B(|2��}z��1�<�(O�:c������a?���G��p�X�e|���2���D�0�P~|\W�2-�.�D���x�u��+��Ϙ�B����y{4׆��z�N�����'�~�E��?ډd#H���i:�R*}���sٛ�#��nc�(~ʶ�2a(k��z)C)�����{�$���:6HO�s�OQj���E��� �+ݿ�|�E� �mͤQ��i�H��]I"���5�Q�5+Ѽ��u!�4Ht�Z�Nz)�h�#	ï=]�=Ⲇv��,-v7�5�g�ʪ���4N����*��`�1���>�E@��#ط��,_���<�~ё�9�I���K�b���9z�뷄rbPc�6g�Bb�r�YtsZ�O�M�3��,��c�-��(ݥc�|�" ٜ��Xۇ<f��8,d���j�Ny7ɼ��
��fVܾxwH�qTW�Hm����HV}՗�3Mf, "��B����.Q��d�ȊBZ�"I���M�*��G�A>�l�R�&�4�)�1������s��B2^�������"�UO���N��'��¥1�A�4o
����2��l;��`���t���S�I4\� v+��CpV:��xC�,��J�fDv��i91�������T�'o�x�* �L´�L�MJ+�f�]O����B%�2�
)X۠|ň>6��6g
�M[�Z5���+�M�X�-Lcj��OCh���:����d��ö��3�\�\���E]���1���W��?`KM'>���Ǝ=���#�?[|�,�x�� ����!�ʊ��� ��9��D��;�K��/� �d�>�x�]F������竹(�V9q��Z��Uy4cԠQ���A���JJ��7��
�W���x��ox(�����wд2zt?z��������{v��hEP��q�(1�B%i��䤝,�-UP��u˄?�DP���o�:�}�S���:�S�g���lW��������X��_˫5Y��)�2�����)�Sr�3S	�gK�.oy�S�������^:�xw���_0#nm��tB,�b��o���Á��=�J�ʙ��?I,�S�JdQ�v'@C��2�4U\+��Sz�w/S��Y��"C� �rF!=Ã�\
,lX���v<�-��X*�%Mɳ���dЏ!��zԀ�
4���i��ڨLK�"L�O��bD�L�i��叽(�Q�W��xz���NNS~7#XZ�ś'_!�B*M�ߧi8�T�4���F�����~��Q�MGa����gn���Ȧй�/pSm����Q���~C�&s"� �|�M��~�r-���L������!���~��hЮ'S�OdecC�nA��&�pR��ՠ�./oEv]��l�QS�l].��Wgk�	6	a�r���r���(�&��#��ɇm�R�ţ��	��4�Dv��v���%�0'��J�e/�$�m3i���pm��B�bg<�8Xn�D�p�_�N\e y ໬b�1݀/r�A�4;��8�tKċ���,�?o��u���/����	���iOT]t�?<�2 _�̈́<j��R���F�u������(�����M��,3��2XF��r�f~�N-��B��]�ת�C���x����a���{Aw��P~�.��*��76&Sd�������Dẏ�X�7�t�"%�����9��wd��[����	�?�����n�1<�ɥ�K\�ҢH(�v�l�l 
���onӜ9���\VF�E���d�s�$�~���.j k�	�+~>������	w)=�B{9��o�Y�*����w̟4u/hi����p���.�b`E�)c@H�7�j���C/��5����&Mn-S�:�02��
K�"g���y<�=SC�7����q=q����a�ԡ�v��`sv��[JQ���u�=/ܑ�t��
,��H���',�mi}*�p�6�wX������=�k���o����!��п�Z���y塩��:��܉ k�9�{�lP#���Z�{�z�T�\����Zϫ�,�!�u�*���)�#�t�_v��h�>�#V��'0�%�I"9���M����S�����KZB��}Mm��˸�w���W"@�c�����c"�t���/�C�A�T�P�����n͹"�蘁X�(c�I��4�X�Ȳ�H=��M���_�<�\4����=s�Lh�������]����KF}������;A�5:o������B"Q�<>�!�2"M�O��WɓO(9/������}	�"3��F�_a�ʺX�󪼼�a�}~	�`Iye3Z��<�},<���Z4- E�Nj��`{G��� ��D/�G
g>���@f?x�LYt��T*zq�fg����G3�*]������{����[c�uä����<�k�X�/������Uq��2��y��������u���
r�n7"�y�E�D7��I��I:�6 s�(����2��:o�3��Lʱ����_�sˤ\Jr:���$&�}{+x�	r�hz,�_��'폘2G��`�a�k��c��{H�mR�rZa��(�hoo@�3��GqZ�� ��~ސ��EW�V�e�O7����'�E�=��ڷjݶ9\��w�2)6T��k��*}���d�!׻U�V��8�+8H"Cs��r�+�_uo>���2��<����p0]< � ���=�1	"r)�
(*�ms�r�
�/��x�	���ڜN���5i-i�w0�͍mC��goI��ُtM�I΃Y����SE�n_����g:V���z��PU����Z��������/)��E��e}��$�E"k@�"n�F���T�R�1z6P�����E�]��5�=#�g�Пȟ$�[/�1���8�{D�qr�MCo����a"U3V�u��qu]�U $j/̖-&�t�[~#����|���/f`�i!$f܊mjg|���<:C/�˿��KP^YɅA��zM3Ju(� n���
+�A��R�nW1�vdk6������]q�� ߙ��J�F6��;�4�w���y�"��ѓ0e/�
^��h�"up����L%܂/�v���֠Mկy��:Hb��I��(���os��˫�л9�b�����	5�2�� �!;A]o�%��]�Z��3�p��#�t�$���6�����;����U��;)�a�+.�ٱ��/�8��f>���nQuR8��o�0���㌊#-q��!�ӟ�|#Fnn-�r�7#UA���}�A/
��t�cؚڗ<) GMC�AW��5����F�s���2�!ɤ;�X�����H���ENU����I�����%O�[Z(L����c��O0������P�<���(�����7�[7p�9K��ﻺ��+�/��PL�R��69�S�DUœs���ē5�K�'��m���b9}G�_�`x��ƒ@��o챓%	F� ������T�����������9b�빴��(�qW��5�Lz�XV������W��
m�[��0��$�\Cw�\x��"N4�Y%r�&��h,��O��e��W��ڌ#m,���������ʙ����n�ad����nb�'�7�6��qHG�����	���P7v2S+�i8u��eD������78��%����ԛ�ޏ�+�����ǐ��E�II��')��y�"�.�.�+�!���[.V=�J�Z�a!��~�WiB�+�s�y��S��M]8�����j �������FgsǗ������EKw�]h�e+����3��\��zʝ���Up:QL�ͽ-7�dʼ�w	0�!����������q�Q�[��-rj�6����.m��(����U/��Ϊ�f�"9𥡻�H�7���KԸ�|�᳜�-�Gc��qk�5��������F���il�H�H� ��@?d&,f9���O��fO�n�m�V.ṲW�iE��mvl$���)!��<4�Q������t-q�i�-2�(���G˗|�'����T�1i��>w���G>{yO+\J4�ccV���1��HLA�B�������X�T�?�uP�o����&�T�L]��F�-��ĉZFǩ�~�y�4���k�Z���U�J$u�MJ�J����̀fI�7�ߠ�gE��'B�y��uWz�ڇ���o�F�*�0+�
Q�ޒ@�{��J����{Fi�@��`25��|������ǈ;��(P(����Lb������$UЛ�d�f�YvM��w �mg��=��h���&O��!
&�������'J�1�3�v��sI�A$�M��۞��� v#�����+t�d�!��3�G������{x�&qVs�TlR��T�<�z�j�}8�\!݆�^*�ؓ�i�S����2�D|3lR��Ta� �7O���k����c�_���c�,`lS�ʛ��W����R�M ������l�@)Iɴ���s��6�d9|kp��8U7Τy��9�g�Z�� �G����'�J]C08�������̚DV����gz^�֪���o�~@��'6�)N�ߝ&�-c
��)X�p��v�m�YLG�Q��:T�J洨A$�K��"õ�?�[�͌� ���?Y�l������W�K���gE8Ѕ��"Q�&-�@����Lj����8z�U����70ҳ"��i�27�7��zL�_1IN��#i�~M$�
9f�𘤎�P�h$�E#���߰G�̗��0�N|w	�.��l Җ��*8��������Ѿ[V��+<_��'�m4C������G����C{��X:��� ��!5�||�_Ϫ	��*�]~�#+��f�����+�fY4���ٽ �������wp�Ete�;��Wb�b��.Y��*|"3aVZJ�*��o�&��4u�9���* �
�ܿ�z����4WF����6�9	Pc����v����Y.������ø������ę�#�稐$���A{`������L7O�4xR�#f�k�|2-�K h|�!ϻ�A���U�[��U�?�÷l�ly�$��bA�	� y�ɟ ��$mQt�>����L�d�XT
%�ZB�3�	����AլRq"�5N\x�3S�\~� �T�6���]ib,M-�z߲��Zy
-�f)�
}7^H函r(I��o��ՠ���#��yA	�iq��R�X��x�AKL+Ib�+��q��ꎭkLL0ǉ���D���!-���W	�H$�WuA��9LJ�L8HG>5tm�_�]�,�}��<_߾�*r��	�Fn\+�p�E!�S�g�*���/N��qz&��_j���x��.��;��-Ú��3�����?M��Et`(�լ\3a�R���zT�����LU^c��723 �Q�X.s��~�>m���!_�H��Isܽ`��LǬ���z�1��1��0�'�n	��u)oD2��A�P�RV�`�����ۺ�ޮ����u�Vfx�\��'�뗓�}��Nk۝�=���w�=ݱ�t�b  �_ۘ��i��\Vqϓ�W����+���G���2xޝE����~�����*�>k4p��?��i��ٛCOfƬT?�-��0���6�3o� �+���6�ƛ�r ?ǃ�곸�G�z�s�Ԉ־���(n���1&r��󉹴���͘�u#�﹑�ا��H~�D욝$Ith.I�*�eX���1ɽN�4��d`LR-�Q�HG�����̏(8�8v�0�����	�0X�Wr=�%:��i�ps4?��R�	�I��GZ��ʬj�d��3�vK@���@=���S�������rv�w��]Nz��8��<�L��>�?Qc�ճ�ߦ�,2�p�Ma�$�k[0��r�Є����Y�Y���$m�F1G��1Nt��w�b���9�/9��N;��Zw����������bz{�Y:8UGp s�$)�+ی^9�hDH{Ӄ����	�^rj�<��Zt��!���>��E�An4��Mo�=�=��g�0�ǜ��*�M�:Ͷ�;O+����%�_x�LK��b���2�r�������Y�J%�����QE�Y%�8��x+R�f��nG#��]=X�V5睾��7��ڛIb��G�;#N�Zc��݁x�Wcu�κ�7/l/Ƭ���k�uU4���-�)��p��p���2�^཭w��v�,$qr��5o��j�62��o�(Y���}�M��z�f՞��W����KӞ�"·��f^��(��L��
~|���g����8~� �q��D��99���4U�Vq=o��U��И�⒇��ф�Ĕ��Y���hX�Q�zo�/��I�k`���[�4����*��[k���u��!�Ɠ��������  �_e�g�z�Y@��k��3������H�1�>����4Y&'��������wC�$�έk��}ى"B5� 1�\�}yh��x�ǸG��Q��(.eV���!di<ӷ�c��f�6���}v����	h��Pg����W�Kv8��������crZj�oٽ��_夔$+ſ��PK   -�OV%H9  _     jsons/user_defined.json��_O�0ſ��3��-����=����� -�&��-�������6�D����=���#INz'�()H@ޤu�6hD�+���ԑ�iw�X��]�ƴj겓kmԐ^�U@@���2��hB9�Y�(ea5My(�t�P�d���>�њw����t����c�B�G|d�}�\5��;��Mδ�0�-�G.�(MiLQv����"����A�Ų��|<�h>��X����7�$ϦQ����ܕ�_�E�q׶��w\/
2?���|����~S��Ӏ�ٌ���&���`o>b�j#m���Wk��#���PK
   -�OV]� �  �                  cirkitFile.jsonPK
   ]�'V�cŌ ~ �� /             G  images/40a6b5df-e714-4004-b865-d48720df955d.pngPK
   -�OV%H9  _               �� jsons/user_defined.jsonPK      �   �   