PK   �cU��	�<  ��    cirkitFile.json�]]o�Ȓ�+ͫ�w�~ۻ�������c�HM��H^Y��l���ݤ�X��T��|�f�]����bW�>/v���^nw}�G�{Xo7�k���]��y�)�Zܯ7�~[��k�?,�?����_�}����k�Φ�ge׉�U�*��hx[�ʾ����fU��-�on��G�dVs2*���Ւ́��j���/�﷛~���JZ)9+�a�|i��4�/X�z���v�k�W1�q�`�):�e��UST��)�j��m����kW�k�d�SXmH���s����-��TV�dTVWdT��/2�cx5����r C8��±��YN�p,衚�XPC�C8��I�p,聓�X�C'��%鱓�X�c'± t��S�c'���1�=v
z�$C8��I�p,豓�X�c'±��� �~����f}�<Q�o��z��3~�$Cjc���01$&<�	n�0��8���ǲ�Xv���N`}eǱ�X-���X�A�q,;V+���wPvˎ��;���ǲc����`}eǱ�Xm���X�A�q,;V�XߕX�A�q,;VWX�UX�A�q,;?��C��̏��������:� ��`pp��������K�pD��*#Gpp�^�zp���I
���Sd`���ُmd��/�G.��*p���y���3�`��s,?���b���;X~���"���y��8����k��,?��g���g=X~�ϯ9 �=���Xg=<�"������<���.X~�ϯP�<ǂ����������������X~�ϯg��`�q0?��?p����_�7s����ٙ��+^������1������y������+�`�E`r��s���̙���)犙�0��`��\{���4�kO�q��c�=Q}�����D����S�1Q�����a�Ǳsv�Rή�g7������kO�~��}�}IԾ�vE�ڗ��+��W�'���D�I��Q��?Eԟ�����SD�)��Q��?Eԟ&�O�����D�i��4Q��?Mԟ&�O�g��3D���Q��?CM��3D���Q��?Kԟ%���g���D�Y��,Q��?K�_I�_I�_I�_I�_I�_9�?Ζ�v�)��Pͪ-��2��Z)\�����8t�����B�ܖ�0��Rv�ٳB6�歪��J�8{������u���M&P��@K���I:���H�x�&�o�\|����n���-\�Ć��5��*_� �b�����F ���!�h�w��I��[�h���F�4�$\�$m'��12(F�#�P7�4T�0�5A!�qa�9,p���� N���A1�Ð�ʄ N���Aq�Ðƪ� N��aA�4V4q��q��(���!������⸀�q�X�	�,���ƚ� N�8.`q�4�Sq��q��SH�Z���޾���y=W�i�aD��R��o���¸���@�o������kXB���tpT�_sp�+b<p���
�k�a�E�����Q�~��5,ˈ���<8*Я9��%18ޮG�5װ�#�����@����z�x�x{��\�2��|�$&Rԇϓrea���E�6Sڕ'�
�4�a��͓zea�0��	�1���'���6RB��m�,�HyI<,p�0�H�H��$bA�F��bY�FjK�a��͓�ea�;��E�6OJ��m�&%��<iY��z�xX��B��,�H-K<,ҷy�,l#u.�H�f�˓�5&�H���˲������"}�'/��6R;��m��,�H]M<,ҷy�,l#57�H���˲������"}�'/��6R���m��,���:� �����zP&�Kϯ��"�_�����g��p�X�;��&Bu �b�;�	�b���%�g��D�L,�?�P'#⩝>gT�D��b0F�S�VΨ��7~F�����3jm".
��Mg�D�u1*�KPW�b����%F��b�Q�ĨXaT�0*V+P��b�Q�¨XaT�0*Vk��5F��b�Q�ƨXcT�1*�k��5F��b�Q����`Tl0*6��	��F��b�Q�Ũ�bTl1*�[��-F��b�Q�Ũ�bT\bT\bT\bT\bT\bT\����z� ��SjuT ��\k���O-szz)�^��A��£ ��gs�K�>�}(������9��J���ҡF ��t(�h,
aK�B���ҡF ��t(�h,
aK�B���ҡF ��ҡ���ڸ����QHO�C1�`��Â7
�t(�,~sX G!=��p��p�(��ҡN�8.`q��T:�	���u�aq\��8
�t(�,�XG!=��p��q��(��ҡN�8.`q|
	P:�:.#�FJ��Qa\#�CѨ@���)
�@���
�k��ҡ�Ѩ@���)
�@���
�k��ҡ�Ѩ@���)
�@���
�k��ҡ�Ѩ@���)
�@���
�k��ҡ�Ѩ@���)����I��b��>|��+�X�P8,ҷ�Ү<yWX���m��+�X�P8,ҷyү,lc�C�H��I�������"}�'��6V:��m�T,�X�P8,ҷyұ,lc�C�H��Iɲ�����"}�'-��6V:��Yȓ�ea+
�E�6O^��m�t(��LSby�'��<yY��ҡpX�o��eY��J��a��͓�ea+
�E�6O^��m�t(��<yY��ҡpX�o��eY��J��a��͓�%�=�t(eb-��C�(��(JG�X�|F�P:�ĺ�3J��Q&�֞S: �Q��&�sJ�`0��uN�P F�Sۆ�)
�zO�9�t( �⩍&��`T<��ҡ ��%F��b	�J`T,1*�K��%F��b�Q�¨XaT�0*V�1F�
�b�Q�¨XaT�0*�k��5F��bJ�0*�k��5F��b�Q����`Tl0*6��F��b�Q����bTl1*�[��-F��bfè�bTl1*.1*.1*.1*.1*.1*._Tqr�P:ʋ�)�t(�e.��C�(./�7�t(�x�\����w�]���\\s~�������]��z������-�onb'�Z�m�M٬�I�*ڕ���k%�mU�:��g����ڮ�rYTΰP��E�J'ж2͊��\�CQ�۫@�aI�/zrqɓ�Ó?)�Lۢ���P�S[��()Z�Um�Zux�gs�Iă"&����0!��Cv�U	�O$��ԇ�O�2����rQ��"oE笝�[Y�b��D�*ۮ�V��ʓ��K���h'�<9�\��Ғ�S�g���!���I9R���0{����L����>d-QV]����zCf���C��:
��'h�0I��wﺥ(��\�(:�4.ݟ�ʒ-ͪU�*$�N>�<�wV�?z���S���/1�N-�F;�����ڣ}��pr>����0R09�PA�B|�W���:d��?n�軺�t��G��cX����~�P��9�W�AF9\v|�N<�!t��.���^ �Ǿ�r8��ztL&��1���N��jH��;���K���|�Sy/��&�^��W=\�@�g5�F\��x2������@O#.��Iz*si��=�jF���3D�]���Aܲ"��j��2F�t���L��N�^	�c�k����M�C���}5:���SƯS�$B�	d !�<�.�z%���� �^�C	�0�����Ը�k����?�A��/��s����~S�('D�h��Ԭ	
"~�
��%�s.��� c0O|T��b����]` A_gy��[A8W]��Y|Eg_��(-�-y\o��þ����ooW��t�~[?����g���zQS�9D6l%� C�ak)��[S�,�l��������tא!�PQ��5S��I:)Kw�N�,�l(�JdA�`c�UjPC�VDpDW�t6ֈ�� DXN����*�T����Q�0�X'��K9 ��1�X���O ��1�X+���[EtW�T �)��厩< �T �)����< �T �)��%��< �T �i�A�.r�8K�U}G�S;R�ٓ�l� {7��>���`~�)�/�>��b�q0?V_��Ã�ˏ���:�B=�X~̏������ ����`~��߈G�^,?������px�a�q0?V_p�Ã�ˏ���:�;�X~�Ϗ��;��>G3�h�~��CxOC�yG'"���r4�p�E0@]@�NNB�@@�K��	G'(`���p�ƇAp�s�v2�&�#��@�-���r4C?���!:w3�h�~��Ct�f����/ڇ�̐��9k�06:�3�h�~��Ctf���Z���)�	t#�S*���r4C�F�Ct�f������s+`��Я�A����r4C���Ct�f����$��y
�!G3���>D�)`��%�3w7kbg�kY��$�kGg�]9��mvy���"N�VNή�A�V*�UY�T}��N�Pn�@e��b. U��V�� T%����#%U��:����O������fʹxT��+��Pu���>��TRu*ɯt�N%5bJjĔT%J�%U���DEU��*QQ��ȽK�U���DEU��*QQ���J�T%j�5U���DMU��*QS���J�T%�U���DCU��*ѐ�l�U���DCU��*�R�h�J�T%Z�-U���DKU��*�R�XR�XR�XR�XR�XR�X�P"gKf;�FY�f�M_�BT��-�~՜N�?q�B�ܖ�0��Rv�/��i4oU�\U�����O�?����ɳ�ݥ�l$��KxI�;!�Ěw�խ_��a֝�P��|��	/�o~��w�k���w�/��e����r�|���o�}S��rߘ���7�=��[o!lo!��P]r��(����[o!���r��-����Bz�-����By�-��P�x�-��P�By�-����B{�-�p��B{�-�����x�-��0��x3��[o1�J7��z�-�����z�-��Zoa�����(�E�-JoQz��7�"%|��� ��=4H�`\.�N����6��K�vd0�s�j*��8��k�ðs�����`�@.F/f��ee��R.FM��2_j���5V�G�}�羾k��nxOQb���_�s�gt8��C��ɧC2<����~:4�b�����Pכն�[?�{��R(U��i�.�`��x�˪_��e�;Ѹ����{�K�w�j�_�)߯�ݒ36��x��m)�b�Zg���dґ0�1J���"Q�m��ڽ(��'�[(�7���o����7��)����ߛ��}>z�������z;�7����s��z�rg�|���W�?��G�׿�<��7k�v����a��Ϳ9���ʻ�|�w����]��]�?��]�-�������f��n��q翥}���fϘ�%�L������K���B�F=�h)�?=ş����ne�p���w�тN�N�}�yUV��#����f�m�z�W��n�nX3�Y�[�w˻���p���+��-��W7RLQ�6f��N�T�6�Mq1m���i�rڪ��|����CJ������j&ڕ�팙��L���x2O%�D<��W%�E�+���1o�L�a���{mC��ME��0�p�|����D�==`�c�	;s�N���'�Ĵ]UN*��!3m���䴕���6*��!����i;�B�q{_��*��JEԩ�6�LD,Q�TD���R��:R��#Ք��yL�6j�F]�T��E��2�5��0�0*�Xèc�2�5��0�0.�Xèc�2�5��0�p�a��(�ؑj��I��#b�FM��dk��v�W�c��u�ح����������7�宑\�8U�oܫ��J_qY�Q���y��ڶSJ�u.��ۮh+�l��m�n][��<!i��8Oح��S��;����^�o�ؕ'��κr���-���A5J�|@���g��n�J}�w?���o��d�P�rU�j�M�\GɴR���)�	�bẁ�`@��#��H��G�����#<j����q�c��K�����q$�j1��Ϝ��T.���O�n��}h�t�?��p9�W��?�-�:���?��C���� ̻]����ۺ���띿�7���������޾���W��^���֛�����#�X��"Pԁ�z�|�I���G>����f����?��~���~Y��~ƅ���7������|��Ï?~6*Y��+N4���~��i�P�Y����%�M�;X&����)���8���V&�H�ٍU#zӭV'Us�$�	�̞�zI)���m�>O/+�O��<�suR�7�!����V�z.�o��y�X��~L�fҾz�Mx��L��3u7�����V�Gc�a7-�O���P
,�S��3���b�!J#BTp��U�p{c�
)�!�V*�;��j��.�ϴ�9��B?�,�s�H��Q+!����V��lV���C?Z���E���E�ѝ)���)��6�'��mi�}���g�m3�"E�;W�H��8j&YJZ�e�G��ww������ݺ��N�R�?���wo6���߶��<��/�/�PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   L�_U�
L��\ �j /   images/5d6e91a3-4a01-48cf-b4fe-ab41826b34fd.png�eP���/:�� ��apw�A������.�!�{p	��!H�w�@ X�p����{�{�ܺn����jj��^�����kj��8��0  ����6 ��  x��>��YO t��^�0_�������5����l�go �-7ا��D?^�D}#ƶ��o~Qѽ�zmL�����˄���Z�-~���Ӝ^����#@�cZ�����tc���:���΢k�^ǯ�+�#�?o#��N��I�ndQ�����.$��>;yI,�l/�l�w��c�VB�dTy�t{��BH�����}��1�o�_ը}.W]7/�=�.}��Y�eȜ��K��s�?�4C}#Ȑy�r�1r���0U���u�T\cL��MYq���[�2��E������hO�oI&��ϳ�2��1J>�����?��=��MLcS5�g�tN85�rN.ճ�}O��JB�XA�Kv��T��?�#�2�sl
��HI|�ji��kn��2�ꯟv�R?�˹�6��Sz�|�W�~�R��c��3�=�����KTIG�tw#i��l����������=���isIТr��!�'åۮQ�-s�T�B.���9��cTv�NlFzZ�9V�y"+��h>D>� 5aZ�J|���m�K;N��^���&�~��8df�B2�g�l2�۝vg�kw�U8�Z��zrt,�$�Wf��5�^��`7|m9���M.~�l�mx�Hi��]�M�Y�M����j}�z~p�������W��/(}�7��:����z��T�|���Y���6������F��ģ������L��>���N��ݴA��Ħ�r=,��^���m��9�T�	dp�I�H��M6y��Ԩ�QףΪ��Q���i��k�I���w:s���n��0;j$������C��B"����H�����A'7�F[�j�H�?�3 ����i\|�5��hﻘ����)z�F�Q�~X�����~���z"���]��z�K�f�ڬ����Q�
�� W��+��f�4�#�ߟ_�G��Zr��c�_��|��N���&7�5���;�+�p �IBO�v<%T�v�6�x�f0P�E&4,�jM)r�7�UA.�k��+�eS���3�ޱyx=r��]�Tw�u�����8@����n/S��Q:GS�:�#v���ٺ�
y%2���(�`#o:m�y�E
D�z�[��@.k�SZ9��+�r5Hֲ��cc���'��fuSü��%�_�\raِO�"u�wI�,�,��$��PO�2m|�1���*n��f�`n���_�i��İ�f�P`�sW�9	�~_l�x�+���u�`m;�u�%�gG���6q��c�%k��9�.�p̣���$�k��d/�J�u��C�Ԙ=)�bZ�L��w�^�Q�46D�Z��H]�ՏͫĖ�CON���N��-��o51X7�N�0�"�����$L��Je~�{�U�y����I����㾑�XQ��������5������n.�_�o�|{��D��������e�n��b�ǕmkJ���Ds$�,$y���,#�K�.]�@�.�\��C�O%�|V!D�f��j�qV�#����C������;�BH����g)������[�O�C�����|x��Ϧ,]�˶s���ov{l/ 6���}�p�^o=ĸ�:l^�U���=\[�F�^������X�`��>������
��q�Y�[9訙��ƺr��-�!����;0ΰ饷���댚Z�<^pUs�;��N9�xT3?݄,�'�������Rb��p��N�w�%��9�����ů!#0S��a�,u�5�7]� J�.t+R��>#�+�P%��8�t���L>J�E�b�$���t��Q�qR��]#���2���m��ڌ���0�#�u~]3�q�t��l��n�k�'*�J�1l�i�5��9(k�������Go#����-������y(q(\�4��_:��2ٻ=0�i��So�Gp��TΊ�an�45T+�r�fW.��bc��M|�O���˲i�n�w�D��T*��|�!m���;�H8#'1����7�b�S[�)�����2Fe�����˝�ď�c�O��<r���\"�Nk����NF����G:˷�+xf�,�\���͡�w�5�w�8*�!}ʠxٝTbu^/���	Hլ����F#����2om��1e���]M	G~B��D��<[/O��5gΉ�\w8�7���D���D�[��C������pK��-�g
!��&�	��.'qp���g�� �	_��k�V���'h=��Q��P5�v��U��? �n��;b�q	�ߪ� ������B?��^wI���U'�k�P�#�3b�����1j1�vF���r��c���oƧX�N��&U+U4 ����ag���*;���*?Z��ݫ�P紥���m����K����l�u��r���^R�g�7+����Fg.�@e?���;�&�³���(o%��U�X�?��6�	դ��kkY���%�Q���q��wu	�:�
���?�L���R�MZ.�{Njh&Q��-EY�Μ?�#�����[%��;+
�p�f��[�ƭ�3T7��.�m;{O"U��dZ�	�8^GF6�|���?��V3�l8�B��C�*C��NƟ{�5��V7��Pe3VkLk��.���'O����ϸ�2U_=&�`(aW]ҭ�'����-��6�C0��I��I�K'�}OU���t\��V�?2��2�zT>�l"z��Q�� O�6�w�9�"�s ���g1�?Lo��(�9ĥ�������։���%q^��[ ���tE�H	(����bc6r�T=��b�1����dنe�Kh������O�xUn&��[���s�k�_�#�{2��^�jI+���1��sQ�ө6�?�+��[2���M�=�i��g:F,��%u+�6��r��x�;N%绺?૞	j
{Lx;��.$��t5�C��T���MQ�;&�r5����ѩ�	�v��`�ieʷK�~�LV�`k$ �DJf���BTu�PK��Wٽ���(�Bir<���� �23��fv6<Fm����}	��g��ˎ����5�R�#�]���y�hE[����P���Jf��w�NbDA~��Jy���Mއ�=���Q��i]�/�\��_��]�0^�F
îǙ�Xʘr�s�b��$$0����i񆃺�tߎ���۪N���W&Dd	�@�7��#�&c�a¤���__�@�*���`�kc�(���k�y�i�CN�U�R�Zz��K-�P���wRi������N���Xt:� ] �/�n)�Mؕx�ً(��82U��H�\]�	�&9�a�6	�{�� ' ��ۈE�z�].�@)R  ZY���׊�9r�A�8:L��}$�9e�㫻���&(�Z�s� C�5��0���A���o�
�e���5�<��vG��N�AAQ|YjG�Q�?2�d�D���s�b*! ��!�~4(8�N�و8Q�/��+�&�"�yST b`s�M�� �*U��zA.��6�L;� E��J!U�5~��:��cF�g�`�|�Pi=ۃR���Hf3���&���YđI���$���C8����j9���%P�7'*wu�A��q��+��,�H�P�5������	����A�K���17+�������J=] ��~a�y�g��<�b#.'��7�<J_�OH�0}��[ަ��Z+o�6W�n���Q�х9�Kd��N:^��6�5�ۧOtݼ�Kd&�v$���A�Pۄ4z��[d�\2��]�qFr`��t�QM��_{D"5B^X����,��9���Fzi��r�n�*GlD�#�ʻ���0lk��9;	)����r�� +��|R��f� �Hܑ.�$��G��3�!�p�־��I�֏@#��{�R, ��0jѬ�(ܔ�J���[^��I�ޤ7kʵ!�*�r�$�q�5��'��`���4�I�����GD)]?���@��J���lQ� ]v���M�)C�c���_��&�qd�&��+<2NlN��UcZ*b2:�Wa�r��S�}��B��Z����M�ئ5	-�C�k�:��*��B+�ͬ7��G��H��ĻE��}=�����,9�rx�3�,'O�5	G���H�qZ%�p5� �.e{���M���v��
!�]RB�����q+J�Iy�J��ˏ�Q���vy�)�]�X��kj�ʖ��Pϲ/��yI���D�j.	�EG�Wh�-�6�P���]�m�7�,�gҾ�b��`C�����pT
i��{>�G��X�~D��a�<��S�4[T����}�Ӫ���cD�Q���kG�5#}��+L�A`1֍J�p�iSz���>,���Ǌ�1Ԋ��Ƃ�Vm�k�kT՜�?g�J�4J����Y�a��"G���O�������a ���O�P��9���8�؏�MFQ�����Pu��k[J�~TS���?Ώ�5o����A��qڞ3�U��6�[Q��s�;a��������=Îd�$��źވ�r!0�E��h6y�.3��fL������,y���Z]J���g[j���A27�l�q2��3D>�����6T.��x�;��:����Z��`+"Ǒ��8��[Z�8YS��������k�}5{4|����1�F���hH�v��T�ı���I�ɑ"����͆���l���5��z�H�̒���[%>bKe7�����(zn��E�՘���W��"��fK���Z�Z��ަ�>o��!,M�y߅A��*��vO��7��Y��2������<�dbNa�	�L��R���'�LF�Bu-�F���[8S���v���wH��S3�tH�����,��e�������3G3T��0-�;���I��3�� UVjjfd���/`�KZ��7Z{�~�3�-�=@�8xO}���Hx�?�O<�¡�0a���JJ�o����n����Y�Q��z$Y;N"����`���R�Ԉ����[_����YίXe����PX��BS��Of���UG�d{,��B��f��_l�a��[m��71~���O����'��u6O(h������$�Mg~���i�쮳�c����5�·��&59<�Bdx��z���x:��R�z�j'9n'���rlu�x�a��HHW��
=a�'W��f�g�m\�Y'8��3���[/Ӈ����k�E����K�U��}��#��P*/������
�׷a�
3��uW�,���;a=T��P��L�)��'�!�aL+G.A�]K�P����I�N��
J$'����p����>�-�M��0؛ܛs�{���o��c����_t�1�U:���SE\m��=s�E����� �mL:h ��\��b7g�����l�����&ԹEΐF�])~?Ɨ+ҒU%���M��<0����ɶ�MYZ�\&Y�M���iUj�~.0�R2���v0��x��3����'O�>�����Sj����ԣT,pkN��GD��I���Tu�C8��];�)�����a�n��dnMn�Gd��A�7��ߑ�IL�m��+��,$hXg),w�4d�:lN�$|-�0L^�1�ZiP1�s7���~����T@�m���Qs+�JAL%7�7���'KjZ8�>��F�`�B�����PLĞ��g��d�D���e	?���l���t(��q�K>� ɯ<���閝�����z�|��V�3��D0��	X�rg2T���%���W��)U4��T��8�N3�}�,�F�s�Od�ׄ@��F�/!��1��4��mr��X�>US�۝��g�����oDz��|��H%�O�����7A�{0R!�,��θ��ΰ c-ėe=�
�>ʕ/̆�<�3'jp`��-��l1U#BwVS_ X{�ud1��%�{���/�3g��-�(��M@����7�5ȺT)�����JW9��c�u���J4k�p��v̗tΟ�٢����!��8QC&������Jxlϱ2�|`��f�܂��nv*"�����Ҡ-����;�e�h���_�N���u\~��]v}p�$��k�?�|%SW�M�����n7�������#��e���PX[�p�".p���2���8w\�[��5�;*�����wf#'L�/�}/�u�yBּ5k�<�����I ��A�$�&-�x�����E?4)&����,O���`��[,].aɚ�6�oI�F�����J�����r�E'�e�ȇP���#��;�d��JC����N���C����������9���}r����s�YũԲ+
R��t�y8�t�"�[���T�R�"^��S���ad�QXX�x���w4�be��t?��#Q��>�7���u�d�"%厄Px�ˎ�ʋ�,��#+fB��w�:ZdZ�D�@4GBM�*�t�ql��nRdo�!��z�B�b2N�	�	^P��b8�IͿ�9.�QJ��c-A���'��$�����"����%��[�N��JMd���1�C�9}]}M�,����8ʬ�-�ŀ�G2JH$���=��r��0�[H6�j�R�1����i��
��f7}.ke��rL��2T��sː��L�KZ��)�g�񋳥�;���bQ^߬uL��y��4�� �\37��8M��5���Y�lu��_����aGb�i���e�T�mk:��nI��c/fݞ�*���>���T�j5�,�Kev�iWfb:ǰ<;�Ԉ0~E�𢎣7�G��K2z��h"�Ș��2h�Lu�9���"�Cl1�Qy|�0dO0�;g��%������Z>DD��'�r�kј��Z7r��W����F��n1#}5?���B'��F�i����'�����R�n~�\��P�
%������\Slb��
 �z1�W�Hi�"�|Ä��=~G;/R|6|8Wcʩ�Ћ��
]9����Vi���"P&�^�d��.0�&�J��`�9Y8*Zׅ�.�҆f��Ss~�	]O�������\St�s��{��#:ş���:���'yh�&���(��ɔB t�Dd����#�+�E����)=�-S�i�%��5���'�ѩ�
0_tV__o���t0�����*���M7١cZ�CYW|yCM�<l�=�j�LaDY�y$z������0yr6�Sf����(9�&E8S�F.ծ�����VI� !,��g��ʼ:tc��Do����K+K�DO��с3��eA㽭u' ��� ����%��[&��� ��?G�S��B�hȨ�nExH�[w��P��XI�Ւ�WPS���Rï;��tQ~�S��3.��"#��H���ƭ�w[�9-�Q�+~l���������oɲ95#���8G7KjJL�`�7H���]����UJ?Dw��&���%�(I�:�jck?7>���w�G��V�:닪5v��j^<(k@�<�L_�P� Yo�����=_0�ɉL��+J�'H;� ����r+-��/�Z+����{is4�Q,rmk�Kí����ͬ�MC�N%I�-f7���B��p}(V�V�"�c�T�`���H~7F���eR��������'$B����Z<;+� WTě�c%I��t\�R��R�J T�iߎ�%b�8�s�3��h��	4uA�v64�_�dzP/	^8G3��;3[yl(��v�yX��Pg^bCw���<��۟ɪ��n��Ã�b=M�Wܲ���:|��&TqH�:`n��@��T��&�(ȧp�b�<(S�'G�g�:K�ԇ��~ޝ*�����ʠ���"�wҎ�ʱ�A��Gn��������/�A,y�����]�������b/y�ۓS߇�r�P�U���(�5�8k.�j�B�8�Kݭ�[�Ea7]�
�6H�ީ9��Z���&���z�q
����<��� k��d©8�*��P�2�h-Jo�׊f$���2����ΰ�W"���6�.��z�ug㮭uǇY6��:�2������:_�М�\�>�K�&ǳ�g�ti�����4R��s������DE�~�
��`�:rn�O2c%v��*6G�L"x"�T�)�����9���ڇj��yߦ����"��O0�͒X�*2���O� X݃_�\ F����H|7�^ �����]fq^
9a�̶_yc{�n�ǡ[n.��"|�6���HH;v?;�@�������EVQ¯2�_؉��<���<�h���0�����*�]x`iG��Ƨ0E���Zڭܢ�.(=��4��V2�5���#F�y��;(Q6`����O*Ҍ6	;jR�9�s�6��͏�)ub9@F���p�	��߈��뫑Ue������*�n�Ք��k�	{��SZ�x_�Ou��:�;N<`�?�:�q�ܖl��^B}B�'~S'�?�������=`w���M��(�|P`K�=�Ko��I���W�w�'��������vc��2�o�f"/���[�9��`����0�Ya�{s�]H#���*/�%�b�mg����wQ߁�Wk��S��-�_c�Xc�9��?��:9���A����;���"�rL�W��bܦHF��֞�&�	K��ٺ2e�'s_�Л���/�=[(���fE�K��A^K����T-�{5�η�^�23�^� �dL*���y�Q�ƃ��b��Q����\�z@�m����+8ȋ�5�1��\S+_ZֵF�����r��uzYF?��^i
)�,�3�����V��L���爟)�j	�&ʉLQ��(�o�S]���6zȉ$�-�G�l�_���}�^K���U�������h��on��~�ɹU�rD�4__�����߇�2T֧��hg����Xs"8� �S�т��\���J��#9^ǅ�Ԕw�苮*>C|�����y��Ȟֆπ�1����|�EU`��4�^>��KW����>��C����q,�\�_u�p��Z�ݰ�ïG:7����$�����}�  !�^V�,+�Ͽ�  ~�i�J�R��:�F�����9�"�@"�LV�A{��#��$|�J�&(��ԉzh$���&(�gH#��g�U��u��w�%��W{��rkm�K�Ӓ�G�|�~���#�&����u���t��6���|����UC����"'���c���s�	���XL�B�%�����ߝ��p3�����	?17[4�'�/O����Y,єq��GV������l,��)�U���y�K���������%���~�C�Cd���?l���5���J�R&u�����gZ��vrj��R X��Tq�c���id�E�0輹���>p`rS�3���D�'Y�:�����kCG�g4��)� -v� �u�t}��~[���I�G�֦�% ��c�k�e��&b���	��ZZs�9��1I?7���������E���m?-�.N��_��&kmg��a���k�h%�����yb�l��9;�x������W����2-�//GqZu(X�������	����ᡕ��y�mD�����i&Nk���&�����������a��-,,������x����w��q�x��a�79kO+{7/{W�9����K���i�O����������^x��̍��������'<��}���'<u�ݬ���=]�=���}�]������_�ݼ=��2n�e�d��D��ă�?D**�C�����n�zR�?(��ml������K�����gK�"��G"r�V��S���#_�je��f-�'l�k�������s�`��������� ��o��]<�`.V�X=�p�?������q�9�`��|p!A?��5/�_���Xhz�?����Z�a���
.��',�a#,`��g�c�!,(������aa�߬�V"
�ΰ�p�;�l���\l����pi��8-'�V�N0/��O9`�w����-]{gk/�r��Cx�y��xyx��H����	��rC8y����?�<��k���v��zXü\=t]]��i�� �9��m����ü`r0/�'�n�/�.���6����]��6��O��,�����=������wN�X��=�{�d���WZ����6��c���-+;����S����u�� �BpK8�0��� ��%�%D���	h��0+^n�r�t���yXK�>���WO���W`����?�}�]�v7����O��c���Z1���?�&���rq��t=UB��������_!��_!��_!��_!����?͔������U��yj�P-U��j� ��oC��0ܔ= ܡ?"f���E4/euy�}Lj<L��L0  (�I��-��͡���q�;*��㝠Šٹι�@=�X{W�6�@Ȁ@�������a�]��d,Y:�E�OX-i�S���L}������ÃV髀nۀ��٨@����#����O���� H�/ưJ�r.�K�7]n�?��F��t$ڍ?OK����R�sӴ0�os���Lb���X�k����"-���&�i�D��3�2`��n���~ QF?�̙��.����M��#%�^���%�бUJ�Q�CK�q?�a�5b��c�D�2 qC�p���(J��o�#�D�@����ôg�,�EG,a.�j���u���!膻�'*���TÂ�蠰*�qG��6*�X�)�=#�����܇�>.��>��?�z%�Q��`���ӱ��ل�-!X�=ɞn�_>Z�yl�q��&xя�I!.�� �������@�����?��9��+���4��̳b�
�ʀ0,yG�!OI�UL⬣m��WfO���[n����L/�z�\�+?̼���E�V���8�]� ��NgiF
�s���Dwz�[����<D�<�OG%���P��l^�VO��l0�xw*k�U����u^��jl�4�I��S>���$�ba�V!���6XJ�>/6��6�����}=�����U¿������g=�K�ݽ�R�h&G� <��' ��S���>��������3=�T�B�&̹?��l|�%O�sL<�iU�kyS� B.��B&H�BČF�Q��4�7!�^���%?�$'�xN�dkf伱���	�j���3�cyq
 ��[T�&����
K4�{t�{R2���i@6o$0"USfe�m�y{��L��f�ئi�3ݺ�����H~Ĳ�\� 9����J�L{|�(�;�Uv-�@�R��-)<|k ^���U=��0 Aq�"'�t�Z��*m�p6%�����	���M5�ݗ�)���ڰwr�r����;糃�4�����|9��j�RF�36ڄW)Q��'Oza)R|�Y�1�ġ Aᵌ�8b�@(�n���.�9���`B	��Ł��Ɂ7pT>@R�kӟ��9�(	0L/�aɇ��7�b�D,HQ��e^�J+r�V�B��%����2��=���HI�NO�ç�{p0�Z�>Ɂ��,���'e�ao.�TX���g[ſ�8��{f�N��#���Ok�@�-dd��$� �&򔱏Zq0p��Bi�[���ll�ڵ��L9-90P�� ?e��n�=�Eo��[M�:S�M���ɉ��95���tȳ�[�F�%���͡�(Nn��|P��[c$];^�>̼��7F�[H}͚����7וHhUQA���vw�c��6�����$���KĔ�t~�W�BW�M��QO��%6���5)���O�`
���'��-�������!��zK��%�ߋij��Wc��5�}���j����fLt�HR�g��>�7FF6EA�(₿���q+Ø��Q����#h����m��^�A嵀4�:�4O(������6�Q)�����2]b��]_����	���E����iT��C�LX��[�*np����#\�XQ&�ZδK0'$�H�޷�C����_�Ѽ% ����md�^�* H�_�ܲeFݑ�6��s�\��1�WT��w$-�Tc��@�Xe���"c���3��8($�O,��I��I.�Eo�'x)<�K*[�_�m���K�d@6��C���^��@_����vV�wAږ�5���Cl�f�Z�6^}dg�}[�e���+�3�鱦$�`Хn��[bE*����fL�uOR�1�l����f�Wg�x!@��_�5÷���!VQ��bKè�A�n�,��(�R[MZ���n�J�dj��Ej�&v�i{���F�0-2�>�$�u����w��-5}T�Raz칶���}���c��Ov�������!��k����c)��QS����ģ��m�������/|&�ͪi�Z��4c�с�M��R��z�09|4�]](Y��`0V��nڊL�bW���BXX(ZC�����lϘu�Bg�'��%^�&O(F�NAr�U?�O��>���O���y�&{�z�B���h[��`�����a��"6�� �*���LNX��0�������zsߊłt�+�]#�,���%�� G�v�i����%u��\�1U����&�"=�#W��It���/��|�f���J"��E��Bc�_���'�Уe�~��ſ�I��v�Ҕ���4��%�BG�:�Dƕ��K��&kS�nx�"�W3�9�>�����$�$#%��EF��<<�w���e�H���􅧦.�X��+jL4�����h�cQ��6z��u�τnx {*���ߎr���<��f-(9�X��e܆��G1$��76&g��c�5M���؞��(� ��&%%޵���<�&-8_�$N?87sY�=�T�y��z�|�ޚ��8p����k��Tlj�K��k#�uv�A}��a��%--��3dO����C:3[9��h���h���a.�i���9���ג��
��@��FfȡS��5�o\�	$XiAZ��R�ʚ	�6Ù�������b���4�v*�sY�| ��A(/7�|������r��c�iu�2�q�/h��d�e��"2q�FE�R��d����S���(E���l�G��Ǔ^�}�V�ж��8fܡ��H<������3�óm�|�I�\IJE%��>6..圣�ץW���@2��iX�n��;��4y�J��e�1X���� ,l��>������/���ߨ�*�=����%�h(_x�]pqb�(y�ʿ���\ߐ[H֨�)��1fj�L��N��L<U+��_,�[n9��1�̘�-�!A�d��TOC9ξOmg���*��$���`���;=���ަ]G��
R��|ߘ������KPd�.W����{{��=��T9�G�Y�����w*e@�@b�11�p jˇ�E��J�v�����KV<4�*��vE=�LA�Pṯ�z�gIH�T�6.SYLi ���Ԇ��R�"kL~��R_	#<CMO�7���^}v��^��t[��DE��������|k	�S%m�y�U< �GeA+��E-���-�&�LK�ȧ�"��{�T���cX-���D� zw2ݔ	�jb��ǍR�����žO�N2�a'�L����+���� ����}6��@���+ŻjQ���{��8H�}>�o�]�F�|�!�:+/>�� lSY�Jn��p/�p(i��9h���!�1\�z0�)�!�ڲ�N�@�L1&,(��U?�YG�0F:�B�c�P�ee�l�Ny!��LT�N��N$��I��AY,EN,����?�v��[D�U���,8t��|�L������)�@�i�D����	vWx���Gg.�����Zџ�Oe��f�n�WW�(F�A��.���(�Y��]�(���L��Hl_����z��/S���)��Ƀ1ld�X��폻�좗l@~}�3)���<��h���+4��ȕퟌ�%�F����K��\����=��Ł��y��?��u�.��}�::�_��A�a�������FꉉA��%u@s�sr����Ö1P���kM��6i�-<���Xx1�iy ?E�9@�ї�=RV��tR`��c������x|��f��K�y���I��E}�L'T6���K0H�,U=R{������Y�>��aO���[e�BI�'�}�������5鯭Ь�2�d�����Ӹ�_��ғ�hD�@���bE�z ��2�rJ��ʙ�8�l�q3"���b�XE�5�uR�=H�s�)���f�B
��p;6b9��؈ԟ�2C�A���(8.��]_f�Q�����`fi\Y�#8JJO�W �Ga��@�+��ߕF���,Ke�+��K�ZԀ=���Z��O׍��k'H���O����6K�}8� ~��\Y���g|�LG"E��ҋ|�y6&�q,�;.[�	w��F����~�0��gM�A�jk��gOʷW�2Z"���f��&�,z�[�L0b��] (����v���ǥxJC�� �Jcxr�av�*&k�%���b�U@�b,�3N���m<�a=U�{�e|P~y0���ax�n�>���>�F�����]ӣ�S�Q
��40tE�5�M���%� �m��Cʨ>@F\�v�1����p	c�O��*��P���_� h��j���q�	��qr�(Q���^�e��V��Y�d��Qj�,��k�;0,���k�}��$�:��u���J���uX�}<�H��	��KI4�F��__j��lGޭ,���!��I��מz#UT�����j@"Й�ܦ�I��@�	����ji4�U*rZn��l[���F�BE�7o1Z��_˽�d��~�A-ԁ���ĸ��Q��;VVU
e.3�̟ɴ����Rztx��e�Hc#|�H֪������M�Pn�|�l�'�F�ᩛ{ǣA�=�!�9���bo��=�y����C5JN�A�4�#�N�����y�h�9��@�I0��ߊ.㕽���[t.����!tI��P`�k�᥍V	�A���ڙ"o&6�j_���p�N�ƾ�4����*d1䌚���)��
BQ�#je�ͦWj����rɬ�]���^�(����/�+���?J�?�8K
�LT����	>�Y��$J����bLӽ�ڬ}��m�RO�岌,��7l!W>H� 6�Fȝ��9���s�_�LW�H�ht2�)ǳ��r���4�Z��y��I���#]ԯ�ͨЯ:˷��l�TdN_�[�vq��r��s�@�w�P��:q쎶�vጔl.���G1)���S#ޱ�o1"w6��Hc��m����9�qɦ�{�7�\7�Z9o�z��I��x����<�~�
�ϴ�գ���̪y�Q7m��r���%�cEӞ�O\��]ܜ\�'�1F:	$6��$vcg��,�n�&:���s��	��$���W��GXd�86d��vT�z�>WH��d���N���p��n[e\�<ܥ]����^r���>{-Ti(<;���5ɔ���t�\���[�Ǎ����_:W]��F��Io���V��R8��O����Dv�����^+\V�hc��.��L��KϷ@����K�I��b�X�Ձ��Y@��X�o@�Xj�13��5~��d�����IhI�j�������(Wd����y�`L���뭠�`� 	��:V�bLy-�O�P���K�����_��c������)o<�r39��v��^7�J�+���ɹ��Q�&�\��d�	$25��#3��فS�0�&Ght\����O1�G�M�Y�ć��Z�X7��@z.`=&C#J&���*������w������gq��_���ҵ�X�hԦ�K����V�{t���R�vQ���|V�KV�پ���*����?� �!F�o0���\��)��.Z�Y.�1L������^���r��qn�v;�e��lebB,A��'�L��⨔q�_����1�?~5�~��.��εQ'�� .vҨ�Ma�/o� ��!7�ḙ�>+*����ąZ=+��uĵf[��i;�~ ��<�:���t��V-�YDZ��o��~��ҶmhR�1�K�y���R�v���6���f��\�i�f�鵌Џ�O��rT�E��~�:��v�<!���V�j����ȡ.��9��_)@�Q�ƭ��^Ex�<U-��!�D�GA�<���|WOLR�\\2alpSH��v����d.d��j��^�,ϫ"b0W�6h�;MyC0X����f+�!�)�#|GJ3�W?1qA�)�1���I��y����.��|Ji�,�h��5�"�C����ïZO͎z�0��y����m+����e�Kgeԁ�+v����&���D�g�>��=�U].�a+�.���}|��\c��|�εO�z�%�(Ú5��Һ���3>~->���]i��K�C$$�%�;T���h��?��|_��;�LYb��|gƏ@͘���Ώ���z﹧	���TT�t��L2�q��Ql犧R?��2�z���b�4v#ҽת_	B��j�
Bz�k��ln��`���p�vfP�GX��;y8[�SB*��8e�����R�<Z���PG�c$�޸íK�H�ѸO��Sq��E�Y�E�}]�f����T�C��Ci��(%�݈���#!����� ܳ��k}ֹ��6#�∛��^Z�5#^6�M�l��K��&r'iS���ՠ�&	Z�?�|�����Q�&-�3iIA%l�g��Z9�1s-��>�{!D�f�-f9����.)���?37'�YE� �__wD�X�C<�cg<�b?�ey��$���&a#%�����t>�ʥ��?�37_�pvq1�Z%���_��\���*�>4�L_���14��8*��������>`�n�ZӨ�-��vXL�u9hu�t�9/��Ґ��5qY�Wd�·���&���Ù&�������Y����f���U(�sd���I�9�FK�Tɧ"�Oh!Ω'ꠄZ���7cɲ�F<u��u>)�����"�/��䟋V�B��K��,�����g���56E��H�1a��>�z�F���A�>�lޥ-ϙ_<NR��ݻ��2�"1*��|�Γ�e��G�}�)m������6ݔ�;����Cz\��{NIU���1H��M���O�M��i��a�(Hᵇ�X��ڿ	5�x�Kp�PB�i �h�%�@�f�����w�ID���<K�IGZ�� ^��-���/7й__��ӱI�_�C��SV��V�*���6�����L%j��é�@�82�t�����<��9�UO��|�O�����=O�����6�V���ܼ����S���u5��Q�Q�B�
��Қ�ᒴ��Z�qloެ��tL\~����Q}U�Y�g�(7� �,<��wv�7:�x��g�9�]󥚆���E��nk<���ܰ�ڞ�a���Mxގ����P���;Ƹ�����ٛ�v����%���1�f�T4VT�|�\�\�{N���(��������������a-�_�� ����KfVVH����uS�Q�7�AA��W4�,���M��~�T�2��P�=9��ޓb���*��[��$q�\EQ���P-��e��4����x��<�{΍ݿrGz+w�u����H�~B��vN���Ӥw�����|°���@��q8������T�i���ڳ�ؓ�c��,{Z)c��sC|TA�8"�إs!�A�u�%�`i��9���a�6�G{~+��Vܼ`l�՝�%��c��㶊���/k����7�j}�ܞ�~)�ˏ�8�e�0_˚�]�����:��,J�J*�m��3 ���W�{�*��z��7��)�o�'��SϿXH��B�I���~&����M%����-�RKۡ��o�9��&�v�}XNݽ�KJM=���"�c+��hD]�̝3`.M
?jQRY�I�{���˛�����[�ۘͷv��^4?�A�K�vB�:�Oj2,��̒�J��Fo��*
+��ۦ��u�C���7�YK(���r"3��~��sk�<&M�M~��(��n`��j�EG�"DZ
��"��RZ������w�TR��[�Y�[_�Z��[!�C���,SQ;��8HC7g�8�ܿ
��2�Y}�.�?}|=��p��5t��M>���VD*Vm%�x2�h�0ʐ��f�^)6��?��M|��q8ooG�};�#U����5�t�Z+�ʶ�¨�/�y�m#�#��O'y��×�@�T%��^�HG$�<��3�y�/C	G��\���R@���ƛ͸x�چ�'@es=0߷��UM��adQ93�m��4m��>u�1W��|dW�=2��<�N���XF ����<��k-D���	D*ȟ%�
��>�\<���0�/N~&�t���g��Nչ����W0�� �3��Y�wE{�@�]U���l̦vD]�#�;�K���rʵ)}W5M�"���o�5�`���2�!!����e��i�/C����� ��yh
�*'�1VЖ��Q�L�YVm���/'ԕxB
���*���R�5p�1!+�+���6�6(79��]H	`Z���u�o��ߗ�R�5��zXצ�%f�:LF ��SN�:nfgz�9|y~�][�ONNΙJ(a�kq$��2�HPzzzV�d�;�w5��R�M¶�H	D�YwC��u��)hؘ�_δu7U$��Di'�n�d����G��r�����p��������B�.I�������g�E�~�Q�߭�(�j���KA�gr�TT@�=��m����Q^�3Iᚑ�<J�������n����^XlǰX\,���ӆK�����kup�P�}�����m����/���I��K��s8͎~�i���:��l$ߧ��������h�p��?)Ԁ����c�2�%Ǡ���E���{�q�<�R����Z �DwNbH���-��@T���a�w�R��,B---��{�
����.�`�k�G����O�]6'���~Ӊ� I]{!�5Y��u �e�[)X���>��]�p���r���_$��soO�N있��%CZ�T˂�\���%`Omy��:��g	x��d��ֆ��:�<��e���f<o����3[`�z_"A�m��>ˏ588HJF�")9�@�x\F��+��I�V즔ڿ�ƽ������9&�����#h��}�U:[S?��#���&z:�2�V�M�����O:[|H��\e ��(�����/����#�����ӛ.磦/���`�;$x@�&v�nޟ�V�n@^���%�B?g����Ǻ2��
GK�-�,W�q�ЯkZ�r�*�{����\o�zs����đ ����###���В� D���/ŕÃ�����e�����(uTe���Y����������gR���sw�(V�yH���AJ'|�"Ĺ����W��O4��w�[*���IǗb������܃��h��P)����j�a���dx��7���ڼd�XFx�O}||���ݼ�K_~!!���?��7�VU[3x
�!�D	j x�;��6�Q)5�"�N�ԩИj�Qר�$�N#�66C�H�b����J��b�ӯ[�*Y�j��2���Xo�#�GHH������ bQ����;^��,n->6!:=)f�ޥ�jǃ�ozE*E��o 998�V�2��r7*Q��M%:m��AhllLJEu�/��4u%�67�m�w)j``����)zpx��t>j9�´)��F�ZR��6i�ROu�k�pm�i��+���|����$f��VI��r����z��p�{��
L���M�F��0]��H=L�&�u����e@w.�!v}���N��[����>�����|}�(���)7V�~�_��ҽz_|��I���$����/"~����!Yq��I*k�Q�ৱ�1'��	�H^3����R8ۊ�i�L�Kk���klN$xJ�L4qg"S&��˂�����IN��%v��1�W�iy-%)��L�Ħ��ۧ���P(Sm��GA�t䮫9V�����	��x�:	��<<=���d��W
<�oO���Ćzo,��h�GQ�NG�Z\_�':�{푹'�M�,ԙV�挍���ݣ�|���oM}�z,j,{U�{F#�@������%��9ڝ�����l��U�v��X�l�هsc����k"�.d*�}}�k  3��	�b���l�TP!�{T@YFF��/R��9��١���Ϝ�u�����r$!4j���t�wBJ)gU=/!R������z�y��&L%)X�`o�E��#����[Z=<<��Y7s�hl{�?G�x�8G��ń�E�P���#��i�s(8�FD�� ���d-fqQ����y�Њ󤤤�V
�HPrQPP�F ��%z333���D��"0r���L�TuȺ��ח��.�-E@�ilA�����u)�5���8�ǝ��O5ֹ��,h 9z��v�ۺںs?��B��&"W��Iг��͍��T>+!: ��V>�Y��%�k��a����MT��c��z�>1 s�����gH��)�nT8��mLh�	�s�]a$��}��p��l���y�y�z0��	���u��P�ʗ�0�]������io�I���H�� ?:}���=^�y� %vzή� A���~�s��*_?ޱA��Ǐ8&��r^^��K�
��,�빸p�^����n��QQQO#������y�t �JY�m�N�8��*,g�E�	'�i��F�l�x;%^:�8I���Έ`�h��j�|4[�7���G����j7W�9�8���}b~3ss���Z�5�.8��L���莘�X�5��C;x	����<U���9Z�-5Y���E\�}��<	g{H�c��$���y��ծ���*ZU{(|1�@���5�@��	|t���*������kOl2��1I���h�G�c�kt� ����a���2Ú�:j����ﾅ�Y�ƴnR l8u�_���-sL�R��jjj��N{_�aJ��gt��eǔ�ʦ�K�S}E��E%���ܯ�rt�Uu�=fIB ��_�.��{H��3��f���w
����c�V�'�|[��N�'/c��g&�[)^B8�j~��}}>]nv �>vx��z��;:R�������i�h�(mo'|i�}��Pk�4�*����D䖶��EζiZ?d� �-��i�����J^��.Æo=FŊ#$*9?�7(@��MqE+IG�a�d�Mq�݇,_�=�<D�T���&g�Gk<���'�6�qD�gg5�^�~ekXFֆ����ծ�ʎ)��z�Dᮻ���T�wh�Oӯ�r�Z�ǔ�/k�U��ڮ�D�t�H��SN�ϙa�V|�zm�f��*	.�r�	%@�G-8��\���#9�p�����͈SϝW���[?��5�E���~�Ӯ%%�Mc��& ���7'�q���~ي�����g8���f(��`-����z��E�!���?������Z$H�g�^]ei5�s�w���~M��l�Y�\����JE�Х�G��]_Q�ay�X�8�,�k���یE����6����x�F�A��g{�d����g6�ݓ1@ܱn��<�%<?�Z�B��]�₞����F��$i7���2(�1���@Ѷ�irCo���~�Ip�< ����%�'=�~����r��\__Sač3�j��)xW�N�I;1pb����������(ꯠi�[J�+�e�ߺ��17�pOhcD6V�#n��\�[٭+tt8�(���F(\hS�%5ʾߴ3���7�P���)'���?�T�'������,��t5S�Z0}�NY��y��2l���V tx|(������5I�n�9��>�2��V[�Cf���/{c+���y�z��R��n.����7/�n�n��(���;5��'҂�kғ}ШtO}ڝ���5�Pd�K�#@ *$�U�刘�����`E�Y�X�]3y���p�<u�I2M|����h���Y�E�6�;8�m�w4��,�&2B�3T1����ɜؙY\��5 z�u�?a�ؘ�:a�����,�x���IӬ�_`�6��æ�W��L��Ӱ����C�1ƞ�yКBo@��,�Y�����!��K�7�����+��L�ix�+q��Ǒ3����OlV�d�^ӄ��H�_��%�����aGԀ��U\5�r\h�&�íB+#@���i�<�A4��hom������Sr D�+��a��¤B�4GZ�i�I�R���)L���(r�5v)�ܹ�`�:q����]4�*:�
�벌� "Ӷ�g*�\?Y��{4��ZX���l ����d}��Z}l^93;ccbc�@g�D���0R�aQ�!��)���1�l�ˏ�\�'��������y��d����ظ�����CaSV@��)P`ė� G�Cj�`������8j�V�H�ؑd�c��@L �������I����u��]CW7�]�O� ��w��2�Zm�ˬ֓�$gd"�`g�P!�b���i��'�&
�7v���ʻ�$�Xk�����,J"�1���7��SrMhxy��I���S	�n.����Kd�,i��2���Z�s=�Y;�bWP�d���P�}�ͬ_i9dd��/W,]�������޾q��R�]���ϩ�����e�'��H))� �r�Sbْ�y���ɱG��Z��A�	\��#��|h"tm{0zQ�%�/��W��fB"��}`����S�e�k,�R9���Y����aHUt���x�&�a{�@��Z-�s}�8di�y纬��gt�(�+��^*���Cql�i<
���)�����?x��sv�75��:�A�&�@�I����G�Ge�N�ەFz����H�ClS?�N�|��(\O��7�B7��k(����x�
t����%��I�A�����<Й�AA�F?��:��=�A�t �V�U�>�6oG��"z{z��`�ǡ&�CX��8r����V�|R?�D��
���܇�Jɰ��a ~��#�g;����gZ�~�'��;��G�f.�l�ݟ���2%�몙��M�4E��Y� �)gĢ�O�>[$u.���q��p�'�H�U��Áz��l��fY�LF,\���D�*HV��Qk�l��QjH#��wԟ�� �e܇���ࡦ�;:���6r��d%LԿ�y��N�Zn6] �Ȝ:��4�2�H7�z�3��Ȝ����]_O89q�6j�'1���Үa�҄W�w���N��AFI���������4am؂�D-=���pI�k즘Ɵ5̐���6:ː��w�]�1lݮi������b��/�"G�į����������1;i����s������L�b�pr�<�B<8<H��~O�9`����;��M5�u���O��A#����-���gm�=�I�5���=�(����$��a"�ş�e��&�P[�Iƨ�@.#&�J4��?��zO��C�ά����S��˶Y�jw��������]� 9�Fl��������4y���#��1~�� a @�cH`��N��h�d��t�ǵ#��9~�s%�w�zY�~�&`g�zp�S |K���-zA���sG-C��vKAi{_� �j�3`�7�q�T,S��a.6'7����a�]��u���X.O;������������c�D�AL�SwU)�dIQj��s�Ϊ�e+�������V(��=Z��.?,;�)c�)E�Oe�_:� ���` �đpQϋ4}b�8����v��� �\U��ӽ%x$�dE�e����T�Z���GU̱5FZ��\֧P�S{�r l�{o�O�EU�;99q���[��9ZA4^�_�IHH8{|�W�Y��?j��&}A��e�z���Y�sϦ#GC�7��⬾�8���M����1""���V��n��v���i�4��?zak���z��x& o�@���~'�[��#'6�vp�o�'ɔ��uU�򞦻(��{��ݬE�>����Ie>�:`&*o������u/�{{��T����?�s�Rۯ�N�q��N�hu���W3��r��-rq���Eu~fyy�c��t��#|݂��8��6a��X@ak0��;-7���ї ���|������!U��y��{;8�iq� o<�
��v�b�h�rH;e�O�x��cŅ189���	��ߪ�ܕ�ծ�GW�X7�e�2x�w�(����,�1U��F[���0�W�S�w�T��~���b<i���YZ���u����k ��Fw��B
�ĭ�Gl��EG��LZ!D9�^����LV��n��J�����@e��ǇtZ�V�$岳��@�s�5>U�.��L�_l�'�=���U0>Z��`�KS�˗'���n����c�k���e������"��;z�����b��B�qK���R�&7��`E:�
���^��,�aww7�v�k�I��r��w-[��B����F$�7�VFl����������1~;I�&�"YQ�W�1a#"UUmԬ�_�������L�@2��#��Glf�^�zٵ�]R )Fb9�d8�`suu�`$�䈅�X�]�����Œ��M�\�P�Q�g�h#QP���7��1�ȐRS�,�ֆt8�
�7�v4T?J}�F�#5,VR��������ᩕ#�5�KJ��2��h�F1�����G��.�ָ~������jj��ϭ[���	Ǜ���!�}���&Ԏ���3y�8}�Qn�ZD3���Y�@�W!?OJF�s�0�Z�s9)��x�
m��%�����������N 
;�'4^r�D��n����^f�;��Ԯq�a���k��&��C�l�A/����"�VQ�~0m������_`�����P	��:�&Y�58~M�\����l?����'O���"�L�>��H��^�դ��#_o�?��2������7-g���Z=b����������+9��XC�4� �����O�������F%�ꨕ����w�ۏ�\�zW��\����e�V G��}����b���������67�X��d�f�e)�B)�|���(���ՙ(N��ҶT��2�mlDh�ا/�1[��vr�����E?:mѵN{9QPP`p��җ2����	����/G�r�>6������HN'�r�=(YQ=�l�����jw��>�:�)�bO8���d-�v��v���:`N]8^N�F�H�äcH�η �q��&j�DePm��f���>!�m�-��*��K�/Kp�t����'V�aa�:HU�qѭ� QAخ#��;W/U���+3����yn#d�9:��;�\���=lE�P<TG[\�#��2���23�&����Z1�w�D�?�Q)]e�L>�[{<�`���5�<@Ոέ���'��3uN���=�L���T
6ĺ�R��4lNڂ_ 0H���f����{*qC �%�R߽?5����Uا�F7�ܥSn�gX�~dX���x����is�D�ݞ	����o�m���֢6�7>������L��|oH�z��t%�a��:��7q	��O�����)+��훚��^�+@=�s��4��
�FQm�r4Ѹ����%���o����DY��Y����~���F���#���`�h@t��W�T��E�j�u�����M�Eс�:_w}�p�g:�@[���,����Z�A�M�F���}\S�l3��rZ"�f̠�CS��IƜh��&\"�~3���/2��2��b�i?-d������f���:���q�n&s�s'v`W�-��2�zCn�T�J)������Hk�ʋ�K��q{�&y�a�ܤ���1~��g�����>�A�`�v�^�`����Vէ�8l��3�D� *�B{|�)�Jc�e�/~�� ��EAt��$��e��WV#Y*�3[g��t�K�����\︃��A��ѿ����ی�O�']yԑ�r�|"�-` �7.�(r�����b�Ne���v��ƃ�K�5S��IRR�r��\���T�V��K����go��Q���B�[7
�n?��k��ٹ1�`Ғ��f���ص= ��G C��Oy(�	c����5�H�N]d�=����'p�-�\z�] ���t��������<B^0w�?P�9+�5���1y��u�$����D�lW��gBuH�d�m_��h�V[��>�����j�}����6?�󕇺���� ���x���O}1��1*���y���γ���+��� &��hA��*��dz��EBE���I�\� 됵�!�C���(inG��o7:�1rO+il$�]s���]UH$����,�M����/Wl.Ӹ��x�����L�����=����zh�((�91����!v�Ɋ�bu�I��J����!@��Vl�kg�֌�ӎ>H��E�.�z����w����|e>8L��CF<3���.s���c|�����1'RX��;iG---�;������Iv�O}O�g(W�FO~ex⃹rX�����d��_�=�!��������]�C{���6a���Q<����}�{�B�xR��K��  +�z�X*��1������C��M���~A�75O�.,M�o�ok�T�\���cK�4���,\0Z2��a�C &f��Y�+�瘢��!@k������|���&j�Lik��D�R��!#:�qrX�nS\�0Qh��#��g%��'�b���Ti?�Wb�뮤���}=e�1�sfn˽A�t�zJ��ɲ:���.��#��xɐd�}��)���d���n���k��$�.��=`����ñpu�5}�˜����yO�~�l��Q�'�N?Cl��_�kG����+�J�=����A�e(�ic*lm�kX\l�ax��E�K}��Ggfg�ȳ�y�;�t�8�֍Sʀ����ZhP^����0EUJZ�l��C��i���,��Y$hQ
˾Gw�ԡ�\�1��M���4�l�������w��{Oe{V|d��/��%XY/�Ee'd�Y�K�íJj�S�R���+��%��������uwS���>�V7������ ��P$��{���K����9����-���n���s�K++��\���sʻ���y��n�Ϸ���lBG,9w�&�8�&tj$��eK4p�"��8t���Q�Y��5�l�D�e��*��̄��X�}���9�zУI�0���k�| ���fl�l�A���͘	~���g�����FA��U��(tm~Я���Ѳ��(�29ƌ�I#3%{��L�lX�:����y���|�0�~j��x�bl<�2x,+�T=�i��ŷk��ͪ�[::Ǌ�ѭ{/��
G�Jx��f^��{�/�A޿.��L6G�L��C��0���`Y����F��|�2�Y̯��C�/��ss��"�,y�}=�BB�~˼������A�-�N����z�D���m���u
v���=Z�pJ�T��Mx��u�X*�*=�S�c{��p0����]�Rjt�b!:\�b�w��c�]E=���N7��$vė�c����d+P�L}m���>J<�c���(���9bI��w��7��0'��^����箸��c�h�~��Z�%Ӆ�=��!��mH��	b"�r��!?z|U����1�H$��ж�q;el%=![�1�3�i���E�{�0��gg!Tie�O?�"5��bg�7D}��	>N������7��P��៕�}"S�A����/�>��C~��ݼ}L��ݼ|������~$�qqpdHEPf��b~�4psS*������Pqa�wL��`D  �C��V��#�YE�-�e�	ë�a�S����(��p@;iR��.�i�gp�� ��D7r�`�����R8r�ޠ|}L.�b��{>�� t;�^a�ѥy���3�3�&
Ќ�E}�}��揦��s�)m�Uc�08T�k���
o��oN�}v�m�V7^�����V��2՜!�
��v�ئ}��x�tG�o��w��V��脠�&z�]���40��]yxl�FR̂�:�+��IS��XS��y��%s����=��$3؜��>@����ϫ7J�G�������p
��縌�'R��9����O+�J�����F�������Ek@ӿ���	��Ǔ�77JWeT
�թu��B&��xs��`����a�t)u���r��!�� ��&�-g�#9a��$-a����Mw+�����ݨ�l���G��{�[*���1Cm�u�x��k�Rp�%�={&��_��o�0f��;n�ssn���z|i���ek����uD�lĤ��zYJ��δ���x� s֘EA�
�	4�Ee3��3\�4}Q{O_)xoPW��(�����4��h>��y�N��]f�1�,������j�c�C�pg�|x �T�f%�I�sA�n>Wh���*��`�㗩k�G���j�v:�ᶘ ���DR��U�<�I�(<�HQj���F�F;��ʚ�F�W��=�t�&�2�ɰ�7�� G%q��2(�0V@KK���G[����z�OV�����ׯg�5?�Q'B�9B$���Ls��
�p�Z}�_�r"�g�e�7�L�瓴��s2�ƶPF� �(�|�`���ǂ��q�CY���Z��F�7j���w `s��;�[ƿ��=�q5Hi��<f��G=����٩Dv.�%�$�'���1|���)>۟i5#��YJ��´t�j�ƛ���rf��;��4Ka��J�0�Շ��*�[�W��6¸a�b��\8\Z|-툍SnRIF|y~���)�숐�wӆ��V����]���m����������]>}U�;�l�P*�I�C^�n�ug�^9����O&~W�HK���J|�����A�şt�z��wQ�Q�]9}�\�R��ɔ4n!DL[�,W�b������x�F�%O��6(����_���I{�M'�Pj��
���%���n?X�v6Zh��֙��4zc��5,�KT�YM��<��6��pr��u�����{�]~����.�g���y��!������ʭ�97\�����
	�}q����_�\�+f�t_�y�5�?���Fj;OB��χ�|ؿC�
;�����>/rF9
��`bbP��n�Lp�[2n���y����d]x+{ݹ����[��u���2bʤ$͍?b�@�C~-��J9d�G)t?I���^�ߜNJe�BG.�W���ll�u'�?x<��(�d2BOg4�Kg
xГ���H(�+�%	�𾩺uX#(��6�V��*�����׏%v�g�����g����~��˒{�e�^ D�=�`?|�U�m��E�Xk��72��:�(�ڤY��X2�ݮPopn���yS�-l
["�3fO�?��֍6Ӥq�`�z����a��Rqy�7&�����>iߣ�M@�=�. �f�Z��w^!%%�c$z����aʄ���f#��]��.{����7-��Oo��pB�Ȩ+��]�{Ii�T����L��*�޵A���j�%��,��gW��l�{{����G�E�B��P��};���C	�f?`q��/�*�g�-&3d��+�?Ȅ����� �@��6�#B�$⦺���:�S^:�X��|_��/^���"�e��O<���%�/��D�~�W\D$��	������o>���:U�?\�R��[��#�Mp�vRE�GJ����n�7 ��=H�5��� Z|<n{8��v��'�o�$�2h��/�98�z�}�xl`��C��fj�Ǝ���q9��c����ZX����:q���%�f���'�z#Y5�j�@i)+���D��W8��I���>�`���L�n�̻1��6�?�5ߔi��02��ܤ�G{�P��	��^��5���������'��Nz>O27dW�j*���wk�Q5}�x��;gy�@�s�'����f�)�H�UC�{��}���3�6��r!f�����.��fΝ,Q��v|4�u�F�>z�yG^�<bM\�h��^��&�lt�	���K�o>�0DT���Q���'��7�vV��={��5�=�����,�q���G�������\_ֽ5�;^:a��p��-.ԟ�q=��W�!�NB������g�JL~@�ZZ��)��LtPeب�����i�
9���N�94�S��I��|��)�vm�4~(��!��p�:�/�N�f��\�t�L�nX���a���\���	���4��V0��W3� �l�*n3�=źɉ[Գ��5F|펴���}��W���o�c �V�;^�y~rV�O��~V�g9����s��8�ɷ���<=��n��:j,����W�����'d%D�4�+t��(�s���x,��`�~R��������������Kj/��o~-�I����e�V���T��j�d�lĺ����>����9�^�W��vB�Y+�
���b����ǭ���䙟.y�.ʛ��n<���2��m>��F�p��_�`Z��A{��]�'y��Y?�'9��vy+�V0�V�ϝVթ)7����9�IU�݋x��R\;N�Rф͎�?A�g�Oy���}xVRug�/!xhiE!�eH#��ΕI�o�
[�
9��m��?ݛ>3-V��__�KH$���륄�I\M�<�c���:�:g:77w���[����y��W |�������;�G�y���P��������S������6����������JҾ���NNt�Vh�mA�{��k8�=��3���<�{�7�Ŀޓ\STq�&�|���#�Ԝ��q;���9ˡ������"˵LgR-�md�q�H\��If)�I�;������6g��(GZ��[�m"7yn����w�hO�I�Q� |�::L�6\|�ڌG�?,L��*m6Kj�i�Ӣq߿�e���#�ݡ��˻>_/)�Ah��/�!�}���F7�(�s=��J	���$l÷�;|{�����QohU~-�n����f���qkgM�2�*K����4T���
~�vJf/G�����jf-sā�xv6�c���yw����҅�Bq�}�����c����yI��[鳚�#�������"S�&i��O7��ð�i9
��X�6���>ʨ!P�d�"�X��jK�C0��F���yL�-�ہҜj���N�*[*4ޣ����Q�_�~���_�T�ڦ;�n�D�N	t�z�7Im����ZC�C�T�6l���Ըj�M�^B���{Q�az ���O����Ha���=Z�D�h�OK��ꯉf��w���j��yK��eI͑�F��(�T<�H<��j˟0��	T�L�>�4�6��͈/ ��gH�]k�O��td8�_�#[F63��3O�7�t[��A���!�q��� �DZ������Uw��D��j�A��a��MA��Ǵ0?��0ܑ��X��W�Z�_����� ��~�W뛥�U9G��U�#b��[�`�w��(*����拧)���v�����V�Q��� ׃�ޑ���1<��Ս��C��fC���˖��}�ϩ�i`�����5B�͂��ꆥG/l���L4� �*qOn\K�=��:��m�8��ͤ�����y�,A�zUsl���,���������nL���I�3@�́�1���vTN!����tWjW$��_a7��y{̶<'S\�#�[����>�}�8�o�m��"�6��M8Ap�ԤU��~�u��`n݇�"\x3��S/|������L!�{�4N��(͜��6ق�ڄd��J�,�X�/1?�����~,;z���KYR7��ZC���efO;������wT$��f[��W�&>v��%������H���wBm��r�Bk�ķ�<�c�!B/�
��ww�/'�/�������3��;S���-.��!��ud|����>�7�����}���/��H�{$ܤ���2h7qy܁��e9�~g��@�������c��N�ʲ����۟4;��T�ry~�{ʜ�>���@�`��P8>�T�YEB�=�^�3z��<�{�Ŭ ��N�	�:�|CE�*���/7���lY{n׵��m��b'<(p� D�̮�h�Fʔ7�+�'���<u#�2��Ga�<3cP'��8=��7?��	���2�9��sʷ�IL�!��F���n��nFGU�RD�
&�g�T,|!�}����x��(
H�_y�4LQ�����W����@����$��Q/#�N>�!���C1Iǆ��oE����K�,'l�^�>)K1��A�缎��6���L璫H����axqGr|�Kf#��m�Df0Q�bl���0��[�q�|4�c�Av�-Ma����k-Y͚�H~q��A��>�-Z�OEtk�����k9��j��/��pl�	K�f�m�E�,���=�!���X9A��le7n:�.�5�g;,��Z�b��𩒖%�>O��#t�����c�������,�lO�k���'R�3r� � �a�S9z^��_�W5��q���/�1!N��rH��l�x��e�G(8�������T��|iY�#\v�)x�����ea�~�/���xw(%��-�/e���'��MwjMwS���pY*=�M1��2 !V阏NUI2��|������Y������f���\�<
;��P�U���G����sf��	=m���_�m_�/6�~[�bE�4�kj�ט[�Qb����U��S���+C���<d����ǩ�(*���)��x�4| H�G=ɯ+�u���	�����i�3O��-�'8q�]�,��""R�U���&U�o�F���T�K�{t1���'��^%�D���:ڀN,���ekg�$��|�$���J�n�"H#T���W-U����`!*l�"X��=�%盝-�r�yj�l�uߎq;ԫg0�>c%v�g3>�o��?;t��B?���a�l1�g����	O���&Zѩ�hI6�M����_���I�^E�$:����)U�W�E	r����j�9��+�>�C���8����Cm������8נ|���Ο˛�X�,=��c��s�˧�Osޯ�D�n��;�4 W��ؿ'�L�zv���c'�e�T�9���zz�5Ĺ�k�?�G��ˎ_�w���rA�Y�N�-�-w���*!�4��?��I�y�u�f<�ɱ���Ta<�H6�Gyh:���C��?�S�>5>B&�4��{�/��Q�/��}Y��d�؟��ɢ�m�"h�C��8Ⱥ�Y�[��f���!�]o��j"�
��u���o����ڍ��m۶:֛�c'�v:�m۶:��6O��������k��`M�����l,i��&�S�.M��Iu�}e��ez?
��_����|$�@,=\�ߠ��1�l��B��X�!F�=1�]�Q��mp��_�
�a6 ���X�b��z�E��znl>5�՞���]���@|�����~�7V]��>e�f���[�*]���]W�(�><<���w\-�2�K���-����ǥ6�~SG9� $;ĳ�ﵾ�a�>/�<M�G�nX-u��i�t��r����KĚnQ�ho���8dw/�r|�899��u�jk�&�Y�ψh��>�@�e��#�Sc�*��0ج2DVf�6/�t/���<gƲ<k2��q��c}�Q��菠bT(Y�$8H)U����L'|��}	���+Q*�}i�r�{_�w7ǭRj�������޾�f�N��\�X�w0��W��ӌ�D�sM_���Ǿ^o(�n�p׍�w|�U743�&�fj���A槫�0[��/S��^�^�rĈOD7������D����|�(�������X��=���Æ��kA�L����x�����t���Vg��S
�p3v�����.м�S	�#�ӬY������`��%��:�(u���C�u>6!N���A�aq'����ף���hl�>��}DM��\�6�7����-)�|<E�֖�s���?1��A]��fJ�C�F�k�/���Ic�e��V
2#Ң+c�{���)"�*�<b�L0��<��M�M�<���z%�n� u;�J��E�g��V.��Z?��lzO�!Bh-���~Y��Ѫ����H����mZ2+mS������y�˃�������
%N�f���[}����v�n��!~'=���O�UƵ�e��*:�|����v"�u�?��Ň�17iۊ~���U����0�!\l]����-����M�z�ڡD�}#��fR���Sh�C�\�߬G�ִ�M����NTq��N	Y��B����l�LBw�9���ǲ�w�b�Ȟ��� �"Ŭ��P��ƅ�����/�(�v ����.�(�6[��}l@��h-��d�x�3�-F}���)Ըzt�\���o��S�Rώ<#{��+G�[D�/ckox���
r�2X'b%wJ�4(��`��P�<�W}�c t�j��$��%�)<;��VE�/�S)�6�S_���H!���Tqo=ݍ��S��B�H���8�򊅬A��s�gK���ϺK���Ёl�c��HTQ;���5�@�d�~����'�V=�{��%�y���J�{P�õh��L8�m̋�)���5��q�[��B��ܫ6�U;�:|�:��Cvd�'��%�q����bޔ����kZ����[s\�����Yb��Z���]�:5�����&ti������|�c�o���M5G:�����k�W�*�0A6 ���[��lz��lEk��q�9[	:��g������~�7D!f��L[u�M��~��~�3u�{b�Me��7L&G�,xk�J����3VJ�4dJ��bC�|>���
6�/��j�J�?т�]i���jhx��Lj�L�����MYF�җ���f�WNo�oͽ/��{3���f�q��5ߜ����2�Ǽ�Ti��� �^�<��]>Rn�0*_��K�}��w'�f(�D�Ze�	�h?�&D��U���y�h]���-� �
��\�v���N�q�W8�������S�S��%2UK�Aٖ��Ԑ������u�Cz�%������&���L��y��Tzk w��w�\���ne���%Dao�v[_�n�V����Q�5�`�6=.����ײ�	�J��#��Ti=�S�(dgS�4֋��j��%~�߇U���i�&�D��M>U+=f�}�U���#3����b$f?
��t�Cn�U��U�+8T)p4)]	S,
8�C�杽6�]:L��q��F��Z��[C���ˣ��k���!��Wm|�+�.���%�i��#�$ʌ��.�Ǒi��jH`�(���޸ٶJ;�T�P�W>W^���B0��񨆂(ݴr��[
'/F�0�4u�{F[���$ϗ٭<r���é���F�ߵTA��#�5Z������v���{�!��x�
���
<#�""��W$�`z$�Dͽ3�&Q$tt挪����/p%�T�H�)���tk:��#������%T��l��GT;��r�O��o��Tŗ���m	�f ~�ho�fC�J,�8���-o<�DD�>����t\|��c�\�����s;+�.�ց�VC{�|v���bv{�fMr�<�wtSo������>�o�����]rٗ���	���&����c^��|8��q�<W���z!Yo����GL��D���C�h�զ�g�	��k��:#�:!jd��!e���<���//+3p1z�Ik���q��R�[���>��s�4�5t�v�_%�p�\3r9zB��
����c�3����7wrD�9\��)����"i}�0d��X��B)7��D��b���/'������V�r}v�eOن>Q�Ї�������5�	�]ae:{�:K4��B%z�][�D\(�~���W9�`�Z�{�zz���tI�m��E�t���c)U�B���<jp�F-F���20�������!��1�>�97 �}	���c.x��RB;|p�_x2��!��l(�������B��/����(��Vd�H������q�C����}��ϧ�ا�+�d�z���#� P����uzQ&��?��1V���@o1:_��A,7W���t���n���oq���N���ة�1u�����P�y%�bW��;9P�>��҄K�rț]t�+�����rM3'�ο�'&�n#��=VS���D��!�Sʎ�4/K7 �N���Xp�B@.T/M6�k���L�W�c��H�¬���:��)ʉ,�f������Q"��������VE�?ٚ}���S:A��Rc����,�T�eT]�c$��&Sh�g�:G|�=[�����	EGjt8���
����=F=@u��ȋ�=�M���fO5o�|�-��]=���>@	�z����Ʋ%$T�ƭ�
 ���#��z��/΋�CdǪ0W�2_:mA(�1r5�¢,e�+w�14;k���_h��X%	CLO'��Ҙ�F�B;�l>/U�}����.��`~7�x��K4�_��k�oAv]�^�a�7�?�F��]�&�Y�j�_�bQ�<�aw��r�!�0�K�^��`#���#�ܭ�#�=bg��*�tP���_���\���_�����&��dCcS�{���>�d9�w/�=����9.�u5��%q�̑���zUHta�_,8U%��%6���[r�ܦ6��wQ��1�o�#���h��'0MX�k�G��~k��5u\�4��>���+�	9�Uap��{��f�$fˑ�\�o^u�!z����F�#�XOPZ����)��ߤ������T�7i|��)�����@�����hp��kV�����I�ݛ�*~��'S<� ?dj���3�@�V��D�G!�>"�mEf!�-!��������|�G6�Xkfh�t��L �=w�W����!wmO��"��v��%Ū��A:�-]#���"4�%��"M;���o�
�{�P�M�|�&����V�O��`l��A�:v�F ���V�l����w���8�nWt LI4V�����{U	T�:4�B�b��W�N"J�Tq*h1���q�E�)Yae��5�B6w��@Z�J�vyi�@��j�NEeM>��Z�s�o�ի��N�	�'���fm�z��T�];iԄ���U��o�ӥ�S�M��&c]��nǠXF�oS�'����0��(.�o��?�g�=�[)��	�~gxu���Y�'����K \�e�������N�xȕ���XFN�I���h��)v3ֆ����+�'�'�Gх?nѹe��o��D�|�ګF����5�����o�:IA�qް������	\��q/�|�Eb��,(E�(��*�t�G%7Ķ*7�QB��<l�QЋ��Y>��Wc}���V����uLF� UU��I� Ŷ���M9:�����7�L��@��T3m܄�Ŕ-t9J�oX
�BV�݌�T?{6��g
:6��׈M��K�
�6�"䬺""u���!�����;���i�,Cqs���Rg19g�[���uf���G�+"sk�8�4���	T�m~��X�z/��[]�,;b#�ۡ���d��柛[$m�T�`8i�9�6v�!DD>��>a��T� D<.W�/"�{宷��|��KB��/����֜F)~��$�&V\u�;a�۠�rCqL_���ד�"�?����:�阮f�\ed{�'c��ϐL{C�λ�q�:�I!�b��[�e��Xwcf�ah\���1�|[/
�F$dhZ�@���U���`R笭g��U{�f��b(jg�o+J�*E}b��Fĩ3�����k���OI�(��$xP�x
0>F�eo���;��>�p/y��ڍ`�������	�[%��Ӛp���ٕ�h�����:�{Bb(�A����@�z4�?�0�I0cTJ���u��(����;�Zx��3W���� ���\	e;g�!�`�Q����.�����,��Y2LPf J]��%N��eh���B�����nc�`��exT���w�#��_��ծ��b�sߋ����ޔem�ߪ+hڣ�&Z�A��u������]��޿�ŧ_`��){7F���{�ݿ:�#��b���j��R݊T{��G�M�زHK+�I�Ŀ9a~
�m��YU:>�����Q8VG�#F�xX��ݮ�&[�m����K����ѕ4�@?�ʈ�,d����ό�1Ohd��-��ٌ���m٬UejP�9��V"s$j�ω�d�.z�\�����U�n3�j���o�r#F�E��Ǒ�r�J�Yo�8m^b�3��z�����K�!����+�Xx��r� D��q=�����=<�6����q[[G=2s��6���c�6Y���B�v�S1JLM�ٗ
�4��Tf�ӝq�C�`�CA��y��*ؼ<;���t��+�4t�=.�䌗�����r&څ�^����3�
*�]_�1`�2"}��"���W{������x8k�~=���tlg�~��~��d)���$���`oE� o��sm�P����l��C�g��t0y<�v�����
� ��S�o���g6�:,\Ys�sG�e?9�ɺ��ۥܔ�؞��*>
�<2�5��C�?d�����F���@4�`� q�6�n����s��2�,O�z�];��Kw=�q�EO�����߂�Čjí	3hx�q&д~e�Ŭ�_1��p��Z7����i��;�m�Wv����w���2���(��܎uV͝��bn6o����D0@Wۅ
+��gT$�'��n�QOT��
�4Am��@���A����#�Ģ߇q��t�aÿ�*�zFl�a��Yڛ����Z���m+u�P�T��9T�$֨}�#��8!���<m� (���]?��?��x�6�\�|����8���*$�>��o>lؚ�C��!�R�"��C�!�3q�b<�=�T4�g���e�0y�Od�3}�..ޟ&1�aA�-�jp7�k���K��Ol9�Ρp�<�X�g􌋘��˕��Q�w�&�&�~��v�C��%�|�+�@k�;��K������x���(�d�*�VL+�}G�	SMDN�1�ȼ`���<�J��2�ܙBU���у������%��ʲjj��z�~z������(��R��	���Մ�Q|�@ű���r�M���8��m�pooO	h�D���]���1J�<�g�h��x�A��^ع��3x"=��q�*-SvS����y�����N�օ�j�������x�s�P������%��ZrJ���f���G�.�Sv��f��;`��t���� -��׮��Q�6=�!,�����6�HQvp�
-b999#�L]����1+����T���/�=o{���$�+/c�.�a1���^̝���@�z20}�"Z�>��#���C��������+%7�v�ؓ*�oť��-@�Y��]����+獍.{0b&g������*>��0W�QÿoUU��T���t�`4�X��i�s�e��Y�ll���eo���a�S��3O����\��|�ц����u.�ߚX��fx�UMM��V�tOL��*"�BFJn�����폦���0Pa2q����ڭ�������s���;��vI�����ll�^Q��bٮ�"X7�F�bMeR�Fc�F�j���#EP3��Ee�R��e}g�B�1O�|�I�玔��j��S�(/����B`3\}����2�X��0=�g�mi�<Y�ľ+Oߗ@BA{jPg���P��A:�.X	�)Q0��{e*UJP�t��(GK�t�,�������Ǩ>7�>N�:����ix���W�v�q�<32���2�yĿXn���j孋��}]���?ju<d��l��(H�-�?�W����H�\���_��2 "ּ!�6��C#�'Cvy�"�1N>��o;�[�a�t��Q��lQ�d�_RE��ج����)�
F�R�m��r�6<�-{�Qw�	�)����Ldr>��Mi��IV����QCv��<�;��t����\�U_V�C�5�6p\���{�:��G�F��$�Ds���7Y<N������5v�DaX�,Y��*�S��KJHJ��/Tv2��M�3)j��o&�f�Q+HQ��w�=<n�����.���-�i����T�[�:���tǓ�ܮ�ݩ��w���I���oQ���[�xE$�HX�X�:��ne*��}n��t�(�`��(z�¡�~|�������f�	J��P����&4k�ʣ}W�؟�ԧT
�{�_�<ʬVe�8�h!J^l��,m`{_��xg^��ˀ�;ꭇ=L(�s��"��Tt��R�������sj����0r����-o�sޏ^��V>��w�4�U$�k?Ey���e}E���2ZN���۾�Ы��z�S��!�R��25+��1���q9 y.	w@�{�B&��#S<�J6���j���������ǲEGc��R���KݥLŦ}P	���z|Ot���}���I�K�`��h;�r���F|�Iz(��ż_Q��9m�C����y٫��D)�\�s��&�A�,�u<�Plr��������Mh֦bc�5F}��h���ι���<�2'����#[��?���2�~�s���p������L�׼m���K8\o<j?űsو�Ԯ/���]�@ہ߻����L�󭠿[�7";C�IH�/�e д0$�s�E����A֘|�x �g��wȩ��t�L����1���a$_S�e�kP��/��U�X�������
۷����H�FmM�ǥﶘ؄��z\�6�����*�q�6������[iߣ:���R�Q�Vnv��ֿ� ����	�X�Ϫ���6�w�Y�`Vn�b���x��??�q�Ԁ��:���$�d���V#,X_R��3�|w��˯��$S�3.۾o
���x�����=��"R��Zؖ���	VV�E��q����m[[�6����w�ӫ�r�3^|�Z��z0˨�^��d��(2�f���{r��i�,�.�1�3�sHQ���~�O�4#.��1 �HW;��uk����\���i�>��,�V��M)*2>tUP�h�U� ���`'��mK�sy{Q����WGfĭ[o��k�^s4�Ê��HgD�2|*9W�o�d�;^��Y����]�.�+�Z��Kjy?��6�܄���S�\�m��J���q��C�Yǻ��LL��RzɤR�=�.qxj��0*�����9yl��c Ll�m1�I��#��g��d:���v.#'������*��x4����ҹV���F�fb�ސ%���0����)kfl�&DɐePA�bJ-4v�l�1��!��!A�$��3�D�pw������0���)߿��o�_o1��h�j+����͝�v���nK��Mq�K��樣f��(�
��.��X���_�1�~�o"#<�xC)���r?9����6���I���a��Z=@�9�8#�-٠t֊����B�X~��5���Jd����Ĵg���){�~��`Y�(>o{{��gE!��w�Ȟ%-��o"����U�*�VY	�S��̼͎� NlNd¡p�)�eE�4�3�������?�o$��E��A~s��+w����/�	.ʙ:F �ov5
p�#�֒R[���0��W\�Mg��u2
��+���V�n�_�X=q��W
�~�Ǚ�ў
]�H�
``:���ä<�Ē ���%T'x}����EEX~>e�{$�/��sĊ��.�H+g����.u0R�Z$&�ӌ��������U���˯�����m,�\�+�r]�&�&���u��S7�U�_��W���ʨ��KHY]���V=�j���xy����:x�7օ�p`�K��'`}狅v#�nV�Ajڍ���(58�|���Y�R��L<j�#�n''mzSO�i�
�k#��<;n��"���y��ՍO���/�FMﻖ����u���VٿDa����1��W����[͌gQL�O�bBCa��X�"l��ƣ���i�rbb�_�Һo(U��@�r����W<��KИ�6\U&��4��������^Ô�	R�(	���������C�Ď������.��N�����%L1�	�&<6Ǡ�>)h+#>�����t��5��3\�qL*�$a��QvSP�G�{��Z��MVrl�.)����~(��h	�>�1��Ѱ��N!�� ����T~����{�e��6���\�|=�\S� �"�:��1$���v+��L�׿G6��O�]_�1W����f����2�v�؝!��`5x՟W��y�𵸭��d���Z�*�1�^����1���a����=��3A��9rS�j�V`"�p�Jd|��d�l�x"�r%E&]�����cQ�J_3� �E��SL]EI���`�x�V#6D�a��{��ۦG��h����N�[u�zJ�3QD�	�^���[���U�\�����ז�3����鬲I�fC�rN-׍�W�T��N\e _�i�^u?�
��8�Ă������{4������"Ԉf"7Ee�ؗ�����>���ōI�}���1���Ts�T|� ��EwF���:"�zoA��𕓕5��{	�S﷖mx���*#�̢>/��4� J�\��K˲���E���ć�%v�0d"=tó�"�mm�w�z@tOy��`ۙ�2Vj��Bu��/&��6K��I��\����֚+�[μ�CB���N�40�%l���i[�,�r$?]�0���>��r֖�@Rkw���ѣ K��B�r(?~�Xʵ�͖4���E��xK��v�Dq��|MM��M�iw!��헤|�ǵϱRC�]�����}EJ�{�TG���l��9�d���˓� ������$��bt$[9`	�n����wu��c�b�ˆ��T��ы�4�hԅH��&-�4�J/Z��|�^S��H�W7��b���+�y�"��Is'����G�
�骘�u�;�@j���?%�G���p���D:1p�F�0���
3�a�_;�d?��b�k:/y�~ʠ����<S ��Ʉ�S}z�T�)�y_t�!�N�t��1)M��x�Rگm�)?���by�k�FZ3��+
���rHj��"NN�}C���z����)���($$a%�T#]�R]�p�o����-�ŝ�d��[��~�I:f�*T����6���fJ����)36r	�v`d������Ӂ��*������i�d'LW�ݰpq��m��In:\��Z�ɨ��K��c��	c���_m�;��޶�<:z�<�P���x
������ox�bۣ$����1��[�X���.�`���b�[~�:_pz:H���] ���_Y盍2�e�l�EQ����պ/݈*���0_�&�cȢ�����Vz(q�v3>�u}�Iʪ@�x0��|.�xu�碮6��$�V��0O��R��1��|�qz�(�:z���`�\�HM���c�5#�?�fZY<�쌌0$}�d?�s���8�h�j��Ɠ�+"�]�����\k%��$��_���w���q�Γ��q��bD�,�m�����$��$�S��J���wC�`���
��PtL����G�]~��+_���*��n#��cV~r�66>Dr��ѐ���t�ެ��5	Ύ:W�*��#�� �ް��Z\܁��M�~Ϻk�?[��HK������/e��=�7i��n�n��Ң(~.*2�4�eTb����F����@�5�w�Okry�%|�!u!;7��4!/J���_���#��6:�Y�ȑ�RY'�F���\�7h�)-�b�͡�?�e8.�_ⴚ�Qa�L��=���Ʒ]T�e�n������q�{�;C�m�?��g��iG[�ȯ�D�3JJ���4��q�Y���7�qֿ��s�q#kĳ0o§�|"����OPwd����rVW59�o�&N�6��w ��Ȏ��ˈ��)�z�F�ךÙ�e�����W�"�N·���lg�u��=Z�������N���TA�p�@�{�����0Y��h��_�"����i)���6$�N�3��F��>�,_>���7�.��s��MK��|?������m;ZRt磚��SB-~BrE��m�5�#�i>\�M==��ߊ��0�������˓��W��0-!���t��`���]�ny����	�5ɘ��n3�U��G����b�Z��Da� ..�/V�@��a������=�4Y4�Vց�a���������h"$|���9�I��a��X^���<�h�˪�	*�@�Ѕ�4��?jU��Q:��r�ޡ�=������mg�(��D\���°Og�$R�!��x�
�C�Ԃ�^��%�{���Y9D-f��Z��'F����;�Ӆ�����Ŵ'�������R�`�C����Y�"��:�K���ɔn�S��I
����/�?��9_Ti�@W���
����IO��݈�*0����1@��=L%ÚO։���\S�rђ��Q���
���ry(�;5�[�*��3��Nm�w�7�����'���x2]29��^��� ���[�(x�_��$.0�[�of�͌���87]�K�$HWm�Z*�铢�1�S����t�ܟ�wR�����L:���ǕLr?$�z楌����.���W�Y����5���@�x��TG3u�� eD�I���@=;.☊�<Ȳ�z\�������r *����vB��Z��]�,�.�WHc; r?��{�����8��p�jR�(����>7��\�:�i'��7{4�����cQR��wP6Șb7�X�8�w�� �ő��mn�[��_9/��5���<w��˅SMaS?1I��Z�n��w���y�uCP:A��x\eY� 1ȵ5EwHY��R��:Q�?�pp���
+�f�2f��%2�0b�I��ʴn3���5koo��b�����cC\3��������\Ɣ�#UQ!��OZI�Lq�9���/�jý���8�q�N�:��Nڭp=!\^��Gj����!}�z�?��*䐏G8|�O"�{���JۏA2����o_P��r�Y�$�{����J���Mp�eO'����J��ϷB�jVi����1,����,7,��/�Qf͗^2n ���%$q�f����� �KypjP5�ީ&�i��.̮;���k�
��<�Bu�%����
LNO��U�a#������W����w>�Bo����g�W�� ^�0��W����E��e��n_����I�0�]��H�����ӥ�NΖ-�;��X�S:뎾O����JK�R����@Z$�����5�93���,�q���u�$�t<�C�'�.!�h���tkH�ǡ�]����ϭ����7k!L����JuC{w��x��� ���t���+�/�K�$m�NΧ��3z7��d����|%t����3��p�A�������/���p4*��d�֬��ʁ2�re?S��b*r�^��e���3>��4U/R�� 0���}��1�-�րnT�l��'*ļ��7�g#hܥ��ʁ#��bR�b�S���#*�`e����������q�E�G=%�<��G��B�6�O�XVA޵[��:{������
ٮ�����6���0��ϫ�~G��tujTuMΰ�r?Wq�9��.³+��P�]�q�|�ܒ�W�V��B ��(^�v�╒��U���9�n+�؎���1�����.�j��$�
��4B:UZ�E��duѓ/<%��a��ļ�r��P����1F=0g��zԕl{y�=�/gM��g��a�{j��D�o$��;������0K	Ew2�b��n����>�B�quH��{A���>qG���w��5�ki����&@�d5��H�o�o:�S��R�#^&��]V��PP��ӡku���0���,���W�kU��Z*�芁�.\WCw���� �"���R�r����ƶG�_T�D+��:�8�Z:�%�U���Oؐ%kʞ��DN�K���r�>'t�ŋ��f�]�|�����x����'�̳/�	U��3�Z��I�%Ϻ���=�-�8bkp�4�)Oƫtۙ�Q����I�Ḉ�;ZR�C�u�K�F���&6Y�t�Ȥ{l�@�o*g��pԐ�M�x�h]���^rD�R����?� �����e˼$ɺ�\9�)W�>ϟ��Կ���/���N�K�]����:�F��V�+ހT��[C�o��ޔ�
=:��q�;<&:�t��'���]r�kɬ �tK$�#�zl������R�2 &�_���V�<���5;j�J*�_S�lt�5������X���Cj�bYC�?q��(��5��E�) }��ق�R[�;�w[�l[�y�b�'=��Vb������?�R��k\X��*2Hq*�f̖�`�cRF�rj�S�T���Q�V���Z?l/ִj\�7U��ﬨw>��,�h%�I�Ѻ�s"�Z�2�ˇbF���p|\=rX"*G�pU�r$��c�8u�!�@�.�W����{���ԍ�_��쀜`R��m�p�'DT�0�Aq��G^z!�f^�������z6$��Q��w�#ء?Cޫ��WU5S��0.�fO� �U��0@���
�eϨĚ�$"B 4#��:i��v�
Z!u�����x�V�\t#y��vgBL�[��*�}߹)��X7g�3�y� ZȵnG$t�k�w��4�hC�7[bi��աVL�7(����?xQDyF�Hބeąx�/H���K���Yk,�����93EMLe�TD	�Z�mI6�ܜ7:�Ѹ�e\�5���p޴T�zù���mBk�G�ke��q���B.7"��͗R��AW3]Xo>�=��z)�~�1�gl�����l�C���"$ԋ0��-wptD����u�ٗ�i�Ζ��p:�Jȵ�
}/��?�o/��j^��STP�]ow
�5���A�	%�EZUش�� ��U��*)`��FQ��f��|���c�JZ��0�O?�>A�P$�"�����֪m���@�hqr������d/�7\�{ZѾLԞ�#4�AfT�OR:����k��?1�,$� �Bͣ��tv-����Z=hb5��XK�,��\U����'����3�L���@3M�_�jp�Yd�ɭ%�)�v=�Eg����?�Q\�p���*m���_h�Ƽ;J�[�&\���v8k��V��S�S�9��2�e\�֭�-���� ��FlY�k�)��m�����[^,>���|��lI\����x����q�����l���@ń�1����?W��q�)ư�6z����G����;�T���E�H�tח�K�ͩ�&�
�-���d0㷳%�GV?�_�*��s�j@Z��2�!������9�:L,Su^<x���:)�ua��-��ȗ,V�[���N����~��{�㎜�6\�}��Y�e
c��[����[�Z���?�el�k_��2�2O���9�֡��@��dC��ŉ��L�e�m�ˍ�!�0��V;�,A<j�M8�
��0Hϓ�F�f�zrr�B �oF5�  Mi�8�~���	�`����Z�a�Y}Ѻ���&�5"����b����^l7����\�򊁋<=��4����X<u��3%��5h\x�4j	oH|PX�!�6-n'���B$�>_9}M�:��n�����D����ɼ� QpA��k�I���x�_�p��@���mRY�6�qLOԘ�Z�����nL@_�������eWC!
#s`�99��.����{��D��`��H��}x��琺$n�q���]!�l�_�����(�L!9�6�2�`+ط���w%�UA�1���\�W�TQ]�Cɕ}�=�#��&������ 5�	]�=�����d��f�0jA�N�/��\�.������
���jH|�t�W�A��������÷�D��yz�ᇐ]7\$-~�'�/�0�}�����}�Kc����}M)K^\RZ��׻`�2�d6�L�V�*!
�Qx��X1<6R�^G���p`����E�}��܏s$����<����(R#�ڔmn����b�����8$,�	���۠��Ip!H���Ig�J��uR��ASqT�X��	>�o��a(�\/�~����R��⬢?^͹�����j4��f�����%e�Y�qfT&��)Sp ��H_|.B��B�@������Dg��V��Io�1�*?��I�Fa�W���7<
��%�h��co�O)�*W�L��B^��WQ�/�.K�nA�����f\,&��h�ű?�ήF�껓��� �z�TpW?:g;��p�p�<~�7���OH��3������[sa?1E2.������]*��ZՓn�m��)v�t�J�Z�cd�08��I�=�&y�
A�~�����p��ub ��� �9�E)�iQl�g� #ar�"���1iKf�ѼLE���K�T
n�kQu޽�5�p���,��0Ȝr�0���:���6�p��s�6����K�J/%�D�sN�{p#2w���b��I<;ܸ�,�!v��� ���)��$Y�]��� ���RT{:M��䃤�����\�mbRZ L�lR���1$�|t,;sмR�n�P���x�]�@9��P�?"j�C-Pq���{��LH:��N\�%���3��oB�)ѩ�]ev"�%�0>�+F/�܃����P�n�J.���H������H�Ӓޗ�{	zܱ���@�8���Y��)��&ɣ$�9���	��i�tv��_���(�8��Ua� :�I~�C����b;��1�h�Q!u�u��t���m��ٺW�]0Q�Tν���T�(���2t��}�:���PѪ��f��*��:�o�BlD8��+@�rf�;�5��w} %c�'����n��� �@�:O����P���I��Q�-�S[I�Ǐ�cM�y.��V;����6�@�ƪ�T++P%:G��Zd���H�O��S�Aޢ�w_���i ��x- z�Ӧ����X/N[Jݨ%P���0�܊����|��~��������6R�A?��F���u�K*��â�G��WHbLW"�3���;g0$�٥~���/�Zs�G�D�r�C�p毹�zMqЧ����#�Vo�:c>���u1s�2��z0�ϹɓB���R7$H=�n�v���Ѿ�@ zև�2s3�N}�]�',&A77}ҍ���~�f����>�~e����#����cR<HyX�X=#��f�u҂���TQ�C�I�u���U}�iϕ�h^��R6�sNNF�)��>��?�1B�P�m���_n�����1,ѷ�.�̉f��7ӓ�E�c�څ>��Co{V�)qľUP�}rAl]ֵ ��r�8���s3��9��7�� �U2Ű����=�U?K��T$1<6c��s����#68���O�kJ�=���� MB"�G�ԡ����|x@�����w����	��՝�De�N��=�&�e�a�+9&�o�T3��p�"��b1�*������ڠ�ԫ�w���ϞY����k��Ũ#@+�DC�Y7��䢅%��#z�{�djK���6�a�܃��`����u�ˊ�����-���|h�F���0o?v28�<ՓYO�Lq̾yYJ�����HHH�&��C '5R.V:�;�����E�n�"�/�����3;?��wc����pHa��d>��$�o���h:��H���Ƕ7�����ƶ��m۶m۶�7�ض�yg�o�������}�s�O�;�.��42gD���.K*YSJJ�q-��Ł+��>��1�Q��_�6z���2:H�.���J�|@��FӤ%�9�x�ه��w^��h/&�.C)O��vo
I�d����0��4A,����ex�jd���M�Z��M�Y��:��r"f}:�$3�'n�d��姄�����\��fzN���t�B!e!!5d��ş�ծ`��&?��F�8.���b��)��_v�޼0�*� l��n�S�	��Q��=����=�mȀ�um��ϒ���5u��!�Iȝ5����:0��mEjS�K�3��������?b�q�𤗢�閬�������z#3^;r?bM2�32�\����!�<�퐜�J�p��/��l)K-���MBVG�
5�
UhȽw�!dA�PvMю-�:�x������SM0�G~_%�c@&�EA:��1b��	�?��9��g��Q�ZSh��x���H| l��w�N -n�(��f���ɓp�����r�:���if,и��C�.��z��L5���;ʫ.��Q�>(�+Ƹԁ׃����ꚾ"l���r�%¶��
�h}�oh��g��{�w�:\}�����L`G-9V�"y��� ���s_��1��+�h�t'����ަ9���Bk��iNK�|�+iL��	���Zw5#��Y�+�q͚dk�oz�ѓ�u��y��x���h�}E<Yť
��Dĸwv�DY߫N��E���FN�.<V�×n�+=��j��S�O�ȤؗD4!�����}V��0O�.��4d	�s�H2X��N�\Z��u�x��2�7�*9Y9r����=����t���t�&uR%��5{x�i�Q�"F���V�zK�f0-|<z�n��Є�';������>H����>��)���êm	�</^��kc��6��F<�y���瓓��jX-.��т��n��x�n��4�N;�A���� �E��L$�E�4C�2M����"�e���d4��\�\��,;l$)���<��Ź��Ȑ�@�Xx��gA:m�'Q�&1��NTh@g�X��I��VMT�[]�_J��c�:O�{�:�����[��8eݑ.:3�6����lpi�\�<���d��1�i�l�����\!E��n*Pt!�=��.8н�x@	�����5�����������j��8P@F����׭
@�b�=쟿fι�-=��ň�4Qչ�����������Da�)���h��h&֬�����MQXi���.<�+���*��u��LѨ�I?���c���g2�	��7];#p�ۆ?I6�;�%k����7��� �ŭψ���!ij������k�yM�̐�x��� �e���j� �)"�Ϟq�v��=:6��[o��M	�L��e/���ʎ0�����=��\��_8��9���a�U��3� U�l6CT�=M�=����� �S��@�����R�b�j����\m�^�o��֭Dgn<c�`2}��H�p!(0� ����AΠ���s�m��WS�`P��� gl!Itxu�5�x�s���ꊮ�O�u\Ӓ�\��N���z�ӱz_�����g�qo��"��ް�����8+I Z�R�
����Vy�j@?2^(� J�x@��6o��N�N��1aG���D��0OR>�n�TL&C���)�JS��h"j�(~�m����q&b"n5��P��Օ�v��q[��gش�yAL��"��4�;�ڼ'�o�s���e��j���MӗVxh����E����đ�Ď	@�.5�=]m-.]g1�+�:��5��(�cȻ�?���Hg�@�ɻ�1Ka�?[,�☀� |�Pv�ױ��/�,O4۬�\,��}���/t��L���'�{�1������m'�Hz3�j�\��Ib�dO�e FK��8�zK�bA�Io�C��TÛ��ȍ��8�"��h�^=��v�F��#~�!x�jLlİO�Z��5֌{�c�۟�s3�ĥCH����\y�5���>��;=��4����i��W���#U�
�\d��E&�&�3�2�9�w�Y$Oh����f�Y���P���/2kC��1�m<TG�w�;�-�:��`q���3η7s���+�S`��i�EƁ�6vn&)�n�o5B�����J�����#�f9��u���p,+ ��ԠyVz�^ax������c����=���V[>>>��?e����
�k+b��2$� q��tec�NK$.)qՍrHP;��^x�8�z+��۹��Iձ��}��3��=������A0�:qR�/W$zlB��5MC��ôr!�y!�_*�)`ù�D�0F�,����G��,sဗ��\�E�ff¤B!x^�@K��h4���S�E�`�S�w2�JW���|���q���v�QI��K&=�K��T���T�fή(���b������P�Wf�� p��HⲖm�M]�7��'A������s�.+��#�{�g6�:��4�Omڃ;5Zm��ld�E�v��g�������Uj�v�&/I!���e,uYˬ��w��W�V���G��)����%�p�"ę+�{=�{D��f�0�u�@���J����3�T:G���ٸ�[�
G*.N(�F� �H���V������0Hx,V�v#�.�ja+�{�،�yV�����&��$�ys�@"����%"}�����0#SBp�lpf�M��f~�n�١9����5��r���evy����쥒�a:���.7�%]8"��Shl�\2�Iz}6�v޼�A#��%uk1C�g�l���N?1��khݐ��0�����jC��CY��'̿@����ʬ�P���t_�l���h ��y�����#Y�!��+�q�cGt��8>���f>TL�NT��&jtL3����<�m����5�T����n#��(���o�JsKF�++a�e�"�3.և|,�U
���u�}�Ɂ� �nUN��y;zC�/L	��J�s�����M.~m��x��9QB+.ݏo�'�s����%��+��P�TXQ��r�x�9LV��F�]뚉�����$,6I!�ً}�:����9��,X@uY@RDU5���GK¡}�-B����є:���T��G%D>�*�7�	�j��o�u&P��)���O�6Kz��%��c���s�zZ�K+iP������� UV��E�ȗ}fy>�v�7��<�����"�Q�����dyp��
���p���Óo񪞹��f��8}���'9�c��ǉ�0�v>b�\r?f!	��뷹����Xqo?�Y���<p�S�6�)M�~��p�y�.A(VV
��X�f�+5��#�����n�qa�/L�dqBB������������D�� RĤ��9��tzr�y�J���B@U�A����DU�3�k��Q�!, �t�{�� %兀]��R"BL1��IU|aH��ϰb�z�ThT1���@���G�S ��k�!�P���$c}�Q�B�r.<�q����|ϲ�Gf2�GA��0����p���䊢dU.M�6��9i��$A��c����d��8�	�RIǝl
��Z��]BΓxmA�@n��&�8Ӹ����w}=�B�,|ԭ�+���|&��'���>���GijQuu�X��t�P�h 5�M�����-qؗ�j(���?�������w[�q��"�uI�՞��ƑL�L&1`��1�%Q�Hk\+1F`�s�E�ۍO9��XQ��:��㛁�)b�F��Z�����{]���:�'}{�Ht�Y�م�� �%U���A��C����b�~�ޚ��`j�#��n�b�'M�ĖC���Z��>6a����#|C���Ȕ����=�N���W�'��m�v�,6���-�*�����t&?2�Nuhs�F^ʄj:��n��hٍ=���@J��DJ������
���<��D�N;� ��T��������@=��)�SE�������^��%x��4�:SP���5���5�?�	���4�ْe���4��Ua*����\����rʄ��S�,B",Sj*-җ x�H����O���>�Bs��e�AF �҈#˟J\�t��k�WSǹ���?�#`�]�Ֆ������mjᲞ�ׂc5zë�{��&Sh�:}LՍ<�3�����0��Q��"�JF*~,IR�+�U�?�D�3٬V5NĽת�N�j���ja�`{&h�k�.��^=�O���MdmZ�,p*�=vPf:�5�-�34�w�y��-\g�U�gU���H����r%؛i 3 6�=�?n\�������|�*���;�!@�j~��Ö���f�������&��7?�lw��z�C����,�Hg�����}��$l12D	,BJ(� ��� �	wsfՉ��U�j0�b/}�	3J��������rnS��*��ᠸ�\�9��0�O�3���$Q��i{��޴�h�~��$�ȣS�t��hǼ͆��_t;ӱf[��f5�����2��Ӆ�a�(RiQ B��sԚ���d����k�ƂD�7U�rUz%͊�b��4�=Z�m�5�����vGh��ynߛ6R�����: ������vs��]�!E�����X!�*[�)�~�xk-������V��
[ZVG���lh�تEZV.Hyf�b�jtQ	��2�N�1TC&�sqr'�Ė�'�<��αtbY����_��m.5�@,�^d������W�E�p�1���/�n�sg�vBQ������a���1��줫+���yͣm�Y�m�4z�s�Qcƈ�"EA�J�v��uU��ǮK"���sQ������u�N�8
����2�t.�R-�'��;�Yr}U��Z>�y�\%m��!���}W(ʮڬ�����FN}�?+�w���u����C�I!ǸH�e���P���P�'G\���T��0�F¨F��
�9�����8�S$/��7APc�PϢW�7z�iR2=��a�a���s�P�$����@貓V��A~���	�7�]W.�/�_/�V�m_�@m���ߞw��q#S`����u�0n�n�a�u��m��R�l)�*��P���f0��N��)��_�D���>��îa����?���>qlؘ�Wg����On4j>��mQ�z��8�N`�?Ὗ��z��(���<8y�v#�V�_$V�~6ϭDkc�ɰ1�3�隵z��Bj�@��:.~3��/#J0���Nm��gAB�I�<�g�>;�z�YvY��Pk���R;8�2�2��*�F{i�K�x��] & )R�[�˯.<\�B]3��r�-����x�CE1ǿ�\=���GnqDl���e��2�8��<ޤ���a���� ��= �(l�����p���e����7��6��iՈ�m��o4^%y'���	2�?���y�S4@���1 #�7�,�_/|򸼰\�W�*=4|9(���*��*�t�3�)Z��מ�����mR�l%@��G��\ؑ�6Ȱ�󿄞�VO%�U�N�ݹ�A�:V|71bL~��,ۚG�h���-�	d�
i�M�T�`�]A���RM�TW�H*]��c��z"�.��s���)�s�HSq�k��P�0�ԝ�d���L�p#��4cκo�ȭ)u
LN�Ʈ�_����}w�È���������(D�8�rx��#O�v���>�p\�VVU�;��B9;�䡦Ģv��#�n�*���tJ�c
I֐�x4{�
��� Rc:1n�u�Pƀ<U�K��>�Nl(�r�1dIKN���ט��i�R7_��Z� �X[�UD�wz��g�e�型��A<t kMKC��=�X��gny�&8�E�@��6a�P�c�Ջ�n�`�F+��l+�s-�^~&+�K�y���Yo����J6ڪH˙�!é9!+��
�^��,�N#��ڏ�/�O���R١�㼸5�e��A�oc8n+�,(�;�.��!�@�`0��!a��Q��l�i�C���3gcB /�z|$����Ɖ�0�~�l����z	�L;�1�@�v�V���GB,���P5T���W�Jƙ��2J�I�B�m�!�V�;n�XEդ�s>ԔA�}�o����9gFiPK���k͒
�C�0Z���+F��^L���M�:���B�jd�t 6��$����\ֶR���|g�&^����-i�"���$A}�����W۾'c��Y=�Zڠ���ҒGTM�b|Gr�;������'2K�`���Z���;���gm-ÿٲБ��H%�Kq�	���徎���(
LT23k�
�����@l�^�}��FWk�*]�p,9��2�<�c��d���V=(�V0��=7��	yn���!F{s���WSn�@U���L�Y9}�
=��3F"��\[gg��X�`"�\	�����4�P�,IxX�^���2�ȌЖJ��ݭ���Y�M�ӖW�O�H�/hGk�H��M���<P ��؄ᆼ���$�>�ayg��&ҙ����g�^hi�X� _%1nT��C0Xp:�-���2���֧l�s۶�����;a�CWWgnuy<�YI���j�Կ���gm�ńM����i6o�??��9r�Q�\��D�6�FAVa|.�������<��׍�G������:�g��0�s��v�5nZ�a�{-����]U��)p[�r�ϗ��o��=���dsN� ��� LD��H[�`��1�����l(��X��k?�C�Ի�f;�撅�>Ep\�H�/>e��xJ��VD'%�ӑ�Au�I^��R��b_[SzY�k��
߆y��)�}Me%:��[���ѥ	�H�����E�1�va��iĳC���p6�?;�+zv���*�G���v�U��jf"`
H��8;6٪��6���Bm��qs����W<�?7�;������u���J��ڏ�����z�~?�)T�^9XP'�Z���1��>���� �9pE����@&9��a���)���
��%��$�X3���*mʠ�ļ�/@��פ��R-޿���)ux�a:�}sss�4k�b���ςE��=��X���+��/x�����OY�$�%�?㮑	0h9sDZ���P5���(&̫}e}��~���1�r\�".���j�c��_;E�w�}mJ���D�`�K�![c�,L^O�,���D_OM���ceec���0�UX��0H)R�"�9��Y�N�#�%���*w�YED&kIR����O�S�=Y�K�}���d��wS��|cs�"����G��W����DW�N�)��r��|��WS���w��\����Ꜵ�xُsc�+�u땃R��LQ�T���7�zW��v����ȏ���V���5FG>t�D�т|��OJ4��Qu=1�q��S%K���A�)e��>)�/J�Z E�0�(mz�U�(We��l�������Ȍ.�k�=w\O:���E��4U����NSs[�o��!��� t�V� ���8᥮�KPzaˢ�&���G6� �� 
U��/��C�S/����a
�Q%>b�+\[���� i��a6p�2��|�d	s�Ǚ
�)!���+�ԡ�ﳱ!n��֠����c�-\o�����{��0]�_�h�e���}��(�Ϸ��w�w�+�tkT7��x&P#��ֈc��E2�����w�s������ÌY'|=�$a�a�-;�%��(��!����X��!4��[��B*59-r�j�_�6���X�5�ٞ{�Ȧ��1���:��*�^cr8��oӤ�7��&znޝ�H
Hĸ�tXU�5�IC#�0��I^N�{?}�[�}���μNxM�9������~��ds6��~G)�a�,3KJ�ݽ��ڎb®<��P	�V�&Ao���A��۟�1d���C@@0~|��r���-~����'�X�&�م�b	-�x~~Ms�ѱ�c��ٹ���
EQ�"6��`�O�/�"R.���%A�%�`��Kո�P�#�)�,��}}�Mᶊn*�(�"��I2Q[&f�G)�ğ
��Ο�)���Rd��~��!��p�$C���Zl�Ù�s�T&#0�������������2�II����&j�0'�J�rK�)-^6&,��������X�j����@	p��).����M�r�$Q�=�6օ�H�|s�Lk�)p��u��4�Ͷ���
�Ay�HH��]�EU��D?��l��!��v�r�e�RݶBp��^w=��1tQ���؉	�R���v�9Ze�N�{{��׮���oZ���X[9��
�b�,?X�@���P�[Xb�(�U�*&)�|�?nެ�)h/��z��z�0��0�Ό���m��%H�
۟�_��bPp�-{mS�b,�o��� ؑ=��]��z�S�I)��O$������ˀ`ڱ�6�+U`�fc��c�.q�M�Z��t]A����9+��N'F��e��M��@�_����"�`4g��Z92n�7����EV�&*��S�5�x+Ú �����&��7u�\/I�eMD���q�vz�b.��|L����Ky�pgY;���3_4
K3�!�
y��מ�s��Ht�� K���D\w���i�1	g2����tf�Ih4'�0cq��u���i��i��R,�o�|&�?�(�����Sg���bI��-��tF�1��,�����<w���!��1�Y�{�D��7@ l¯>�4�e_�J8ٕ�ВLվ�!xn`�k4��[^^^��ߊ��V��L
,9�A��U0N���`�1�pW�����Š� `�w��XM��n2E��V1�|���q�M�S���9���r����CF�$qȗsKm=���ߞ�詀r��~є�<����Q۸���m�.��]c�E�w��@�����(�ǌ.G2?��/��O��% U�
���_��RV Ʈy�p7m���Ǻt�0���l��ԈŠ�\��Ν�)�����HwN�_�d�sK)�aɂ�&P�N�V^qش���yϋbs��T��I���'�q��Q��S@B�-K�(h�뢠D�Sƻ,�S���!v�Jӯ�J&Q�7[��:�pݴ�����U����~;T���r��E>��G<�.ء-ֱ�kȲ(o�S?�0p�f�IV�dΰ~{"����<jS��\�L#�5;�M��2���`5�����⑫E��V��ks[1��An��w��8�3-v%��V���R��.�j,=X��w�����;�T�
�Slx��O��7>VաXz��>+��:���o��Σ?���s��X��>��$������O�=d$�p�>ɐ/�؃�D��K@Ǵ����s��3�y%��m!�� �D-�Jo�J��X�e��i� ���I����.;���t����M�N�ЙЛQѺ�|:u� ~���KMklq���ȋ���J�"��� �2���~o�e�*��WO���(~#���4#��V:`+/ ��, �n|BsȌ!�j#��گF���~����8�A��L�/����@�*N��_h�@�Yfr���a���>��9B������Y������*$ӆX�ϫ�I�->��I�[�)�ńP�8��,��^��P�Ǽߩ{������/밻�����\����`�
`"k�݀%CuW��f��[B�Y�:������g���2���ͮs���Ko?<OOO�
;fN[�]�
A���:����9oO�bL�n2!J(N{F^�|"8F�?�#�^<����=~ݳ?q:�t�A�4
�qݥ��˴��S!����2+;�X�ʀT;��t�$�'��>k\�,G%����;)A��]�<�L�ܰb�W6�mylU����t{�ۏ~3ӟJ��J�
��|t��^ ��ݻ�A���8eS_�Y]Tk����,d{2�6S�j�Cv��/ ��=$,��I�!5ߊ[)��iN��:�)U���g(f��_�5R�)g�ky�vT��Ը�۪��2��}��	���-@�a/J�WbD���sB����gw[Q	m<-f�	܈�!c��(�K)���3���߶oR�8R��ě��@�A������˘߇��`)��j��'}8eR��~d���f��a��k���C���rH:U�2�I*֣�a¶F%�4/2I�=F6�9���]����N�OKʧ��&�a"N��]�R���Æ�,������ey>���(�s�|�΢K�
�"��'�m[�����<
�}E�T�C��0.x�r�.@�^k4qZ3k�?�X�E����P��D�9�=N��̰��<��*wN9	PcIC���M��WPA#bUQM�����LD�%մI3� �J�Ȑ�0�}6	�\�W
�&��iF?�VUE�_dE�u�$""���D���T�N�mjP|����;�,v/��A��n�s2��j�ތ ���.�X#������X_ݦgo���eS���D	��� qqN�F�!a�c�D��9Q2�3�,<�]-��# oV�כ+�}�z�w3��c
� ����~��,ZB�$w���� 곉=W�=AQ��
�D�b0J�~ �(�:H	�)±,�-���Cq�B�:��'�U�����3�ުT@�YT�j�^Ѳ��@�k,�}���c��h!\�����R+�O}�s�0�W����vĕ�Ƌ�*ӡ!�ܦ
{�x[N.�c�uD	������4���X0ʧ��}'0�*�3���T�b�wSɤ��Q^�{������~r�jP�'���l){�E�d4x"���!��~�ު�h���+��blZ���Q���fks$�jP�N��7�up/���p����zs�q��8Ǎ�t����ZW-I�&E��d�ߊ�Ø/v�h2ݍm��f�'ȓ=�	�쾴ޛҔ�`����W@+wlf�0��x(��<O	�N�C���+O�y�+�W��Zc%��'����(�`e��$��y�	��ݳڤ(�H�Asg~�����rz��ok,z�a��zL����e�yP��b�!dK�����E�F��K�,F�1J��x�H��8N�{�Ϧ�k7��	��P"	ݪP�߀N	O�Xlэ;!i���R�M*{"�_�h� �VU�a�c;#c�o���a5w�6g�g����p��d].�'�q��U=��n=m�*�J��IO���p�#�/��iN����1:��=CU�i��¬�K��$��A����ygl��Wϩr�Ade��@i:���|�7VZ�[��h0�\qqq�Dt/&V�N(ٕQ�?LT��m��*L�+U{� �$�� .,��J�+����G� 1Z�֢U]�6N�J����@�z�T�]hĳ�b	���S�7�q�"�Z�6l�F$2^��v�6�N���BL�BBB������/옑�5Yx��c�DGkq>w7�ř�p'�Bu� ,����iQS���u[۷���9s�<<X��P�<O���1�@�'�$.�N�I�D�D��A&\��!�/��o��
ʒFR>�D��}�0�]����-������_
�Q���Y�sH���0�8��DΣ�,h�j����Op��HIer�y�
K���M���qp�9�s��ڌ��`��~�D	/��C�N�hаgJ19#�u�IrĚ�F��_�4)r���>��!̼5���0�3�����=��/GZs�=pɊ��DY�� D�MK���%p��Qf�~�t��[^���`�i-g�#�6�	c�D2�D2'�X�bC4�bOR�D��c��tf���?�Xi�D�'m9`��߼��|ŏ2�����zK���P��X�{\Rf�;M]��(8W����8�̸��^��ⲃ%o��c�FUʤ���%g��=/�>B�q��>K��~�i$¹��(?�e���J~���tF��0��"�a�h�d��Q�99���m�ȸ�\Ʋ�"�������dk�m�&^��^�p[P�d)�n/?�.�����6��l����cI&<�}��*������ꛭ]AIn�>��������"�B�YE��S�_��./F�-m�g D�*#�%��f���8e66`F��ͺڹ�ѣWָz�N�&?����IĤ_��!������Sa�A��a�9�����8s���u9�_�s�/�����fO�M�߄j&��7�c��c����8���	O��>?����)d3��]�I��LQ��#؀��Wk�%!>'�e.	�QY5HpH����F�@��T����7���q�����f��%߹�7n{�c� ,0�ʢA�� Kt!h�5�ݵY�A�q���Kڰ����|^��}��r�J���������H��D��b�����\"Dn�_��cpv�DI2����4�i����8��pݙ�>���*2�Jj3�|	��d���;�F�Q�>v=�q��H~s/�PG�0t�f.�Qd>����*��`if�RXz:O�寣y��8=׎���Uu&㉗!˧bB��*\n�Dl]+D�3(��TW���n��8J�բ+�I���0P	����w��vV3X:�,m�"d���8��Ij����8s�����e�	�ɃR�{���&����l�7d����@� Ud
�f��Y!�B);g�
��|�fV*���/A��f2��z1Hn�A�	�wG1�f[$؂A0C��t���9&��l���؅k�k`��p�EQ��~�5��X7l1"$=��R5�i������xA��W�i;���ˉR*�@B-1|ĸ	;{f��;t���B�t���ӪQ�'v�0��~�k�J�8��%)�E�f��i���71
�s�������@(Uq�OA���}���!B�x��S�E�z�r��j	��3��UT�k|�.&��M��S����y�6���i;���e�����j�TYIU��TZ?k���G�����)���Nc�i�d7��;�"�ӥ]��AS�@-Y�d�����J�)ǽ^�Dfذ�=5����>�o��y��bFNG�)�[�:�����G�0%��ϣ�pA�]�H��S2H�����(�ҥ��Z�V�j�N���MC@T
s�8i� ���l�]aUY�7�)��t(g�)RV�Ѥ����p����I��?��r�$� G�K�_ ���%ȵp�j����f�YM�,g�Pen��o���͡@ۺ��MheU���j7���6Ř�	����&:�~ߦ��wV��w��
~���ph56�M����S<�	=���T�.�WR��@�j���F�E�[��<��x�v����j�R�O�3A�k� R�a�G���wϨ���[o�������;ҢJ+�:t��&�gt� 4a�x�z��b�ʭ��0t I�i۲�f���!�&б����"��>{������n�E�~ʅV��P��$��8;�]��CC�㍫�e��8L� C�<	��;��Bz�b[�9�P��Ů�[\�U��R�3�^<��am��M^��t�� �l��!β����Bە��X����Q4�'��f�yr+C7k�>c@e�6�B���s7]{Œ��+���G�AW�I�۟6����Xܧw�ʸ����a�3��F���Ukw�31�}8><>�X�Zh��eG�6ӑ&���yZ@�P�,a� ��Ȕ1��A�]�ZG�M=��i~3o��?��B���AȎ�9��O��>�ԓ����;�5sksiN�ԥA��[�Y5.dp2t���G&9���j;+M�r���Y��K���]ͰN���!\���0��!k��\�>�vi��e��3QZF�D���!^T���i��|"<b)(�����jhG�K�%h�����:���p^6/�{��=<BvԈ�{F��W��H��@f���@�G ôvOzf�ɛ�?�h/����U��� p��Cu �s��.�Z{���� @��r~>MP�EO1t!$H����i'�n2�SE&��Pa)�c�f?�z�У�<��{���ַ;m۝�z@J�O��F��	N���lb�G�� �z~��᫙?�i�Ӎ�����ߐ�]�	�I"��}#l�#{4O���@	��,sX�܁Zd�h3|`Ȟ\�t�T%Ӻ�� J�j����D��f�o����
�����ͱ5�sҬ	�����s�����}�ɛ�B<�{��l-99�_~�����l3���E��י&��1r@�AK�iflO�s��qmjn�;o쿆!I��#]��ޕ�2:k��V��.�N�a�:����U�JHxN)�RC�`���|j�ka�fDx�^��\�3���f��?���ǽ1����GxV|��>v��yS�~Ќ��!���X�Q��1$�UO���03�xn+��[j���&_?���.G���T�3���h	1V�]�~ٕ�1�T.D�[��rG�ʭ@A�B;�.k8y�W=���	���s��b��v�3�9ش&~j�����U^��t�3�@��p���N�5��Z�	�I��.d4�[����i�TX���Aq�!W� �+f����u*T�Wm�k�:I�v=����Q�*Z)2 ��;��[�REe0y�%�KK�s�$v�E��N�ei �eO5���t9�
`�f�V�g��n���9����\L�)��h��?K	�Ci���IO!�O#3�C5Z,U� uɛb[P�%��Ba_�	i�C��x<8Jppq�׮��|ي�J���~���Ͷ��_iSÀ��8�(W�AJ0EQtA�g�C:��n����
��(*x�����?�;�)���QG{d;�~�<�n:���#=o\)�Ti82�؁�@���n�
%Ȑ&��$��4�4��ܬw���26І_�^��~���=^�@E��4�p5���9A��z;�p����,ҍ��S什+`%+�d���`Ww������`p�d���/�߀�!E�LM	24���P�!���џ� A��c�d�ő=t�s:����\Cj�m|A�Á�'J��cq����>�F�z_^�o_�W2�>Z���w<~'Vo���=���T��w9���ʴ������w��DQ	Wg��5� �޵T��d����gL��b�Ђ l{�wׇ�R��k� ���b�W���3���p"����ug}]�P����Pw,����(�����48,Î�,J��ѹ(�Q����l����o� ���<OU\~��ϊ����%����� ����D��&�f�m�X_�t];B��W�Κ2��+x��"8����?_��n���+.w����VL\�;��ۧ�#���&g����Ѯ%����3=�h�@����G�Eߗ�Ԡ7.�hq%�C�F����;�� ��9�w��m�zP��{$24XJ1�OF�:������͗�c�����6g���H�k��=����Җ��b(HE���%"*Q7�&�Em� #��b��Kp=qK�h"Q��;ȋ��( F�iL�?� �[�wu�ѪU�!M|ڽK�z��T�~I�q�Z���nd&�(m�X�*_��P�BEk����ű��2���mE{q��������\/�'�kJܓe��u�>:�9���n�TE5�m�(e�� v*�V&�pt���pm.c`�?�9�V��K�����}��{�h�(H��� L�U�F��z{�R��܊�\��hH[tN�7� �B�3�5��$���!1Q�-4�̒���L>o���h��͇�	?Y�e�zc>??0�y������K�����7��-z�Dm��$j�dC̑�N��ffu�����S����H�b$2_�6C�� ]?��d�p"b�x���߯P<�����;^�~m��E麝崯`
�����'��������I�[�a�_�K�=�3yO��{J\�;�w��v���A(�]�-y����~�j)7W����31@K\�' �L)m��R��Se�Pn��b��xq�����ﰚ��������<a:h�<���N��&僱'�L#����fb�yXH�D^O�,ix��ӿd��xOG�@A=]�����̕Ec��lY!ɐ���:g�J���l7��JKh[����x��� ���W�!M�X�~I�r}�����"���70?p^w��Z~�-V?�=��۩�����G�V��0�X�Ą
��3X��au ��R(ծi7�x�(ɘ�����|;O��o�����r�Q�w:oU�d�w�V���\?>��[(��SY���#����e�I�r<C�0�;�K�rq\�/NO2٬�_��K#CH\m7Cտ^H�e�,z=�[U1���h[{� �[fZ�Y#�|.�8����d2=�ݪr��r�س �����w�����6��y(�NTީ�bv�r�n�.�q"M�Y�ԎTk6���HAv�]�����o<*�)EKǬ� ���s�.�,C����g ����N��%�$��{��,���my[�]��c0�E�n"C!#57����B*����42ٜ�G�~a?Yevl\�R&�~j��S��T¼�$�!�}Q^{��8����dC�mӅ�~�E<$�iom�/����f�ZPw���t�Amu[4�������ݵ�S�	�n��Z\Zܵ/Ŋw.�o�e�a�'s�>���֖s�m/�뷺{�"���B}�p��R���Ԅ���02lw�V�ؠ��Ο���#���>��W-Z�8��uz�ؖ5{<y�[�G���M[m����~��|�QH�]~{	[���@so bt]�|s����Ԫ�K.�9������9�A��7]�����>u��{f?���U�9Ý���Қ��M��YkW���̛Au���7�Dk��?��=�l%���������7���pUr����59d��(�"C��MDk�/���j���(��s�̟1�6���u��g�(�-:k�6y]�o'���[���b3�m0!#��l�W�C�-����XY����=���BG��_Ř�@g�R,��k�4�6)����K�R㜺8�~��-�$}8˭�m����w݌����L��F]S@%˞c>�?�˄x��CD.�Ŵ"���)�0�58��<u�m�U��:aMs3�j��_�#!��|8=8���m���u�@z؀)7��3+�9S��.䧭*^E~$�_��A
�2c|��(n\���1�&h��(��*��"8u6ŕ���z�p LBV����cB	&���[Bg��B5�Sr\7���Wz�Of��L�	K�AH�+ߗ��(@��mfU�`�w��.��|�G��,�n~�:�K�݌��3�����is� ߻�h�I�~�i���'�<�PoȒk���9\A�kgT��M��ׇ0c��dÄ�j�,�]��8��-�<�-����b6mX��'|_��<$�Jua+!l��ei�����P�þ��֡S�Y3����~���DlXhT��s
�:([Ue'L�LS�C�ǒ7rKĬhS�-�/��������/o��K$dDe�L�8@�p�.Y�e�]y�Z�nR$L��,Hh,�����>d7�_JM#i*���.J�m��ʣ����+]ƕ�X	��H�C͹�����P�s!��e?�n�(g�F��V��m�m_��e�u
Ow�:c��t�{H'R���u���Ѕ�ܛx>�l��	q�3
nH=r9���6��w�*~�� m|��K��j3���Z�4�r�<��S�o���4b�u|�����e"XF���}ՠ��<��;����w1C��}U|w��F��k�/���;2,��;p���#�o�80ԁHyx��=�
����<�S�Ja�,���	U����M�<��O��Ơͨ2��C�ܪ���`��D���]ލP�9Y*ItX�b>�o,�����QYŴ�������
�\n'tt�n䰊C5_;m�V�ZD�ƭ�N������-P�'���W��zV`��_|���������I��<�A��#�%�1���מfo�8���V[&�e	�m����]��xd'���G��;�s�E�y'��?2�t���=���پ$U��ǼѤd�3{dk��4�5-2�]��57	�#�В�*���67=3�&~����h��o�g��"��Qߵ(hH+~�a,+J�v\�<������-$$�e���E9ָ�&>�N��R^^R�����W0mIS=b�՛&��8�B�W�,�Q-8�5HѸ`b`$%�1%�%8��Kپ䨳*H<��^OV���RRdh���� &��U�K]�x�gg�'~���m9�\���kL���[m��h�0f�:⭅[q���^p}a�O��D�¨U�l�^���a/�2ɿh����'UB-?���?f��Ӛ��f�w���/Rdd�'m�QF* �o#�Y9��m[�dw�Ef�����)�o��(�S��.'��7����ѣ�5f|`2�.��JF: ]����O�[������H��0i+'x':�0� Q�Mza�w�"@��Q��=�a�Đ���6��ax}�"K���Q7@�4i+��N�6�O�yP<1��^,{p�}�߿����1��E��s��+U/���6�va9�	ԋn>��c\0�;KJ�n�ќ,7�E��h�����.��X40(�sDU4ƀs�p�^_�9b�bЇ���h�U�Y�
:��ꓟ�̅M��b�,�B�!\����vJJ�6����:!�g�s���iY}__����~�)�2�R��
�!�Ah��J���p
��J��ñ�~Xk�3�V��B�h�}(����������L����8QΖ2% I��	��e7!<�2l��X[�g]�)���?�܇��7粮fTjB~�S9z1�r�#�H�O�:e��G�>s�7g�G'3������f�[�o�8aX��d�!6�d�4*��\����4�j�%��%QzH�x�^B&�]�C��	�H�x�lΌ��MLL�6��$���z`6"�w<w ~����t��!�,ZN�VɆ��$b6��y���D��o�r��k��ۓ�c��q�WS�T�>��\ڷo@1F�y�K�WF�K���έ���S>���wݯm�(�b�#�O��{��1e��y~��*D<�����V�.��J�o��?�(vK�-\X�4g��˼x�O
5:l��f��U{����ԣ��Ê��4 a����>A�ݤ��l6�ti[{�C/R��3���>E�~@���Z�n� �_r�q"�E/�+净�2�&�zfx�S���a�	��̥Ƥ���m[^�q6'�:����t�����K�N�S.���׊�K�SK=6���4�
�*����jP��;�P�����-Y�u3U���!yK�!�+�����`�f��E�kY�s����ZЋj��oK�p��S�e�ۡ��+h=����j��o����A��{��2��[NA�w$���Q��,�-]Ob��s��#VE��Zt�&-���՟�f;cc+Q(�9��� z�Jӱ<�yU7�3z;W�V��H�I���ls-�!�pz��������"�,J��7g�񡇓ݥ�FO!MG?�;%����
��=S��P��]�/f��:��?C�?�h���φG���Y���B��6!>XpO�"���t�_Qa%�r�~��r��r"��.��i|���w�Jzxz ���{��ՌO��]�kiz�9J���e��r*�z�愑Rx�H���v{C0�igSe�p��:�N划�(�m4fۜ��N�7&������7@� �d�����dD"
�~�]mOg�\�[Cѡ�3�8i�;\8���ͅ�%Y2���\W���Vn��/z����y���TK�T��z7��0b�����w��Y��N�����__��e*%},�
x�u#��e��y@��%Ã��P�$Z�!?m�e��z��/?��.��.]�<���2���`�;f[��(1)�C����wc��GKZ[��M|Hj����G}����ѷ`�+����my����_����d�`���f��V!��p��=q�)%WQ��]\�u�������; R��9��]x�?���,	�'vHk�8���)�R�?ͣ+���Y������I]��+e��؟��iI��7��ȰPxT����&�G@�o/1�`c&H ]�M� ��9)��})|Y:���uNt8��:ǟ���!>��D�GG���� �G����]?t��u�^��6'n_�0׾�מ۞���އ��mz���(�$X���fFP�f�rߏj��ԁ�D�\�/��^����ѷ��;jy���-Ö�Ig��A2_��o|E<��o�G��6��D����v�Z���V0:��h��5v&h�IS�$u��2\�P��hȈ��huV$�ݲ�V��n����#�/��3�d��|3�R$�|�R=0���R���X���Iڐ\=�;L��Ң �53��|Nm��|>dT������F����=�7�Pz��~e|��/�B�[,�x����p�68�?s$<�Q|>�g�3v�k�&E�zj�7B	�D�(�R.�{���߂�)�[\�kW���	9DQR��h�-��Yso�}d��!�ΥI�Z�g���mRs�Y��z|t�N��*M Jq��n�2G�$ne#ty�n�鰼w��I���q�����t1�۹���("��b���ye���m����v�&��]�xS�TY�_Uk�����\o ���u�:��*
NB�7��)L�^�Y�?]��<fF*����Ŝ�qX��Wg��`��ϩ���QTuK^���CE%v�~�H��|C4mՅ�b����h�Iº�S�M��d0�	�6�`�3_|�7�`���7n`�Wz�I06�����4�	��lȊC�9��v5�t��z�|`B!���5qå�]�<��jo��p0�3����?o�s��V�����z����K�
nCyJ�fy��g
"Y�!;1	�i1��=uQ���m\�J��뽕X�����:׷���ȱ2t*G�����Q
X��0��P6�v¤��� �a֮��2r�&23�v]���G���j����Ԕ�2���/�W�5�U"����M�4�Zj��"���	������7x�V���)!44B�����kH�i2�o�r�����aCY5Zz�5aJ�6�_J,	��M�.3�)��@o�m�[mq����������,��U� ��r-����S|�Fg�V��6(}#�P8Y�g�]Ԝ�,��w]��n���0a�\IsD儩��0&����p�{�Nap�)3�Kvv��P��a<�Q�<�j˳����djư��z���v�8�)Ƴ~� ��Ū��	����ᎣbL�B2���}���j@:\��㊥��^���������i3��,�Z�]<3��eg�m��:&� z�é��r���2����|ۮV;�~Ћ���p�YǱۿ��N�p�Yȭc�8ݍS��_֟�*�!�)IǼe��p}�)b��.�j"������P*��
�
��X�&�ou���Rc`멻���2j{�0ql���oC��)/�
(���s�Q��69��,g\xJ?��k��[̨ߴ+-��	�6`fnn�h���o�b��[����A-_�a�,��J���|p2��%`�����D��������.kݕAIp�mL��� �t��>�Vm1�*�w��ݏk[-e0�s�A?-Iq-���ݝwo� ��22��X��Ġ0$�Qi����zx�R��T'	���eOJ�a[+�N!ů"j�/^�����ֻ IQ jlt�-^��P�<�@}��eN㭛"��)ܺ~b��P�@�d�=�\yj��l�1W��y}�lo	��z��A�hn��s]��,��ml��c����e���j�m�R�������[��mw�p�y�(��*����?c�d��)GR�a��4���kI�(�?��l�LSʛ���"����='߿��&�/n׶��q�&i�UѤ+͟��_�H�(�JN֦∧�wX�Ů�1m�����W�]�1"�I̖W=[^b�|7w���|%�����=H�q�_�K@ V�!��	3J
f�gW	��TBW��F
��Sl]��3,S�Y E�����d�æ|���\��C�=/�'�_�y�C������_�PyM�ø�j�o�0�k0��	g�A����MJ$���QM�&:`֦W~ڮHjT��cb����#;�mw\����O�1�O;��1��I	J��K��>�x,;M�:�1��-����x�5!��V8�օ�2�\Y�ܶ,kL��R���mt�GxK�M	�{y{z�J&�h�\#�����֫T�����[���E~�A�)�v߇H.���=rKخ��B��)j�o;�NlE�Ն��p���&���cu��Ltk]�"����0�ZZY��F���'G�X�Pʄ��kC���5�C^D$$���F��d1֐�W����m����sý	`�9_�+��0�����#a;��9r��\�r
g�K\�����87L��0���"|y�����{gN���n�e�,�o�[��Qý��	{���F��:�l[9��A�*x?�l�,v�;V��r�a�Y�:��B����������ǀЍ�IY237@W>�Rx������-��򭍋��wL��֘��or��O���̣]C_?J�6���b�.�A4@.P��[q�����{^7��hgN�ń#�"��:���v3L��a��������Rc�3��~"n���h�c��\����an�9��\��^yd�v�������:��l�<6j����g��?_/2���ƙ�qZ���5:����t\��p�kcg^��5��.��.+�D븚�l�N�ݍ�o��QU��1C=��L �}�K��AX�W���,�*��g�=�%KO6�4.I9Ձ�]���[󷅌C�ayH\�`����Td���\hA�6<u4|��s�g��%a�,��fi T��=��7z�*��q|/���΋�U�l��oR�r	:j�ҿ�w�,8�8n�Dd���a``|���wVE��׽xz�x� �`���O�U܂Z����+�>��{��{_���E���%|3����EqUi#?8��Lr$�-��?5��ԡF���/�S���%�R�NQ�P��?��Y�Ⱥ}V��������@�ۯf�J�(�G���kT��n��N�c��b�%.����3�B3�#�P3��H�`�e?�l%`9M8u�r����K6X���v�?�O�EZt=U�5}oi!<m3�i���B�^���Li�j�i�����׵�oD, /�O,\ʤcF��SU�|R��I�K�H���h����f���x	�~�v�_w���=Rez��Ő}��KW��B_�c+�r\���M���ЮT�\j�*�a	5l����Z�_��d/s�����EH��yϕ����]�y��)?�7d�"���.��S���������C~좞�Q꺢��xBd3C�w�%�G�	�*�,v����*p�,V�%�j��S�_�o�^�����tn]�F@#�0{�1���`�?sx�����RNNN��fm�t>��1v��h��bR��!11z��Wm�q
	�V��|ཽ�l�{h��~�� }1�O��#��ק�F�ۿp��6��k��9}�� E�GRIN�G\�u���ֻ�2�I��G�$y��/0��R�=��v���8���^<f_ⵣ�]�qb��9�Mk�T6[��:�d�+
�BZ#�Z�:����oB�3��i�?2��1��_��[B�l7^�j8�&�1�Jf�ҹ�I�����֐����%
�i_��A��[jNUUՠ݃>��\��N�׉iEa�G��ׇ�m�(���uH;�έ�D^0L�e�[[���:N:����s8�s��|�sj����u����������J�E�ceH|�� ��w�%Ta."���Z��ޥ �0�K���·K]V�G)��$)��3A�偁��4�Oe�/y�:����������@>�����
������E��3}�������:��᝿������l��r�U:��Ũ�U�Jd��`���W��ת�����f��8��vO���j�\n�u�;��Mķ��i}����7��. �>�x�v�C�c���h"e-	
z��/�$��
��(��k_.�x(;g�[Ӧc�^ڌ�*�|��rVV�69�]q�⚴|(�f�6@�s<>>~ˈ�Cub�h@�ʴa�)O�
[.]|)tOF�1�,������t�3�u�E��mΗi�w�J�ʍ�.�0���2^�<*����m�	������=�y}�E�C:d��FFa�?�nq��T�p�S[V��{s�t�VYƺ�[�����T���!��o�"##r9\po�(?O��3�feA"�������D��;�%/��&�uk<�b9MN��0�����	����B Q�}Ow�4�sw��^��FH� o�w�����I�Ո�m����ƛrx�0�$
�)�D�PS2V1��ϟ��*9OO�
�\˸�Uz_����%8��9��B��0��'���%��(�3�ɛa�etYHy8)�sr��BF�00���5�5԰�0(H(bs2�u����.��_��%����/l��m@ඖ��2a�����N�ԓ����ߝ9xĻ����ܤ�ַ�$<x"��潹�����u��?�j]\F����a7{������qXEȇ��f��V�?:rP��ފd����_*�A���%d�r����Oۭ7~/\�&��>�<�$4_���1rf�zOYU����	y�x��g$2���0�Z3����z|h*�eZyz�7{!(��7�.@�r7ޚW�C�^퇨��cp��+�I�+'n��<����wڏ��q���#�ڐLL
�f��#�$샻��ܞn$�և�<��'�r���3�G�/
����I�����~�Y@����g���3�<���n�m{t��j�T�pj���^�_�R����7�����`���jAq[j~ΰ�	�m�%��)�H���\n�+X�?N
6�L{�\`��S��nB�Ô���.B�����5]1| S�%�z���ћ�J��"J(9�<;)� �CT���r��.f�4��*/�AG_���%��}�o�Gk�L�q�Ȭ�k�H�Q}�����_*���F4��C��m�L	_~�{\��;�T\d�(v�
����.��lvҲc�;B!ƶ��t���:����2�iƬ;�,��ʯ�z4���7��9�~?"�.�R�^R`�,a��u�o)\(�C�cŮ�Pq��բf%7�S�fԛ��h��%��0���P��vYdDK��=�x}�+]����o�=P20�������_����ׇⷌ�j!{�~�ү;X�j�d�U�Ю�ݭ)�3���F��#��G��Ɍ���x^��+�[�	�J������ﬆ��cH72T�n~!
����bpt]���2%S��{	�n��Qc�M��h��F�R����c�E�$�|�ڊ������xӎS�b�����ᡤ�@�J�2���\�V3iq�$��s*hDG,Kɔ/ȟ���|��۫��g�f�I��=�dAR�y�wG��$���P��coD�<?�c��Z������nn�{��^��ub|T&خ@���.��F'OU�������߿�#���v�C&��aB[_�� jq���ߣ46|ӳ�����X��B ��(�p�̨.���N�J%�q�1�M��[a+�$$����MBGB�bT��\�����7Ka_��lJ|y�+kn��}}9w?Yj�υ�E��}��� Gț����?t(��nfrܗ%k�89��?���6)�|��
�8�U���'f�@a�[J����ek�;�܏_^��փ��y��S,��}��=7�|]�}r?��ӨǛ�G�ojQf@�a��&<��>c,?��O�by_��.�f3l��T+��h�A������Q��h!��!�P��v��ٿ��M����q[4O34@S��f&s��lx�p7[%LB\p|[����(���&��N1��(Sp�)v�4�h�sU�.���w� av0�U�DMm�GR>�%�b�����o�4w��8�j��"Җ"�/׶��f����o�9��LC�rC��4�h���J-����R��G�2.��Y���ڕ��B�ݨ���<X�e`��㭋1�fz'�����h���6�vMl<��è��͏�oOٛ|[K}ȋ�q���t�c1zWĞ@���-a������y�t�ѡGĭ��4�S���Ƨ�����?�
��Q��k������3�������;��"1!���ү�
M��#�	��Ц ��$OV����s�oۅF�aH���7����ת��,B�A3G�HWB<�O�fO�GGGP���Y�Њ�kg��1d�ל�6e���I�|�?ھ�\/_R;ƌq�q$�~O-גV��ʛW㮵�p)@(i��� �3 B���yM!���p�=�z_��C�ف�_�M���5y�"����	��tZ��9)<����魅AZ����|�TVC�@>���-��k�ȅS���mN�=6� �h�N"�5��̊=|��R� �k�)E:\�򑼵'{Ɯ!�8FE���ov��w��c���?��6ne�R������dO���i���y]�2DQN�a�#���c����J�
>�
aQE�>ֿ�˛4��7�.-!��Hjdh�wr���A9�ǐe��tV���Sڦ�T`'��e�3�w���V;�u���:�lp�LI�b�P��:R�4���LSPF��Q��}ZU��t{���32kPBF�����n�Lp���۸;}Bс�m�%�e�Yd�T:�x�5�@���*��}��-�)�2Q�	ծ����|�芏�D=�6�Y�������׸�������k�u��ԟ;:H��
4E���Ht�/ZVd;���(j4�*Ԅ�ԤI���]7���Q'��K'�(�\�M�,�m^Z5��@C��]�5���'�"��?4n��P%���p�u@�Z^	egl�kkI
t�k�N_�u���4��1�8'�� �4�~��7V��m0^1"��"���~���:���(AY{��#�9C��nZ���gg%Қ��A�>�C���D�@�oYu��=�{d@�z�
�g��t��0n+>8Z�WZ��.�)>.��)�5;�z>����>�P{����V`�֏�b�ǹlZ*9� �������O��)����(�i��X0�������)ۦ]�Zx(�r�FQ�Y��>� �[������	P��(�e-8ہ���0�[c⪣��ϱ/��ڬ�-�����b��v���z{TUaR����ZkY]�߬1z���Mu	qzR�~_S�|4����xG[ŋw�VN��0�I���	���X����{�P������w�Rit`D������kW|����>��j�5��mZO���i�`�]KE��v��=u�d���M�֓(;H�-�dwm�+��], 2���QO����GMZ�JOZXӳ��@��D���C��O����+��O��5+K���$sP�'j|�ݸ#�L9���P���K�L�	���ޫ`/�ɝ�n٘�-N�����V�[e�#-B�"S��՚?P�*T���}:q�)���L���z��1Y�Vj��燗�}V�0e���嚄���8� E
�XD��ݎ7i�%�U������/OA�0@�p�冉P�|K�.|uP���.�q�1:�o�����8��B��6�JZ ��tۊ(�V���d9�ߕ�ME���^{kb�Ă����A�L�����SA&�xI~��y�4�j���j�q2��Kjs��?:�R[�R_:7�"�g����t�E�Y[���ƭ����?%�ll�q��
�h�9݆_UHg�v�"�2�J<���D���渪*Zʔ�F�������A,��/)�;`���oDJ����oc����t]�k��+2��b��]2�P���mT:�۽f�g(�I������Mi�=ՋG�3���}{8M�d��^��{G�C�?q�hh��\���[ m���<�ug�=�ڠ�i�!3Ѡ��/�<S�'u�sߒ�U�U \��D}���_���MfJ�կ`�8��Y�쮵��iF�\�FE_MN��3i�q�1? Q���q?M���S��J�s�{BѪ����� f)�EӽN�	�=O��͘v���!�:Ș�D��Y��3_SA��-B���4����L�\>��"��a�_�m���a~zcL���C�链����<s���p0�s��/�
i;�������1~�U�~7��;����@���3O�Vq�d?�}f��~������z��D�Y��j��n���)S��ށ�����4�P%D�#�53i�m���I#�`^�m�I��-씽VÚ�i?�Q"'ǰ�M[���4��
�p���������H˵>�k��.�	�O����0�	f� �p�Q/���pR�M�
uy@�/�ư Aeg�թc$�1�VL1��YVX#�"�KP��~G$.]+���Q��Օ�VT��Q�}:Yh0�_��4�g6L��1%:�%����=m@�5=ɒ�(r�ګ�����_�N�|X�������L��Ӑ����UҘ,�lyn�^���{��ty�s'�ָweG���]�G7��1�4�����E�j!����ؔ��Ll\���&����i���3��}%�N7�e���Z�g^R�B��r��z}���PG7�'�ə�X+p�>��	T�(��#�|n|�{�Φn�8�	��gw�-Ox��'e�� ��=aC���O���s1�����x#�r3[w2�X[s����ʕ�w�@����!�x�lv���fq��s��}]`m���[;�տk�wk&�*��fj|<�I�>��t�����L>T7��s/<'Zj�K����d���%P8o�J70���	��B|�>�w�����HF�m�y���G)�.�7U�k �c��	f?��!!���>�Z������Co|�3LϠ^�B������/K���n�jU�|�
X��P�{��^Zk~jX���&�j�r��f�$��ZN}u���*� �?���0|�OU8�~1��U��
4�Zu��ѐQ9�&�dxP������	ù�i�\�ڣ��iQQ�[���ͭ�3*�irwĜuf��I2�i�m+W��}��V�D�P{����9PIEe�Q;]E��s�8`��5[
u��k�1��a+�N�R~�t�ÔD���K?�Yt�;s�:���X���i�Վ���r�5D����2i�"���9�Qn6�.R�_Y+̗������ԯUR"����:,�'���S̎�K{(��چ����_�[�ą?����V��8�4���$�J<d[�j��̢w�|�R�KW �T��v�
�G#�$׊�&4A%��׺��TV��6׀�5��.��M�u7����gs������&%˸n`{�� ��*Υ۶U�}he�)}�ÇY}xo���Q�`�G�rP���W� ��\w�}�k[���/o��Z�i���ݯ�h3����.�/0k��ya���s6{�EP��HN���'�X�~3�2M�%[=��� ǙZ��ca~��$-����9)�6�y��u�*SLf����f��Z���h�5wh�}��K�Js�ݹ�'�v�$o0l@M�e�'`�����8R[��<f�<b:�6~��N�*�q83�B�(�#��3�j�LP�}`$��7�ZP�uVc�����.ǝ+G��S(���^�P"��,;��wo�J����k���|&��Q�A�1��j�XO/L?���=�Ƈ�wWt�֘c@nt(�Krd��D������oT�#U����	�SP+QH{+�8X0G��?9�w���k����J�SUh>y�pE���Όsǻ�
��
�,צ�o\̏Ϲ�?k��A�UW��Չ�J>8�Z͍���΅h8j@�JU�v�Kda�Pj�g��o���ϓ�{ѵ4�y�I⸌\�1ԱH�^[5`Ee������m�
�j�,+|#�ן�M�����C�FԖ�C����Zn�ٰ�S%'�a���P7�>�$G��A�2����&��I7�d�l+��ɞI�+]��Qp��ŵd�0�y�v5�s�vљL|v�e�v��Х/ /
W|�(S�T��`v������e����o�}��Q����d���+R/'� ���i0�iY�*�8#��hi�#�W�k���@+����Z�<�ZI�Ň-:s�P]�o���-���co�m⽝������c*���* t��5U�����4��fӠB����H�x�rw�K���*Kъ�#�"a��0@"W��Mr���'!��lb6�.$�$ڶɧ/'��rh �(�3�lM�LI�B)�\)�̦K��*
�?��CwK<��Su�_���{���m��Tb�H�ʑ�t�[�|�#ά!ډ��V��c�����*�xq���Ҥ�N�u�[� ������5�jۻ�P]��f��1S}�N�]�y����� �����T�c�62���R�mc�vE�F$u��y���4��{�};��m��'�G7fn���m��a�������qJ�lu�Hۘ-�7�O���ۍ��s�.�*��M�.I�(��B6�n�'�~'��*Ո��R�T�qf�R:E^!m�OS�7,r=�뤦`��gA��x����M)dG��|�.]����W���P������<%�ԝT��H�ʭtT���%z�S�՛Ĝ>)Q�y	����iR�]��R��^y�*��2�*H�2��>S�t�/���I�)�k�5#��m�'��'Ce�t�� i�'$��,? �oU��9�~)u���Zɣ���Ċ�i]%i��+*?�ӕ����'�%�u�8e��m�Vi+�.8���W6��K
e�Q�FS;M�q�JꒃNwt����N}p�NZ�x�%8����,D_�Q-��Ά��r��3�0W���*�Ҁ�|ْ��TY+��pI6�s�d��M���~ʢү���u7J��}Аa��\�$d�ꈧCB��G�����{�s�H����7)f�&�&�H
eʱ�fc����	���H��g���Ѷ9�<"r/
�}60�u�_x�T��t��8������4�G]Q�;vܤ+s��w��K���L�y\����Ǯ})w�� f/�-���!�����2��#�v����	C�kX�Kт��F;��.��*�����'4���q�)��Ҥ��6���0iF�̪�?W�.Ua��/PB�oIW���<+Q���9��׀~Q�xh��{' ���\�p�F�˴��l�,`��S.8���Wa�s-CE����M6�`��ų�'qL���J2�~���gț�����\'�!�K/�c��m����6��r�|l����?~u��8���qI���v
��v4�&͒Y!$�ש�8�x�gw�>�E˴hx]�h\�U�"W&SB�G�#�j��^�?�[����Q�ץ�1���"o�L=l�KѢ9�/�5��z�)5L�%JE(ʚ%ɚ6��Gk$v�aEa+��fw���*_���F�Z�%�:iڌ�P�/�u�V������#����&�&�*�?jIZ߯l/�[�4(9�
��+F�.�����}�-�����M��H󞦚a$ŕ�����r�%�m�F�Y[��VXlh�9�a=jt�a�e�9�G�HJ�g���Y���=�1è���md��)Oൂ�諰�\6I�����3�Q�#�]�PC��$�G�V�%��0�N	C�5'�eeD���z�#m�rzK���?�5���hX�^�	g?�X�樷�{� C���w�����/+��<����nr�Xj��)�V�n�ٹ�9a�9M��N:kBqxIn��z&ͫ�W�%w(�(Vn^�-�50�ޥ��_{�86�2����A߷F)�Q�ɨ����K����c%,������Y|���1�j���N�ײTy5-K-�N���o_3�})�Ѷ���9���k�dp����<�q�J;[��~�p� �C����*"��x&[�H��:M F$�����ds1�zLA����]fۖ�߿��6�58(��u�F8nW��D�O{���7n��׼�q膳<��-��M'�v�$�w��FW.)�ɟ6���05�D�jm�I�"�3YvL6��P�y)��ٱ,o��抵���\�a1�z��|5h\�2�P��M4�t���~�wVo��. C$W���:t��$E�ԓ(���k�K�$�l��0�5�n�����E����O����7l�E3�ڥ��X�Hu-�i�J7 �A+�P�˻|~�_\��k�l����j��L�ڡ09C�]4�F��(t��7q��#�����>-t�m�O�}��<�s�R����<"�<'[`�us�/�Ǿ-I�˺ο�Cl�1�Ěc2��ƙ+�N�k"ky��O�;���s[�Z5���+�k�.��N��l�V�d�� Q�b>\Ge�,\����gG�?��1��/0�_�ğM?�@�٢��]��sc���|�{tC���/w�΋�7Ia<�Ozw�&a�N�.�'s���{j�B�vh�r���\V������_wp$��T�j�T~/X����<�Ȣհ0�����:mF�W�Z�����`�x6��-���q��,g^gzMܸo�8.ˈD�����{N��|۸�[G8�緟{
/:M���8���Aɧ��͢�	�[�ut��y�*V��=�708���/w8]^���}dhq�ɿ4�1Ok�hU������p�c��xK���|Fo�]s.a��ȹ�X��G��\=3��+|~N�+��Q*��3��Zf�tr���2|O׏XF%�X|B���?	b接�|\�թ+�5u�ِ�4+Uܜ��̒��|�����dUddP�[\?�M]�Dj�E�~%ݸ]�XV�+��u�!�@������c=kC�*��|���3.�l���K>���8[9�+%c���y1����M����f�4MT���'�
 y�����4�Dl#~���ߎ)�eT���p�� ��x�n�-,�0���E��y���j��ָ��g�¼�1{N�߈g�g�:ӠA@�k�R�C�.�Ѭ��[T�>x#�~����G?�׻1k[��Z�U0�4�� G4J��$9�[ɓ��쓗	d$e��
�7d�6�DV���ލ��a��ҲpYpVD��	6نz�ۿ̽�7���%��q��n�O���*\&����B���s_wzUM����hQ?.{����j��fH	H3EA�J	� �"E��CEJ�һt�"��5\%�N(^��G/���Q��������zo���?^���9{�=�73����3�:>�Ѿ�L�6,�/���c9��:�$I�Ǎ��i�]�й���;ڟ�z� �Q�*�zD��	���/+?Z>N�-�T��[��b46�y��K�4/3�T��8�<HE!.P�.ɒ7�T��^SdC>NB�$D��p�C���(YØ!�����<�Wc����u	q�6�� �'�����;X�U��E��rr�CƉ��J )N�1�A epo�>�6��m�U�T(���+�x�jl��9ğ�b�z�_�+z��T���f���g����Ҫ���&�#��Ogr�����`{��h��4�#󂛳����W*�٩��*�!�Ï�#/2��d�W4�]�r�f4�Nm"��s�k��agljz�e�.o� 𧱱�o����e:X�*�w�?�ʪ�sI>hg�!�,���V|���n3������ബz\˻�����]�e����?�5L)+�l�!�ޥ��8�n��-,g+Y���KzuK�g+�Wڇ4_�EN
�|0�j����Ȅ�ՠ���L�dS�P�`�{��Nt1�:ud;1V�(-&t{s��-�����XNQ�NU���6@�k�Op�i$tb+<[�ӫ�׾�z�dU����?6�(����$���2ll�
G�{��4Rٲ[=���59���[�8P������J���\���	t-��3nг�n�s�8ߨ�i���ɝ����X���������Z����1M��O�-4Z��y��i8%�TE�����&�a�֟XZ������>��}�+q�~n�p9��"^ jdYl^�#wG뺽Ćj�\����vK��A�œ���h�PB6�9P�C5^�x�N*��]���!�gT�`�i�@��癪����k�?�(��S��s��LW��$|��ك���K�7���h?x�W˟^2�����e����8�T�Z��։t�?�`��ف����m��	cG;i�Yi��5�?W/�>s�j� �Z���T�+�	�D�*�����M�'��҅�s{��7�	�e�tg<�pM�U���/�V!5#���9{t��\V.+8k�A8Z�#IՍj>;�er�(�G�БNٻ�'Ɲ�u�4��F��}�.��S�tu�������2R&\�3�sǯhӗ����<�څN+��@���|����h�B�ہ��Z�NΕ��;���.���� ��wɐ�C9级�9n���`����ۓ��P��~�l���ɞ�BFh��2nǩ���f�!�- >��4{h v���v�dl����U;����WA���9	Է����a��z,��b��4�D�߬}���4Z�Z�ٷ��Ƶ�nw�~r�S�oO�{S&�>3�:�Ɋ��g����}���'�38`Ig��-���jb��CЇ�5J��
��I_�%��1����IO��|�W'�g�d�S!���f~��w�w�D�9g��s�a�8�T�72�!�?)����l��u��o�X�sE�d��x�;�t�m��.�]ja�������5�+��WB��B���x�pn��@��Mݾ�qH�,)�������;Z�xjg�war�k�"�^�Ie����m����r�PS��EP��	kB���+H:i�lv�J��;!u�W��=�QХN��rq���?��|	�D�vǂ��;ѤB�C���Q��l�u�3�C��Un�755.�D��R�k)��:*�ڴ��P��E���y��"�wԭ~��)�<��Io=�\�"�~�(gɇ��*�!��Y�!;������)5�w�|t�!kq58�՗���X�l&�S�K�κ�ry1,�ޘ�R��z����1sp��<QSe!j�D��t���#*�oGf���TKD]X��a�T�A^��?���Q�ᚄ/.���B����. �	*��k;�-�z4R�/ gv�E?V[�h�wԬ��a���8�2B�I���I�×���L0��޳�nnچ�TV��Y���߿K�17���5���/��,+��r3�����6��v�Z����Z|���'*�erز�z�h�N�`�s�ƙ&�6���+b��9$D��WA˼��Pp�Ä3�&c�Q��s,�_9�f�\]�����&*�4M�"Nޜ�կ�UW�۝7WoKfi���h�\HG3l�I���Ӫ'�L��������#!EWZe1
7x�[������M��^ET�2R�Ԣ�&	�~��_�]�O����t�d��ߚ��-���T-�WQn
f!��x��j~�[��A��oDme�r-0��[|,f!t0f�_������z��1��L�q+�{�bƛ�yA��u�{,&&r'klS��▽�a���p3ւ�3z��Z5;$��f�O���� ���ŧp��Wsᦈ2E*e��L�}����c�f���M��@�Y�_4���I= ���Y��SF��ֺ���^����!p]��ɡ�kpm�[m6^x���i��
ip�W<��:�O��	Mn�>�y��C���np���\���Zͼ�J����F�;y_�{����Zg��d�\lz�L4��]
�`.��oVF봿�}W�aǖ�6Yh�~�u.Ε�R����"�~���k ��&塑�C`ϧ�1�P��ǡ� �=�n�7gN|�׌Z)�m��,��6¬�{#�Q�ܯT�kԽ�m� �Q̩r��s�m:�w�c��Ӗ�-����ő��}�A�O�Sy��_>�U���H߼!��%���a���؞�-Q(ý�gr%s;�xzw[��\���UH���HC��S�16��q��>EX,gy=�<�8Og�rL�+;r���ScO�GGd��$�3��{f�Y[��g�
$\̭��k�������N�o��&�x��A����Z��a�y�_џ/��AQ,�>�y*�`~��>"�*vG�xY���B/�B���Oa�����Fn;q�~��o��%V�����ɽ��?�<�@��Y;& �v&��}�pS*_�����E�62.��S�:���7��s��c�N��� y��Q�Dk�y~�<�hT�w k]�����q ��$:��uE�U#�Ե�~}[W��@e(l0������p`_Z]z�*��������j�lF�5<NI�xb��X���Hi�受^�HY�`�>������V>�����c��Ks��]0�wl;W�ͭ1ZǛ��D�������\F��!�<�G�f�9��<w� j���;����8*���������4`k�oҶ��{����L�T�����l�!��%��ψL���4�:��嚗�&AH߭2����X(�?�yM|Y����Sn��a4���Vu��#�9Wr���֌��X}C�1�p:��������ف\�
^eFWWW-�ބS�B��찒�2KB'A�ׁ�ze�샑�:%�e�^e��+_�b'|n� �I򕱝5,�������� �d�z0��l�����Ej�cDBBBP���!��uu\9$!7�I���AQF꧗{�s+FٰK�r���]iT_���BG�{A����:���-��ǣ%�ȅ�?���wqw׹�����ޝu�ihfffs�4H��@v4�*u���JO�ZF�O��n&��˻ٸ;�{�EW���"�W�,��x8���p�Ѡ���)�95���i [�Pn}}=��^�ttuu��	x�ɻ�O�:v]�Z� Ev\S�IGe�p�:�7��s��5�j�yꉵsA��?>?t_ �{-2ULO~�@���{��ӧB��҂�gOO1�:\-L����'�͓���DvP�(�6���� ��ަÏ#7ۯSz�%�\�*M�ÓCx m�3���+�'�?�s &0��*7���f��v����#��Y�U������{���=$��h�q���ڨ������v�H^�]c�F?���|�pgww"��gOD9I����K�%ј���04U^������YFɴE������B
<�&�|7,�a��+�Y�O<z�`���'���
ϕ����Jɋ����$�-��{��ѝI	�I��XȠNj���'��K
I9���iK`�P���ߴ��e~c9f��]�i"9���E�W����(�@s����Q��s_c9�Iھ�R��)��cA�����/���=�dQ�&�U�>>��"�}�:�1�5۹�v���~��gaՙ�u٩$?2րc��(�n.��C��+����ZHO�۶���2R�.V?���l�+�?�$�,ٱ���w.�|`�Η$��,���0��v���MbEA5�o/c�4���I�`h����
��70�W��sh�|�@)�~�M��
��D ��`����W����.����ؕ���|��&a�?��A���n�ӠT�;�|�	�"����5�
����6��P\)��[N��9�I�`��=��C];��*+g4�,�G��ضQ}���F�XO�T"̣���;nx6���m�B` ֟�����P���枞�"��� *��qGGG-o�%ν(�K���T��p��p��L�§�v)��e;�H���ֻ�b�/�{�R�e��bK�`6hp��_%�m	����իV�����A,�-�����tG(�E���8F��cf�KU�h��S�b	 �L7���A�x�D�*�&cT780ͬ��b�Q��Oin�@6�{{{�u��f1/�����xGznn��C��Q!�C@�,HV�����[5̫���u5�i�A /��ݜq
��[?ݟ#�y�$�a��XU��"������><;I$�)9� ���J�f�`n�ST*��������;r��p�{�	x��z�m%�91]����:���?�QTQ�-��(/�p�����dn� Q��k䳖�}�ݭ-+/�||�yr���ID��t��	%��lY�A ��H�	a�{��j#�yj����&E��Dc�(�a�A-� f3e��yx��t,�u�~����C _�6Z��V�G.G��7�vŨ���s��Ro�5}ͯ5�#xTLQe�]r��U�"q8[- K�m�?~d�?�5�"b�=T__���Ұ4�1�Ez�ܦ�����h6��K����J\��Z�R�أaDMUVQA��1>>6�jDi�<y��)C���UT�sPS��k�x221���2WWɄw,x����I�[�O���ԋ�i�����/��:D��.6���]��OO�P�J�6�? PK   �cU�rH�  �     jsons/user_defined.json�_o�0ſ��g�� y��6UZ�*��2EƦ�D�aU��:YZuh������{|}أ~�i�D���ҵ�Z���Λ��A'1�?� �h�u^ܖ��f�֞��*{}ߺh�g �+~�2
�4�Rq�0IT���
�<aXs)���T�8�̹tٻA?�/�������[w����;{u��׶n�r���P�5�n�6p?D�Lp�A�r�n���Y*hz�f1X�8�{�6�3@��A�M�yc؁Ƃ�,���g$ ������A���M)u��C�g2'�1t]6�{{�����O������N���8�X�ڙs�߲�i�ج�'��:'%üL�YUc�k�K�IF��Z�G8�ৄ#�Ӕ�|��<��<e��A(�:�E$1�`�Ǘ�jFD�'���l��Q>��'�����|v�x����A6����b�o49����'PK
   �cU��	�<  ��                  cirkitFile.jsonPK
   1�_U���R�$  �/  /             i  images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   L�_U�
L��\ �j /             f?  images/5d6e91a3-4a01-48cf-b4fe-ab41826b34fd.pngPK
   �cU�rH�  �               �� jsons/user_defined.jsonPK      <  ��   