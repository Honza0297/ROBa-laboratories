PK   �I�U�G^!  �]    cirkitFile.json���Hr���@�:4��替����-p��m�H�2;r4�����.jfwF=ꭧ�p�|�ؿyT�)�GvW^�?l���a3��9<�����R�,�[�?.��nw��q?|{X~�n�����8��qS���z�Oc��*�j��b������J��VR�U�Yv]hW����x����oW�B��`UCif�*��23X��V�0�f�B3�U!�������`UCof�*�e/�f�D�J{�{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K�k+-|�
����������,�:l�z�5E��U�j�}��)�m��m7�fqsi�v˲J?����"�u],c�m��i����*]/��5���l�D� .p�5���l�D��3�xUJkJ��}Y[~��h������Ua�H��
�D��U�%����,�,��2�,�(�%�,�(�%�,�(����]�/����~�m�H��i�H��i�H��i�H��i�C��N�D���N�D���N�D���N�D� ���kg��N�DP3i����h��f�Da��f�Da��f�0���i�H��i�H��i�H��i�H��i�H�1{���,�(��,�(��,�(��,��^;���^;���^;'�?n�a���zR��q�<�?������[���t�҅$��N�ءt�҅�dcW��C鄥C�Ʈbc��	K�<�����.]C����ءt�ҥo{6v;�NX�0�l�Z6v(��ta���ul�P:a��г���ءt���$H��v,��|:}��.h{�������O����]�'0�N���;�O`>���v,��|:���8X>��tj8?�u�|��v8~��`�����p�`���	̧	�̰�`��ӥp�`���	̧�(���O8�G��(a�Q�����O�����'0�������O`>]���,��|����?X>��t�?��|��/8~��`����i�$��|��:8~��`����p�`���	̧k��ѳ��iV���`�Q�����O׏����'0��|����O`>]���,��|����?X>��t�4?��|��
o6~�,��|�6��?X>��tU=?��|�i? 8~��`���Np���R�D�D��|�i�8~��`��Ӿp�`���	̧;�������O{�����'0�vIa�W�����O������'0�v�����O`>���,��|���?X>����?z�9���5�?j��|�i�(8~��`��ӮWp�`���	̧���������O;���k`���	̧=��������O������'��en;q��/s�yo����M�r�̰?o�9��wg��󦛙�ϻef?os�9��?en�X�Θw���r�3o��X�xc�M6��o̾�&Z���7�@*w����o��R�xc�M��o̿��>���7�S'��˘�}lr�[�x��W����7�e�����lԒ;ޘ���Qr��w�!I�xc�N6�o�p4��ɖ��/}���g��E�xc�Nv�Ƚp7��d7������점;�j|��;�o w�1�&=�s��o�W?w�1�&��s��1�_cu���k����1�_k̿֘�1�Zc����k���Zo��5�_k̿Θ�1�:c�u�������_S�m��+��"J�,��m_��1��������=߫��G?�}�,e[lc�-b��[����&.;i���~�_5|��_�O���9�\9_���������~�������-�)����7t�� 
#�
���!���>�`� ���R"H(���
�ć!���>Db� ��ϥ"H(�.�
��3�DrU�+�X��pSJa|r1a�[��M)��	'Ą�o�
8��'�V�+�R�CLX/�:N)���6��]s�X/�:N)��4)���L��Ƅ��r���-'���X���8�b��x��qJ)�3/ &��WX���8Cb��x��qJ)�3Y &��W��8��)3V�+��SJa��1au���8��)HV�#V�)�0N����:�:N)�qJ����n�cu<bu�R
�t6�	����R��ALX�X���8�z�����R�!BLX��:N)�q�$��=��obu���8�ƹ�V�k��SJa��
1au���8�ƹ�V����)�/�>_s���+�	Uqa�0����U��z��k����`\=XŅ5��pU0���|�K\�;�1�`�t���cL<XŅ5]�����Vqa�yo2\�������g�
�ՃU\X�p��W���*.�:'���8.Z�չ�>�ur]N���w�����B+>�:��'�>�˅V|huμOl}����������0Z��5>��qb.��C�k1|b���\hŇVה���Ǒ�Њ���񉭏+s�Z]���`�Ǘ�Њ��U򉭏/s�Z]s�[�'bN��||Y���J_�B+>���'�>�̅V|hu-�Ol}|�����D����2Z�յ�>���e.��C�kD}b���\hŇV׺���Ǘ�Њ���������\hŇV����Ǘ�Њ�������/s�Z]�[�يN�}|Y���*_�B+>��6�'�>�̅V|h�ǀOl}|����j�����2Z�՞>���e.��C��+|b���\hŇV{p��6��2Z��^">���e.��C�=Q|b���\hŇV{����Ǘ�Њ�����J2��d>�,������\hŇV{���Ǘ�Њ��>򉭏/s�Z���[_�B+>�ڋ�'�>�̅V|h���Klk_�B+>���'�>�̅V|h�ǙOl}|����j�6����2Z�՞s>���e.��C���|b���é͇�/�}|Y���\hŇV{���Ǘ�Њ��d􉭏/s�Z�-�[_�B+>��#�%���/s�Z���[_�B+>�ڳ�'�>�̅V����|��m��Lo�L��n��*3}�3Uf:og�����T��n��2ӏ:w3yDe��sn�A��d�ܦ��2L��m��+�d����2L�m�+�d��f��2Pf�xn��\&����̕a�xn��\&���5���e�xn��\�R���Ӷz�MMse�,�ۼ.W���-�re�,�ۈ-W�����re�+b����+�d��n[�2L��i��:�,��9*W�����re c�d���E�2L�m�+�d��&<�2L�mu�+�dq�dqݟ`��a��a��a��e��e��e��e��e��e���n�1Y�2Y�2Y�1Y�1Y�1Y�1Y�1Yܽ��MU�u:�(c��(ͲX��}Q��Я6�n�����W��z�Bߗ�R��66�"��)��J��nⲓ�i���,W��ʲ]Ų�*)�۪+bX��2�}�v��mb�:����,K��s�/��p���q�x��W��M���~��xX�=��ߓ
�gE� �0>B� �0>kB� �0>�B� �0>C� �0>OC� �0>�C� �0>�C� �0>3D� �pz�ȔH�jse�ۂnJ)��2LX��xSJ�� �a��`�R
�G�V�+�R8=4g��:^bu�R
���w��]�cu���8�N�&���X���i>Ä����R8��`��:^bu�R
�9(���x��qJ)�f�0Lܝ�V
V�+��SJ�4	�a��x��qJ)��'1LX��:N)���)�	����R8M�b��:�:N)��d3���'����x��8�Ns�&��G��SJ�4ۏa��x��8�N��G?X��:N)��I�	��5V�)�p���0qO7�ǛX��:N)��U�	��5V�)�p�<�0au���8�N�z&��7X�S�_�>�@������*.�a�tO�U��z��k&�hU0�����I7;Z�����&���I#;$����\�:ib�D��U\X�5�K\'�x��k&��hU0�����I�:Z������aҵ�V���*.�:'���8.Z�չ�>�ur]N���w�����B+>�:��'�>�˅V|huμOl}����������0Z��5>��qb.��C�k1|b���\hŇVה���Ǒ�Њ���񉭏+s�Z]���`�Ǘ�Њ��U򉭏/s�Z]s�[�'bN��||Y���J_�B+>���'�>�̅V|hu-�Ol}|�����D����2Z�յ�>���e.��C�kD}b���\hŇV׺���Ǘ�Њ���������\hŇV����Ǘ�Њ�������/s�Z]�[�يN�}|Y���*_�B+>��6�'�>�̅V|h�ǀOl}|����j�����2Z�՞>���e.��C��+|b���\hŇV{p��6��2Z��^">���e.��C�=Q|b���\hŇV{����Ǘ�Њ�����J2��d>�,������\hŇV{���Ǘ�Њ��>򉭏/s�Z���[_�B+>�ڋ�'�>�̅V|h���Klk_�B+>���'�>�̅V|h�ǙOl}|����j�6����2Z�՞s>���e.��C���|b���é͇�/�}|Y���\hŇV{���Ǘ�Њ��d􉭏/s�Z�-�[_�B+>��#�%���/s�Z���[_�B+>�ڳ�'�>�̅V�����{��m��Lo�L��n��*3}�3Uf:og�����T��n��2ӏ:w�wDe��sn�A��d�ܦ��2L��m��+�d����2L�m�+�d��f��2Pf�xn��\&����̕a�xn��\&���5���e�xn��\�R���m�re�,�ۼ.W���-�re�,�ۈ-W�����re�+b&���˕a�xn��\&�����uL���+�d���L�2��c�xn�\&��ʕa�xn�\&�綺ɕa��a����O0Y�0Y�0Y�0Y�2Y�2Y�2Y�2Y�2Y�2Y�B�٘,n�,n�,�,�,�,�,�,�^�⦪�:^�1�E�fY,�۾(oc�WY7u�����T^=O���e)�b�m���r%E\7q�I�4��u��T^eٮbYV��m�1��b۾h�uL�6�_��r��s�/7���tn�w�ð[��x[�,~�6�ǻ��f=���a�9,޾{g�{�8���^|�ygR6����<c/~zv��B><��a����������x�8����o�n��E��S��Ε�ڒ���V����1�v����<nҷ�ӿ����'���i�^��l�y��>X��.��#�Y"��(�f�0N�0R�%�8��Ha��4#�Y"��H�f�0NC1R�%�8��Ha��4#�Y"���X�Q=��	�O
�]#�fY9�*@�k��\$+PG(�v�p�e� j� �ԮN�@='t�����z(�%P^��4�����(�v�p��v�.���㜹3,�)���(�v�p��g� �o	_�F8M#�r ŷ.f��4���T�
��v�p�Ji� �m\��5�i2����PO��4�����
��v�p��j� �i�]#���Z9�z�zj��I�V�+q�����v�p��l� �i�]#�fF[9�z�zj�����g@=��zj����V���@=�k���t+�Ȋxf����v�p�bo� �i�S�F8M�r ���]#��X9�z� �t���Ycҹ��;��0�	�'0_&�Y8=$~,��|a�t`�����|�a����C���	̗��IkK��e��K�p�&�+�����/]�񛴨4~^�O`�0L�QrzH�X>���0�8��!�c��ä�$��ď��O'5�д�	�&�	�tq��ڇmD�v"0�Є:��!�F`B�	u/Cڑ��B�d:��+�	�&���tig
M�����&�P'��1�
L(4�N��cH��PhB],@ߨ�}
L(4��l�cH��PhB]�A�b�?2�}JI����)0�Є���!�S`B�	u�Cڧ��B�:#:��O�	�&�5Rti�
M����>&�Pצ�1�}
L(4����'��>&�P��1�}
L(4��g�cH��PhB]�I��݅O�}JE����)0�Є���!�S`B�	u�.Cڧ��B��c:��O�	�&�u�ti�
M�k���>&�P׫�1��O�	�&Ե�ti�
M�}��>&�P{�1�}
L(4��g�c��D����>%�>%�>&�P�b�1�}
L(4����cH��PhB�GBǐ�)0�Є�K��!�S`B�	�Ú�)0�Є�Æ�!�S`B�	��Cڧ��Bj� :��O�	�&ԾGti�
M�=�����e�O�i�R�>&�P{e�1�}
L(4����cH��PhB�QFǐ�)0�Є�_�aC��PhB�Gǐ�)0�Є�׎�!�S`By�0so�I����ބ��'=sw5���D�?�e�9~҃4w'w��I����^���cN@kN�d����t�\kN�����t��\k&N7��0�Bk&N����f�t/�\k&NwO��f�t����4k&Nw�0-[3�����e��8��ĜnC�+`M���/�K�Ĝn��+`M���&��9�N$;��o$��gM��F��Ĝn}�+`M��f��Ĝn�+`M��
��L�na�+`�����L�����fbc���쪭��X3��fbc��֚��5[k&��Ll���Z3�5��fbk��֚��5;k&v�L쬙�Y3��J&6U�������.�4�b���EyC��Ⱥ�����j�W�A��rYʶ��f[�>6E�\I�M\v�6M���Ͽj�W~�v˲��hn���a]���Eۭc
ᶉ�j���zi��K�_n�����q?$����ϋkN����\��W�*���O��4�O��t�O�ǌꑢ��+z��Ѣ��/:@tD�#�Q[G�:����(uD�#JQ�JGT:�qtD�#*Q�JGT:��QGDuD?���:"ꈨ#���:�����uD�#��C�ZG�:����htD�#��FG4c�tD�#��VG�:����huD�#�1�:�����tD�#:��NG�_��3_����d��d�����)�>���~s�tқ�s�!�[2�~]~���S"yA�D-7��|��`�iʙ�^Y�l������8�-W�;͆i,�}s�;����1�%ӷ�ǷJ-s˻����~��vG�U�M5��>m�_�p��Ǣѯ�M�*)��U�������v�/۪�-�v�M_��_�w���Û�q(ʗ/���>깢q?<+���<.����o����q�+����/=�)�������Y����ݛ�˻O��P�z}��%�E������?&��ۭ~���������nu�����?�����1a�S����S�H�O���k �{FrX������q��;��)�
	͛2���o��}S�p*�ӰE�mS�MQn6U�ץ���2��Z�����e�I_������k�`o��.���f�2#�����n�x�eY��o�.|�I�����җ3o�s#��qnD57B�F��;����m9�F=7"΍(�F����������o�������8�zS^~��9�?;�)Nڙ7ʹ�و���刯(5}}�g�ޘ^�~����`�^���z5s��$�^�t>ߙ���Ӥy|c�f�oL��i*?a��!~/�މr����F�̼�΍�fF�afD)s#���9K��79O�_N���O��i���k��|TU_sTy�V�L�����������q��j�x�9>\>��.߶3��3�Ǚ�˙����g����Kgvzԥ3;=�ҙ�.�<����������q��j�x�9>\>���N_og��g��3Ǘ3������~�I�kw����z�����p�\�7�&��o�e��۟�)�v�Ͽ�����:}�J3�.�,��Z���ҽ)���%���ή\���ӵf[o��$p�tɳoæ��mS�7]^\u^u'����zrQ����/
�/_�u}��ߒ6g!K߹}�Y쟂vSW�M݆�/��=�X�k�u�U�J^'_�Y��U�bW��^��V5���V�y��ᅘ���Y �..�eQ�.�ʪ�ky�Ǎ�ݛ���v"�^����u6�M����[�E��u2��Z������95�d�nʱ*�g��9�֒W#��z��~=֞�>��.��{��3�+OXz)>}դ�~ܭ�ߩBHW�U�C�ɿ����8��V���|��/��>�������x�o�����6?�g�j�?�O'�nx�x�~���8��~q�>U����������-�=�Qps�� �}m�:,�˫|�çU�^��s�'�a?�w��o���F���߿_�m�?o��7�2~<�o���j��5#�:>��n.��ώ�����KJ��'��}������!�'�6��39�M�x������6̈́����[�\w��5_����jM�p]�\wX�\���گs9U�U_�%�*�K���*q��T	�)Uꗙ"�K��Q�b
/
ĕG�K�K?��Eօ�N	��K���?o��<n�d_�Mʱ����٬���������x�|���×ŗ�PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   �H�U�T�S� a� /   images/dd298255-0ede-4bb4-88a7-459da88d83a5.png�eP���7�,8���@���$�4�@��N��w��!Xp�A�����sϽ�μ�·�������m����K��()H� �#BAA�HK��@A�lCA�J}��cb�%�^��r!���1�X�I�l��`W�	���HA#��������(RL�V���D�*�)g�.�Xq�FO$w���e���L1�b��9����î��U���3���W�m�I6#O�c,�j��w��͜�==��3�Me��o=t<^hꩿ[�w�'�.���3?��. u=m�]94���n���A��^z���jhه9}�`0���s>����8]��ͽ��2���[������7nayfhs��e�~��Ův� �����^��8�NwdS6$��7[Ƀ�m1��m�fB[ŗ�K�<LpK�"�K���'n�^�����Za�>�d�gI|��h�"�����(��
b�����3�����<�b���������b��y��r���'|f����)��d+@5�u|����5�����G�~��iL�i�+�`�;��/_��K}��3f��K$納1f�g�aޜ�n����+AP�������>L:9�6���K�!�Y�c�8�;���*)�d�]֮�Mz~�z�%��o����h����W�-LF)M�(����WT]�����NX�mL��i�3�źk�Ų��jܳ�a��	��}���� *e�=������\�S(Ls��c��j'X��VM�̍��Qk�$����̽`�gU�l�����Qx��]{>�|Jp�>�Z5���;�}X
�!���
Kit�;�}s��f����˔CA?�|e1��=�z����S|�� �[��C���[����L�x��-M��l�.w:��Q�ޥ]f��"�|(]X�
vx
�-@y`S��ȴ��dd���%�{AUto�!��A�CTf��s�U'�cG�%~���#,��RZ��}X̋�ĕ*� o�J����v��ǸW0�3�^���o���#���L��E�6�K���p�O�����咳�-ѹG�=��FT8u|n�m �LHiļDq��T�]i5;�nA����D�)����7�9Kj�U߯�Nz�&��^�����X�DPG�2�>$�����'} �Ϝ��0�0vX����/T��|϶	���xwT�̃m)�8���bi��jrѢ�&�5��,��R/�I�K�5��-����Y헭I�sQͷ��S���YYw1gf�mi�ph�$e��7��2���b��a:�%�or"��ƾG!D����b�&cw�W<2�W�<����/�ԢBbZ��^�VN.5"�*�J�_9���rպ����z�{�%�S��C���G=g��#�)�t���$�q���,/?���}sG>�����S�m���}���ʺ�LP�e!��P禨�>��M���H/m�h!�܉����gm�3����5�Kv���v���pA��Z�?��UQ�|�w��)��Z5]����,�-�[ND�CC��*0*7d�kl)�1�/�_����c2v���1�X�<����Ҁ�t�~��w�m�M?���+�R@�j�ESyEPkUG���[�[E���Gtì8��_�*���RIڅU#��m�^�~3e�u:����zg���s!�R�h2ו�jD�EN��5=�q9��j�(�>���+���ȡ�����?��p��B�F���/�8��{��6�)�Bߐm���*؉մ�ίHTI8]Z\)B��W����W����T���N���A:ڶ�#b��ô7���R6J����O��i���T��3N�ڣylm�Σ�A�̲p�p���k^_�N���H?���6oz����b�F�!�������F齆ufNX�&+�whf�h���i:]o ���R�+�N������e�/��Cf8�2H��Q�LoJc��C�YZ�h�C��q�`�����ѹ�\�\�%��4^��cG�N��S'r�����ORO�Q����R�h��򍓦�W�'F1���]��]�ԛ�Pt�@��� d���fK�G
�r�7�4@,9aw4�W3�����h��a�<bF���e�)9�ԡw�h<��&�؛��Jz�1�4������+��PHd���?2�ڭ#��f�K����Z�fqN������*})�ɄR-�c��`�J֑�`ċ�����G�7 ���['�h�)O=y�0Ӱ>w�0ڤ��M�؀��1�*綐���ѽ�k�9
验�O�8zQz7�m�zL.���MDu���iB����e,�K����X��JP��Y=z�Ͼ�+�K�z�P�6
�P�\)}%�s��Y��3��X�����f ���-��쫶�m,�U������;nW<���[a���kl%��C:�H��$X=n#�M�}��80��B���>�[RcJ	���)����CD�/�? T�ûQa,?C��q}𩀕�R���J�{���CJ�с���{P� z)���Wz�!���\�� �%�}� n"�άs	�@ߣ��D���T��9�-(+E���Vx��]q�ÿ�7bTu(���!B��a�����cG��=ܕнj,��YS7+���
E�|;�|������ݲnT٦O�$L�o��-.
[���xH��A����)���h�;cc�N'�9M����{�\���"�u�)��!h�v̷:>v !�E@]l"�Uie$��%��>oY���vA�p/��@�A���WT5{�6b�`�@o�y�>YG�BjNܑ.�Rh7�F�{���w�4�&L-�Pd���'r	��]��u�N�trɷ�'P쑒]���x���I��}f3�B)�����z���f�X1�����MY���#"�HD*�P��
� ���y�c�U�.�Y��kH!���DX)�[���O,�K-���́�����6�U���{���|5�f��vE���j��	�m��J`�>��B_b׭YV���U�@�����z�bQ��W��X4m�#�J�
�H�<���A=�r�D���x4c`�׋���:�Ð�6������Q�^L�a���Wu�tl|(W<�\%����@��έ���"_3[CѮ�+7V;_�7�D�vƤ@�������{�A%�2���}C� ����6J��'�{0����@��l��.��b��K3Q�q�v�V|?�ΰ�@���h�ɑp'��r��b#Ub{}�/�"��'1Vp�����ҿ.�S�}��I��BKC]�������6�\����E��uS-g`�#/P-!�-D���M3�P8`�Nּ�m�o�siA���Hcx
4�f��ۭ�h��Gjeg�3 �����$SM>[0O�oI�	��~o`I$��8�o,��#��BF5'�q�w��v�a��d�u��t�W�W�"{Cܵ�X���R1�g�ii:��;�o��v6T���yW�<� ��� q>�eT,?���U�~�<������O�VR�����wq�ppK�-ﹶ��V���:�ZLD_�2�oL�,fq�_e9����ے0d#���t݄ �Ԩ4p��	E'�b�QU��Z �щ:B�D�A�fB0%U)g<k�K�$��U~�y��)8^.�����Z���U���	�M� ��,G=��Z8�G�a��ϧw���.:�b|l1�K�[��Uݱ>���TUAf��'���ё���'x��+��r4��W���9 Z��`G�J�l:҃���-��@R5.(���{���~�P|Oǚ�t����'�o�|鶧�F��/e�g%��&�	W�DS�r�_Lq�����BUZ����Ѭ!�2�ޥ��5d�S���\�$)&Je��3L;md4Y��?�����/v��~E҂[�Z,?���˳ߌ����C|��O��]���P(W��CV�6�|ӡ���D4z6����z��W1h Jh˟�4�J��N+sL�83Q. C��
&'��d�(E-z��',Eo[$� �h���JtH�o�ɕhO� � ���W���J�g�|Tm�{G}N��()�H�?��ߦ^��u.�:2�|y5j�J��+���u����-���/��_�q�&�@Q�
���c��S�~PN}:�I�_큁��M��m��^.)�.�]l~�}Z!.�V�ثjN�-�o�pȨ1_�����ǃf�ORn����C� =��{Eô#;�K<=�!B����H���6LLs%�\�j�ۊ�sQJ�{9��	���/�t8.��&�^GhXi�m�q;�|��"6�m���S�$蟙M�G�����Ljʷ��2�
z�B{��9�p�U��(����i����x=������׊S�?�9I�y��G��7�/���-(�~�� \�^�~�ZQx] ���EU3�?��R
�"p���C�^Bki�(|Y��}I��Yo����
j��|��(r��٤EѤ�P�������� �g���1j��H?10�M(�5n��P�i�7������ݲ��}���ݟ��B��N����[
p��V�	9��y÷@hu�G�����'��#����A��ǖp7SMoе�B��,+4�}W�� �%��������$Yn4�.y&Tl�ӲC%���7ɂ�;G�-��N\>�K���<�>���f^E�PPЁQQ%iQѿ�o��\Ӽ��Ku*a*�֊�퓮Fg�h�a����t�@�kvN��ƣ����|pJP���x�W�~΍��	�s�W1C_��:������P�6}��>(E�j��F��.B�L����h�S}���c7�)��U�B�6	�8��A��ae5Y^v�"!,M&@M̹�����뽦c�����>5�:-,�)�9)%�5��k�w"��vڔyz�Q�>����	|�W�R�p謻EY�H,��U��v��8�������b�^M(xMr�Q����+b�u�]'(���4j>{yUiU� ��f��t_K��v����=氵[[�_�G�s���d�ր]�N=m_am�.���@ ���j�FE��� �{|�����uv}�n�2|���Q�pԐ��1��b���\�l��|�]mAF`GRC�)Ě������b�O��.���A������
jF�F����|�<� V`G������+?�.���?���/S-��5�HEm���@& �Q���J.�H�gol£"&�/��?����-3�������)37773������y����#ȕ������0��F�[G��5�6���ɑ���y����Y�������_Rx��+Ȗ��	�le�����Ύ��jn�`f�����X�l�����F�^o�do��3�l�<����HJJ�+��L!V�/����_3!&&����y������3'/�_d�#fc��g{�b�����A�y^~��p�q?�����	#lf4�2bedc34�d��d��J���dm����y� l\@VFNcncF ����݈����Ȅ��dl���E{ȳV�,���?P��P�� 0'7�1���nM��\�, #Cc ;'�А��؈G���
�|�+�)�����e���y�����Y� ��Q�9�</x��������� V`UG�y�pp�Xظ8@�g%�Ϥ�`{�g]���`bc}�s0�yf��2��7�<��`�������%?��?+�=,�lP� G���
`e�aa�p��y @Vz ��m�!&n�O���)�_b��8<�w{��˦T�v��jZB�j�����/@�`c��22Y������C�7�`lf3aa7b42�3���`CvFn6 ;77����(6&�. {����e���/�"���Q���|3��_B`dae��� ���b�����1����ׄ��?���_���2���K^������"�C�����!��+"��)������s�T:�\f��J��\P7��>�_ol�4�������v�t~�Dp��G�D�K�I.�E
%-&���k���uts�vI}��뷖&wU8i� a_����P8�f���nL�3��Ԑ�$N���V������V�:2�h��Ҿ������-����2٘Uzf��b�Ǟ0��rx�BΌ�<�/�|�^�}B���	�b>}����H�?oP�� ���;�M
��w����A��ߣ�"��|��^�#Uȉ�n�!���ovdN�^�x1F�M�ܩP�����J�<V���Do���\W�8ɲu�I����<w������}@����as��I��S�|]]���!Z��?!F�.[++;*�����	�asafc�	�-CV��b�4u�s�F�������.E�o6G��P�p�tQ�x0�hβ�"]���V����P����ӜY}�*�h��?� ���~-,ϑK�j���S�cUᒙ���-|�^0�t���*���9���g��ʲ�`P�} �ˠ���c�>���ύ�<��ͮ��rk�}�Q�PaTߞ����w=�o6i��/���e�؃@}.�a��ׯ���~��Z3�|�b�����Tyy˶un�ݕs);�� �?&��N�xx� (�U�r}�'���1l��,k�n<�^�0�O��Rw�?,/hQ7Y9Y�;[���� ��`f���R��V����ށ�m�q4�8�aBɦ��H�6�'�~�$��[Fvt�_���r<⿕�D�g��E��֎uy,�- JkK��`�FEW䳏�,w���0%YRW"�̎#�L8&�������+��|P>4!b�;N��Y-O�N���&�s`�EFB�E���)C08�`�2
�p���/(dcKV�ԗ�Z��^ҡ���u=ĥ雍������+� ��O=$]���$�r���:�qq���*aoG�-4�Ѻ�zl9�O�/Y�cl�3�~�{A��:!�Dǭ��V�ހ�]�Ö�X��� ��8�/��P#$���X����ܡ���RL^�o�V�M�=T��ї�R��0�x��19�=��:5�������1=�j��@��W��-cMx��R9r"��
�T�|���_b�;�͛�I��ݓ?c��_L9���}�e�J���x�f8�/��OX����������Z�g�_� 3˜ڣ/���ŢV�4�2
���n�����`@jSk��N��T18�|IE�q>�D𥑷�C�������0�DBR�%DcШX�G�Ca�Xc�)��C���"-�m��J�7MM暁��^w\��Cn�e/ʥJ,��t��rr:5>o�e��s�����zq\Rf��̏�g�ӵa�w>ᾱ��5��ѕ\������au�]�ɻQ,[�ݞ_g&�}6#��Hg-	��u ,��sو����M�k T�D%mC�QgCA���+4+��H�Qx��S.�>���6��UR*$�q�DI�N�lA�M�ԫ�	�����V�9���I����������]��i$�"a�è�Bd��Y����z���ko����z�zN��9�)��<�U�c���Yf���������M�3��b��"�����R�a��*�����ɯ�PY�R"t�μ�R�2�����N��� xA��z�@b�� 
�����,jAV�rS������꺃��-!�%�q�:/�M�l�Q�������1;˃$�1<���{�2������I����o�R!���"���yfF�8L�l%QFN}W#R�X��D���G��ܼ�N���D��(u8à����.��#�8-&
�[P2��[$+� ��?_�s7=�<� �I$gAw��4�s��(��J���&��v\�-����9��F�&��#mhɇvXg���l��xn{\�u^����6��F�be�w{ּ�N�Sd�\���xX�.!�kt��?��S�{s��W���=��-�L����p�09��8ڏ���=(�|��*�{I�x�xk֋֙4�P�c�H����6�
 9�v}𣈖����"��W�/-���L��Q�:b'q�u2�]���b��.bZ�NR)�UҼ��Q��<��1ZaLt4<�ޘ1��#���]��%B��E{�%*�So}hh=::Z�ٟ(��K`�+(�H밲�J�j�������<�I=�:{��	��y��;ɔJ䮬�Z�����U)e_�|A�����&/��g'V/H���ذ�-�[0�P����J����
 �Јe�♕VZ&I��YD��TZ�\�ȁ��Qx:Y-k����f� �� �K�y�_^�c�=�\���*'�T!�dk�n*y{Y��3�~�ܡ�%��9{���9ϴ���XZ�u����$�0����EՉWBa���)��&�L���k|>�|��Ax&�=�S*�����sݜ�g$W���x(s;x�"�c����W0UB��I����H�M�4}�ི�B�e�-�RTUw݁��]�JY�r�:��~T@#$�N&�H��I�Ty��k��W��B��&��V��cI�t|9B�}\r�0�����*���v�*y�%�3E��~k�Z�ۜ�|s��5��U(˒����J;�&n�ǒ?�n�c��^�����d�������N�$�fQ��Z��$=\h�xǙrx��/C��ӻp	��h����>����|�[�� VZ�;*��N"���g���Qv�"�49
��~�$��?���[DL�0�������b`�M��b(�!r1E@�#���<���}~_�#�v��z"��.��80joԼ~�%�c�k�3�`E���g���fS?�����DG���қ�%3c��{��O�o�P����"��s Q $�����0���y�U+C$��ڎ�,7���I���໫q<4����/�N�Z��K�N�7�<d����V�Ћ ��yJd�z�&(+"\������ h�5@����1;\�a[&	��g�_�t|��m=?}��q�ޫ�Z��=u���yQn�V0a�T8��B^uH�,*�����0�k $߿��G��e����Zb�j�k�$�7���02�`Bb������J%~���T�d�kG�ېWȼ��z�(�Z�=��FE��ԭ:U��5=����3�������E3��d��)1�jDF��")��CR�{��	f�Qb�]����Fv���
�l�gvV�H�r �X��TۢI��t�+S1#�MޤGY�c��r�B^�_�<��6��Ɵ���Ѫ��T3���}��o�ozXY��5��,�<�?0nq�������2
-|���O16���t��Qf��<�V�����[�A� ���~���;�ߏ��~���^J׈������-�a�61.<��,��8�������M��4sV�r�13���L�0R���D�G����O��dJ��"5~B�z�Ӯ����#H�y+�t2a����L�����yV��^���`J줅|�y;��i�mφ�]�B��-m՝&���(M�]К�Y�,�U ��aD唐aP|���Ņ��Yz�|ë�3��[):^~oO��I��_��޾���0��6�YS[[��]Br�}��?{w�.���b�"�ש��W��$x!��Irﻥ�D�N�H+���y�B�^u��j��1��zʐ�p�|�Ir��ظ&g){Ľ��;r�(�Ț�O�2D51!�iR�U1�P�Ֆ8�6�Z���]W56*�m����������#�O�j�ġSEQ8OPYW�s9�o�E>�/Yj��y��Drێ@��s�b��s�#�{���<ԙ7d-z6�RJA�e�x���w��ī���̔��{�)�	<���s�Q��˞MɲG�I�ʌ*���Ҭ�9��C�`g����Ϗ�bhA����6�ju�C���@���Ha�E����ph�]B�#%��[&F�ڡK+����L�����Y��Ǟ��'!kI��P��Ej_K�z:t�[���a;>SHu���E6���i��])��V_"��e~p<�G�'�?Ηr�P4�䌸��F�U���⏽HzO �a\�y�L�\�jG
۞�<�NT�0�{e=�������އJ��y�jkk�796�(Q�S���\�E�i$Dh�f��L��t�9�(Vz����t`��+I�5�z |�F�,�.>v}�W�_���Ͱ��>rz�c�;�1d�x�IoϬL����s����!����5saT�eK/�}���y��A�@Un0�˘�sX�a�z�(�\�LX.f�%����V�w˅��:�B��ad�1n��kH"9f�?0n;�;�W����|T�2�-H���W_ɀ�[W�3�Rɗio����t �Z���H��5��|�s����JP�R`��?!B�1�B@F S�^�������Ƙ����$<�d��F���q~��;�-��<������%�2�e�������P>$�����I��A�o��М@BU�;�.���\��e��`B�B����n8����R��E"�R�E�ĩ���8����ω���Y�=U`��p�ˑ^���j����������	S~� �Y��q����]�Ѣ�l���~��N�3ʝ��TeRAİ�u�@��)�}��ˍ�K]~M��s���zcE�v��No�W�����}�T.�;pR�r�6��ϗAafŏ�Z�Sӯ�O�=�,���:�VV���kXN��z��J�G����/�^��3?o� S �戃@+w��U��d�١��
N����A���t���<e����o��奄:)������j�s�T��X�nteK�E�UƧZZ�-8��ߜ�
�����R���X
߾�v��?�q��r�۶�&
\k�$�@�_��]!�P� �RѢ{�U��9t�f��z�]	�"����hh��8"[�t�<Ĭ��ϵ�e�V�O�73�|{��eo�cG�<r�P1����s
�л�p�8�t���^rW��fj#X��].�BmL����>�@%�=�5\�X�0I��-C�W�FK�^�~�y����m�Y���f5�ח{��j���e��z��tn�d�2u��p��_;�.+<F���Li��UB 5�Dt��v�"��	o"�>�m)�\9,iP���Ѐs&�AhZ���K�}��{i�F>pE�6��X%�/��n�sU ���P$���Lrn5W�%ҧ$��D,����l�h�}rH��s�m�����A,�\�K�-��ᮃ�����B|֪��ZUK��3���q�i��J�CO0\�T�b��}�䪋�k2���IV0����0�BwR��m���Jt�,ٟ�x_������m�
Ϲ���n`��g���P��eo�!�LǱnh>w����mI�F��t�}��F���Q��^3a���ݶQQ"�i�r��A�x���ލ��i�V*���6{�#�$��[��u)gAc.�˽����:����h���ߢOJ�̉_��jt�:�?�tu����ɫZ�'�>�mvB�[�E�Ͽ&���,2D�~�!��Q�ZuBo����Zb^���� �OT��a�k�����6/5���(���o8�2�O��O�qw��U+�`Ni
?f��b�!G�3JJ�|O2y�,�m�$��q/�R�����0�Qvm�a��f(+0(����P�EEEE��)Z	��>�vT��`��Oy������j��f��>�w�5@},�#�(�2��D���\������6�_Lk<8uk���I�]S3�#����rMU�oM��&O���TGF�tz��$��F{�L�
*Y�3`-/T�}i�k�b��n��{�8d�?�������P)k�����`��Q�PV� { r��P��*}��N�?�J9#*���Ym0��i\�yn�=$�xel8�Rᖭ�4w"�{v���;V������Y�d3��DH��C'����ot��\�.����'��j��Z�zI��;�Y�Y���dǴ&�|��+g�L|�a<w�oI�bp_��Ou����� ���	�N{ J�S�W"�n��N���?n/%�!<$&ܿ4�A�H��cƟ�#E
H�������>n�®��EjY.���7�Tl\GE��G@���vBD!�]CY�F�-Q������F��Cj��@wl�L߾�Õ�r�Q�۝�^�50��������8r���p�L�$�)agߎ��������[�u�~���rD(�Z]9v�8����KY�^`OOLSQ`�����L�K@'@{w�*#��U�L����vW��ǖ�o��_������aҹ�
� c���!�:Q U��*/e��=\����|�6�~��ѣW<7�.m���+F��ʖ��I�f��0����f�C�O�D���}��.��V�nӏ��_��}����������r4m(���.̾�O�E8�Co�:�C˔�NK\�.W��D��ڟ�Z���g���a"��"h��%d��]�
��l��Jsy���+��җT
@쿵��C���@/�x�%ϩ31�{׺������j��a��$��[���h�6�J��{(*� "���*:�Տ�[�r���ջۦ�VQ����c�L����7MVj�_,P��>�%�8��Ƙ҂�7�B���g��A{���<i�A�R�G�� ��Oqß��Ӫ��w܋�(�7�ͤ8	ǭm&������sv�깗�ro�nhl���cXr�p�i�B�j�I�Q}������K'M��՝��<_��tK:&���q�Al+�ԌZ8��yq��s ���{�1�����id�y����i�@�?�ԙRB��9�'q�.�,�xx�z��F,��C4@/3����0�ʌJ���3���Ơe�����B���h��i>CV�-��ѹ?O�6ks��î��Ue�[q�<�RL������_��V�р�vj����j���޹������W;j'c�������l�-{F�����΃5�e��20��	(4_$�`��S���*����W�t���#�U+�.Z3l��#�ⴛ�r
t�SW�g�����픍�z���ʾ�z��p�B����M�ď�B|#�g:�z�#�4
#S��=�ˏT��i��KNg�S�Q|_��e*�1{i[�+�W`�쾻= ���ߓ.�֛��x��`'�׃�%[���-WR���X���4�P(zcn��J?Va��r������t�_���?���y�yM� P�v=7�f��m|F�̬�rI�H�IT���1X�Y��W:���?heV ?&� �T�L�r`Ӗ|��F�qO�|ƻ\�z�x�cԛ�'�N��E���&]������1볌���si{%���z�p�P���R�d�q���~*űˀΊ�����g�4
��t^���8#�� ���W��a��|Hx���������i��]YC�M1OA鶵M�ZR�^س�rh1�w~ұ��vk��AՌ���=�U�#O$�u�3�����C��|Ų�����h�ҟ?bu>F�E��g��V��#�muzja qS8j;����Sq�UL#�4�-U��%,���t�r ?���	e+e�����WX�.;�F&΃��쿖Iz�_�<�_��넺�V
{�e^��OlX}_���)�S�����!�R!��:����0B��+�i������ckh�vzc���s�q�(�m �~����O3,�b�d�\�m� 2���üd����B����Q��a�ԓ��_���nWc|T&�S��0�[ZLln\�x��w��-7 >J��r��� b��Z#g�Hl3@cD�cN<ո3A��XYp��п��o>�K9Sg������A���]8����\(�#�b�\J/�5(n9����]ƹ�~g��%����Vb����Q:���Z� Nvm��~D�G����`���E�x�]v�F�x�>��Ğ���/mu.2t�N�m�l5��I���NV�t���]g|�3�CX X�k�`�����g-ZjW��}�2}���G�|�3x�H��>B<K4�ﬡ�l�%#���	~7��E���wb��B/�}���E���徦
3��W����1�a��*���X�f���Rv-�*�创C�����ə���w/ ޻�pzpq�XꡲÂʊ�,&@���P1�@<~+[Y=x� J*��.B+�xNW�O�-I�x�p��D/!W}��<C��Y<C��ڪ�z�2�9 q���'Y�����`U�_�{�y]5�N,�VvM��Dy>�x��u�I��u��	T�B��̊��O�ē����?jV�W�~k;��m�Y;�D��D`p�#����T����x�ގ!��9/�`%2��	_4H�3gBC���G�\�G�/)FOe�rMTn��������
6��� ��b��VnX2N�SS�=��ޏ��.�~W�\m��ψM�pluIJ�Ax*�3ɩ��:LFs�Z��dԽ�HߏǕ��,�$��t.�·��s|�X��y��q�d*�|=+ �h�V��-�����+��<- �S��E�s]mC�'�V(x���s�i���1p�;�[>�����;�� ��M���.R��P��99;��[rXcz��X��v��\>S\^ZMŭ��j4�#w�w�z.V�HÑ��;D��6p3���^^���q�dK`�"=�����W����n�h���Tx��8����a�[�^9�S�� ?sF���W=N�?��D��7�x�M��G���q�;��R �G���hЬݢf��MSq�.��tk/�d��V.���\�Nԛ EY���'��} Cj9X��@x�����l]�+���_��irۛ��\,z����P3N��	�t�X4�*�8]���5ਙ�j�\��Ș�����üW�qH3Z"7���@����Crۣ��[l�f��2����9�9 �<�<VM�-zQ\�4�eX���g��>��}���GŶ<��6;��Z�+�z���m�b�����:~d���tZK���d5���IL��K#�|m���o<�N�$i��������cfJ_�N�<G:�x r|��)9`v�����g/�d�ozN-x�SF@l�L�,1���	88����u/�CA)��<��R�R_)�M�v�=X���.�,����U{9��Դ�!�+�j�S��	!R���S�+�D]v?���䰎���?��7����e����G�c�+J*V���\�������2Ƕ�.��0��x=,V�ɨ{r$�8��BƤJ��*�s�VpHv�l*YW.	�K��׭�!Ljne.
Y��N���.�L�����@�%/���Ϣ����"�*�IF}6��o,�����F�_
hA�"��
��'�ޮ��/I�]pT��d�K]_Zio�\RB����T�k�Q�-�D�6J�c�.�|����ɖ����g[L��=���8���5f5�搡�Q8a]�꜡W8h�ƶ�Vj՗t/A�QŴJ+_+��ޝ��g����zc9ޖ��i7�Ƕ�Xg�j�u��S`g&?[�˃��o|�)
%o$��_�_2i��JFN,qI�"n����;� ����5C�Q�|kњD�BGt"��^mį*��yPj�7���4��_Ș#)�"g�a�����A����6�.��i��+l�ۯ1���c���f�}��}��N�������4olo:4ͱ�%c^`F*E�߾�s�)�}W��K<��t�a��b]���ȑ�,�Ts����Ċd���vTn�!�u��s��T����6�Y�����V��������u��6uDg�v��CU�'Ȫ��z�5�TK�h?0,;\y"��s�$'/���xL
�L-�!�I!�����0B�Ğ|��X��;�0��Kbq�_
�E��#�eQ����*����shH�4ގ���N*7N��Ȍ)%�-L�����Pg|�}�~�t�R#c����Ļ��qywp����";$-��ʺQ�Q'W�lMq�ၱ�����ۧG�Ky).ܧ���	v~� ��]x`��QLr��e�gp
^y�$M�����I/I�ߋ�Q�k�=7q#m'��a���c�!U�`�6^�K`�8U�D���r�����`�:���B�O�U�sQ��Jܸ���1���k�
�yy�$�>�M�I���.A�s�57����{/ٝ1��z��0=��;ak�Z����|�/�vv�����v8F��v�N�U��*�l}q�Ү7����"�F�\#��x"0A�5.��b��SZ\����.�bC �Jw�ƨ���y�ZzI�n[D'���l�䡑�;��/��[:A±�wߑ��I7@���޾F/�o�������z�S�\���j��F<���*C��y qAPH�d��.fg�LD$��E0n����K���q�������\�0~2�l���I� E~s�E9훑S�^N���,����|�J�ٰ�}�3��b/V+�ެ[yn�|��t�ly�Q5l/��n����.)�
>_[�L�X��^���W����r�_��O'�܎�h[��-��F��!��nvb	��]�49��~N�$�:��{�A]�}&���M*�v�lt:����ͷ�S�A	zN�pت��p����ˡ��G�
o���9]�FT�qW1Nwlv�Oc��Pko�"A_>y��
���L�� D`&�̀����*ۨS�QU�pZr?�sP�1ܭhtt�o�����|/7��g3�mF9(B+'��:���x�zd��͟�[9���޷���.���%���Z/�TFY6�����{���+\{�fN��,��䴔���M�<�.��o��߅��u��{9��c������er��	T>�A��Do���)��������+�h�f��t��IpwMp�@p� �ww�%8� ���ˢ����/�y�����N���=3��ͥq�0��j�w�~�͕��ó9t'��U:9w2�'��&�V���.u�������ݷ�� ��-Gx��?Pa&k���8�X}���OKO5��A�&��Q%�tT7��K�,�pس�,�E�=qL�������゠"S&�D�4$H��5�u�9��g�Q_�A��;8�w�%���Ƹ�����h���x)b:��d��IUu�5&%r
�@F(rC	�\^#����
:��a�aUŪ?�T袄Iy�4�D+7i�i&���F%�'��d,���M���^	^�
�Ɋ�S�>>�=�?o/�wخ֧��"��bb��s��� �Ԗ$Z��/�^`>~�F����|��/�����Zq��byeZj�~�
��W�C�/9:a0k_�����%/���N�����O����wpϱ:Q	U*�I����::���冺�ؠv�`z1�n���VWO�J����|������qE�W�6Z:�(2WH�(��-3���*����2@�jU�h����}����)������|�,##���piDx/ԙ|ƨ+B�2N���۳��\,�pX�|y�Z�U7fb!= C�XR<������s���e�P8Q���8C��������?x���^�^�ɼ��GP�S�Se�I�@Rx�`�׽������Y`TbԠó��;��j{\x�hU��n������ꊱeF���P�]l�N���g��4I3t��<���a���Ĭ�w�R�p{��A2�W�t��PV�S��~����Zd:���TkBL�����{�/G=�_[t�n����γ�S�p[�W�C� ���n��E�`���^�y�Oq�`�C����G�{y!�R�5����H2:�`�l_n���+�\��\y`�inRhdc��������\=e�ϺU3��)�ɻi>[����β�c��O�߄�^��Mtٽ�	V�_�T�Ld.<�{���L����ˢ�U�֫]���URe�X3�2�H�>%�Y<K��i����qb=�f= �����NN����Y�u1�E#��� #�Z����x�6Kh"(��h����C��O���6ٛٿ9ՅU�.����*��(x�Uk��	�|p�5Z�.�u�ty�7_������U?�_���]�>C���a2~�I�#J-�ʆ�mJ�	�I3�/�f7�:�_�����S�~�F������U�`~�R�5�ÃH$HԆO��O>е��8�WV6�v�X�$��O��i�d����,�欚?E�-T�i٫5��*��ML	����g��w>�z]�Ӿ59hI����.�{@�M�j�	��x'�0�|�"�����8�ׯ�2B��vL�宭11��h��=p��'�#Y�@T��V�C�* 꽉f'��Z)(����
5��K-�Κt]!I��.mοK�3L�����;a2�':d�������lS�`����
��כ�5���0 ��ڜ�ʪaB��Լ엲���3�)jI���3���q>��$��H�� C�};PY"��Zy�ns���ϭ�Ͷ=m��o��ԳW<F�^P������=[Ov�D��?������/����߳�1a��b��  Г����;��kmHe��tѫ�06�_��f�m[�I|S3�Cl�t� ��J�86�Q�eL�^6�L��Mii)�6�P�PղBʴ�v%m���G�q[[�"�u|k ����$�!���BL5{]��,�O-s�H2��~]����w�\o��)O��N����C+Hv,=)��V�杕d�A��G���^�r���q�����(�H����" [��P�����T1KyLX�=lZ� o�Lb�%!�
�����ɦ��W.s�\R���k*ޠ�ٜ�"BM�G�}<E ������Љ�'���RH�AW[��x0�t̳�f��<N�B���b�9GxI�7���s~�����⧫����DK���x�+FB����]Q�:_�����*Ӡ�G���,}��)Pr�z���2.�$�&�z����m���Rl�ܟH��.;����%aG'��ESK��ӈh�qL+�H4o�|�@��E�F!:���=���7�����t!��İ��v�YCI����j ������"[h��`i�%���ɳ�A�����A� /���fdt��S�"b���E�;�n�����֙��\կ�e8`��6WL��W)a�@1��D��$��/��ݝǂ��P��b��-��uA��pyp�Aw��g�.KU�)��ֻ�Q�h~���4Բ���3H�Ѱ�P��^�g���S�?�Z�ȞM����+;^�}�"��"/_�q�d���W��;I��#��(��^9�ި�?ot0m) �<��=׵uE9^�����F��\$
����'�-j������9����wzn���3�k��+���v������3h�� �$ c�J~�X�ƴ�m�����EՍET�!ƋX�x����k7oo�4]XX�ݤ^�����;>�lfn~&�c���\�+ﺿodL[��]J���߄��)|$~��-V�w��C�(M��z��6&���[�U����X�/ރ����*�O�^L`M[����d�+/m&-�%j�&n���u��?#Y���K��(Ղ�OX�v���h��b�*_�[&���c��Mj���������)�#V�A$o|�3�:��7fd��d{n�ymQk-8O0@1�!5�m�տ�/�<�e�~�Ҳ�wڽVuB/W��$�ob`b��.�4��~%�Q���I���e�PA����>�[�L#?��U��x��D*YDM��n�mw�P'x�M����F��M��,��VEE��D�*�H��^̞J<�Nk��+�z����K$��!��*���h�f���ȍ��E���uĜ�(�c8@��jt3�1��v�.T�$Z��.�����.�e��D��t�YJ� =�$ P�_�N�>�E�!B��_%ް.��]`4 N�����\��`�+S�����g��j\�R����\DF:��i�$��s����s���ng�2�+�vh',�� �P��B�:do��T�}]�G
H�t).�e�S��rc�ex�ձi�~��M}�ɭZm�c^~\��(Ʋ�X�Su�S�"�JЦ������׶��J#[Jሂ���O�v�+���-!��r<����C_�������}'^���ϓ���қ����󾏼�S��/��ٽ����`�G�%��+������Q ܆3"8C=�@tdϑ��ga�
N[_ͺie<p���.�"�����H~;��X<G��
�OӟD8���ftp�f�
E05�6�m�g�[)�L�E�b��#�rD }�?~���\��23@�|�!�!)�gx�ku��?��|��.���У}��pT?�h1����C�|nm��x���ЋY֌"%��K����"���#�|�Ო�0��Fpݔ��aJ5>���A����{F1��£��|v��a)��.�t���ל0�x�	.}�r#p8��tG*�|�6�+��F+�����m3�K䨔�+���<����#�&ɬ*t�u���$y�_���Som���QW�s� ��5�|��.���c�yn{V�-h�|���y���?�(/�s$�P�I�A�1�P�K����-L�W�X�H�C��U9�m���[��Z��e�N�c'�>8\����9?��0����*`_��D���Q�K��uM�­VcM��!x-�Q�P�O��3B�X�r)�x�q̶�띶ؤ}BO<p���᲋��!��A�ӏ[�5|?˝��S���_�y�~<�%����u�>��R�az}�L��(x�4n��qGȆ��{v�<
�4�� �������<$@��9|�7aJ��*��F�U��D�X���@�>��S.�M�/������K�NL����iAJ��hK�m�A~����d[
�����0�8(�,I��j���BO�Ͻ{\���F����pw�r3k`�R}���o�}X짊
�O��*Q05jW,j��ß?����6^�E#�Oq:�d5��sWHb3b���L)}��ڕt�+0�d?�,V�*_�
,�t&	Č����y���UG�?�=�P��{����"��������>�_Yo���]�W�Ҥe�׶=��e>#k���T�����93��x�X=Ӕ�B���#��ݑ]�Vk�\Y�*)��Z2d�T����'��j�W��x��ܚ���bcPxV���c!K�=���T}l�1]�/�Aޤ��I�͒�c[SO�y�nڂ35D|�A\��36,���$Jcln�Z��j���"�豀���r���|d4�n+P$��-��[��թG6�j�F#)�S�r���\7�d��s��{1�
�\���H3��C.+|�>�^���=�ۣ}�[]ٛ����V4h�/��YaQ���{�fz�'��a���f���^W��Θ����$$LCA�8-�+��� 5�^�T�8��9���.KP�b���x���m�n�qmқ��uS���g��sc�mSp,��[*�;�Bk�.�*���������@��������e�<�`ފl~q�C�R�&�pA�dBBBj���lR�eL].(V������3k��-��NM��>!�e3���;�֫�l�W�|� ,�&S���{�����	y(BS?��󉯊q����5S� �ߓd�)��/�a1%�=7�_1ȴ���38���6�SVA*%�;���RA��T�R9J����QӬڜo�viдky���?Lg��aso!-O`��b�n���T�]aX�j��ͬ�W@��
�QQg��?w\B1�@�v>u�@1�+K��f��
q	1k
��WD�G�ps���ـ���\����߭��v`��2�̄ЅG���]�-�*@��`!	�!
T	��n�յo^r��$�+��|��[��6N�`)`��U|��N�Gm[n����T�Z���G$���S��6����;�,�xa��~%��|��.`�`� �ݧ|��Β��RXT���jb{�ȝ����x^/��t�s���i��@A����u�C��Ð��x�Qz�������g��I=nx)7my�N�c�vN��yv^!�>��u�t{r�Xؔ�Sq��M� ?6���-�����xS�d�	����㪩o9l��ҽǛ��s}�5,o���)���s��*�R�T~�� U`$�7�k����Q�J?�9ǝ���Nu�:�i��vy�_�l�<	���\$� lV�*]K�",8:|I�tN�533n+���C���O��9f�]�洣[nꃓq�3K.Ő���{)8qWg�!� ��5�>�m�o�?��dؽl�|���<����RLp��¤fm��Р,��F�d5I�:ԝ�;?ĥA
����Sl�1�y��ss����E��)dgg�i��h�=�݌�;L��-�.��5�D�Y2�����sz/���r���c����E�eJ��-�q��,�G�d�tp\�Js�r*R�N����-`�rN�]�E��^u#� ��d�>�+J�Fn�l�V���sBT�O-B]�!HT��0(������#�QLЕ�L�>���K�v�ϕ���m�7c�^�g$�t� q�Hi��'�0`��	MzW����
��FP�ªEɞ.Jj�z�p�9;+Dۙ~��2�S/
caa咮��}g�����߉�0~ܢ��_�:<�(���7w1J^��]*���Ǎ��䠒5�ia��ϣ�����y�����sg�������^R��#��`���'��SJsfKJy� ���{g]��VZu��\��nj�J� �+�|���
�Zd��n�dFrZ�&�0�Xq�-,���K���(���T�@%D�~92�,���Sf��Β6=e7y�7��g�zvF����2Ψ�e
!�[��dq��Es��s��	�٘l����Ä˺��{�i��|P�r>�r�����\,C̀��A`��׽aoO�������M�L��<�(����æʺL�z� � �{q�wL<�`�=:Y����󬯭���
�ֻZ�.���iLɻ�>lTd�z=�2j)x�E�@C+0:���s D^D�I�^�(����uvr\eh48oyB�݅���L��#8 �%�(�TF,W�*��Kz�x��f��v�
��(����/ZYx-�	<�y�a5�����	�l9�.�q#���)�M�� .�#��c$��4ʝ@i��x�ʯH�
�J��p�nxX���gDKG�4}7������������y�&�=�>�5$��^:�k�%S�@j���?=�Nc|!0�1{�_W���o|�E�g��ވP51�(=�;�ɧ1��%��yFNcr<~�v4x	\�ma�WPp8^�sHP��Q����E�D��7-X9q���R�qc��V���CgV���ץ��]�kk3��ݟ��r?�����04]��(��N!��9�����7�j���y�	縆�M$��I� ���qҘ�T�q���� {f�ꋺ%��7 �z���c���ΌG�﹐�Kf���#b?��{�К���1�n>?���n�ލ�}U�>ሎ� .�@�1F�r�� e�H}��<��1�.�G��jjfV�t����IZCXگ�������\��PY4�VhO�~LY����݊��#����k�W�������OݖU�v��o3�rQ���U���(��""\���	
ً!�6�Y:�p���'����I�G���G��bJě���U���d9��4^���z=u����V<2g��OA�TC�N�x˦�����H��Jݭ��.5�̱&��Q����I��X���(�M��y��u�^���t���a����^�E8��R�rwd�z���o(��Y�K,��E!���dd� r�5ߴXp%��?�h}ν��i�"��D����)���S�;F�d&R��h-me���}���i{�,+r�5\4L�*~^���V������9����A���M( ���/L��@��b��C��Ǽ��X��5~�G˱y��*| &��Jv��:���xӉ����V�@���p?�Q
[ݶϸ�T���NV���s����f�j�j�Q�����b6AVK�ЫV��(T�sT����ƿ���7���"�j�C�n@�4zy`���=!�q��j����Qe�{��,�ha	����6ͽ~ip�	8���
�Ox�Z�*n���ظ�����%�t��O��mW�O.����I��7/���UG'�>�ɇ�e��2Z��L��,Zi��2r��{eu���+��׷�:-�"����t���q����񘦬�=����07�z�īk�L~v�Wfg-�
н:�)�����ֻ�uxڢ�KN�s�d��⋱%��5���nʴlK5l�CXE;r�K�xл�buĊ&�xPA y��Iv�:�������s���ŉ�͊��z����n��<�������-b�|��ZS�ov*؄����e|b̘��1�S�.��_fU���F�	Yý�����o�a�u�
g�=ͮ���!�����1�KSv3���k���ιwe�?�x�E��:j������:
�P�����KC�|ɯ��<7<��,��j��b�N%�@YNo�G�7�|T�}��8�f}5�����-u��ˤV�+��)�%5[{�����(�ry���H��sv�� vK%ɻN2Y⓲x본{�rѻW��t7#Vns�F��X3��]�y��-C�[ְD-��X~+���f�X��>`(1*۩���*_Ǔ��H����^'���x
ˁS��BA��7��D�"S�/���GZ�1-)ݺh6�<�D��(�Yw����0�������t+
A���u?IG��;�G������F$������<M��,�1D&+ww�I�@��D��)���I���878\q*���0��g��%�1��nL$��9!ѕօN^��s��t*~T��$����5�=��qE�;z�$ufoBs�!F�.��ag��:}^
k�1��T�A�=N���s&*V��4��r�I@so����!��Y��� �V�U!1�Xs��<?�cf���û���>��ubs��&k�m��n��t*9�@6�e�xZ^���W�aWpUj>���|���Dا�"U����A�4��B�0�I8m2S�ChE�t9����_*�Q�Oǆ㰵O2!�H/�:��Lw�oi_�w^�~Ie��~�oari��~Q�M�o�7���J��Z��϶�_�
��O�?�� �P��s���#n �c�Ǝ��g4uW�!h������wР�϶�L��r�!�m	��e>�_~�\����Ǖ@��k�v\��Բ�03��	�!IZ�D��u���+X��w�h�G'O����|�D�_˿��h&/(�c����b�b��o��\��Q�;�b�sK'�w(6~���b>"c������;M���N�UN��©�9��r�Jc5���a��k@�-���9����o����N�`�s�s�vr���m��
�<s6|IJ�4_�T=��X_�R�)�^7�.\*�m�!�p� ���[�t��w\�w;�ï�?��.��}��C �!�Y�'�r�ӰJ�vnT�~��b��A��x)�i`p&� �VHeK*GB)O%N�X34�ï�7�����)�_�KG��0�|�*�U!�9�L�x�h��{H���6����9s�VwI��r�P�0Te��j.j7�����)���3�1_�຀�H�>Iq�1�weà�`� [���4���Z�0�Ѷ������_r��\W�\4%l��S�B^�M�cA��M�x�~�����C�z�w��VQ��I���� �@Y[g��Ҫn��#��΁��|��ǻ���Z�����`V� '��	D����a<�C�K�qN T��B��.���u��!a��:���$G�&/"�}"&"vpW���H��pސ�v�}��B�0I'���Q�T�� ���CdX�)?�R�s�|T��Q�"��v�ז�zE��ݼ����_�Y6,��X�䭷�@�j0O!�2(p ��E^���W��������Y�3� 	��Ó*�n��%\��˹%{����g�͢
g�DG��OM_j�Y���8tϯV�%�F�ھFb>ɏ-ޥ:j�W
��{�+�ߌja���R��rCxg{~�{ڂ���I��;\b������-q����}j�ל�Zy����[���CS+�`rD{�0VxC��'�h�B'L�|%Z��tyE֖D��61`,rd�TT��Q<���:A���`��,OS����Z���#�r]����i�Q�;�2��Ҿ�i����Z�&Nri�*@��x��F`�-4�׭��)f���"@:������a��D�Yu�F1��P�G�_���ptZ�̾�b��pʑ��a�����@�-!1���M���ƃv��U&C����������QA��KŪƅ꦳d���*�mmJu;��TD�W�K1��!I<_�T��.���Oe���nɑ�����y��N���(���ۓ��So@�����Cw �j?�J��Læ�L���_�5���-x�K��S,�h"��r�����gM��BZ*��f��v]A��|SC��=_��KECk�`���7N���@�D�>�'�HLt:\h'1�'D��5��Gl��l��	�x(���2QkѶ���b����ж��Ux)z>Y�zҩ� {n���c�D��@,��ꦻ����[���=� �5�%u�h���[�D ��k�@�9��$��ؾ�Ǻ���˝���N�c'���'��ܥٶ6q���ᶰ]�8��Z��p�e;2���dM�51;&�v��C���b��A:-�Յ��\ e�����"��aXT����ףQק��z�R���� ��T�ʸ�o��=�R���f�0�:�Аk�-jm�ْ���tV�Შ���L�`������(B��[~m���祢�~ܘ����pH�Gn��%�y�����)��'�6��On�"(�G�/�ՙ_ͭ��/إp&�jT`Ā?~p�x�l`,C�
�G����][���=.��u����h|���DT�	"�M�@�o"׈�8����8G���e���|�^fn�+�=o��=KF�������7X�����sU�$����gf�tr�U^!SEJ�(@�r��:]T2r�H�%��)J(�A1�<Sy�+f!���5D-���P���a#_ ЭT�	VO��G��8)i�x������Гot+�WW��gf^̂���/Lz�Q֯n�E
V7�
>�c��w6Q^�8��k�@.V��rЇ���hc���'9��U��T�x*�������
��N�Y�b��^��~;TD ��%IP�� X�@-͖]��(���R���f�L7ϔe��ه.��j��S9}�:_]��hJ����O�2��&�!��,���Y��{{�_�ɞV=����؇�K�ӱ0�}%��%��.j?��Wz~'C�`t|��U�#
��X��7�3rt�Ə��)��,��D	ٰ���������54�:;����J���T�H��P9g������OӔl��t�C��������`�_�Ju;��{.s}���Zg��
��y��e�&i��\@T�g�9HN�ʈ����g�R~v�L9�Xf��S�B��+�ǜ[["�v(�`Ok��T�0q�Ŵ�Y��^/7�I�^6	�s	��MDSC.�a0f)�����#�Cl��.�}ǽkxi��%�of�G|Tҝ���m���ѿ,�߉x�n�!�ǵQ�4O�+��ƗuX =�	[�K$�Fi��x}�����l�.�����bG�57!e���H�Z�G7�=�X��3�(
rn�51v9�����ɓq�oJ�0
ټ
��	s��-�ht�ҕ?�����N��5���vҾ�:�&���鲃B͕ܩ��nYEU���mH��v���DV�YՈ��a"
h"D��`9-����$�D�+Y�����u���t��W�R���J�qp%��#�Z%JX�ɫ��`�!�����:�*��9�n����"�@���4�h2Н�����^����-�Y�C�X4ը��J��+="� ��.^@�UsĞ�Q���Ӿ!���0/ps�R3mǦu�w���l�;n;1 9n���"+���P���:��#���S���H4%j�����d�K9��t�p��K���H�o/��nSp�.�s�+�Ns�`H�u�� PS��+�Q��?0�k|B��j\t��[!%���(��e�����ݕ�щ_v�-_v���V�6ȷ	�l"�9��lJIQ��`��d����t�rnh� ��:XƉ!I�d����j�����G�ٹ����a��՝��k�fx=�9�I�!e�&�7l!4��j�,�0��z� �瀽/sm/
�޷z�#1���}�����),L���� oS�ϥ�}��Y 9�ma�a�٨�M��Y7R�^���W�{ӈ�,-�c�h)��8����D���&V�t԰�F6Tv�Rk�lS��_[�����J� �S:<��ih�>zu�ulᗁ��0�;�@�j��?�盀	�X����X�u�HV\�pJ�k�s[��Wy�;���h�+��X��:�͸�Ợ�ΰ���e�X-�2g�*U@#/*{.@9Ė���:q�H3��X�Y �v:��9��Klm4��u��O9�7Lv�.$����p���޹IQ��W���Dq����@�+��˚�&�eH0Dd�X�p�@%����7�T�>-�ut���/�|�J{Dc�Q5�
���<[�m����0��������㥵9�����k�< ��^p�C�� �.@-�2�#��X�����[�eJ Df�i�$�Λ� 9FGϡ�����C�a�h#�P�M�	Pe,�����t���%�M��U��}���������}=���wt���[�:i�w:����3�{�W�R�qP�]���bg��P�[X@ۿ�k��6̤��F�G}g�~�d2
7a��:B�*�U
�\G�d�g	�d������YSNY��	�"�-��5F_ȝ[���&��[ԅ���,1�c<�J��`m�I�(��-}�+`�W "%fR�XU��hG���������7�=^K�ٖ�2r�{߾(����J�����o�T��[�;�_v(Rl�%�8de�m�@�9�m��䰱('am��KA5 �:�dxfR�gw���68JX�w����s;I&�4�I�UYk�A(Z�,6>�����t��d���;f����C�w���_���U�c>��rɁ�{����8ώQߘ�Bwu�2�s,�������g8�_Fڟ�����o��u��]���I툢��Ƙs#�5���,*�|��p�N�A0�ܝ�����v�k&f���`\d8.��R�_��;��B�i����`�}�p���E!-~��r�z�-���`9�t�3�->� I93� �[E%k��+6�X�fm�j�D36_>����B1�ŀ|�������݁1ڦ㿫��em��w�7�}��xk�e3�t�|UG��l�=��6��9�&�0i��0�Ƴ���%�����(d�<fk��ڻ.`�Aѥ*�4}{N5M$�FP� _D`X�����W>wf���K( %\�_��+�$z��r� ?����Ġ���$��?:7�,932e��WL�[U�����d��ᴨA0�V��̿1)R�mH.;����.����ţ��&����Q���P�P.���DL"�:S����|GV�����|&���ø�3��stϓ�i�Gt��v���=�����=�% ބ�036��q*j T--�@�sWt�|s��Jt�,n�q�	���B*V稝�r酈02�p�Bl]{�7D���Z�A���)P��)�����h3��B�����fj\�e�wI�7H�)��?�n4.��Cj�������Xm�a7jyQ�E"��) ��l�֟�'Y�H�m!G�8H.a�X%����b�]
JH���]�M��q4@�@J\��� �yG�Ҷj���bųa��c?�����%�~��X�`Qk�̣��"����	����Rc�@NM���ݨ
A��>��鿀n'`��`\W��a�ζ�g�^�x�ǢPK��&�C3=�[��mo���1H��Gz�RȬ��5�q��y�^����x<���ސ �|�2����I��!���c��m�R'ՠ#A�7�z/Fd|*��*�1��r=�Z�2��zZ�ST\P8���4n�%;��g2��9a���Z��UQ��.���"sS۰�0�����O�����t�%���`��d,�$9*������{(W��d�w��w؏�Jԣ���?�"N�ND�.n;:<�dH��7l���&�W� RyX�������{�ׂ�Hݳ���U�J�iI�|�Y�b&w�����yF[��-�?X-p�Q-[�u�3��)D{�����d�	���R9īG����=ԏ7�+�~f呣�����ѧ������7^���B�˛��]}��*�]����c�ڳ'�A�E�x������U�R�h{F"�<��p�E���jW_*ʿ=P�Q!��H�+R��ƃ�ş��m0�`��6�d�ɛ��7���=^r�\�=�
?z<
�����uEBz�rBd���8����ڨ/�)̎��Mwc��߷_z�������Và��eZ�� )�xr)�D�?�Mf��/(������K����Sח�\cH�X!�*��)S�����E����K�@�.����oV��&�_��!�)>���?��x���g�Y3{����9X�F&�a {y:^�H�n�x��0�"� �"��mm�@��k�=�}�R��l�8|q=\�TC���P�����#%|P� �^,?a0�^�n۟���'�nR��ۚ��7���������e#S�����_e����Ã�Ț��P�gߛQ��~fZ�(��"D������p��$���x8d8,�O��h���q��e� �O*E	���{�nl'2��w2�}���{��Y/��[7���9�x��c3��
�a�����7�V%*Z� y���7������R�]��VpήT:5���u1��/p��@���z�	1�/D��5� ���>B):Yl�Y���n1���s��}��h�'k�T�v����pT�B:�y�0�H%>!Q$�,0��]��;(��F@T��e�/�9�.��|>�o�u����~c�8���:5��XP�b��>�H�$��5R	9����x�2@2m��6�ɵ�}���j꽭^S��>Q

�/���5�in�_�
VN�w��c�����v�t!����2�y�{D8.vbH8��f.��E�����}ai�I����IK%U�Ű�ؑ���6��o��W����i~�P��vX<��c��s��!��/��-/cP�Ff���m�5"�����B��C�Ѭ_�o;0aU���*P6��0t
����{Y9����b�$S�R��f�u9�ֶs�9��g3��;a��@�5����L�ĭ�ૂ| p&��H]Dd�k�/�20y�Yb����1�*NgR���q=��;�'��BHvej*e�	�Ҿ���Oow�ZDCD9"�a��1��E�e�GGb�j,j3��Ei�x=�R����AX;[���v-�i�j�tʓ.6vu�`4�6�NKh��}�L�����E���X��5��L��Q��c�=N������~�'�wK��c�@M���+�E)m��avx:��#��^���������ԉWY(N���I����_%�R�5.W\.��	���D��~��SD[����m�s}?��JQ!�󔭗!>�U�X��z̮9CGBn��&��#�i����~�R_����?�uî���v���9�v��>��7��ŀN�	B���Q�0U�
�_����&�U���n���yj��=n�X�d����;���d����_�<R�z*?���7��D��Q��ed
r���4v�~ڜ�5c��n�D��݊I��1,K��Ͱ��e�ո�W���.ί/�nln�h^i8Z�Kks�B�uj�uO�	r�Æ��R��������U0vH�&��"��C�r���-�eg�D5�}���7���C���\��Z>�%�3�N�+�G4a�q%��+��8��}�Z��JL倥�N���n�P�������0ܗ�uZ�~!�a(V� �ڲ�g@5���ғ��?B���?�����΀�l�j���G/��;�@W��������`zZ��$�q-����.=�����������S ��f��P=E�	���O�ZDI�+��B�ΐ��
� ��d�O��h.��4����"u+�6�~��8�E`gG�:��6>[ :������kE?�l�I��Ս��y�{v=��a�T�q[㻽�_O�))SYe}�z[��/���h�^\d�>��:�_������d`O�:���#�#���lټ�Ӌ���бK�3d�y֐d⋉�� ���vټ}�[�/]��W[�+���`>�ȣ�"��^�u�&�Oe�!��*�t�)o@nH$u��*��g|C��Z�G9�Bf�8��U�R8}U��vOI���{�ʪ<���Ua�>�(�4���w|�ir��L��S�竮����z@�o'0�J����j���l�/�8A@�U��?*1ܢna�he��#��E\�he�bV�ܷ,J^��l�	&d�P�3�rdTd�'h
1$D1�|SG����b4�Or�x�t��#_�f2�8��!4���h��2]���5�'f�W����u�W�&(I�H+C�h�q?r���D(�#��7~�E�������E(�I{� ��:�.1�q>��r�I����rg�A'���(��n���D	�����"�|����JtS[��(C�&�Ţl��I���!�H8c �䩿�t�
3��Jd�9�SV�w��}�O�}�?�=]]���16�����V�L�Ϟ�7ԓ^�7G��o����z�8��l&����)	�����ʅ?4�sy�(��e�Ѐ��N�h�� B]Y�7_[}"�t����gg �ʿ\�x�;k4��3P��D\�m&��vj���]��D��s�	�=��[ �e#L�6#t�/,�p[��v���4]���l��c¢�mWG�m/�mCz��K_�j����(�0�)�`�s���Ȃ�����Ax�W����Ͳc?�%����������B=���=��O&��Y�F$9H��� NE�e�'��'�ہыÁ��iX=�Q3w���Q��&B	�y;����q�'I/�1�Co��2TߒK� ܤRӖ���bX����ʋՄ�,�)�/u�92���S���;�*2�YV�ez��ګ�3�N�7��8��3��B.2(���L��2Q>I�f��n�{!�}�X��[���]J~v������i�	�Ԍ���Y�c'���I<6�:[C��r�H�#d��A�l�]|8��G�YF��t]��=ap���!h�w�������������#�����굺w�s��U]�1���l�/�)�F�R�A���<_v�Ȳ���qn$�tZL�m�*��ۯe�j�/X�/�A�[g�	k/+k[+�Hج"u8 ~�z"3B0s6?�D��`-q�,�6�,�t>���^���5MIʄ��w������*�[�O7�<�`�|"�lOMP�(.�_n������w����|�3����LwoH�A����RW����~P�3w����9�M�1!�5�Z��nt�������a������9澍6x�
�8��ä=�џs�g^7�����̋�$o���KE������hg�U���7�j�j�k�r^�_��w_cwfY-���x��t�Q
�?dDs��y��9�[\��ħ
7&M�K��d�H@E�Xs�h��^��:�K����� �0��h�Ty!�~ �*##�n��)OT�,�w���BA7��R��P���7�竵b���Ҳk�������A#�Q�oy�
�-��TKB^د��d�Gq`�z��"n�i�s�EE�����w��ӵ1S6V[_�,Ȍ����@~D��j�\��[H���k���	��8TO���_��q~���[w\/(�����D�3�i��J��x����0���A1g�}�*$Z�����~1�
T���]�����9�4��	j?o^_o��6��oC/�S|�v�-�׍���b*ũ��
��E-�򤕊Q�G�����x$���L���s���8<�R
je[��9Kv-1��y�h�c���y7��jQ ��9R�V�5�ϟ-6'��^L�:5;'B����=�q���}�85@��93?��t���3�ۘ.ܵ�tWTc�k�+����ۯ�:ne�p~	�u�����%�b��{����&��i�`&%�+�p�Y�@n�8�x�`vBC+S���Հ�նT�By�@�<�/��G?~#�MI�+;����{��c�oG���f�y�/�g�7�r�O�.��1��S��+�OҐp�h?��1�j�g��#��Ih �Gb��hCX�J�sp,,�4�=��G��B����ntS[SG]� 2�:|���),z	-�����m��$�`&R����{�l���9�P��xE�t��V�ޛ3��k���?}�b����q*�s2G��uѐ�1�i�ͦ ,vn�����z�Qsr헾��/�S�����͍��'����C�&���7�}H�no��3i�����W��H�ﴍ�]��|�/�2��E�-�6�-u��h�{�η��÷<�� QIB�����D4d�
��~g�g��0@vQw�'q�>�YP��(]FA�I��dA�eJ�h
�M�Qɓ��F����XEʡŽX������le~����O��'2׼(H���ÐЛ�i�Lp�Q|����d!�WSm=�b)��;���͸$�G^�u%h�Eõ��_��i���%�:��AC �_�紾b���ɬ(R��Pɸ����kV�<��޲�͚Y:�ٲM��2ڴ�*���iC�1�p=�ť�K�k�{3������[�24s����d�{v��I�͌�f4�+��������OL���$鏺mv��q��_�L>��ɸO�c�����%���:M%��x<�GyE�<	N��
�����v ���~X�h����g׏�l$��b�a`X������S�zd��v�k��e�*��̟ơ �EX�46�v)ZP/��7�A]X4x��6��x�f���Fqf�F �ڞ{��W�Wtcvv5b��S6s͎7�'��}*�X�Q�2���
|��`��5)��F���a���H`��.��s���DU�%���MY��ѫ��u�A�R��*�u�!���!�B���}��əf��K������k�SzVA���{jI�G|�mJ�b������h,'�U(�i85o�����?%۽�,������b�C+J��rT����d.�C�픎�b1;~۟������u�ˮMn��I<�S��n��_S�
��i�^���Z8��ގ\z�>�R>�&���_��E�W��~ߠ��x���:o�X���`di�}���ך�Q���%�������\C�:�醣��hD��袘t�=0'�0��3�M��GL5ٔ�>/��~�2W�T���=��(jj�uel���cBw�F�4��4`���|���ty;\������~���]槻c���P��)�Dɿ*WY~�W��*ǐ"�T$�d�M ����'eZ����,��p��oy���|_O�>��t������@64p)�\+MX�`�����i1�4E��p�5�@9_��P�"J�	�N�wp`����C��so�5��Q+�NY:���_���s�D`*���y�S���eD�*e5@x������x(���7\b˫��/çż:�}��=�)�mg�瞸㙁Q[���_v�}�����L�}��N����7�]�z 0�'� �R��3UQ9��f�+G�KG�qkUK"�(�H��Ð����`��4�c-FAf�����>�_Sw\�l�a1ϲ�,_<J��t�}lj��v�?��2�0p/�:������6���\�1h Χѳ�CItIn���I�6����������;e%�j��]�Ba�s�2�Tr�a `�A�62ͅ����'����=�4u���D��P\vB����R{�5��|Q�
��LZ����ؠ]��b�JO^��Rd�h���u���>�ǋ���T,��ED3j)>H�S�W�8�P�>q5jj��ݳ+���K������Ģ�4WM�� T
ię�����?�W�s>�+Sk���MN�A����Յ��4���0���w�qQaX	[�B�QR�)٘q���X�`��(�N���_�8:͐���[�@Q��)E`���`6�¢���R宖<���(q��
u#�<n��6�����w�A	O�WCc>)a�K�Y�++<���:<H2��ը��9��4
$���m�Ý��)Dи����������K��ڑ��#!�H̫^�~�� Bh+���a��w�����"�n������yqS�I6~b�m"Φ�3UKocU��&ص;}�"
P�`�&I���X��e��J��~�9��[,��q�� �OYE�w�5"x\+ �Ɲ-]U�aP8M�=�솯���;�5�m0�o�b�9M�Ov/\F~������&�{��J������"��4�8mc�~Y9{��[��l�)"�����aד c�02�%�+���}ާ�FN㿼M
�PSO����OI/P��������$@�j�~�zX�-�(�������#�����S�����/s�s>����Q���<7�	�2q�F!,��C�س�v�����C�J$����ԭ5�Yj��fs�D>��̓����$|[Ne�g�do�%$"-�6zor��U)�S��������c|R-���8YE�~8�8tY�}��l"u�
�����R�%���!� �BR Y>7{c�{�%'O��L��˪�2�&Y:�	PMZ�7�6�\R���n�ѭBE�����2^{X%�u~+[gRt��ϐ��d��_�GΏ3J��Pk��YLR�:�_�m[s��f��4�ܢU،��!�.d�~��գ�Zp������Ğ�f�cW������?1ƃ(��7Ksh)b����E3*�)Γ�"
�<�Trr��CĘnw1�0�ןt\�;�_�C\
�lm��9Ӟ.ﷄՑ��>���׎	�g<��4����*����(��bKHf���Yx$���@+�����[�44�2>hhi�<�莽�����ܺ_19 �ֽ�h�#Q�%?�k��`'.���"��i�S����d-x��M�.m^�+pfi��B�Z����GR��i�c�M���`�ۣ�(�s8l*�o�Y�����t��4V?��&�Ea�T�:���R�dѷ	`j^�1��9�^C{��ipy=���v�&�4�R6�)"�A�x�D��"XJ��[#���<Z��w��:�F]�-g]>׸�b�8li��$��>�Ћ�I�?)ið{�ޟo��G]mLL��s�yİ���F��aXY=K查[�¾l`�'_ތ5�r�������|�I��"d��pd�=�hUt���e&�
��n�iNJ
��2�(4�����<+�@�e#ϧ���&@]�H���Y�(Qw��h��%�c!f)�V{(a8��֦뮞�����B��qg�6�M�F*=Y�����K^� ��{�t'�%R�����G]�Kw��oz�w���F'���3ŝyQ��i�d��+��/}N�y��}ba����^���	Ƌ�h!�=Q4�c��)؂3y�]�#O$��M)��U�d�W���h&掘���m��>��������8X�9 ��O*���W[��gn�m��Lp��P5��Wy}��e���հ����ґt1F_�j��N�z��f�qۗ�� �X�2Wܯ��{ȥ\���@E6�e_�=�I$���k�)q�)Q�\�-0[�%��b�5(��$�8o6��SWl]�%�^&G ���{����c�fzl���"�:0FHv�&��<yPG�Y�//��s�#���aG��M����kw���=S���X[\7�Oj/I�_�w50~}�҂��g��Z�EfTmb����o��
�"�H��E��X�M��js�8�8?3#F�J��s�sFpۆ�a�ё�~\v�H��{��	���l����86�\Zr'rtm�`�
�-�%+a;�7�������_��G�1r���H�|�>���lԍ"A��O�!������!4�5��~0�a9�����o/_�Nʻ��隐��{�j��ܒ&p'�H\��*.W�n{d/HT0[4q��Z;�W�X���]|�����\����ϣ+����o�=^m	�����B���bl�����AAl<����?L�F0&��<�f�+���p���!�!:��#ڻ>(��^V[����8���p�B�h�٩E�]<N^3#�q��-��CK2�	[��y��K��ۈ��HE�ֺ��{�koF�Q�w��xM���b�>W�\��T՗;��%D��nO8ߞ�v%�����p��V7O�.�t�I��-�U6g`�r���(#�T���߲����`oBH���.��/=��!�7�d�!�9���J�Բ7axΛ��c���}����:F�rW�K{n�I}4���4��$�����FR�����m�~7�*`J�/4�2ղ��ed���~�Q�~��8?��X�Ej}:�M�	A�Y˵�� �&^��EK���s�%dB��u7'�ޙ��%��/Ԣ0*c`gT�{�҅�S�l��[x�-��fT��C/7�G:���?&z���l�4�M
�8��",Z�{����wD}s����\�����AF5jp�������'��&�.�7N��c�@9�R!��8��8�P�.n0�_'}JJ����aw�dF����{�'''�CNNU�*�y7@0��*	4�ؤy���G��~�������� @�Rw�x�v��#i		mau޸�Y^y��&�NB��%'Xse�X˦�ǇjiĨ�1f��(a�N�9>O���춇���`61��E�	x�,}>����6Kg�o9����7t�b<����^$�,��A	�]QLJV�DZ@[��hoW2fD��:\XR��g�h'#r};r�ng�zM]#O�PŇ�=th;��f�"��/

9?���:�!,�$�U``�0���P�2��R�!-!}� �N���w5��n,����JV�h���O�Y��D �����`h�rnC�D&�#�D.dKH�(�cH���Q��,�)֚1�Fq�|u���z�؁�XNo���G �݉��oG}�Ѧs
�]h��y��Ӌ?�����b�-�B�*?M�U�$ ��$�H�&�O,�w%�K�1zL�+�.���DL3�OT����J�Қi,�]�D�y�`�6+&����*�w'�L���IX������&� %��;��B%�^�]F^b�$�Ic?���C'������ '��M�yjUf�ȁ*E�>T�����SB��H� 2ገy�=�oЦ�[i�J�ս�y��X����um�r���G�^�l�.h���l҂B�	Z�%"�pጤ��Vx8�V�rq��<)�i"�j]���BDz�n���7^1�����pE�0��R�O�_�C����핏���Q�Q�3&M**��e�`c?ۋ�d��}����X��/N�;�j�i�Q�T�{��9Y�[��2���"8q0����N��t�K���B4��/)Qm�$V�����E&r[�1�]���������g�܍���w۴ާWֶ5�.����0���7y"���~��.����K���I8�+ëEsE���#��Y�0��o��LY)��{x`}�~���`�X)��p0F�5�^wGͦs�`�>�C�k�W\W���q��A|!��9 2D�N�ھ���[��`�l."%�3�
��f�u��l؝��6y&s��o->�pr:�E�ų��+X!2��	���"�2�����,�Ne�#nd���'���6��':�T�5����%��_lj�#�I���e;N1??�I����H)�3�N���}��`9��:z^#R���󱾚s�N �.�"�/K��*���(�e�ޏ�".M����'/�o6�j��J����v�����C�2��u�cW1�ͮ;�T�Pà�p���YWe����aj�m�w�o�����<@���,GqlX��3b}:�&�Q���UA�4�� ���o�څ��?Օ���� 鰞�?�x{`#a�;CY��/�#7,��$6F�d
:A�2�p�8A���vy�V�c�HU{���,��8��	�P�pS4�oPFo�+p��Qv�O*`n�t�
�ͨ���ə�kǘI��|�s013�dHJdL��`���-b��NE���xA�'XQ��jX�@D���+ꆈ8":��V
����T�!�]���Q�ѯY0�*S�����4J��?$~٘�h��ـԪ4P�y|��]��3U�%�I2f?J�SC��S�!�ne�ܠk�c_S�rBU�Q(�\�j�4�7����D��!�jE38�}�A#�C������K��^��Da�깿
B�����c�ϩ��
������wv�4;��`�'���v�7���;�l�>3#�ȗ��5����V��/��W�����|�A�TEfJ)�f�}���;>�JG��Z��Qz�V�sǴ8������/�Lb�������~4����rmR�#t�w��5<�fe*j���0i�IwQ\-��P�j3��g�w�"\+B��*�&%����=�NWZ��>�:�A��E�����l�g�fN4����K�!�Ad��&��8�@_Wh[/��2묆��,�KUO���q�(����e��a]o����Se�D"�;��N����	(,t1�nd{��Qw��Ңqې]Ɂ�W<���O:�쪦���+dRaˠ;T4�>�R���ꛝ�|�g�a�.$ڢ%��=W��5������Wի����f$�;�x$�B
�Ǜb$��q�T����T��yZ����<�����jW���������ʼY"��.��r�������m���y[�FA����oˌ�uX��W��П;�c�&n�y�^ ���5~"�k2�v�i�\O���8�&-}��jf�|��=B��C#��\AͷZ���KV�o^��g[}�n�r�����v��4W���&���"����SಋT��px��*N��c1{�F?\��UQ�pRPe�	�����ɒ�}���E�،��9o'�5����-�?�F9qvO���@��ڼ��Q�K�lx���4}'�� AZ(�P{�WGM]�����U�:� I\�,��#A��g�gn֚�?|Es?օ}����T�Y��wWT�=�g��z!({*�o(��}����ol��j����!���$Y��{�#{�bR�p���´�o����!��i�N�d���!H�"cJlK�ƚ��xe�<HfLv�T
BbWc��Og[�I�b�j�2*�u
���`9>�}'I'�*���9�d2��Zݰ��*X����.pRp�ѥ?Ϗ:���H���{Jh*�.>�(jD�ڏ/V�OV��"��aJ���ʴ��Rj�oIuh3 �q�N��LG�a�T��^,���{�xN�S���կ[%юy���_ם��������~b@�Y.���Kaؘ�_�3���h��/���0��p��>���"B��H%[��|�겍�� ��W'�J9�qs�)"����Z��T�|��!�p2&b"lԣ��<�>�,�)�3(x�/�A�z�ELa���AM�x�.�Jw���3x*G3�i���k�F~9x�� 咄����PA���o�%Y�����e=~7מP�r̂ ��*�pF?��J}��8��?�  ��q嬦��Z��`�����L�*��M�d�u�~=Dc�4��� �$Ӗ�ڤ����Gd�z�[n�7��[��܆ޣ�K��8U�;����v�ق@�i�#~iΑN�T	ƣ�05�?L������������K5��%��&���*��-�-CI))��:W�ā=��zFO��Gy
�gt��v�=�N�FYK��a�)��e�'�j=��vC�Q�G�3�B_�5c�Wb��p��4����`���L@��߾h����,^-bc� Ϟ0��X
|�ѹ�&*�W��\�W�͂�>P�BI0*��w�Ar��N~�Z������C< �!P����`>������8�>%�=	��h�֔�Rn&�Dˇ
�r���O-ϝ��� ��f������{ߑ(��@�{�B�T�RU[{� Ζ��=�B���M �yמOԘ����Uy��B�V�d�rc�Ŵϑ_��Ԃ�&���n��Zo��n���Z=.`2	3):�L懷�t�X[\�R�<0$�\\?�Q�����$S��1��r,�plxU���v��q�c�h��F�;�����#����(�H���=�jK0���=K8�i� ��k&�4,� ��� �IK�!�ٝ۟ҟ��J&�8��Ƒ��sN�y���Ƅ৖��^�|~�}��?<����4Z�Qr��ķ�d��oB���|Ɉ*AA��]P��2�a�D��я��jX�7�I�a#����a�n�j,xnot�2� �w���]hw��E�xH{�Gs"hc���`	��W�6���"�*�&LB��+qc���/�c�!Hrz��[����|wM�g�ȏ�M��D>Z��I���,��ۖm~Qs�������+ww����.ªR8e�%���7���6L�Ƣ�	�v�S؜���n%���W�������g�㶃J��Շ�[�O_\��<z�,�~�ʚ�Uc��@�r;�|���z����l�Q`�O�ĭ�E�X�A&C5�����5�j��:�I��l�(/�� 9�I����Z�#U�#<�x�y�$�hyJ�jם�4S=\1��%$S��+�>Ĭgh�|4<6bأ������v%����u���ﮢ�s'���.IcaJK�8Vtc�}O<o)�������7
q��0���V6�j:��f��3�yX�sDQ,b6�(�e�8RXC
51�nVI`��(ȩ<�~oX29EA��H��_�=�2Nq��%��4�a��Q�=��T{CѠ���Q�� ~1~ʪ$���4��Λ܏#Z�X���>��
�XhDe^;{(kޯOz�W77#&�{((>+`�J �dݬ4Mq	�@E����1s�Y�Cp���1����'s���qo���;�k�@�pU�����F�/�:vwxY:_���GƱ	-,�,Lq����Ӷ'�;���ށ=I�e!.�6���%���$��$�J�m��N#k$
,Qى�ˣ3��1l>[h�h�0zxII�fH�W*@ ���$��煭���VLfj�M �|�XĦ͋e|���á��Y"�I���}~����B?��UB� �����A2�co��G}�v���P���3P�@AF1�B���	�Q�|'�t��8g<=W2�I6�5������Y�ܳB��b��à�5��t�K}Tm~�[�r��w���|J���zdGbK�÷<bJ����Lg�57�7&'�&-���pm�)�6�p'1�*�~��U���(�E���w���E2#��MK��˓&
)ؐz�$�=������j��l4m㵛P��39�t�<H�k�>��Jx�vcGFk��d� iE�-�J�yc4�?�BZ���
��sF9���lV��\_��Q*��K�ª���5���ԩ�3dxFx�]���rdio�؏	����o�X�C���z��3ԉ�(NȐ
��oa�9����B�>>�;�Yށ
����H���m�à�"���(!��p����
��`��k��nXƝ�������pį�OղQCO<-�E�osM^�� �ZZ��0g���
��H<�3�*eN��A�so����h�"�x1-7�*���D_q�_��~e���fo$�FbX���|4ѭ��~[�!7Ht�w�7��^w]7߮��>�������<�����گKf����/��Im�㒮	�
U�'��d�؅�uLI`��p�]58[���uz�҆�f63�C�̸�Rӌ�>���Jj�}���ׄ͹�3-��w�w����K;!��p�W��5r��"��=9Ҙ�������a6��������G��^�g-�b*�i�+���,���]�Y�����bT)����Y!�8�,'-�:�0]L#	�za��z��P͕!Z{�2��n�_�F��a���aU�i�(��eB#A2vY��T!���ׁu�-�M��eb�&��9�ڈz5�!�O��cvE#�3?���X�X��ru7O&�/8��y3 ֳz���O�F���{�HT�c��Q�!��j4��R�N��Ff��3<�V�˖���3�_��Ϊ��̐�jF�	������-�~���2*
M0��܌�CDN�/g2��{��Gd[
L:~���4���gd�FZ��y�*��}2A4�Jf��Rknֽf��z�׶��0�H$�;�e���9�:ۭK� �A>�����'��,�Z*&=����q����vǠ��=�D�e�a�]�7���d�_]ҝ���$���ӻ�ҁӰ���X�ҚƤ�f-+�R9�z�f��9*
��7����vg����1��9ac�7��
��'�o���D�wGчa�J��rY�&I0�ҏcSZ2��8�S/������y�P+��1�߬���"}�!�[3G��.����;���Up��U��yy��h�Z�Ţ�<0���?s�wxs������zE�/���l�H���N�EZ�og��w�Xo���������+�u�nۗC�t���|
��l������N�Ӳ��_�F���ِ@2,�W+ÿ�y�?�($������9NȒ^Z���f�cO���Q�p%�A�A�K�Pd":����I�2����������?|GKC_��F���._n��F��n�&��ӕ���>�`},1�8�mqv��9C�w��{z�t���2����)"�N�	����)��t2��%�%���6�.���W��1��+^9�(��/.��,+�Ӄo�,�Ea�Gzb/��X@���`�R��$����ڗ���An�n5Rg���X�ad��l����`���܆|8T����R�Ř�y t�6�����Ɋ^}��f(FkN����i������N�ꮹ6���|7b��a`�R<�Ed����ay�̍i��^B}$P%�
h);9>��xh���xE�6b��dx�Ԡ�"C}A9��Q���}t"�R�Hʿ*��h�3�hA^�b885e3���o���Q1s��+��08�^@,)ڳ�y�MvMy�aG�>A���^9�Eq��>�w޾�m��U�<�%���>����t��+x,+����m�����Ȅ�m3�.XHHX8K���ݍ�Ђ\t$�y>�� �b�ώ��**|�cX>�іA��*�iR�a�z;Ũ��k�H��'���]1�~<k��
�����d�n*EΩ^�Ww�a��ˇ��Ƙ������ՙ��b�$���N׾�|���X�ž 7x�P��QE�{��x��w��F�q(JT�J����/���S�����禭�7��g�F'�|߿��(%R`�̙\S�A��b�tA{�Pɻ�Y��?�8�|�t�p�Y}�U�����Z�Ŕ��4h�~V:r�:��_-Y��Yk���m,����/���V��ګ�OL����'DMIZ�y����/lTIn��=70�$ �9�2Ȓ4uquKf
�����A[T\\sIff{�{{)m�a��$�j��}ݖi� O��x|'`��cT�$R:cj`]���M���Q�)�������ߕ�N�%�?�S�����"�Ha-���GW��;
�6���UB��U1�2��� �s�GD�("�'�.-rd(�[ʗ�$���h,x����J>�~ �6�v�%4\9I�}C%�<	us����S
(s<��〻�p�G�Q� �(�P"�	S|�9������Ի���V�@��9@kT�
δo�EX���9)�����'�0�n�gr��Mͫ~B}���'%DN/�lS?����h/!A�}����'ϱ���v/�z��& ;ʺ�m�*�b!Z�UL��NWjNS�M�8CrR�	�
�!.[�ݙ��Z,��1����n����������A0�D��X��͆<o{�W�@�9(yH�����
.����s̀淓Q�>���DkM�X�W�v�8Deg�ةa]q{�l,F�����OO��<q���rD-�❣�fߕt��g��b	��LE���*�~��V�-DQ
饮�'�$�egZĜ2�o}e��	6�ՒY�A���� ���f��+�[�_s�L<��'fR�x���x6��/��=�Wb���)$qYQ �;��vb|�aɃ�J��v,��?ċ*����aK��ڷ��O�o��r2i���|8*t}�*Z}"2_�Mf�����"NV\nC�h7ɿAp�H�UZ�-��e��ƅ����[�ӆ���ٲ��_�,"�Д��.�~ݯ��/&�N���/�!jr9A�|��ou�\��n9k�;ef��n���l�����-��yAD�yCW�<��u�%K?�|Q��<�V���u7�~�mzHJq}�¬��u�çO���f�K8n���O$H~7|�dp��w:��W��+����ѯG+�Ĭګ�]450�����V��F��l�E���#��� .:l��^�J*��y��)�����f��{H:L9G��Zc�b�b]�&8C2;(�f������گe�X�cٻ2�
�v�L"����T�G]��-�>��KR��t�Ynq�B4`D�4b�o6�I_�J��R�x���	,�tR��эXP�"�}lt੯���v�2���f��Z�^�U5�����(~��R����8C�՝�P��>7y�1���dT���Bf���q�x?�*��!sZ�G��TK}Y<$�����2�������>��UU�d�+��^/묬���_#]m��*B�>P����!��υ�߅K���y�+�Mz���޻��lm��>�x���t��K7\�-ק���˦����L d��[<�<<H�9EJ�_��n�wJf����� `b&lz	��o�Ti��CY�z��v�����$�;9Ŀ����#o�-�&/����� �å�Ւ��65J/������?+�ؓ�<7j4�� �d��3�%�`J/���h)��z�>O����3yF��{lW:��-W=�"�XԆTpb�wjb/�7�/G������m�K�ɼ�����U~��5�(UX{��~~{&~�|cKW��;�WC^8�M��߽�Yz�3�(���Ѓ�����E	NO�b�������@�2��3~"�9�I�^�^a�"!3�0�@�*�|l����N�#Q�W[���v�K��,��2p��M>�A7�V��4���g�K�������0 ,H J��Kr�����E��$X����p�G������덹�u��(��Q�_yw��pn84F5SF.��ܨ�.�k�偭��~�)����Y�}�r�����'�Q��*?"�W�.��gL�F��D�=��΅��h����6�J'!��1g�W�M�����%֣OG$��j��L�! �  ��՚pe��z�3>s�G��C�t����}��]�0<��ITd��~V��פ�	ay�Y�֙%Ӿ�*�bg���@$�ZI(K��3K��E��K�ʝK�=�=���x�����5|_��ҷ�RUh���wV�U֕�Eg��U�j�\\h�Rt�9�����	i��,��^��Μ^��J��	k#���կ�_$�V��d�.���u2���?�w�`Hq#?�O�O!�����I�@~ԬikY!�����.���wrj	.>�rn�.��y�3=�El������)��Vo�*�lc�/
��'Q$UYU�qT�i7a���8�y<�=�`�C�E��|��ߡ�Ă��2���	�[�-D~%��ⱈ���ˎz�.�F>/�gz=!\�̦�e��W�&�Z,�r0x���s���;U��N㱡�����$8��>��w���P�Q�缹���Rޮ["����&2G���dB�k��X5p�\�K�݂���	����m�y�<t��ck~�]�vs.�v��Bl	-x�U5����>�;�+���.;���n[��&��e�����*X�( �q���&�}�W���`�K:����������^s�� !݄	�D#&�/#�mewL�jᳮ��Q����6�����#�GN�p��S~��4$4��VgƋ�ŚH��VW����(Sp��Q���X��N����'��C.@�j���Po�0,è�d����w;g��1Պ���:P�t�r���/��Py��x�>�Ka���%��G�kJ�+����Cч�+Hx�5�Z�#Gl�X91#�6V%��Y�3Ă��܍�gn����d�}w�~�����E[5ޙ������Wj&]�+�Ği�$�]��(�Y2���3����(��w��
?	��0ҮE��uZF���o�㵻@�B�1�ZN*��~^ s�-� ��h��PG���3�M��u^���Q[�[P��IZ�<��j:�����j
 N*u�L0Ep�?��w<�4G�����Lޖ�_3��m���|�Bn���c���X�
\��hJ�j��+-W�'9���O=[-�_�u�{���T[��ƹ2��-Xm=6OM�����F�o��-|�$��s�l�ɧ:��skzr1�i��,�ѽ����4#�7y^1��"aJd�?I^�v��	0���tTݏԄc��l���ڑ���{{��w�f�T)���B+e^����oiB�\nG�x��Vd�nw]��`#G$c���3�@P;�֧=��hQ�4�P�X�<���HA޺�⢒���k����4A�N>����E�T��yvڈH��W�=�\#;Uh�iI'���N}�ҙ����S�2����
%�iT�t�!�$n�j�`�ߑz����Xu�}*��y�Ec�,��Gf�b�t~��5�'.<Χ�TI�cA?�qζ���	I�	vS�v�>�'E�v�7?�pQў)*qjH�f"i~^I��/Τ��rě�ڙP+�jwdL��ť��>W�����J�%���-)��Lc��b\�Tc�v��Ã�s��~������F�t�W�ɷ:HN*���O�m�����	��hz�\	M|
����hx�խ�M���"2��/�z�����Eǃ��vQĨPFjb���R�t��x5يB�h��sPLڢ��\�d��a�������+P����|��$ۿЁ(���u���T�<<�11�����C�g E�T�`����ddh�o?�����q�bZ�ư�ȇ^8L��U���+[�Z.j�|���8�HI��P�xe�%�	Jv~�SWv<���[����i�1.W
���ib�P���T�cvJ#*�f|�-�z�*��L,R���D�aŭ�A��r
��N�_���F�1���HC?A� l�Ǣ�Ζ1�Su��ɞ�oix�����ˀ	%�<D%l1L˘�����7�U��å��:qU[��������GgʨR�&a�����M�>< x.J >�a�v��=6T�/W��9��2����>H*�v o�K>`���J��C�@Xz���o|��a+ g����2�����P��
Ņ�٦$=)����3��E#ڴʊG��I��@�.�Z�cr�=�P�������~E'�v�ױ�}�+��������B�����M�$L9����?����UQm�]�X)V��[��^$��-.���][��ݡ�����}���&w�{fM[OƦ�:�WTZ`=��/��/�
�2 p���C�� ����W��D�̓�6����Ћ�w�$�W����[% ?�94Ӱq`Y����mij*ټ	��4���[Un�-�ѯ��� ����ppS�,t�&@(��f��t��_r+�T3�I����e�F���\���|3
4$m���v/V$9�'�n�IZ�*XA �2Y���8x���J���k�3x�w�x]������5��MMC**����:)�C]�fϻ�b~Y�,�Uw��R���:f�~���v�w�� �B{�=<F(нrG�$��տ�Gq��c�m����M�����a¶�M��7�8��������ӿM����k&'&����������h����Pt�q��0���Њ�;��x�,����xv�1�D�=�^7�_���*��rT�gݫ7�ʑ���SV���4C�xg)��t��@���4�I?\\AI�(�"�R�1��������� �F���Dd�����,�[0ME���H�����H�x	S=�@�� ��XA��r���՞[42t���ͮM���&2%�Nd���
::4��L��,|���<-����'�~�`����0�T�����E6�[��&�D��6���
Wla�Ck�S��X� �p>��@��?`c���f�G˫l�}���?s.���onRO:���)I����|X�����d��5G:B bN5����u�g�-�g���EUU�}-�'G!�~�J"�E;9ַ6o�;i����D51�d4UVw���[[�iw]�e=i��g)a}��Q����*S'/u	�9QV:��Ů��Ȯș7�u�1R�������1�D�L<>���X����6w?���M�+D��C�hll�����i��㯴��Y�ma!�#�pE��p L�Iz���cJq�$	R \����OaIt&
�wg�9��8�����=��8��������K2^��]�R�A=U_x;�a#�$5x��]�2�@5���P�&R��r��~!!�O�js��V"o}��@ˁ��G*�D)�C� sy�G\�z��D���5�7�a�'t���3����������`381*�]��I\z/���,��������oC׷����Ym~�[��l~�G�D|�[[��f��Ɂ
z6���~��F����Y�Ѕ��zdN��\t<u���N����}�Mp�,(�8�,���r􇇞P/�ҿa�)�����[lC���$��|������vw���;Kme`�ơ?�b�`{I�]:F11��-oP��:�u�d��|S�dv�d1N���uQ�Q�`̓[�\����L�绘
��
<�����,v=X��PI� 0�aʿ������X��)!���H�a�%��t�SD�2�z���Xk��=�\J3��yU��MH5ri	��ZC���st��ߑ:[��EaiQ�j�\�ą��/�j
*܌Ӝe�Y�S⤢�B
m�A���`�Y�2v	;�*�Y5H�x��\w2R���{�<'��j�"
͟G��o�>dv؊�WV�F*�K�0�����)V>�	m����y>���r�K;v���/��E�p"������bBZ<\�+++���h�^���#��ٴ�����&f��*Ѩ��(�p�}�X���\QB�)��G^��e��[�����%�$�a)�Y��AEY;�$�g��!,7w�	8�c��E��"����f֞�ieUo�y$WzB���COQ��6��y�ŏ�����?�F��1�J�# 
<yp����0�L����_�21�,�O�NL���D	�8.�z�y�ļ��x�<�iƓ�0,o
�7o�ܘ6׶lo�'��ֆ�	���31~��fF����0DwT��)S~
�
�SD���SG��X"7ג5 *��EjZ�{NB���8��+A�`��#p=B��F{��Y=�.J�5�P�5j�s �N'n�#���������M�@b&�~��u	}R�5<����Ŧ�z�"��'"BY 8���+U����G��5D��s	{ -�:��90���[���^^��u;���,�+�w<����w�@n�X���¶� ��cF�K*����I(,�������AI���~��i�/M��&q^�����ߧciniQ!K���%u����rY�"��{E�T�T�nX'���ٯ�߿�d<$t���B�.��S��p�d��_��i<��>7�}�&�������w�ׂ��?���&k���7_̟]�v޶�7�R�x�I1+���C7�\��T�=�W}&l1�]
$|,�g��qɵx;�\`���K��/�~��P���.ȕ�h�F�s�w�|(��Ji�����ޟB5ڻ��a���qpP��d�����-=a���B���N�R|1\Bj�*��oh�|���.9-^�S�-�X/9Ԛ0&3~�B���W��P��E9���� �i��Xc�+��e��po��"&&,�KI�T��ز�!� sae�B��?����˹�^����R^QU��8|p@���)2�Cq���7�����W�Q���c8�?�9�@,X��pՀ�����b�]l�8C�"��Ԕr4�T��S�K���a�����b��Np�Բ���J���T��������/҆ݍ'�AC��N����-��.���~�l�r�9I���ǘF��ui�_v@���#�������y�vIA%IS>��4}2��^!���VP����/p%F$e"@�d��S�Sā)$����H�wWI�ĤӇ����]��s��A!P͂�jh f�X�`�hm�`�����k[�H�0r������)EX��4FLnL� �����$Ɏ��a,E2�g�ԠV�4p��9Ua��A�)�ݏ��N/��j��V
m4�0�0P�����'����TN6�\��RqߑZ#��ZG������C"\��E���i��?�}��6�ʍ�$�򪪛�n<||���s<�$qM������<k��2���?6��
+'>(U0iJ�͓Z;���KX�FJ\)�`y�3�&����kjJ�%H��y#����ѿ���Oo��ݢ怉"�
��3X���o"�X L�zE��~j�y&Ssk=�W��	'����Ѻ:�q�:���*������ј����Hİ���Z�35)�<�e��Ƣ�����'�L$?���n us�)�%�>eB�lbe6ξD�O�jt�U�> �F6&�V �l��C�ȃ����?gSV�}g����}F�M�rA(5o}����چs�@V*u>��O�ۋ6�S�v�M��⾸aUU�D�\a��$C�0�e�j׃eS�����la�k�C�J�p�8���gm)���kܣ� f<ɷ��?�b.�IpKK9�H�Ƒ�M�Ԕm�Y���:o���.YZZڿ�\�9�8 ��{��B<�����*� N����2V;��a�h�$��ji��hA�ZQ��jb�5�(�?>K��K���ٺ�[����<b�Q#Lx���s���s���ڵ5�rP�E?g��툆�1#0�hk�5��(�B�����N��3�(�WX'���;[��
��X?ws��V��m������#�a���&V��b@,����7�2#�(4lk�2O�(��'y��@��Z0�O�;���+9��wEV�t]#U�(��Fu����j��B,�w���j�W'��fl=8���P�~v�z\�h�5໐*W�Ph��KNF"����+E
U�[����S`&��3����q)]~���m�.�+�+���8R��XC�J5o�7C�ũ�C%U��ZzCw�����Dc��|��bVo\�@�m������B�q�ݱ(����Ɔ���ϳY��;T��w!Ldd��"��k��3��b��hV�L!	*J�3&�M�Ob�>϶���� j*]8��0�LI��q�}"J����J�r����a��lr�r$Ch(���	"��D�W{��V��}��T��@�+U�#�uM����}v��;a�u7t���_�ٰ���ʂM���ϷD���݁^�r�}%��£F��S빔v32��nLxu���x�o�m��d=�?,����2LuU)�Us# �e�䄦I���C��|�p��\���9�6X���g�H�@"��P;C{����|2me�P0ps�^�A���gr�an��"���#�Hn��nY.��(�����poy��d�Oo�PH3[7�|y�@O����e�fpK/G�::�����>}��7ifbyh@M��t�B)]{5��a��]���������|<.�k�� llt~����>�[_P1xS���]����W�&��&�W��V]&7���Pmd�:s2���)�9��Ʋ�Q91��&�֕'L��lF�_��mu���ժR�-��*��e�#y�8V�r/��3���(��.��BN�J0*$���p��rɒ}V#��G�`V��
�����{��7�7�·�{�Ub�)I�\ѪE!��;�'��Z ��	�$ֱl�b0�<����
]����t,a�&C��Q�|��b�p���٥���L֤�7��`lhu���xl��<�%˒�x
i;F&�(�����z���!�;�n�(�弑�m����՜��*���]��~3��3�R�0>>��/�&�va71F��O1 �nd��~�W�n�⮝���tN���졗i�\Tu,qrV�x��EV����� ���LJ�b�i98����}W������W�����!?A
%����hdd�8m�˭rT�b�W�3Z�٦�(9�͚����̄���������q�����6�fN~���|��J��b03�d��q��أ��}ÝS��+G?V���?=�"���r`q#j�rsp�A�܎#��4�|��3:����ч�u��;I��L�6T)����ƊL������GRE�.5|Z=�q��-E�#DU�8ȇ��֕H����~EI��m����mP�hL$I`���I�Vx{1�LI&�R���╩�یE�yӪcۺ]D�o� ILE��b-G���;6o�B�C��W��s�i�T�<�$!)��#s|˓��o��gfБYg)Լ����I/�h�zS�� ]cG\�oL]r
fc�+bG+�O��Dα�p�҄M���.�Ͽ�%g��ϋ]���ןu�����\��q��=�^\,֘�b7��/
�ڍz�p�d�q3��hU�x�%���(%��(zqW2rR�Ň�fT��>���r��'y���^�_����ɏas!�f򹡊1��ɱ�T���6'P��l�D�( ���g�Q+�1�����	��j<����g���!	�'��{���g�]�W�WĦE��a7�Ŧ_�Zًim�|]�z��e�eH����� m�J�V\mr�j���DC
[�9��fB5q"gJ#IIR^UM��LR��x�y<=��9��G��ԑ���Z�WD�9�5J�p=���;�8�ɖ��]����Q"��I��4�����F~��/�&Ƴ�k��H�"(�O�P��3�1O�[���dee�ݩ�<801oP
ͬ{kAG����Ӕ�B�����n4�f���W]�L�0s�_�h~k�y��3�6������q�e���A�BGu]�c�Gz0<8�I1K�S�k�>Նk��� ��c��@"��V�9���a�	`�ec�0m�A�p�8_����ɤĞ�*Jˋ�L˗�h'�Vԙ����=nʺ�yz�������W���}p�����~䚺�q�}{{���w�^x��3��� ������1�q�T�`�iuG�c��?7�Z�(�+e jEh4ka��w�,b���2�7�I���]�ʯ6�qH�2Uā�uZ�b�3�\7��,��<��D���c����ky,.�����]ʅ�Fb�~�ܘƝ�Zlز�~oo�Y�փ</|�Ǯ��ÐwL�󐷱�ֆ���U=?�����{m��`��I�{`}��!�_U�V��4I��Oo�d�67?��R���?�ì,�^炁^^i��gk����ۓ����"��@�&�[|ғ�0@��ɾ�pT	�V'LTa�+�'��,��O��/��&�������Gj)&b[W9������3���dZ�:�m�s�H��b�{<�׫:�_��2Ɍp���\.&	����ͭ0���DPh.�w��ٱ3��H��76^2^�TA2�/4հ^LDr��8���SD'��.//?����F�����铙�iS��5��g�ZR�&�fR@OZυ�\�NR�9cYB�b��o+ȁ���MBM̨��N��	�\���-sbޏ-�Ls��GH�?qk�ta�u`y߉��:�s`qX6)�R	�i���z�Ԣ$�v���FI����vELЄa��2j@x���$��jʨ�zSQ����2��um���s�I/��Q�����d������o�_��B=ĩU�"n�k���7<��G����ORs	v�$�u,liKC�'I�MxP��>o.��Y�:�%bF#Sl�7
J�Hf���
眢�_^��cbhj#�d���&����2���]f]b�r�HcyN��)ET�b�xd�]�~�E)�ܨ���b��ǿ���Ij&�WYմ��i��σ�!�Pn,� ���:+��mA��܍{�m�ޜgg��_ �f �����=�Rv}L�@�딇������?�\�sn�ɿ��7��~yw��y2�TY�pU��t���w�+�,�z,B�H*����@R
��OI�f�YG�Z~囊F7��`������_F��[���XftCA��-���������yH��i������+UFC�*��7�K9���'%'��*������kJ�[��f{��ٲ2��C^�J��&Y7������
�g�g_���Ya����dm��q�I�}h��ڝ��i�'��h$�1��(� 5��D��,Vm��=A2��sPn%�q�(�wĶox�WB��u5�t���/�d���s���x/m�H.��uG�Hf�"����ʪ��2��D�s�� (KG�Z��c�K\5|2C�ގO?Rg��f��9ٕp��1܆������Ɲ��ͯ�=`�}^�ο����˥G���w�O[�<����@W]me�)����kl��y��lPMGGQ��mt�d�f��|U�HS�S���ņ�;���nO�0��Շ��R(I�۠I��$I@�,QӔ8��{n~�t����{��Ez�+[������Ĝ��d`s#��[�@G�Ȁ�����IFԖ�%�5�s�8�X�}����x���AA�O01��Xx�%e���!�S�.�,�fE��mM��-/><�ڼ��A��䟧�w�r��z㧯�I�K�� �hk-v8�~���R��?��Sh&�������V�%���b��@���{w��V�jx��:d��)�V�H�(p��A�=B��m~W�ײ�O��Ap��8*�e�53'�M�PQ�u�ˇ�H:O$I%�0`Ρ-��4�6::���̊_�BYz��p���<o ����������������B̏?�40��X�<٪���,Ҹ��Z.{n�?��˪�ɽwԹx�'����NG~�*�c�˿��dQ�@�h���4����3�*(5�2�M�聣�ƚJ��M_p#��Ԕ��FLA�A"��9�9V�-�9�����b�ä�|�Ჟ-@�($�H%	=SlD����"@?JUr|C�cC�t�헋7�:h.^x�U
'�X�<bw�M_��؅c�z����-<�{��N��3��^i���?:�nDds��R�:n<��z�UMP�h3��I~599E����YDo���0����|tU⥖����$H��>pK6��t#�L"�'�ЋGu�����?��]�B�
�����2���=|<�c:ieob�a��/�����0�h�Q�{Us��#����#a#b�->��*a�֎�8Oj@��>�W��c�+�9�������ч���]��hy."y���\`q)���/ 6Q��b(�)�r6��m���pNPV����+d�v��|$��;f�-o�S��I>6��'r*¤@�"p���S}T/i
!���[J+�uS����Q��G�� �t&ob\Q�g$u�����J�|AI�������H����bL����Dեϳ�[z�����5^ �p<�BU��??�Hiv��`n�����ƐP,�a((%˄�g�쩡���Ӻf�����/Gu�T��	;��'�>,C�Uh0Q�Ț|���C�2w�wR�5]VM�<�y��F'���3M)W$Ȉ(���3���/r�n�����-X[3�%��>ّ�On���\i��r�of��wڋ 룷{8�p�g�d��@,b�a����{���޲}��5�ݛ���d�4��|�0���{��U��.����?3jo_;�D*�Pz<-?�݂'��pn��j��B��an��<'�T�7�Vb��2��*��X�>)���H��0k5 ���?�3���,��T�WV�XN�g8p}�7�HA���m������k��ղm@�W�́Q���J,����m�G�����o�p��9�E��z}x��s�w3����#=�'�h�]�B+i�LA
�����;���ٲ��1Na�x�Q�ZD!�J��$�V�L�p'�'2������'[K͏����p��ى�8	�0dsuH�9���\}s��{�l�
�[�L�j�͟�R�-���m}"�/<���kc�����6�X��4.hhj
O�(X��e~b���0�@������vE�H𛍸��Q
	y��=	I��I�o�o�Ā������(|NT����?Ǹma�#,C� )�M$���c�GĚ%Ed�V�N	��`~�0��E���I����[��ϭ��jX��Ga�7�:�������B,R8~�\��I�X�f��.��g`�I1��<G��0��w��i���!����V�(�0B�� >~�Zz�Ę�r.m���Qu�./ŵ6�7s��h���������;3�pv��s�HM�y��wIh�؝%�q�
�i�"V����0H�"��IpP�����9��r������w\!����/.� ���Xb��]�N�2�_�������:�F
FP�FM��\U9cEYN+�a��sV&K�ds�Eþ�R~�q�Cjg}�����K��M9�Y�P�?�4����V:oW����p$�~kH�"K��c.>����Օ͉���L"�/�n"������\ڹ@)��Emj�1�"?Q�zLL��U?v�8q����.Us�r��G~C�,r�z�|s��Pt�*�	�,) �a�����n�k����X�(�F����t9�Rf�2���{{༂�,ڹD�`L��ed�>�W� m}+3PP፛���XA�����j`��Qz�,�h&3-R2���Hi^��%�����
K��S/��P�S����w	��tps��������d��{��;�KC,0�t����%,�K��|�׸��9ژ?��j`��w�ȵ^m�G�:I0�-�{\_����_�)`���Pj��ު������F��+7��E��L��ɖK�����B�P刊D�����j͙��[�ĠD��0<��3'�����>a�a����;8%�"�E���(�x�$V�x��|{f� ~S/׮3.�I�E��s�(��J�Ʌ�i�PO����г�hX���A���a�gg�+���|��j��0��Q��ь�(���O�_��4aP�-9Tйr�^ZٮB��[���(�4��c@�.
<ۄ|?�'U�S�|  ���N�Eg���)#�������;��H�>�r�lZS���<=K�Ld�y�J=rJLD��^gi���ӛ2.[�Coo&/&���#C���GL���`mym�v���u�b��!o�Vw�I��v:k���|P���R���P۞=��m� ��i}-kZ�����.�ܛY�e��t�`���ۧ�Z�1 ��N�@�MΨ��`�4�J�9$���y�6��he���>ɤC)շ���D���CP��d`�I�����R����E���{(S��H9�X��d:��i��	BN��5� ����犄;j�
��}��9C"ݳN��y���nFFs�{���������J\&-m��%tP-���B��;�~�_���i	�|vqqӃ<ɜ��n��c��������
Ώ�M(�vʞ�ԕ�FA�Sl��#h/u�.Oux� �ӊ`��/~
�O���1⾿�_X"H�E��&�Q�5�Ut���iU�R�^��i<�͹��.���,���q_�]���$u�}�-�P|'Rt[�)kϟ�Ȩ�Hs��j}�ݸ2�{�$6p�=��g�Z�����������U���G�d�T~����Ll�=�Tu���f��c��3�<�|ހ�:f�_0pp��k�1���]�4�(G��X��� ���|� ��ā ����|9>Ha�i֞��GRr��B�ӓ�%* �~�c����9��hNX1:@��ptr�h9h�Su邪�:>���I�*�J������}�(Pq)�'����=�h�R�Ƚ�
����.6�s�LB¬���y��l��,+�7yhdm���<<�]�-=�A�����WS���s9�� W�͟���^���|H��������֓�rŲ������|���_����+ױ<��x����V��*js��"5r��z��P١�ı��]C�H�QRp<6St���8����e��g��Bu�A�!�O4e?t-׿��A�.��|T:@�w��$�~%5Ո�6��ia�-�p[��uQ��m�������٦�D�_6���^�y<�;��B��
s���WY� ��Z�"i?;�5�LQ�}��G�]z�dE<�;�;������-���[���U��e�W�M��C#B<�9�"�8'a�H�����Ā ؉�e�\��8\��F6ը!���)�Ν�[��/.E�q�Ӟ(�Cr].*���M3�D��Mu0�ŉJ��?�+d�J4�G�KF7Ҁ��E�F&����&��a��S�s	j<M��!�5^�k&�vV�]WƗHۆ��D�̃���Y�>msw�����|c�����_�}�����2q6/m�et�]|�������3�zs �������u��:�飌�2U��[��"�e T�J'R��3Z{0f�X���Ƌ�!N��TKr0�@����#��4ҷ�Y��;�q��_m���hVwk�OD_U�ihP!,�ڨ�M�|G����x�V�[�Xh.��e���ΊHC��FL�K�Q*t?�7:4�?���	 �;����q���r��K}q�n��֯2�2T�u��K���?��f����k����羐��&ݮ�<�{�6�lx̼��W2E�!<
M��,��x�	ƒ��ɚ�����=��6[��rR��Һ�<��uۇ�����ă�q���Kd��t�ܯ�X�^6E��B��?��f�J����Sb�M�h�'bR��r�c1���KC44������@��A��}���7i'D霶7�1,ɏy�����g��Y�蔙U���HD�x�̈C��(�,�>�G�o���/��v��z/+�D�S/\<\F|�9�Z��ր��|�L�8�'lֶL����O;c�F�!���YX-A�Mz�>%R�"��Q���b�)0Z���q�[����<�8��Q�2�{&���u&��v*���-߷8n��^K���͜5_/+z��!h!�~�#� �����?Q&u�v��ڛ�v;Kc�H������ǆ*���1a���
�%���7�'�oW��gI����ڳ33J���_��C�v��ea�}�^Oy��AmI��_S7���*�ʎ�4�a�ce���a�ɢ� ��-9�FŴ��z��N���wDt�2���%BΰC�˧�z�4�y���F7G���c���!�8	#�"���In�@e�������E��[����r�Iꈛڏ������<s��<8������̿��ս���"e������g�H�6������� !!s�ڜ���qk��G?`�A/e,3Y�H�� b�O�W�}�ݶ���b��*�(!y�!n���%n���p��j�RY��a1XT��MDd#������V_�����/r�xVW�[��3&�D %��.�3�/C�8+��s�����qT�X'i #git��
�!�oxC>������"�)��a�U��m�M9���2^���FJ�cجd+��s���$���v��=��l5����o�#����ת*�k�L}'�sFO���|8Z��0ˀF�[kq��.�� �����ۼU~#!�8���l���pL�9�q��o$y��B����3<#�YO��Ũ��7�tS�d�Q��&���LBtb705�iq�X�z��-6�c��w���$cBr_��8j�a7�Y�/�(+��U����k׳��Q�O��Mӷhqq�Ӌ���-�6�s�<�h��0~*�$R�s%��e�� ��ѱ�۶C�*�7:\E���8|C`9RAf+]@/�OY�`���Go���$���U6�n��XL�@��I�]��)+��X�1��T[�P��4<7�((�
S��˟*Yаp��?�n�}�O����s_��r.�a�4���0z�]�9�:�0j��'�dc�abH܅�?v�>;xn�
�����ww�O^N��S@�������\B]H�H�M�O�0��;j�XL:�z�8ѱ�I�c���'Q�^X��2+�V�&�� 9EB8�_]��%�r4�Q;�l@N�#c��8��	��2�K�x���� ����.��)8����
�����t���8��x�2{{{&P�|�mЕo�)���=ֽ��,r���5�X�� ð��д�f�9LW��3=��>��>o��y�rrrJ���J�X�iJ㢉"B @+��TA]�R+��� �U]_�32B;::�"\ή���VH����Zʬ�������T@jl�2n�\:�!��oVaf��*Q1��/5q���q���[��&7Z��pO��'�69>���e�@Ϙ%�-�[����3j���t�C��:<�¸�g_5q6M���io��w�v+��y��U�O1��0�|��u��&A�!���	�ط^��9�.�*�ͶR.d��W4����sj=��Lf%�iY�0����d��t�D��!Q�G�2
�^q
����ҟ����
<��І�N�f$U8Uj�m?���C𴥕yc�(a�B�F��yj����=�Ed/�7�:�+|޼e��cQe���H��o&�p������8�s��*B/�k�-����{���[���<Fq�Ș��ϲ阺���(� �`q6��un���l�P�əc$|�����n��0�Q}�xcM"�O��F�J��f4���v�#���߿6�������JE6U��T#" ��E,�oV��J�.�!.A  i,R䴄qu�������3k��j秉V��.�T��UM���(������<����]�ZV��rn���4��]���g��!e^�[�+� ��JZ2C�#!���Fs`;��4�0��|�`��B*�wʕ����n����Q��$�'%��v �r�l�=�E��G4^$��-�7��>j���+)C|�������I4��kF,-9��UW�% ���l9Z��[v0��1kV"�P!}�T׹� ���}�������������n���`<�������2Ŕ���j��&���W�1?����[0���J�n=���vNp�5��

�"��?H�1b��[�;�ه���Вd7�;�:|b����Ԑ�zݴV^��z~�:=�L��:r@����0@��\��^�g�t�2u��y�u�5W��Z�֛7(h�s���mГb>&���4φ�OD?��n����bŁ��Z|��\�����寨'��+��P�U��%#���"�(�2�c ����)����n�7b�e&��R�L�l�3q��X�&��s��"�����d;�_)"�}�m�����������ט�+�<����5ӺM�h:uM%e����5���E7�=xR�D[�Xv=��<ǫ�}��E�U�[w$��Ah,����ѵf�ݭ�
�2=��w�����Ń�P�3����^b�@��"1��\aq���X#�#!�@���'�6�ᡆ����(%�������ԈM6�d��#���	�ʟ��P��~;��L�/�* �H���%�BA�bf�����ei'+k�؀K�Ai+�8��4.���1�����	����OF�`�x���f�C�9�<i�5�䥥�����a�c��ە@���~�؎J����_6e _�e�� �g����%�k3�,�J�]Z@!&��ę;�N�A�Db;&ǣ8��5�a�������@�Y�{Vs��7��R�ME#�����'"����k�rX3YB���}d� ��q�XLz���m����0��ߓ��뱦�9�踾�ƹk#��%Zlx֦�Ñ�^�*4��7^K�[ƁY���7�����_�)�����_��������n����������<^{������
\�D�&z˗��A�?���$�o����\G��������?6Z��$4tXᗖ�������f���dh���:%8��3c|���C��bl���H���ʓ���"2��,A�ì�6Db�ىb�Q30eXڵ���wwZZZY�3�#��#��i����Z�E��
$~��	���@����h�B�#9��O���������G�Rg���4��t3}�'T��HzġL�az�R4��j�J,y9��:%�m��0ҜSZ�9t��0����B.OE*�m �&��-���v7��&��~���6��z_���y�tv��jH���A�zGǓW�ۻ�s	zp�/��V�{w��}ͮ��#��}s����ɸ�.��{7�W'�[����v��}�ۤ����*�饩�~����[�p0RR�����r�e0"P|���,	����)J�nb��U�F���߄�?�bQl#��*�d�!�{kubf���"�4k�E���TN�יִ�rvq��AJ��Ri)����r&�O�L�0z�4^��P��l���ø,��w��:c���}�u�S�����ZY]]=�Zuw�{�i{��w_�m�n�/g�L.��kǕq����sc�F���Q�k�s�B��)�r�T d�=�?&NEk���.���w�#i]F�2I� ��Y~"z�Eݬ������Z4	B����Hn6P��ʦ���7O}R�聜�5��n��dQ��8�>W�<�y{ӎ�;�2{��qxÝc]+�KGrCK��j�J�j�v���e�ߺ�R����x�������0��}4��;����l]�o�@�n����%P�H�#a����"b�	�E]�u`x��ˬ�nx�{7}��n�)Β��Z'� ��~�O�1*�V��ɜ�,�e�$T����l#�2���g�h�eO���2�yIzWh�6g5�A��XZ�6�k�j[�{�#~r{ܝ�6Md�}l�����e�mmm}~~vvv;{������p8��������cf6e
�Z�d����ηy��S*b�c���o�8}�5#��MlQ�t��Mtm�f6`X.z�������լu33��$�=���{�o� L�����q��*�<1����v��^cF�������e���{�B�q�@�6P�Υ|@���%nYcj�dp������כ0.�k���6��!2��o�Di�.
��<#��
��/���s_�����#�xI��߿�W�c�|�Y2X��L=�C�SW�;�)܍�ق��ѡPR�
��T��~���7k5YǙ~*%/��l�ҷ%�E� -ZU&�W���Y���.��P��\S�#Diy���t��'�mí���`I���%��V������ Pn�r�?���O�&����j0]Y�_���ȁ�ř��~�w�������6���S�vwc�r���_��6������{�	]yt�߿��:��G�����Fb���'r�vF��S4��+��%�Z!̩3��\IG��J����ym ��RJ�.��/%���8�)E���nb��c+�D>���.�|]^�7�.�k�2�u�:
� ^�!��"�H^�pK���R��(�@Z�����LXWRX"z�i�*x�b{���a�;:$�+����es�"��$E�hm}5��r���usKQ�2TZ"t\TL3�~�Ch�(�g�Y���3�_w�m��lb�֛��C��Y��rd�{KӾ2Z��K��!�����nɤF�6�
����	;<�> ` G�!�=��nڸ��2�����ڭ/u����N)��$-�I댍��o��;��~������&�����<.�T���v���W�¼l"k���㳋�����ʨ6�`�B�)^�8��[qw� ��{qwwww���+R�)���sϽ��#YI��Gf�~���r���o,����W��}����nn��7�^O���/5���|T�DXpb���`zx�;���j�Oi�0�� 3�U��+t%V��"U�y�"Cf�e�ߖ���T�f��6�UU��g�O�9���Z�����4�[q`#i�Aǃx�[��7-��w�ܟv<=o���j�[�C9��Q5��+V*�	�G�Q�Rq6��]�hu�g��i��E��+.�w�E��G��!�	����D�()�}<X2�����܌�q#�EQ��>�K�h�%ť��{�NBfٱ)
��+0N�nyq�����3ŁX�zq2��1�Snf���:i~R�y��P� ����^qr��0��--[x��Dg���7�Y���fq)�x�J���\7}b��{xx(�8\\n�Ă��Z��1\�
��$�\74Y��.�A�[�'N��p�%<�Z��VGՋM�W��P�a�;�3��)�uY%�f�@��T\�1���C��sz�8�y6��H�8��%侓���7���#Q�L�^?�q�>�wx��Mڀ��R`ά��4�S|��c�ة�+�=.�Kb�.z�p�����ŹhqnT�?93�O�q0�'zL�5�)�*zFI���L������Z������s��[�AX�Cm�*[�Qh(D��G^rD�~�� ݯED��0�<���m�)5Sڠ(�|������X	��;�z�1����R��M��~�D�c	��o���,!� W��Ɖ�����+3��N*����Ɯ�rmY��Fȡ��R�,��B�/��/��)sT���Pxd �Y���@V��ɲknx�s��"BeA�6�p�%,�Pl+�������=j��I5��e�O�3�,j;m&V��E���Jkv����20���5�E��<�Y��A??k�H��}LAZv��uWH�_j���J�h�OC:_B�N��FQ�'\������j7D�EX�f�:FYB����n|X�%��ƛ�x���U4�ƺW.&�S�p�i���B �_=Z��[wו���>+�$������}y��n%�������~�6�Iç������&ڜnlϷ���!Zz{rT#c�`״�?<"sՔ� Q��zL2�w�*4�B9��b)ߒh�6DiK��i!0"���#(V_9[�o-���(�C��@���۷}�C��
翬5f��V|�����d�T��Pi����`����(�F�X��X��di��6��:���|�91#%U��R�8|��	�~��N���G�5�H�3�<�q�Y%0��lv�V�?%�.n_z�1�������X�,�dՑ
ٕ��> �q���E����TR�::"���ѷ��ِN�Z�LIb��!F�����C��]r1���F�S܎�������_���^s�Q���TĽX��?��*��Z���){�w�,!�NY�[�A)��}��Lko\Hʼ��y��z%����h2Y�Hؘq|'0ci>|"q[����?���*���%x���J�{���䫁��rs����
�G������*U�dz�i��x��e3J4T�_��p��{EO�~�}+=R"�/iQ�j��ZhΙ��6Je\~q-~�2	:M��>#���cR=����lޡ��J��Vǽ	j��y[ܓ�9�.�WFֵH�ŅwQؿ����r�نLd�H�A��f��W��W3=���X�8��jp��7S�#�<jA�b�%3�睸%�FPUu�tkJ3��<�l�'�~g���}u����w���k3���P�P��x�Q��z*ك��b�������}f��p�` s'˙'�������Zߔ\h:љD��jֆZ0@>�����>��n�;�\ݽؗq���,-|L�H��<��lv{3g��X�Kl�L��C�(c��()��*(:�'�&�ʙ�GK��[�J�����K(G�� ��K.��d�E%g��UkU���	 L!�2�+[]���;SH�%A.g�K�5VYV�ԋ�!BB�@\f��$�|7U3\�F�m+�t�����{}7;�5�����-gXF�s��5�fGo��F��0��u$X��	)��*�D�e��y
�W��h|�i���]zj#Ǒ
 Rd����?'#4Y�,
��v��=-"P�c��|�t���U���.~aiw�?C��SsW{zZ��^����(O��"/���w!7���4��~�Pd'��=&�[ٱ��5�-K�����)�'a!LJ������.��:���G�3����n�k�U6�U~BFQ��R={!=���`8B
�@��@\�l�CL�=&��F<�}sJ6�ck�?�U6��y�5�ԆNY�,��:^����[N�1�I��5��5��{��=� 4��͛����ŗ1w���4K8Q���48����%���M���f�����<�LHI�R�'7���Eu5�̛.gT������r��ҩ�y�*,��2K� Y.��)&����"KL�f�?�Q�T7�;��D�����穳��'�v��[8k}�_!�����":D�hmjc���R�ckm�X�l�ti�nU�w�Ù>����띝�:L��_s��E�N�p��lUH��q_��"ȶ�f,��W��6Y��'�	�W[��4�Q�N�EM�Pbx����Y�O5�zb(�ė���')�Rj�ė�[�L�hnMG�]_��7~y��ڬ������ѵ�����%��nM�͍L(�g��y/���S�#ZN�.<x�S�Y�#$?
!.4B� b�g)}Zf2﹠շ�lv���
u��K�/���j�,����w9c8GGT݆M���O������o�J�+���@�u�%-s��ZԒu�]�E{'�O��W���Im�a��EJ�8ͨ 7�|%:X��8�f���o0�ۑ$��Z������x�#22r㲎�@\���Y�h�w��lY��u��y��s]��LY� M#f�D�y�4ܪM&d�����o��*ť�$Ƀ�����v����my~�/�#:��sM��Ň~��K�dW��U�dx�~ݾ{�~SWw�u^ ��g�U�RH���_�3L�3U+�K�i�e�ue4-"��RN�L�3��^�z��Wvm�d��g\=�v�ӷ��{�+�ץk{��gX�ti~�
��Y�|ċ�ݕ`�t������8�('���ٝ�E1��ks�ÆI$�-:8�ܨ	?$	��2H��0�w�L�۞��=�
6a�,o�ή�(Q��`ļ������V��x�OD��+��e�j�eE�M�x�I㥅� OnID&ː�\W����Ъ��(������u�Y䌶}���mTZ���d�Έ�r�䠋KQ�эZ��V~��X��D�s�4��(����D��:����ͦP�ks7F@�_`�#n;�?D
{����kI�����{R���nI*�����F�uR�7�SWood�C�?z��"� ��$!��o�d�a�]����%�	�yF��\\���5R�p�v���0������.��aLUg77��ͺ����{�!>���:�R���c&��@����}����[���ѫ`�ۆ��J�l�ֶ����z��^Ê�E%B����<Y��9�B�s; j���%V�o�~��tVj�.��@�՛�̢�����O��'h�����n�x-W��^�J�K"Jl�-�N�?�b�i��f�b|*���R�ь���4a5��&�%�|`����.?���[��!�pGb#55�s�J���\�VJ�䥦���'FKh�IC �����{�jI�$�U$��cyZ���, ��t:D��-�a�1lp�q.�	k6#��l���y�;ZPh�`����5GYd��|�Y��~L�P$�/;�å��a�z��,�&Q�!-7��: �1��I��/�d��'� ��SV�ČТt����ʷ���Σ+�Nj���z����7��`�7�)�?��- 2�y��0f�
V<q��`�kk/O�3׵���5�g�ܮl�τW��g�\��0��!�U9g�'�9:ۃ����u]����mB��OC=�=�t�B;r�� �dY���H�7i�/��7�1U ǡ�#�z܆�f�ȸ�%f8�",�#�'U�J�|���zy^L���Ǭº$d�t8*�>>vr^8�n>⭩"�٢�Y�=�O8����
F\�����v)&�E�E�J}���]���je:���ow�f�ϙL$q��>'1yZ
�t���{Sx����Ɲ4K�q��l%M���r�*ܴ_3����=��G���3s���l΃����E1���kR�&��c"�PE�a�O��s;6D�M��z�$7��N0LN��Bס���`[&BQ���I�_	 �z�,I����6E?��v�w�����vТ���m�������4�a�Q(��]�{�r�oZ���j3���y�"~`QL@/l���rI�-�[V��eԧn��}���T�`�3���dEF&Վ(��ݺG2T$GFFB9$�Ǐ-M��m��~Q�FMM0��
��Y,ᴇX�}�V}V�|վxm�{����2�c��7f��5�x�a8���k,�<��$#�,p�������������gܳ�*��p�k�1B��EDx5G,�-��ǐIJ�W&	��/��/�_�N
�;�ϻ��{�P,���Ί�����
�䲉���?6����<�����F}zE��L
�HZd.���%g/�k0���Ͽ�(ө�m�J%I����z�M�Ե�_V^T@)���ߝ����2��}|���3���.���(	���?~�X�' :Bt��ܮ��KJp�N��p3�*Xʳ�ƜzK_g��}_���|�SM!U	:ݒ��xd}]5�~��ݳy�~���:�2��q�yK�bp�z�ǷZ	J�2S���)R���ד�c%a����97[�����,��,���$�2b���w�`��L�)c2	坯4�����}��7���~���˕�Ъva
F�®����U�?x<�U|	���"�
qlY`_�����|��݈(1���k�%fp����]p�O�%4~Yd�5>F���s@����캖Q�E�Ƶ��(�&/��Lr�|�7V��8b��3��`�2NB7�@.FUd8��gSpht��K�
��;[����y�H;;}��w�e�^P}$�ߞ�A��%9��&,m`o����}��5���p�냻Ͻ�&��a,��&�:Fz>��X�yZۍ�˜�����ל]%�A�y�v��[�������(�Xf�>Uה��wĜ�R6�}B���I��al��Ȗp;��G;��ëQ�%�������*��Q�H�t�k4�M!�(*y`���>VYY�����Pܬ�\uP}�^* �4�?n�Q\�sẌh+�u0B�U���5��H�b%[۩X%;2;���Q�F�>��~��E�P�!��<a��k|��#�A��s��AͧpK�9�h�iC�k�����\o�q�x)8����4&K+E4�4`�фz�Lb�ū-*,&(k�ǿM�x{g??{���,���yz��������_0�#��bO"5T�gmt��yFi����y��7K�?r�!��(G+lK����������z�\<��~a��R�i��ey��%sW-�iE?����O	g������D!� M�X|	�g��O �SB31��	�eH2��U�slas�>|�5���Ҧ�>]r�N^3�-&�W�,���������<#+��g�o���N�����˝�4=�Z�q
���J�HHQ��@5=_Z�x
�a)�������9n�9�|Z	�%���P���O�����QA�K��%$ �!�������N�w�94�t�M)�@<��	"Y^�4��fE��Vw��ŗ��Z)�%�ȭ޳�������=�&���L��k{֡��Xύ%�G��#�$T��K#4�n��7�FS;7��ݕ�{��%��# ��/$FnE@���Rp��Jd�����;��rX�t*x���9�`�gT}����4� _����$ID�1F�m]�9��$��*�}k{�K�]�QƆe'�n�Q�}�Ҡ��O��"�x�[�O��9D*���S�n7���d:����,�˖ ���K��r��!�R���͞��ȣ�2Ŧ��ߏXViA�����a�7Y��l!n��U���`T��}E;���?�}\��>��z�V�K�&��:��#�rҬ����v>?����߿�Z�|մ|c\��ĚZ�ƶJ�F���ֵs[Y�M}�o�"�>�!�=L�\^�v�M_�w<����8�T��8�-��ډ�iV�?����Ȯ;���r���`e<���2�۰A���)��.muޱ�c�yc����\���{?��G�":h�A��s_9�_�~���M$��Ѐ\<?�1�Iw��f��}�w����L8cOpgY�0cǋ�*���n��1nY�M�����������m���|�f	᳭s9 o�e��uB��ܻ*x�+�ή^L������s���=mm�<���*���e��4de��=|SH�^c��5�M3CI���{9f&u�1u��yx�,�X9�7���p��A�&���v'��̾���ǯ�\a[|P��j_��,��"�-a�	<;�����	g�7E�2@?!u~]����P��q�/�9���Ú|m��~�{�������%��wa.����&���D�/F)S	U�áʹdJ���S�.�s�]\_��@4TY��E��C�z�?���#��u����ƴ�?�<]��c2��'���t����c����넁��ن��i�?M�ZI38J��V��m�䈇����qz��}m��A��M�r�����,�"�����K�	�%�:S���<��&@����^5NҞؽB�"|f��t*����!b$l{�'U���.$��_nIl��c�Q��8s����Skm��~�~h5}8V鹨�#����g�O"�M��BdG�<�	H^����ސ���-�bi�b��IB�Dx�[vnh��`_O,�b�{)�u�zm^���pj��l^�D�1�'
���954���pĕ�sB�/�G� ��7��1.�X� 
1!Z�q@���T��|�\FǞewsw_߬�e"ɋJ��m���7�-z����{V� 5@�e�ޓ��Ej�(�������ɟ3ȿ�vd�"i���v	+���n��� �؍��~-��*�3k�������_0���D���d�48a�*L�Ww/wLlt�Cֺ���zv0 ds��[Z�k���i���:���992zu�w�(�pJ1�:Ey/ߊ)d����/�߅�����/�	�5(�i{���$��#���Y|�yz1KI]:^���o�(8!�~:�I�2b����a�_�~�s�X��&s���+fle���_Ôo�z@Yz�r��G���������e�|��'�������Ko`h�"��9{�S*q1���@�-����M(�2!۲���}��q
nu��n�vd�Gf���W�G>����3I�=cv���	��w�}��w�5�/K5��Ϙyʆ\Zv׶95�=��!�u@���ˑ�&��?=$�Ҋ�K��T!�����K�Ÿ� �	�+�ld7S	����у>$)-$*,��+!�MG����wP����;�Uh/d�����{7__����$s��&�0�D��r�w��P��6�&ЌcL5pUi�����*����g�R#"<.3�f�&4�]�g"��l�x�@�^�n<��k���U��Oi`�H�!O�T�I}K%�4�yPv@�����g��Yrll�om�md�����3��Zz&��MN�+�a�_�'�"\E ?!$���/A��ļ(�w�	�:����dD�42t�by����jz�����LX����Q�x�g2���GR��}?���ܽԗ-����'�i��	�
���YW�d}8���`
�	�P����|�	�,T@Lk������g)c���!9D�0����T�x#K�P�6������Ŕv�`M��o��(���#�a�f(:�_� G����z,����[�$����f�����~gz/iq�qS�.)m,�X�ի���v���^��Ƀ�z���]4I��kF�oP
�G�	������X��^�i@�¶x�9	��O��m7��^�zG��QM��5�\h�����|;�@=��7U�h�Q�|t&B��ە�vX�&Slp�%�5+,�EF\1�`0��cR�����y:N5^U_���� ��2���8�3)�ָ���l�>}�"��t�'���Y�g���⳩ޒl󄔽�]�O�t�N?$|��
�5,h&~�����mz��.�B�q��ވ@�w���#�j0��.�ha8����X���40�B)���1�?���h,�]��B���6�%��'�|\#�X[Cu%Y)�e�c�<h�`����02<*��J�� KS<%������ Dc��b�-ʯx�C�"V��ml���i�oQ��^���C]hae�aE�e��*�����qG�I��i���x��ǭ�գ7*Bh�oe5ڌ�3,��.۾� ��Y�ߦ��()���.j��7��%,.��.n���V�'�J�8`�D�"�r�1��V���?��ۑA}�_Y�)�`����~�i��;>�ݱ�>�h5���X�ƺ�?m068���of��5�Իܵ#�TV���_�u��t�Z��AT��e��S<��s�	�ɥ�_u��<�N^jǅ�aY䈅����͗�=�� /����b���|���
�����6����A�"��Z�c"Yv��Z15�k���{A1���M�ܞ/ڍuo���҄�J:�O���zw�!HdMf�>�A����
E��cI�೙ގ��q,1��E����N�{��```I�|��4h5N+ꦙ�1Ѣ�s�.�>7^��XU�F���!55cpR�*9�t	�i
��
��GMq�4���*�H��t)�NV�@�Y���H(���r��~�?�M�|E|9{���`U+kh��ђ��!�"��뤷�Sj�=�̺Vm�@���� ��V$V�rǄ��K�d���A���^�V;���\0�ۙ��Da��V�j�8� ������(i�"��"�B�����NZ���c�1��3V.<�/�Jڞ���&��j�㉲��E�ۄv޻�ݴ��HP���m�#��f�Q���+����򛲜
���=����]�����0���A�U�X~����vw����M��!��=�<n�r�����`C$/��S�σ�'�*j�DS��T��QUO�Ĳ42�/㴣��-��N҉_A�D����"q5͐�S��Z�'��.d�G�f/)�V�>5�t�M� 2ϛm�בL�р���}b\׋��������{�����S�.=�������|P��4S���ע/��_�)���Sj+@��a^���,x���4��͹��@���!�I����,�YX���Œ(L(T��^��MF6�Vj���|Q� ��S� �綿]�����G/�/4Yi��gI�Em�X��x��}S��A9��'_�����C[�7^�X�\��tU�t����YCW����Q�݄�<,�%µ�+9��-z_ѣv<_cnaX�p��Qܚ	���� 3/o��!�R��d�^���-�km}���G��*���(/��b��N\%�:$��i��2�,"�&>���!àd�>ގτD��:�:���&:J��9~�? �b�?єD��l;��;�F�  �xi=ǘS�v�[x椏ؕGW�w\��P���,n��b�﷞�`���`��c`j�0�J#$����`�$��U��E�K/��7;Ȯ|�^�\�lyq�N��qtLꍧd:{�����?�r��4���wx�S�)�u4����=�5�@L���9-����3�z�,"���n�c�8xH�Y��NXm>IMܚ�7�[�����2�5�I ��ô�:JXF:z6	R^^n���$�� |�kT��pp0
�lvt.�(I�%���!_�!�n�}�A]����_5��Yn�����g��B�|D�Q�����edƋ���/	�r��=��- `3'7z鴾���A�,�y"�[$�|��85?>F�N�׌�JX�Ɍ�erxt��B3���%�K�s�7���PY��������lv�[&;q� [�,�a�ڣ�w�7�eÓ�2)8�6�#�&�ʈjVN�/"��E�ܛ���z�����R�i97%�*� H��G6j�b�]���ڶ������Ӯk�w�vt<��nvol߿�-p��|�ɫ�6��#�����tB@4�8v[��R6*� ��j.U.��4cY��P ��f�^ž���8��1>��A��O'�"�������G�r������?&����7��=����G���|�;��x�I��"��h��ͯ����TN(P�?���!�`�#�Tt��
c���a�/a9k�@��ZV�^Jg���5�Z`��L��]�^pr��]����l=ʩ�$?zqDO8D������Ą�W{�kT������X"���K۰f1�0T����<F%/.�k)�g��I�CY�]>S9/���D`-H�<�6	�8dٵ{�t��뾫��T��^/�����:����Տ��Rv�CCA��۠*Cg��l����?8	4&
�g��\J�hx�UȔ���D���ƕp�h���Aɔ�
�
-�,��xV�K�(*0�x	�����}��F�G���g J��!Fƚk�O���/ɻ�d�<��)}R�,{���i|G���<6E�w�pA���0���y1;I�3�'1D��d�.5��0��,,-yX��оh�A-����阙k��#ԇ�S��}8>��Z_ݜR��$�Z̜��4B�ڋ[�(2TB��mwp�C3A^�A�HG�blM����i
1Ry�F*:���(1�3"4A$����kv���>���,	����K���A#�����BϨ!�iv��Z ڸi%�Ŀ9��u�]�ο�������H����;��V�?�3ߍK!׎AQ7�6(M;П-�L��05��Z8i���3;��	��#U���p\������_Sȫ���.�c�L- o�p�+�L�#Y������Vqp����_��<�%�)}��=(@Ɍ؜ �����[D �t�J��ٝ�[����|�޾�ҡf^+�����k�,cщو�:�'*{�����⪧[��m�6Q�Erb�q'��h�S������=� �$W:}�_�@T�R�N�¥��<����}�\�|��ې�{1���=�����an�d�����y+� ��<ߵZ����9����GR]l],�!��wauf6�/��Y�Ȑ�%a���x���1X4��^)�c��JYb�Љ*�6h�\��E>�tlb"?	�W�n�-�,w�Ai�@znn�G:"��"�����{�%g�.iv'l1�)z�)�ڏ^csw�B��J na��H�A�g���b���CI�k'C�,"-mH�6������q�T��(�2ѿtyy9��_#ܗ���nR����߈��	�7��A6��u���������CS�t����|P��FY�Tjq��q�fD��f�{~D����'���u?g��64H��<�Q�d��b%��a��qa��T�����'7��i\�Q�W]o�E�+���= ՍD�j��҉KbS<;�y1�T���l�2T�7�|�˕�p_#��J���紘�h%�����JP�3,�|�V�WF}�<(7�!,힁Y�4�z�_���:q���,�EȽF�A����U
��DD$�N�TOא��$�4@�?@��A,�
�A��rb��Y �_�<�
Y����O4��2^��'r�_���.�'''��x��\��C���cGaA�Si�\�vk�`��a�Cgl��ؘB�͍c��� �k˛��-�<u���N�^���{��:�A�8��6��Z���Pz/���˹�GB��E��+U	�B��P�(ˆ/��
�M���鎐q5��I����Kg����yd���I��ܮ���e��R�� H JC��Gˎ����!���0K�qp�V�5�N�n%�H�p���=҆�����+ot�*,iXr�����ӊ� L�ϥc�8���0 �V{L���)`ޡ��,�Ư�|(���v;�u�x�@)�nd�ȷ{��s1���k���L�|�Ko�*��v��v�[��-�C�ahV$�Ǎw�YrIC��f���A�DN� 3�;��i�=B7���-���E뿹Am�>��]\X0tuM�X��<��@��ؤ�E~��V���"ݘ�߫J�����-�WNs�S���R~0�@^t���K>� M=�$�p}�b�\A�^r�@���
�A� � �a��{�g�A<F]�P��L�����w��WF�*�#L�tMCd�8�r¦����.!�cbݭ��L@��)�?�
�ͯ�E�v��Ξ�[���Bs
��r�D�,���G�����?���&s�LL�[RԿ�~ʫ���ہM.�?C��������˓l�!hz]������`��o߿a�����JU8�Q����-B�ĪTC!��V]{tu������������������/)����3H
�c�,�W�K�݃k/~1�E���<�@��J�iz�#'CZuJ���o��SH��Ĩ����&�Sv�(�AP��'"b#�M?u�v���eW%�����G����Ǜ��U EI�z�K~�uF��+�T^8���]1�Hu-��d�r	��`x��4��\}���I02.������Ӥ���J�s��g����'�������D��!l�u�ZZ�3���`�,�pA, �d,��,K<�[��~_��`(�3��$����\ĕ������C?���y��j��||z:sv��ťoe�������J9��]K�M����ף#�9o,?�s�N`OqЛ�� Zl{��`N�gs��k�`�����CQ��}�
��@8I:+�&����\�9{�_K~�HP�E�>a\K)�,|7^}c�/7>*��J˘V�5�a��k��,e�����?|���"ȣ��[&;��<�����j�be�#����W��l��}S�j,�g,�R���PR��x���sZ�7v?ӋӒ��g�o#�hЀ�g���7|�H�����D�&D�,l(R�a^�����X۱�n��ލ��l����+~T44|�Q��Y�����,��ߧ�i���$�6�[���J1��N\b�s:W�i,�,���9]�H����z e�\="DIx6.[S�L(����.�HT�_��BJ��M�aeyD}m����\��(�e@��T&�|w�����BH�M��J�O& Gv!����5����SCC�Oe�G&�]n��x�9=����w]��wF�N��?�]z�������mhlF���c%�jT��.�"�Xl��ٿ�U�yt�-��ܬ��zF��LNMat�����3oml�mo�VY��9��h	6oU�k�f�W�ͧćq&#�By��,3e�z�M5��R�YPb��W���Y��5������h?�t�Py�h��T�L5��9N�����-z: (Ѽ���v����v��%X=�,&��1�i����=n��z՞��!҉���,��	UT�LM��K�;���%�K,��3u ���7��{)>�%�;`08�j�UPG�6��6�+�F�y�u���~f�.�l������He�?��27
�J`` ���۠�\\]H�X	�hG3
�0�ɂ�ҵQ.�ɠ����,��=��_d�9Vm\/9H�yG�Y�iE�r�c]��Ӎ���¥3d��2G4!�	�F����v�'�0,�1;D�*HY�z�f����Y� <�� ��u�R���T��S��:E���T>��0�\R�K'�E�#��[����b�4^�$F���-���3���ɱ����z��΅Ck�	�G�-����N/:�x(�A��؎��uBY+�7���E��~3>��[��-c���23�W�������v�����/;���qS��|ĜX��4� �����,G:O.��D�E�S~ߑ�e��c��I������q	Q�k�'I!J[J�c�3�����[�&f���a7?�h��)�!I�����q�C��h�#��̄�4�hD��,p"JQ����:[^B_/l��^�ĭK���6����7����)`]���k5�̜&�h�1�4�=}�mo��o��ӻ��_cq[�0[����fa�oh������r"�ʩϨ������f\9w:֟m�����]\nW\mc��]\3u������J� X��sN�O��x�[X�~�l{��|���1���6�l�/�k�E���)	�a �_����r�Z133�����$7���N.�+�U����*����y�+D�W���\La8$T�x7x�b��i"Y��/��n��W���g��@��w^I̐a%���p��6f�=X�=7x*۩���c|��Kg�J�+���̉��|�F�#� }Ù��5�p�	[�S툨 '�1kEۈ7o�$�8��ws�533��Ro�xrLt�X;o�����^qe��� t��l�+	�\���u޺f�m8��x �]�k"�|�*+�Ep��Z%�$��вl��2"=_�uhH���J
s���͓��N󞽉��8�$E[7��p�n���_��!Z�C�P]:>e�w�),�bR�&���y�,4,�daPD�V�����'�;�hD� �\�����T��Ld=C]cc_�c���x^��ʣ�ȇ���h.=MM���4���;������%��9G^G�2_����y��.�X���ԇQ*I)�G��m	)��h��dQ�(z�"މ>q�p�
������?��99ƷFd��N��N�1���訵�:������yE�]�X!>~����ٞ6�`H��;Ƕ���K�6�|y�-}앓i����j����n�T`��Ǆ��i|Wo�t�lH�:+;{
�;�=�I>R��E�P2	
H�6���5tK�Y�AGʇO殡4dXK�:'S��TI�dR|�f6k���$Ag����[�Ò���5̌�+Md��D.���ɐ�2m|�k�`��jB�є_�h7<���(��{�_$)��)���w��BB�s4|俜۩������"�f*-yR��0�>FW�/k���>�ǲy�~������q�0���+:�77rT�WrT�#^�"y��b��^QR�:��i
9IRE�X��|�l�V"zn;^0Fx�.$
+�w�_�u�]Syo���s���99u�����pX�
��,#k�AT2�q#����ETR�K��C���Tg��N�M����V�����D|�q�Z���#��_Jum)�J��Ju�Y�{<f��3eԔ2`���͗{��Qd�ݧ��H)�m�>���01��imh6A�G�.A�_	^�GL���cT�J8y+P�c`��q�*�������k���������!8���:����^��~:4b�/���׈��[D��/X�1y��xs����4{Y�yTzZ�}M~��}���T�Y�I�|�.--��ah���-mАam�9� �H]�m���[�1M2I��'�!�g�Ũ�6�Q�9���߈NQ�v0٠�ƷY�h
C9֌�) m/�8z����I�ّQ�3`�o�������������r�*T�7����}�����n@9�u�;��9�֊�N#���_b���S�.E9%"��S=��F�P	n;�]\�HBB@�HJ�i9�f���kX���-_w����#U�;[��;Cv��̾s�֤J���&�q�:\;�&��!�Z�R�|��BT>a����Oy�쾸�\��a3
�w?��q8����8v4�3����]|�ҭ�s�nw��mE.��j=��2�=�'CI��_7lĖ��^�,Ѡn���(�,�k�p���8��}h�ɋ9#��gTw����ʂ|��^-�2�h}�Y8��+��`Ay/�ǌ�/��P�Z���U�UU���Rf�GJd�Ē��*���Q���^��9�0E��� |�I�U������%�%���������%$�|�w��<�q�-��4� �2�E�c\5U��	�g��3��2G���v��S���`l����"�r7z�pd'�g�k4#��$r�6~���$���y��}�H�����?.�l�O��a�]�H	�{N�/X
��Յ���j�`��2Jّ��&��ۧO!�Hu-#���rm�B�>ďA�'s��8�u��p�1�����͹��r��Yj�|G�u�0��1MTi(%��_���T(��ʐ�>ME�5K���w�]s d��2�B��0��{�ݠ�R����BFWG����U�]����󷻆^G����r'�� �>��2>���x�+���3���.^ໞ����n��a��j3j0�.ٌ���[��1��
��
S��c��~� )�"��9�ttԮ�l��W$�aQ��r�%^K�����-â�va�K`�n��z()ip$��������KB�n�.a�o|�y��|�g�u͟��}�;�Z{mc�L��o|�j�Q�mp=NK��ﭳs<~�p���~�k\-�Q�k؆E�{����o�a�?Cz
A>G�1�Y��/M��X��"۵V���3��9p�/����*hR��	6�!�m�`{�c.�{�=��M��rW�v��}0�gڴ���91�"�p���PB�Vpm�XS�.N�%*��k>����?dF6ǃ�������ȫ��y������۫��T��[�K$�?�-7�w��5�St���ФO���v���t`�P��b�_���/���χ�X�R�/6^!e� F������W�PV��9����[O��G���Dr�^+���s�#`iv�Dc��q�)��R�+ٳ�D�z�ߞ��晥4�\����JdLm�� �>O1���d<'+��ژ,�UK�{�Sk���-��S��5	�T�q��F���QV�U�!?�{�m>�߭d��Fa���I��з��^����D%$#�E(VJǳ~ه�]g�Ev�/u����)��p<��w��ظ'���sy|�zm6l_�p��i"���$;;���a�aZ�*��t��c�S>xd���?cB|D�V�18����I!�����%]2�9�r�o�(6�aj>=�փ�ʧҿ�f� �w"ӧ԰�Y����C0v�S�1�_Z��{�z�9�#���ɨ����3|D
��y/���� ��o�� hK&&@訕?8O�>��ڭ�ŀ��"��/�9t�ԧ�h�e�^��} ��t��#C��bv���Q�� J��C�uJ�pЙ^����L��t�T�~��SA��0��%M��{�2�^R-�n��k�Շ��0Ҹ]"�M���.�[�Ӥ��� ;+����|_��k,�
E�=s)�c`fE�P�O��jb��s�C��y隆<;B:/��K�P�W��sQ��_����wc�u��Z����K�Cc����փY���r/'��/�e0v-�y�)�ȑ�>�V5O6����q�u�<����~�V�Y`D�D	AĢ�گ�ҋ ^tڐ�&��4U�3$�0J&��d�Wҕn�i$|�)���+A��G��ǃ+Y��oke�Q|�l��ǔ���W���u�Jh�[kʗ�H�����f��e;��V������ϵ�])��ҌFop����&�!�My
�XC�j�{�Il4@v��	�K���گ8C/�ALJ�$5�u�l���Z��8��}�3��.�5���=��_���R�����Iۘ˸�iRp��3ԟ|oM ��SZW�O)ks���)���7Vןn�/�~=��]F�,�&e�hQ� [��d�je���"��s��t���,�u�ge�^�P?4!�� L��#��ٿ臁#�eeq	C�s�?�No6DST=y�H׉�6�'P���忊)P<+.���[L���Bo����?�D�w"�-ڏ�ȋ������1��IJ"%$̆�4�5��麶��d*�=�����7_�W+|����C��/�P�������p��{#�?�����67J�&]�d�zs��fp,���KE���Ek���ד��^	k��j�b6�,�dfL�_��o� ������!���e������0� 8P���2�I�������mn#svgVQQ���V9�(o��&�r+h�X��b�����.]���G�e���ϯ�k!�*+}��`�b#��Tp�}}���1�)����ߋ��~'�k�k[��9;�]��Z�'6b((�ü����B%��[���������S֋XG�dШ$�����S�U�fFNCs=6FX��	!�Y4�AQ��&  `�ha�Ue���i(@�sue�'�`哎=K�x��R#[��n�;��(q��)%��E��q��[3Nw�SK�6(B��}�?SpxF���aN�μ6$�A3��g�
��V+O��T�ZwK��� �f�g^�pe��@�<g0�{��:����t��ˌZ/� �����+D����b�Bj�C_�y(i�=��xG�x:�A�q��W��d��=	�������3yWGu�=�s���7f]���8��SԻ��Rk�qN���bq&-cz�غ�Ef�;��RUJ�ؠ kur7L%{���)G��[�~XELq���~�gq��X��#����%Ãqg�Ld�/roq���T�A �i������W �Z[e��P������;S"�澑�����*���
nl�,�������q�T��^��Y�_P�������N�Mm[����y�
��}�Ey[h�[�K�]�{���/#�h~����l+T���LˢuEE���KQq�ͳ_!N�St���� �9L檐�Pw��)jP��L�G'�T��K)&q���ʧ��L3>7����X���s���@�Uᘁۙ���}C^����i�gP��v!����e+�A���k�A�Rx����oy�C����|DD"�.O����ܙ4��W	�Os�RX�"�姹�F���y�r`#8�H��s8(����h�[����ͼ�E6�S��@�݇{�[s ��P��If�瘘X�ږ�Yl\�)c������n�z�/����F���|ƃ��D3F�V{m��T�`0�@|�=J��HV�E��=�B��wd��{�<b�� �Z��w!���:��,��NذQ�Y�`D�+g:qA��`]+7��o�ߥ�C�]���-�wv�|`�3C��~\�
Z����������u$+�]�tP��{�G���j��Ԟ�jf�K�O�)��O)T�^�̎=	dPi�.��Ț 8�$���58.�.k�H�1��(5�S�9��t���J�]z����J�E���F��	W//7ǀ ~�w�2ߖ��9�%%W�		��W���i\?Z��Z��N��1a�1��QR���]��p7�d�g02Ɯ+�Ͽ�K>�ciCn���r��n�-�$666���&&�!�?-� 71�g��^~�<`�%�U��ux�
���8|�g��)Ff�?u����u�&�p�۬@�9�ɩ�����p�����|I"�# ��O��Q Y��Qϛ��w P�NH�E���d����C�c�{�y8h��E����>3�]o���D�yƭ�|��n�c8�������s)3	I��THUG�d�-]�{�b��wuo�2R���\���R���)E����(8̙�U,���j�|�j gf��ޮ�{q��wK�I��ϕ(;���L4'�K]�a���� T��3��0]^AIj|�%V8	5:�R�w^��+�i(��C�J�11�M�q鮮afCJ���p�d.�"b5�/����$�em��s�# ��`H�v��)hN�� �Kh�rIQS3na�J +E�����~��� �#�B� v�l�זE�D���D���۠��B�y�Y���$\%�L5ߜ�k4�����iϲ��A�����΁����?u��6���?9Il��e��@>��WO�TƈW<���γ�c@�HڕC�郬)���s���4����+1�Y��L1J�+��=���j��7�ޚ��k�h��j����'C�k�<�P1g�v�%�~�ER"�VA�,�dR�ܐ�.�p��W<^�������Ƞ@�t
�ɾ��'+����(�*��*���Ąv�\򼁿N"�}Tf������C�l����N��*H������K�DqZ�U7�#ӧ����X%�,�  s� \_�5SӪ/J�R&m�������%!�������������P��e��Oz�ߺ����`�c�:�E����<�C �É�F1\��恠W��r��50�j���h��_���g��c�����B�W}������|�]]ʺ�
8�� �;�qg.{}?A	/.ݩF��D�zO����/�6�J��ijѡ�J��Ƞy�G_ 4Y���j���{W�b�d7{7��t��?����j��y���>���"P4���O���KP�Lk��vXP�[S��1N/^s�vY�"�~M����v�|wY<va��Q���]�[���	�#�\[)-5fH���7���&��|,l��`���Hꇃ���ɳ8T�
�x�J}B�ܳ�bU}w��jTTK��ڹp�eu��0T�m�T/�eO"޲�(6W,-�q�P���_6^k���lq����3�Uׇ9L���g��f߂j�n��s�7����R�*x腠m&x>�>�� ��*/*Q��n�ї�|�ˤ���~�����09��I�����o�}��-���K-m'G�Ȁ#�-�խ��j�3%X;�[�W�6'�aE�w��k�]Th��� �����P���R�B�C'��k�C>����U�0�e]������+�c��*ǤOg��4.��מy�, X�������>�5�WX��U�Ol��y����j����j1bD4�>u	��T�Op~Y��l�&��t�@���F$e&V�gj�7-��Xl��)m�71`�`�=����Ic2ے祹�x�QZ/p�/�z��s��H��6��&['�GC�w��v�-#=��	�U/��x5��_�)��T���W�1t�[��kx���w�m�8����t_O\"��������8"���?��1����S�j7�&��m�@� l���'�B�sN$KlUgQ�֭N�8 �x{ߵK��o^�J�������Dl���@K��C��II K�J�ty��o!�w�0(�տ�%��
��9�A�f~��a?m�ga�\�qC� �b�(�"�F��T�|F�K,�rC�S@[AH�������Q�L��������	���j��,��)K��������ͼ�_���
���R*�g��ח%;j�\za8tp0�:��f�F��g��*s��«~�N&��5��$���#��C�j��=��s/(�_pүZY�F'���	4gW��7yV14iAw�h��y2�0���}�/z�W����wo䭠��.Z�,��X��3w3���Z*�"�n%ܕ2s.�ț���חh�.u��J\����z���P�Y�+���o�}Z7�P�������l�3�mk���X=L�~���X@���(C���G>���BW�Ș�D_��t���ǿWŏW]��vݑ6H�s���챈��9S�3))'���_n��OW���}$'���A���
�[㺍��ب�wO��#R���!��C`����������׹��)�m�Ta��Va4>������h�B_�11��B�|���{ӯ�i����O���1W��)����:�K�胿����D^��|o:��l�Zʩ�����h��ݭ:T+�;A�X�	���%/���L���|�KQ��Gi&Ą�̓lJ���+'���F$	8h�%�ĳ�y�t�xnD�a1������dn��>����o��S�<���k�����5\V!g��ƅ��;S_�i���=O��䓼ɒC�x��a۲n Y?��Ԅ'���TY��y1-0u������������޳ut�{��I�ߌby��)U��:zg���n��˾�T�v�y?;f�@��l�����Z��@Z �BMMD*T~z&F�:,o�6n�-D?��z��U8u�ʣ������CC~�s%E�#D����%�ܢn*�ߢD����ڏ�O��,Dq�HO|�c�� :���퓈�Ãϩ�8aADȦ� �ǉ�c���@<Z/P�ղC�ܜ��������Ǡ�������8�6��9b�v��&�+ n��q�w�����%���_�9����
��b��B�L'�;�$�i�?�\��x&��DY�c�ax"��c;˥�Q^-N�Z^l�Y�W��.@��.#�E+TOO����82o���Nzα.�@����t��1�U�b�M$�e-��(�L�j �����U����y�q�
��z���Қl��C��u8;+v������w� ��k�+8�]S�먔p�?{����XT��3�����6ֵUdd���
%��Y���a��h��.^�x,�}�~���_i�E�9�r��r�v����wdi5��%�fH��O���@���B%�Գ�ӵxB���RWZ����\Q3؎\?���2#B�{�ʉ��20�nA��S�8���3�:N+W$���0-BN�&�}Y��o�OM��
S��"�J��{�|����f�W�dճ/���q�7^2H ���+�V���W������5�BD�y�k\ieI)� h��G\Y��q������,g�!o�!�eL`%���ctp0��6��� ^A��V���?�GXG&8Q�����M��8�T�=��1���B����_�we�S�AJRB;:��-���cK��f���!��Q�DH�	J�V�u����:�͌��Ғo�8�9��ng*l?fP�I����ık����i��Tś��N��Sz�n�H�D핉gR����(��۽^t�����ړ�Ӝ軵G9�Sm$xEV��2�촶���[�G����{��M��/�ဣ���E���lpn���ްFV��K�p-�Rw�e*}��A�TLc��(P�Ocl`�bq8��zUPM*:�Ӑ�=�#�&����G��H���St;G�ǉ��"/���@;gl�["�b��}A@�M;k|7���U���:���P)!f����;��K@����x��#��1*�������_NϮ�I�p���"�����n������t YQ[�����W)ۋ;��pK��j���D��L�O��Ob9��֣sB_��+�ڣ$����fz��Q\P4Of�7�yX�g�dע�A��.�����&[��g�� �ȼ�a*C�1�FVŒ9���z�)6���OK?����>�.�s�Ev��Ĕ�V���P���PmOk����P���V����s��e_Ә3��������&�u}�.6TXj1O��b�>�E嫼�V���*���͊놧�rU�K�WP\QH���_�w����>���릔y��	���ѣ���Z*uj��3�_��殩��/�p\ҥ+�K�l;�"�XS��'g걪����tC���ne�W������8��(��·����".D��R������S:����Op"��Ɉ�F�t�b4���fat����TT�n�L)�KK�4�:$��*F�%��c8L��zI����yp�Kݧ����IH�'z'8�?�(:��}�d��k��%d�Ƌ�$�$���ߔ����S���p!����o�L*c�@P� �S��� �ly�fIq�Ƹ̩_�8�j��,��3�3k�"�$�
65W�5���N�3k������oGx�0d��wx_��} ���O�����3v�O���n�\f��!j��������;a��m$e�1�/�?�:��0��Q@��u/�`v�7M�gtYϭV-uZg�
8z���@h q�~�����I��Zh���jDf�|W�9D��c��K?=Z*C��I���N��X�&4�)��c�lI I5���P#�C���{�I(�����/��{ �$��K�G�|�y��uS�k�xȥ����1w�߄� ��V!�!O�t�Ll��m��f�Ə�v����-3�3Ien*/�4~#��R�	p�ތ#����9`���7���SG#��|˻�����F4�������%ex0�$��u���֏~���_��>������~J�|��o�I!�6�MQ�BL[8�)�w'f*�s���ݿ0�ϓy.U��lň��ֲ*���8RC�M6/������m��z��C4�����4/lGX���^l�P�s��>|c�fF�N�N'�z���lحUq�PA�e��}: ��l��//݌FS���טL�a�xZ}bZk�^���F([��jytV��֯p��ϴR|x��y�>[U;�?�!���7�U���m֮9�D��ʜ�9.	�q;�C#�#Y��8Y��i��3��+ȑ�|��i[��������ڱu���m�
>��6�K����@?e��W��Qr-���avM[[0 (��g�[�H�u�����]C�S��k%x��s�� :��������Dk;�����Vv��c�y�$n<�/F��3�)'�~DL�}�3b�넵�ܮu4Q�~SR'{���ފ*�1%/�)�����X�8�f3���e�ŧ@+`g�U,��@}w����K�i���7��C�]�J���P�JF1M�
�%%�~�-�Y���ز��k`�����b��>Jm������Q�ʧ�@����Ǒ��+%�`Aj^��=xi�ѱV@�nם����jwս'Һ�7���1TYՕ�#q��#l_��yr�Sqa�����J�f?�f��?�)f6������iol���<�g�u����D�KF|�ˊ8�V��"��;�xM�Ex��3��N%i�3��03K%]�7W}�Z����7%�f�D�%��^TV�w�Aڟ]uB2kL�~�
sJ���+�C��qd8l	˘@���L�N|�jL�4��u:����i=�$,Ƹ�[a ���B5�����3���Sl^�ϩ��_θ�Ru@�v�?��)�y�l��
Z�iX��
y����ƪ^n�����J�3��1�j��ʅ���W��r��* ]<_mG����=�a���,�/��OT뗓�i����o2��?��HR���`P�Ή�/Bz��������JA�����.ףl{�p��' ��2�*���Y��ٞ;�H�j���*�>�,N�c/<M����x���i*ԭ>�Y���pU�om{��ᇍp�*��$�l�?��J�ԧv{@4[� �݆�0�HA�-�����k55Q ]0~`J���饥�~�+־ ����W�����#�^Y}��
 *��8<��T�M����S[�!�ʱ���Y�"�?��a�Fp�P��}!�B��'S��s��9r�%~�� Kʣ����O�gI*�O�m��k&\���\��R5�s.��B�- �4��*^��*�@���^7Ӛ�s&�w���GZ�U�M]�P�Q�k��>o3?�q��9�
�e?�aҢ��Q!g7;N��J��\r��MWd������X��+S�ߖ��$O~��5]���)#���p0)rr����(9�~h����Zk������\�Wd�2�
���5���=��씱�:�ƭ�k1�+U�t��P��a�z=�֨�G�k�V�pڥcUG���S*��0
�k�EzM��!�2��S7�o�[d�mQ���I�bi �I�Û��F�E ��\\gV	t��4;ᬳ{`Ϩ�%۷���ǖ��c�oj�S#�MRȢKN�E��*q"@�pD%�ѣH�nB��$p�Q�N���m�������d��HRýi�����[s�_��g!��n��K^ޝb7�\\�D	\�)�t�p�1������&k7M ��z7:�颍��&�u%F���x���h��ܹz�ʹ%X��η�����Wnf�U��j�ǌ�]	��ix�㿽���N��#�'M��	��g��R�%:=m�����Ȓ��=7H��)�,.�ޮ��U�4�6n��$���;\���f������~�	F������R��7�����-�f"�?���{���) ��k���Z�$3���%����2SX�����J�tw��#*3��~-��n}���ې���` ��!/["m��e���ȧ� �۵T���O���:a~��v�sT����d��ۉ�CU�D�x�}[+�؇+mߣ)\��[�2P�`�b�������z*u+�k?�;*�{E�V�a4����e�lK4��5�_��p�#�@�~��Z�]���їٿ�F+9��x7�S�Xn*ɖ��[��J�C��,�)����N���<[��	H�=�����r
A�t�m�=,Fqq��}�N�!��-x��J�;?�m��$I(��0�T��2���f>G��ҥ�=%����٘�-�1,���UZTD1����<�W�db���4|u�\����Fb���=:6�Yi�1?	WS�]���)d��@ǝ��� ��*�ͧ���7G�j|]26�+�f[����NH-~-f��S\�Q�m�X��&/�+�ǂ�3����d�n &f��{����e7���k�����K^���<�A���TS���a�'J��CD����l&Cc�n03!��R�Uϑ[6ǥ�����@�v0g��e��vN��KN&��JW��@��H+�t���O)iV
CE`�F��,8W�� ��,�v�T��f1`��L�鎒�~�cU��}~���F:gKE��R�;�03�M^�,���hlW��
5�t�[�ѹw�Iw>�ѥu��EK��ᅾ�b���Ա�R�O�����64�&s��9�5�l{

�4w��uut�#�	Iض�)u���Ր]��kT�h����F����},p>S�����<j��g8ă�"�y[��Jaj�U�^�u�+��������=���se�ڦ�wrR U����6�Z��NӋ�<��'e>9K�c*��|'��4O���c������2��2��4�̲��p����r�~Q}&��� ��$+{�	�Fo�8jYE��o��t�?+�
�G@e���JLq�PZ�����zif� �I��!\�DɊ�.�C��6��j$� ��:�SoQ�(�����;��*,�V6�Ƅ�Dmo]�a冓G%����
HC�Ҡb�� ;=�1+����n��[_��\�@�}�c��Rx���9F����ǭ1'�� Rh fs	Iɷ2�Ok�T�;�+N� H�]H\9&�*+DV����%�}}��9����'"�*ғT~<+��9$���ù�#���"�{��ØG�)��4H�匄�\���|}z&#��0�YT�0^�EI�N��;��m|+��;���d�R3����2.v���ђ�q�D���)@�JXO�/�rv�rrG�7�R3V�n���o���^mw��?�Y_��3���d���%/�x�&չ����+����)(9��C���6���h��|h���M��[s�9FF��L&��xx
^�`�xx�[v��%[����db����L�0�+��S��P���*д��6�P�Rc۞�����jh��]
:���Ȼi�&�e�d{��E 0�x	�*�*>"bB���������n�Τ��a��T���;Wפ�Y����_&I��aH��ѧ �����Ug\��Pk�}��W�,#Ι,# �ns��>/`�$ڍb�3��NC6�f����x��ܩ�0ù����|a}ųJ��X�SUl��%�e�ߝ}�ennN�� ����z� ��M���ѯO�v���Y�?0��W+���ۓ�1��p����HTH�QA����/�{�嵩od�'�e�M��)�閛D�(��=<<�3��H�ҐO/b��w��qۻ�U/�u�f�o�*�S�VHHfU�"���xD���$�<\6�d���f!��{�c�bm˱r�ѧ�qvM��p����WF��&�W��O~���*߶�vΥkr0x�f��`��I��sb���:�&�|�O�I��7&��i�,�٘�.n�} �����8�⨻ �
�is��1�x^r���AD�T,*�uxz�}����|���o��:?Ft����ci�B�P������1,e~>�<,��A�Z.�yH�uL�E/���CU�v�9y��u�rh^��"8q�Wu0g�<!�����jTh�y�N���t��bC�eg��y�N�V�$i��y��>����ᙈ5n��Z�{6m'�.���[�aJ�j'����;oU���h65����u�k�5����5��DG���Ɯ˫�?M��O�(���yJ5���xY�H�F�=��R��~ہHu��QP|�Rl[��R���!b�j:�F�Q�6�� �#V�S���3_t|���i�m�Ο%��>-��P�S�>(�cH�]��܏��s`���;Jql�d(���:K04���x��� �%���[�)�A���x���:q����P����sd��]�������#WM7���ڪ�٭?c!��`�kx�YbS��:o�m�����f�����k~����i :ʚrS�K��Q�F5"��e�Q�N
	�PNű����֜6l��V&�
L��|��-� �v�t&��T8F'>yv����ނ��M#�K��b�"PT!�t���Q��T1}�'j/���kGAژm:�.u�3�h�g���~luzP(R´!y�ݔOm����ąA�.��--��=�X#������G��~m�n��ǥ>v�>mmmd
(���1�}��ퟗ)�w�!��yx|�m��&��Ԭ@cObR�R3����������|�2� ��*�G6_um��aV[��7	�9*�/%Ȥ���I��1�I�)qd��qk�m՟�H7X�!����·���b�w w�wBY��Տ���+�6�|��x�?�#h�TB��ɞ�M�B��'<8����z���^=���R˓8C�?Ċa��	*�1�������H�er��k����7��@����H D��5������d��Z"�J��%	ƨM
:��d�b`�3�	q0(P@`�I��n`b��+5�D�
P	>�j^V�{m` �C �ќ�?z%|~�r��Zڐ!�ʮ��>��?͹�G�8e�Z�+�V�>:99���`qB��^D�p�W��V��h�Krg��D��K�{���T�2!��}���c�Ԯ�;2xtW�:���lv_��x\�9\�n$t�iox�6�EWJ5z�5���X�w���Y�1���
���L�a������~�K�;":�Q�ն�Ȕrb�=��]R�r��D�M�LcE�g荬��Hd҅�f�h��tqB�u|b�SS���.�n�����HW����o�w�%�Q��.c/��ޏY�+�돼{Q�ߧ�GL�q7T���k@d�EvS�7-��m��0��7�s뭷μ}�9^)�>�yK?^��^�]����K]� �0���\2��-lw���z8����9��\l4�Ř������M�P��(�ҌQ0��>�KQ�!|'Ӯ�YOi�IPֹ��Ნ��6�Ԝ��j���~m��2W�C��!��'�'�9t��/���w�>�y���y�N��Q*t��l:�V�m�_}�$�D�|��=�_"�U���G��i���2�	���4D\��Tv�.����^<��f@�]�8�"1�lض�fnj��S���rz�����L��}�KV��N�;.53
���	���P,	�۞j.�%淛��K//ԬAjw�30���Yu@�����:aU��Y[J=V �R�1l�>����ِJ���v���iW���c�6�>J�g5�8����>�Tj�O���gO<h��y�M��s4����:����ۥ����) �꾿jr��6�x�)`b�h�Ӈ�<�e��B���_�<��~�m�@�u?8zxN!�-Ln�Qf��+޳�뾧e�N�ͱ@Jי1���<#1�����ܴ���r���VE����z�t�1���q�e�S��hyE<�Ĕ&#7��(Ӟ�p��[������m�wuTS��y��g?ŻBU���b��%�I�X���*��&r?ނI[>��c���J@~����i�+P���͗sO�c�eM�����"J��PטۣD�[GY�=Ѽߗm�g��o���]7z<�+�[GM�Y���I���.�m6�}ʥ?̚e�-�q�<�@[���Q�W�]�B���ᢾ�O�}ψmi�
pcE�w�$���)���k�ʛ�-��gĩjC���<W����s��e��gmY�j={h��Z�%M#�k�aAs��ee,�vK���x���������t��ۼ`cf2�h,L/�+H�-�����%ÀKxhhĠ���|_�B��ϣիLt�����J �>���-��o�ℊ5��Z�b"F]�gE��c��S�!�z]4�in���PE}�%emus��zbP���|'HT���2��g:\�����ٚ��¶O���1	:���'�Ƥ���e�,�Q�!��//v�ŕ^�ҋ{��+�1	����R��!^}���گ���O�s�v�OQ�d���߻�������ZUs�=�A̵v�堯��_��);d/���>�yc�aIg�%���8�����S�w;� '�=T���!F����s�z��Ӣ�K�5l��*�cF���o&k�(R`��,�J�#���>�jn�Q0���oQA���Z��Rך�]u�~����e������&�/������l�5}}N�n��-�x�3�_,<�*b�4��|ϣ����F�dD���Zf�^F�)lESŧ���:,��T�Z����J�1
*�ڭ�pB<y���Q�O�&�9��?ܑ�h��&�s,+F�{o��n�d��_��@�����^��)�U���Ѝ��Q��J�����|�8z�AG���ξ�񾏢�J�O��Ũ	b>���/�3�y!\i�<�L��*y�7���a�7��:;����A�<����������{�ek|Ѵ�]t7��^)(����f���T�ݦx�M�г�Lm}0+RLHb�&Z�ȁT�f	�*�TV@]ܳ��ь�SRS߻����Ab�e�u=����襔��$<җ�������R�EL㔰�m���x�>w�W��>�Ӷ�Z^R���L\8ӎ����f
d㜖��a�G7
jBT��`��dw���(��D��F�aD����*|��."�]�Ф��_�kZ]��w=����f9��sfd.�),�F`�^�"-.��I��L�Lq�D�&�ڦ���H]�g�R� }\Oњ��6d��oB?�㪎���[6���b�m/6W�ԅ�_���y
��5�<$�^��z� J��O�w�G\{^Ȑ-���٘��UO>�mRn��bkd|�Z=O���Ƕ��e^�o��G�?A����0ʂ����(TYU	d�w��>]�$��bkL,��ۆ��ll�{=$��lCQ�ʇ.��hσ��fe�"-"Ra�a�V�\�b¸�i��}}�mz��]�'<���?(�WJ3{�ׯ����p<�]��A���ڬ�?y]�z��/�}�O.s�8\�ޥS�&��6�V4�ݷ����V�ѿ�J�M-�\���o��r��k�99n����<qtTc����5�����[�{2���i���K�Li�ͻ��?kж�w�#�=u��ҋ�	I�~�W���=��l�bцld��f|;�F��S`'�Yb<VN�y�5�sM���(&����w�(�*�iI��^�J�̪�^5_Ԑ#Zy~��$��E�l~*��M�ٛ2S;�N�1k[#����[���E��/��.��[��K'�'qE�}.�b��! (RH�$��[�Nh����m�z��zf��Z���M6�-L��mD�Y�~j���rб�R���G�����u�%<UU����� ��W)¯!N��v6��:YS� ��s����x�� �5�e�`��O����'�7��*o��Qe^��.�I��DKO�~�<'$��O����a����X�7��/� -aI��ȋ��4�u;������$�5�Y��B���c̙�^�Ҳ�F��@H�t��T��YUY6E�p�3�|���{�E�������Q�l��bCٓX�9��y�;��r�r�O~s�m>ጢFJ)o��v�;Y���X����ȊH����Ϲ�)�/���8k�21��R�>�y�t^z����4`��e��W� �k�j�;7��l]�����HL͢�R����h�>~�%�4��C!�t���My�6?ܜ�~%���:���9�u�9J1�\�%e��F�{j.n��h3��Hr�T"���xÃ�Q���ɊE������B���!������翚��J���3hP�ӭ���O������Y�$90I�50���Oj�`�wǥ���Q⪈g9��y�34kk�*`�$p�����9�p ���Y��p������\q���\*�I}�j�}/���3΃�E�����Ew��:�������j'�a�E�����
��
�!� T)�❽�m�=Vʷs~n�! ��8�U��<�E���wpp���T���V>bah��*O����y����������?3A���R���G�F���7��U�=�M�I���i��{[^��t����a� �䬣fE��O��Oًǳ�sjdS�p��^�59��_ϔ�j���1S�J��� ۏ������7B��?�J�dl�e�]�`҆l"�s?[��*z-`��V'+S�+3���k��
@dY1���:�<7̭�h��p�UF��-�`^}J�f�&	��
�`m�S�@$ik��� [,�_?��91��<'Z���iBo�a� ��ռ��%�aXz�;���w7�^���~��H���>a6�żi;��d�u^�m~�Gz(+I�6	��y6�WK�S��a��û`�J]�}:��sc�D�'�uIsHҸ�F�,����%��A�D�D��K�!��f��1oM�箫�_��[�*Ο���#Tm�Z���x#�������bC.8�z�H�v�fJL��L��;�iؕ��{9����|�"r^9�n��|�lv٢�<���:˰6��m�w�Bq-V��;E
����ݡ�w߸;���8�	��|�~����'p�̚u�u�Y���[�
�e@W�����;�7q�8�B�C�[9Ch��A2������6��J(��F1D,�Rƙ��D|���w�<�U����&���� ć��E��2��P�dBNK��57[��k(U�6�`K|� X�L��\�i)P�fӄ�VHO�3d)����>�\᭛w��t�
�ţb��H����4�w9���Z�%�p�R���Q�\�'�F腽�A���7���:vTk-��_(ٽ�Z��T�-�;]8�0���î���^�?�<�L50��>��<Pk���i��쉾Dl��GǻԵ�i�|e��!�\ahhPi��Y���a��DD ��bj��\ܳ�%rA�#�z~�; oR{��>k�v��?4T	�|���`��m.�M4|cb��6��$A*�F�g�^ �]f{3a�nov1��F�F��}�	tz�4R~�}[�hQM!�$�<ɵnڿ��z�K�jbhѪ,B�}yѭ�*r7�w���i�8����Mv�_8�\;k��o�^��P�	�N]W5fYw�Hd���8�q�c%??��C�Ojړ0�S	M��-�vނ����5�>/]P]�cu|Y��b��)�_@�3ǡ?����&��l�L	?N���z]U��$}��!�E�3mQMY��W܋YG鞉����85ᇶ7'X^�����ٍ]7��]N{<UͰ�N�3�;�%*ӣ�`��F��3{�9��c�#g���:����10r��\=;G5�؄�B�Kk���}XV�g�nK���9T3q���h-H��9��e�������hh�R��o:�dY�������"G�BkQ��p�',�;8����z-*���BƟ�R�)��I�T��M�'����L�>��"� �z�*P�ʢH�~.��I[.����;D����Y0���Sܦ|��W�(y���H����mN]��խ`ߝ�ƙt���u����Ɩ)%l	�@�Y9�r;��4g�l��)!�I�ӓ��n�E��^�܀/���^���_�E�6����(��u��+�K����R	��na�_���yN�y[�LzػR���z[��m"qQ��7Ũ���8�BM����[]X��YB:��2o���{�+��*�75<<<<�s�����K�k0_�s2(��u=T �7��J���������s��:�b�U%�3τ��i��q�q�O�d+N�x��t�O#�%"�$����jHj$��y]����Y}�~�(��������L���	��\�k�����8԰����
��[%:9�!��$�'���"fg�l����'��U��@@9�����YR�ٷ��=}f�aC�Jj5��|��D�4kn`�����g�����L�%� (�NH�s���<�Z��o�ک�g�h�X�yOX�z����[����;�e=�V���2��~�J�>G7	j'Y�Ε�P��pf�54̮@R���
A. �k�7 m@�h4���OG6����v� y�3!X��G����w|cc���皚�DF�+L�\�Q��|���I�^��nE���쨨i�]�h|G�j�+onU��b���ę5|�&}�yq��,�{5r�ۙ�2��S�>���^z��[����N�P�l�&^{���X]�aSM�m��i^{���iHk��e3t�Ӂ{��}!���̀�-4c,���y��h�yw{�����w~���/��Ч-��òzժ����7	�Ч�	�y|5�?6!��<DF�w���ve�t��dx�J�NƟs�[=k�g�i�J˵~�����+�jkiY�m7�_�ZŽ��������TU��iP
ou�]�/�{�yY�w����1f��l��j�@)�8d�S����ﴩ�8K)6��zϐ��;z5AoZh?V>�@|�!y�����ɭB5h��T���n�������Ã���u��^�r0��~.d�F9EB6-C���o�m���
�v�f�dm�o��ܬW���<��i�?�W�T�r!�B͠{4,ǝ�P짻{���2�)���%�����й�^,/�ڡ��~���z����I���Y��7i����Ŷ�=�.����V�;%OEV�4g�e���A�R���8��K��,��(k����7SH <X`˕�n��t�5;�ʰ������f����hM,�ql���:o��2N��مL����Xihx����V\Cc�ʛ���7�I�ˀL�6~5�S��T^��%���;�8����|t������2̓J�W�w���5ϮOo#��VEm��`��KJл�_)����f�8,��\샯�#��x��Lq�H��ۗ�SW����zz�s�QQ�����s<�g�/ٱ7sBw�U��0�%9�P��1֖KU����������0@��qr�ӊ�/(d��
��$��e�i���0UV� @1bo��?���l��1�$��&R��VZnJ��*����Z�V������%�2���|�b1cf&�����XS�l:_颮��gG6yܨB~�G0@D�I��4W�j��Xp�h��W�o�R��{gT;�r�I�>��x�D��C8?|��{IO�/l�],+�]�I�}K�p�/䝸�LŌ�!55�C�16|��j�+5���!���ϖ�������Y¿��m>��Ω�+�F<��B����SCך�niںڐ�r���u �w侎�X��x�F�X�h����;{{/K�vq>�T�ܲ����t���y�;�"�k_��8#�u �������� A>��N�_�ܴ㜗����;�:P�z��JN>)��m\�щ��6P�tI�����7��q[�l��D�Ե�-d6��'�����$i�~g+$��ӠV�,��\-���Df�WH~}5�1�1vx����\\}׵ӯ�b�.�*Uu�s��s�=���ގ��[#� fzcw/���b�<����!q	�I�w9���{��������sE���QH>I��r��P�o7�ì�I��a�W9.��gϩ�K5�=��Iյ��}x��8�u]Q�<0���w{ƨ�̈́��A�u�	P�>��;8xwz|zq�j��.z�&�̴���t�JɴZZ� /�ûl�?Y�0q��:t��6���e k��^�sب�عc�			V&?�L��雪��hCjkg�5J��P5�j^����)G��`�NI��/���,wI͑;��B�Wם����u�F�	��#��̣
ӡ!6��TS\�DHr�?w�Э2�:!�
F���S��T��u�����E���Ή�?��"1�
\Y�	����Z��?�%�3F}uY����J�h����I��n/���(�5\�X��1$}o�ׂ%�9z�/���<^��}�j�l< %%M����y���"��L9�t��pq*�p�6>E0K`I&�+�A�9��[��r�����}X�u��҇���N��G]?��~IT�	-�I�qXu�y��w��l}D�9���ws��\5��_�^��%�����4�(;���*��x������V���x�vh2<F~����K{�jw�m�yH��=3���9�����TMf���٧���$ne-�U3��/ک�~z6�̨%�e�n�4���F��~7��u��l���>RB�T�9B�7�����d��S֤\R(�1I�I�wli��&�K�!���&J�zy�>*��-4�{�T��]x$������Q�K�47�I5���H����_�4���G���XzZ�M3��_=�?<`���=c�'ѣ(��zD��8�\�7.�W� �������7-�<]��9Z��82�O�R#�}S�S��i���>���;4 ����+Q�m��'�iU�d2�
���,a�b)��y��l��[Z�{�ێ� �{`��(�R�s��Ul���cs��B����&��eB�Hˡ4G	,<��W2�0&��G#c��W�q8{�j*E"Yh�/>���]}�U�* �|�R�����[C�t��j�,8N_�I��G}XTC���M#6��ZX^�&/���Ρ�Zf��=����	^�+��b	Q�9���,x���S�ǎѼ���R���W�%�zcǾ��G�k<%�������_7(uu\�s��忇��x
�'2��1��;{�ꑴ(P���=y<�[�N��4��_O^k���/7^{+�fW9g7ʭDBfW��/�(�1���
mOc6/*/�*� ��TU|������P��˂�9ƇN���B�	�Z�/��諸��ʘLt�-UN��څ���e��e�ݲ`��f`��?���'���rs��V#��%a !��߼�*I�|�$f�Ja^<j����'�T/Rk�ꂵh��xҊ ;�zU�R�@n�J���B���W��Jf�
��v̛����V-j�C������|�V���/W��k�6��A��n�q��}�P�j�*��"���=�lP�`�=�j����p��f0��I�,��3�_>���NZ��_�t_��uv��^ЉҖi]5w���-E"�A�g�}�P��4��)u�Iܩ���ic��~����@ǫCv�S�k���+����~��FS��)��Ňـ�@	ڟ�F�b��g'a�Dz�+�lԂ���=����.;�U��h�������}�����̵�]��nd%F��lױ�.��/�k���Iب��`��e%dvԔ���+�L���≵�fk�4�4��$�K,]5�k�F��3�+��Ku��fUuc?��}a���UC�[�3ðĝ�	NI!H�.��a�$����K1�kT�Z��WcL Cs(�ouz!a�n�;ˈ�p��[A���f5�����xJ1�߯�y��./-Q2;�� ���Q5R��%Ĝ�����d�!��H�lN��E�/i�S}�G�E��݇���+��ט��F�D���������K�Ŵ$�E	[RJ�Q���������k]�+�U#Fi�e�]l����#\��CKϪv��]O�<e�@�{Yz�W���P1�0l�`o�t�uly��koJ�j�8ns�9�WA��9&NNWң��衝�~Ȑ��I��癵��d�3 n$���iECc�_II���2��Cj9f�Z-
�\!`I�ru����)�Kͮ9s�Zp���c��f;W9���ִ6��?v�+��1���v;���mE9�bM}BZ+��D~�����an��A���az{{�N�b��cR�d��)��I�P��c��Q�G2�t��b���BZsҫ��xl�0���r�<��F�x&٫n_h��sf8y�E��݂���1�;?'C�!�1�>O5��L��G��V���m��-�E��>ց�� ��SL.rg�7w����`��Q�2RL\$^���?��D>��A�(��Ӫ/�:dZ=x-�M#��=3٬dFs#78q�C:�x�G%jꊬ ^㻸��XҌe(~���R��x���b+��R9x䝯c���Q�MQ�2�����:F1��΂���
����r}c^��@��Ak�J����ĝ� �ʜ�\�*�ӨW'����N����]u^�Y;�?�����B���O�[�Vf9���W��r���WA�u��|^X(�6xln��шn��b���H~�v�m!��?s�0k>Œ�.im�F2�9s�y8Ȁ��3	!���1�����u�����g�� A@ڰ�@'���t�e����h/��E^Eu1ŷZ���M`aa���Jns.����]�0��g�v��v/8����&�ݯ�t�e#G����96�������W[���ɣM'N��UD��C�R������ᤓi��L�	ӯ
��kt2V�fq���sڜ�����eSN�D�'��r^f�i���>���&}�:0ڽu=�;�t��.���୦����%��eZ=_��N\���u��?� F��$��4)�J>���x�	����1ò���kݓ��2�*L��M�#��.B���ض�UsG7��t�U��\O�¾2�c��'�`��*"K��H�O���Y#Ggg���)g�ټ�rj�<��0�gQ�,�,L��i�ܽ��-S�ܻ�X��=\n�E���>^�[�L���PG���s;p�h+��Ba�I2i����<č'y4�������;)2Q-�'$�����3�(�!#g(`aƵ�K�?꠯e�Ӆ��Ho&-�{��b][�� _����9����Bf�;�1��d�U9�
c�p�E.�˦��!�j-(' ᐫ������O`x�5��)��o�V�꿻�"k�~s=w�WRNiʭ�*��e�ܘe"d#X0R���%�	��ٞAj�E�50�c�Mx~	������{c��˫_��د��p�=H9+Z����zz��J!
e��qM=A��u[�9D2�v~�XJ����st#��ِv�!�̣2�=�\�7�i��P�� m�#o(O$��2��8�:����-�l�u�瘓��r>?)�w���t|���&'�,ˉYX��B6f�S����R+jVQ�I�J��-�i��}� ˗�f����d��.X���3鑋f��_d���_�o;�tf+�Q�\�s����!wu9Ҥo�^��Y��I�o k\�GV��@��\�X�^�����)�ӋPe���=�@�l?SE��v�w�r;|���ۋ����wM��(evcF�h�o��>S'Y��oT渋�lM0�E[B%_���^���o��>���Œ���1񴞂M�Hԕ�U�n�D��A�p��߫������z������^��UVg~�d!�o	���R��3�d���+�WO��%U���1+[:i�~��i��.i��-���͒�Pv��y��T/���F�zS��&X,�9��o<���̝Q�N��o���v3zuU�B��7��	�w��(X�혊4�c�>ONb�m������e@CC��pn|�3��SM�X�%�9c�=��MulS"��K��7�~�zJ�0�n(�i���|�C���Q��R�h� fM�/�1�*3lՁ��o`X/��9[�%��'��нۇ������'�W'�\x/�D98�G�噐�]����t�n@#�iH�.҄6;	�#ل>U���W�B�4unp�S`��V�O7D�,,HKL��T����wଭC�\�k,��a��y�k�+Q��qt6�K�n�C#�]��S\Q�tXqh�e��Oiq��\-[8P��#%6�͛f��Xe�`�b�_���t����&��3,���6C�LM�����e{6vN��&_��d�0:j$���釓�}���~���T�F�|�\�(�g-�z���������#�糑vEt��rc4�z�,�����8�P��G`[I�2�_.�Ry�K�
�#wi٨��Ǵ��������~Z�+��D��a��N,�i�)E�r-5��^�K�ݎ�ݺ#���k	U5;}Č�����@=k؟Xn�3�44�ⴱ���Q�Ll���M�Rl%m����]�Jp����q@����g�z����D�E�>B-�dVDf ��2W��6uTw.i���#Ù���>��U�y+�����L�f�"�rr�`Z]��}A�+�`NB9���-i3���G��D)��s�d*�Ly��ݳ��`�w�m��Ԏ�N}�?Z�'ż�F#��Y��	_[yu�*��� ���qD:!�g�2��f)�O+�f��3^�1�aI�&b�C��Q��1�4Q,Q����vщe."������O�8KhTzXu�\���2p#�p`QN���)����G�1�#��V��*�:��~�n��=��I1rq���!ƌ8>>v�d�	���&+j����ݧ/�E�����,J��P��d>�F�����qfLf�U��LX4R,����b�Z��#���{���Pc�����;�i���{�oY�l3����tFJOn$t󟊨
Js�aze�f�&���?\L=>�'2tP�C�za03��%w�p��^�iA�Ʃ�槧�'a�qtr�1�-S�,G�&���\���^F��a?/ӄ����X� �����G�OV��4�.�D�46�����^�fU춞�͝��O��5M	����ƹ����Rz^��w��Oώ��#�����[3�8Llw3�٘;@��^�ˮⰍ��F�����s����3(��P���z��p��ˍ1�k]^\��y&���^����ㇻ\���4��9�]\_�;��'4n�иMV�7��}X	���w�Ŀ+H�)l�4v�J0�d�єg�V�>���4?ۋ�%�b9���tD[K#s,?��G�T���ْ��������{R"�s��7��5pcu[~3S#�59�����ԏb�`�A5��l���<��o����s>Iт�f������E��Q�e��^�3�,=_d���z||4tC�y:>1b�9��y��@@9��BB]��e�6(���b1�x�+=�48:�Lm��X�m��9�����;Y��������5�B�Ƈ�,��G�-SC��JNZ���Ғ�����bE��-�Uԋ����qؙߙهy�Z,�d����l
�:��?���p �#�gO埐������$Lr$�V�jJ�P"Ұc��9(kP��A�M׽bƊ�{��=���Fi`�Q<|5|��2�bL�t�3��4�b3��2 Y5����m>T1�F�V8I�~c款X�&ƢCP��sJSK��ц6�b!�>�E�z�����_���Ek��l����[�C�E���30�C`�|��RB��;JJ�C�R����D����s/���Y|I4c��.�����,�r0ɞCRa4��B�2�a�+Hk5����b=��lt�2y�5��*0�h��|���S�fM�r<�_��_�����;n|x7��GG��A�xCɦ��uX+RKm
;�<<�T%����L�����Q3�"Q��I����E���9�>EG+r0����ydPWZ`FV�&��n8d�S	*��gV�]\���_���Os!G�.���5(T0�g�����
��lq�[
"�s�,�	�������#��Y������x�L*�:,�Shj���E����$]�G�(v7l�/<L#f㕙<�ɉ��;f�	$ChXy�ö(�(�rE;�A~�����P�nf�	d��,��uUk���D�ַs�<<B��%����`Rw��9�=0�\�M�#�ũc����SL^7xf��E�4�y��@�޾o\F7���y~TT�g��R��1G��k�흑iX�t}�b���rJ쯨��T(�T	����.���L��v� 4�`��7T��ξ>��+
�[�uz�&��S�bz�����U����� ��E5��A��R���R��?[?���"�@�9���\gu��<��G�)��i��sŎ⫑D��Je���H8[�|���Q���k/��۲L�}�vJJ����^<�	��~�㼈\C����ģm]����� �<����O,�$Uv�w�`f>�}���I�,��yy����5�%��z}�a�P�����bu�M2�!B��D�Z��Q��g.W'��,�,�.q*�|���*��P�����W�C�������G��)0u��;�|̎=�@�:��+��фb��F��+*��]��j8;��ϴX����`�"�����}���?(["S��{�S��/��[������8�u�3g��]w�f�3��D�n@>���%Q`l`�a��m�G-2���
W� c��f�~�4ǲ���~�,�V"���gvC��'U�f,�#Q��۝��3�M����+���3��pg%�맸N�4&�8?�g�J�p𖣜��by�8b�ta���0�^�/���W�P#�5��S;��h��?a�ү�������Y���e�	M2���]�����Ǽ��r�;�s*�% t��_��Vo1�/Y�p���2d�~D�K��^�pqIބS�����zH]�x�|�^�����k�)��5�$���<��%��(OT7�i�g~z}��eQ;���Ŵde�e��j��������՚�uTE��m���!d��f06&���Xb���W����w�y�d!2e���9�x�HE��H�w�c���1���৺� 8��1��E>�?"˿��b�-�0���%6%�@+m����ڐ͎Uh�q�!u�wv~Ʌ�Q�[eF��Ϲ_�g�
��?���� d��~�������E�Ģɬ�/�+��+k
��MJ��-�5tw�cl�oU<>�-R��7�{���r�1m+���l�H����}���L�r��Q��2���8�ߤbS[��n�o>��E;X�<�M�?�ɑ�[	�z[�/�)���t}�q��� ���,���M���_԰�ӓobJP3��檯�@*�F\4��_E^v2,ZPihđ��n��9�B����J��>�g+�!����2�_6����mH s�A����9�қ����:$��v2�Sl���v��ڰ4S�cu�J�w��߄��$]�f�0�E�I7�η��կ�n��oG�sҳ�+�轤�Σ338ò�?�P*���(��v#�1c��}{��E)�d�4���16!��|�&�.�Vmp���2rnC��[�hqkA�NWI!��6��Ct����u�w�|�"N^ֆF�g����6�.X��χ>s�cV�BM9�E4�t�+	�9��2�[�[&$g�Sr��:�L�xsd��1���Kd�A�i����. ��T�3<˿_t��U'NNV�\2]|\�X�:D��bS��b���]���X��;���.��h���i�M�ǯ�G��3�����:��S�5��8��=@�y,V�l�.�������es��d~*��"%����+��nV��c���(,��r��GM8a	���mܑ]�WS��߂�������%:�2��gK���=,����0�� |�J��Zo�b'���� ˬ�GQ�1n�z���Y� ����g?�h�51����j�Дia�2��˩�ꧬ�:}$��􉺖�j]�J:	&�h�DȲ�0߮�M��F1YM�aV,��2%т��T?	_�4�4sK(�I��K�lTW���]�&���p��H�����|�Kշ�8mZ{qs����8R�hNNN��'G�	�zP���Xcöq��!d���F��R;��~�/�m�Ɯ�Ղ����{~W^_��Һ����r�nϩyPI�m��}r{pרI��@�'�M��Q���J���{}�АԵ{�U>�82܉���j���B�A%<�WmB���A���Rǜ�>�1t�p O�ix�eS����Hl�i�	)��*`
���0>��s�3 ��ը�8��{���c�G�I�tE�%L�(g���o��,�7��Z[&��Q�>F\^2���ILA>�9X!��J���Ex`���z^�h�{L)�R%~&8;f�lg�
��b��	#���@������O�2��U`��*�$��W>D�.r�x��R����m 5v��tn���،f����$ObK�'���Tٍm
�뵃�ٻG�� V��V#Mv��/�B�E�"x�7��XHHP~����aB4�F���k������m��`c}�sTiW��%1 	��Ε8�
 �Y?�"8_� VCW�Ci��cS�Fl�LUZtT(�4x�������U���8��Q��П���RQQ�q&k8�|�(��1�[ݒDw?��2�bJ#�7�8҉�73G 6�����IѓX��:-$Ydvibh�ߛ:;�pS~б�-��-�0ɀ���0�8��N<m~�d?n��'�m`\|^@z�X<�rP��0���<Z�����\���m�W�CĽ�4g1�A�Gf�;���ʚ&�a�A^��X�����E_2�c�E9Bɥ{��>�3�+�UT�8�P��'� z��>N� 6k�k�c�)F��d�D�'��?���DdV�Hj���bZ���V��5��M9t���3C5�-G:.�� r��	���-��[	�.f�2GAy�� 6%�Ι����_�2<K�K:ӋNݔ�?��%=�6a�(ag��)+�N�.Jyv�Ia�+���|!)�l=��cr�b�!+�������"U����4�v^K����ۧ���8�ne�&��y�� E��hT�y�O���k��%-��*��<0���
F�x���2�C�%��LOt�&�!��A�B��|�]w�{���^�9Ӡv*���~��`LF��^/�c��o�?/W�^�����zP�=}����-�>����r�jTk�����hg�DR�x�Rbcf#ˑ@ۛSC)�E��&�E���D#N��~g�a>�q���PxȌ��\3�ir��' 
������K9�Բ"�y�h#b 6\��6�
ܑ)F& ������XMyG*6\�(�~�~3��E�@����F�
CGoxk6�@�D=W?	�c�������=��=QGvNg��z"����C�}�=�K���R��x�6�]q���f��Y��M{�GKa�+�� g%"/���"����.���	|��D��-�@ P�{AnA'����&�u�+��i���ғ������0���[�[�z���o�w�9�*P���N]h�ۘ�� ���.���(��d�r�����}:%��
��"W��#ƌ���+D��@_ZnP8�O�\
�Y1��#$[Z[�}nm��^��5�B��H����������js�Z�'���:�Y���X��p�6Ch�|���]�=���ɤ]�@-��atDS��j�n�7�z@oU�%�^Yr��y�\B����F����42�m���kͨ׿ǼX��En�Q�������uG��Oj
�*Y#�XDn�&�/L�,_R��`����C\&�B�� ��n��r�=[����$��A�B�i:���םT�1y��ѿ|�z�]�Yaz*�����
�q�5h����O(�����z3�nN8��(^pA��#��IK�|p�׿���q�g�{DVm�Lb��0\g��>�����6�M-,���[��HG��_,L3�W�Ƭ��]�,�e�Đ���1(��d�k�M�X�pr-a[��2q�R|)�H>�Y��lƾ--酉p�eG)b�����y��4��F�=VU�q%U�a>�Y��KJ�0J;n�;*u7��sk�=�̯zO������0E��Z�srb�w��}�/Kڗ$��������*��-����124��x���BY��kn�Y�(0C�������������	�6�	�/C����x��$���5�oT�8V��p֗%�;U@��x���~;x �x�Yb��C܁'l3U�����m�&d&���������y���%��b�TZm)ܣ��*�Ū�q�A
��T<~꨺�r`�0u�Ma泖��uD#��=����q����&��� �Y�ȅ������L�=��
���v���wƹ�������Ui�4#�� (�<��	��_T�@�:�ܬ��Ǡ 7��{�N�=׹Hfx6���A$o<�������y�n7t�D|�;f��iko?4�B�?7(eG�� �Q[��If{��Ő�9ً�K�C�<
��x��-���������v������h���Ex��L㿣M��X5ԍ��6���ۆ�Jh#��+�Y҉1b:���U�2wK>߲;��-Π3+u:�#Zv�X�z�����>�ڸ�C������²��(�e�	��+W�N��{k���ս̵�EL8��j?�o��Y[��K/�M��9���qX��pFY��%ˇp�{�4#�d,���ixI�����h���f翰eo� N9�]�=�`��z�0���l��[��A�����E7I�.���P�Ó��Is�T�A�.��~c�z���o��d�s>0��]c���E��|y�?�"��͐Y��$����	�b/9ϗj]3�z����z�#++�h��$**Z��qʥe�4�M��mt�<��c�=�͛"�R��!
�9�fCfZ�8�kτ	G�c��I��N�k ���j2��i�zV��n.�H�-'V�=.�.P��j,ǮW���*d��k�\"ߞu������[���bq�1��D��;�Z$��ade��0�ESN����Pj���@����"�x�.��I�?c�f����vݸz7�b	��9�xi�L��[�Pl��#\il��:���'���UmD+؋�	'aln>�(�g���OC��n�L��vN��ƷʤQ[�E�M�����5@DJ2��RM%�b&�\N�h���s����By70�w���w�I`!�(�R�f)�+-�յm��2Gt��Z�\{��N=�wL IMs�7��J���-]�g�I����+ޗ�<��cZ��LS`��c������TB$���M�n�������I�#-��ح���3d!��d�'
����M�``%>5���Z���Ѐ�w� �s.cѨb�lP`�eg�r��,{��~�/d�5t�K�v`�i���*�鍼��y鍻����_��{��G�~�ϒ�%͖XlZqq��y�(G׶��^�E��|"B�U_R+����FY����^��^K���T�?b���E�C�؟/���7�U��ݻН"������>�e.C;t�{�e[	}��v�ÏA��D��̭�Q��9ʃa�|�	Q꺼bb�,�U�\�/��t	�J��Z6�K�f|d�t�[ت��X����*'$�C9��S�9V�:�<� Z�o�;�����.6'V\�|Eʪvz�l9W��B��
-AE��K�B@_::��aك���ba��h����:��~����pj�+H5)^蹭��<~L낲�39aoQ�R���/.��#4�����׋W�+i��_���������Z�
��H����-铣1!>啩5�j&M�y~[i�[�Vt��E0Z{�(�|��?��8]#���pP�p�8��0�h����!FE}���5��R��I7C�����PU��j"���h�� ��_?��, 4�@&2�&~puy��+Zu������n�� ����������<
�,�L�l�lwꤝ���G?/��G�+�^2K����R�̵sQmL�tR�8�'���Ҝ�+#t~�Hw3ϦU'#dk]��T
��r�J8C��^�0���?7����)ha�������%���W]_�N�������_y/�8,���Uf-%��}�@� �*S(��"C�.��,�)j��V��$r�s�pUK�v��(����sg2K�h�% �2yt��s&��?�1xq��s��33(Wˡ5V��h��B��٥u��	pb��HrzzqX�T�ڄa��nf���l=�;N^���y�dU�����.td���}hv^l�v��z�Յ癪�V����c�����(�Yv�ن��נ��_ƣ�����S��*gb���P �u52��ʝ�2k~,�]�@z~53�|"��T�L�NK��_:�_��q�hd(�h{�f0��������q́��ԍ�hjs1��aU|��V}d���X��������/�O������A;;��W��D"�e:5#����cY�B7�y���պ��:���9��B^�\�c��OVDW^@9�;�f�V���6̚e(��RPyh��A$O=#zׂ��J�<�w�)��6��K��p$�ܮW�|r���+pB�7�����LQه����<��4|�a��|�{�,�(Tu����`dJ�*ի��;B蜼�ƒ֍��HCc�*��cU��7kos�6��%G�03�bi�B�PGL�{�HC6cɴeʛ�ķ5"W�SBP��l��t�?����]�i�B��`��V���#�)�3A���oRk��k�\[_����b[Gdu=��|ם��qON5H�RGUXO2����:�y�
����m���f�ſ�%Y��qK���Ş�� j�<����>�9\@]\hh���(�K��z8;���֯��S�ŢU�`>i�^��N2U��8�H����x������|�(N����NLz2�%ȟ}؝��EWWwW;ϼ��B&Dv�C�Wn�uf��e��k��^�}8����ce�K�za��*[���-�e��zC���Ƹ-$]�=�MI%���0���k��.44�5�49k��2f=�.���m_�&2��_3��{����"A��B�S���Uz.�����n�����ϐ){��>iΜW$v�ދ�_C���Tu��o��b�Po��n� Sr���4޿�S�yp��\m�Ц-��蘛<�~�c�F�%T=�݃4֑L1�� [ww�-'m��y/�e��drZ ��2��m���aч�<��E�P�bQ4�ҜT�AjY��o�Q��� ������S"��G�a'�5��9��3åP��Z;W������&dm�ngsr��6�]O^eǨɣ�͙��4���zp&^0��C�mD��s�F�1O���i���C��u�|���6hNEt�%���7�`�a)�ƌ�9ͦZUb�7ƪE��D�?��:*�{$��F���N	iP:)�n�J��A���!��s�z�ᾟ��>��X��g�����׵��KE�����/��r�ⴴ�26���=��7m�u��6�uE"����R�7b:��a����O�
"(g�V�V����u��,��b�5r-����m;�}�]&Y&���Ug�&;�	��o)G5�i�J�� �7��w�0c�.(9�W �쒳�8����[�@�f��l���
NrD	$��/���%�j�-���SǓ~��V��HKH  �-T���}��Gu�t�L&�ز��O�@~9��E?�6��}~N��t��I)����uYi3D��/��U�汽Z�6iD�j�~@�q�G�Xh�Y0m�� [��$�7���<e|gt�)#Rʎ������yD��?S��$�ގT�itۉ�\H��Q�?�ʎ�=�����r'$�^;�g,y�����öGf�6����G��l�ҹ�M|6"}�`�Rm"��ʸ8��8�X�������K��J��M�M���.�*E�5�Rd�ӅU�YW�Y3�2�]�o����"�2h��fa~��=
�F5�qa�.�P�8L۵l�?{���=�S�֐�D�Oy*3a���e��y�;-�P2�Z�-�T	9Jx�q2�]���B�B���.nE����R{�By����|�!�'�B���;���U�-c���Ϥ�dZ���Zlz�;���u�#�5-��S�F�-n}��s���(�߅����<�n��q]{�n�1겲y�X�@��B��B��J�ͽ�rK߶6���(�� 4k��͸_��]���B�͌��՗$�;`��HW'�He��Q�������^/j\4m����|&���,:l煅 60��H����a�9�E96���I�ȟ�kx3,�xa@��v�-�b�~r(�AU������A]3���L\e�y�����_jO�L�����&�f�ݝ�`#C$$���)��͠;Pb��=�0�����:���]y3��1+��
`WmGm�Dь;qgV܍�%8���)ۍsGǡ*Zs���H9ʙ}W���fk{z�a��m�o^9�t��>��J]=\��_� 0��$NXD��q���yzm��A����h��xg�R>��|�Z�HAt4�����D�����In?'�F�q�Z�2y*��?_�x�j蠄��} �l�W�a@V�Oɫ�{��~>#�]��f�6'\b�E~���@7Ѝ7&�x,�8��F:6��j�T�zn���L���" XO;�!!���ɍ�B����M�ZI�_��@�-���l_�o겴�*�����lv�;�*�T�o��IV�Y\y�O��,�a���S�7_E�?����&�~grЮ��=�'F�w��{%ty@ҡj5�|���Y�2�R�SU?*��S�u�+��E��Of�Y��dt�u1ͳ)��UƳ�\�"J�W�X<Ay��N��P��!�O���:��.�>�͞��\�K�F��?���L��~k���ˮ�]������b����2����Nl*&�S��Z{�~3<�WsT~�n��b��]�ΐ�H�����7pӌ��t\.j@n0:B;Z�i��ç8��`�w5X^^^��`ߓ�EeF��Aݲ7�~M����dԸ��9w\:�˰D_^}d^�ѧ��o�Z�1�����Jn���G���$Z�V�K�Z�6�2�LH����S�(	m����S3��#���yɇ��ZslY86kyU��=w��8]��.�����۝��y�_,cҿT�V?�J����T��oA?����P.��Z��gڮ�泺g	��+݅ݡ���{\�s�J"��lm�gj]�J�]=ɞo&5���5��;�D���Y��Z��s�������
yS�;������YN_l��٫��qŜe)((Z����+z<�6Ɨ>��w	�b��S��ѩ�5��ɕ��{��S�<�g���G~@�z���͉G�ߨ���6�����ŀ�D1=�6i��h�ݥ�]{��r�.4T��ˡa{{,�`E���sw��Q?��a"�d.T����{��Vy�$��_п}m`�ۧY���a�^�s�������'����T{��<������aaaާ+���Fڼ*A3_m��0��X���"�0L���f$��W�ao� -
��.�g�A�<Z ���|��>$t�3m��9��*�9�H����� L-R�l9� Z@�=��������#x�>3��xy/��AG	�msMg�y
d�ih�f�)O�>ʸB~��O�����b����&�����)�{|�ҙh�|��.��E��A���dV/n�%YBf1x���GIC^xb�Yr��m�|��Mt�[y1�S�+������\1NNr��������}&x~W�$���Ŵ]�9���>�~I��cmO��u)�������|ա[�g�5��A_��{YL��x��~7�u�G��E��J��C����֞K���(��"gG�
��1�j��z_d��[�����ʖ�l3�fB/�,�U�m`Ժ����<������㴏�7�D��񛋾Ь%]�i�q���Il����L�§�f��Y�5�XvS#�W!���s ��+W��}��Dq��.���26��d?�:�u?�(,��,D�$��Ehhշ1�l5{�.$��g�$�%��b_x��'��D//�vG��� [��j���������ȳ]��nm.��
������J���'��\� �����Y
+�;K^��M�$��l�;��72�R�̷z]���l���!�<�����e>�F����pd<�w?*a�b�gO���~��	$�!��BL�H\�w�k�?�^9�{Y�� �ǰD��͔�:Vz��_�}��
���o@ڼH��
,�"$���\��+_��gRPP�p2��v�:Y�/,�ꗥ(3"����{q�ri�Z���=glƕ~��D���w�3���f_�	<�M +�Wd�T�`�E{������8��/
3޻��d��	R��d�D�(d�׊�+zgDD�q2kX��I=��ȁ�8BTE�g����pv������F|�ł��~D�۱��$+�L����5�oj�䝉��*�i4������+\uDЂ��D��/t$��}��(��ES)u�u��"�esP�D��Ri�>A�DK*��%Ѡv��k��y�J҄�0+��Ҍ`[�eG��X����{k
�uW6�7�-�����EC��sn�m햚�8-9w��U�dnm0��(��B���|��o�B�N1��䦟R�����)�����+y���޻8�7�n����
ˏ�Ŕ�Dq}���B(�c�t�o!��������Vw_�����}5�ا��^�C�E^I����^�����4$�O�3X$�w�����'�T[�3�=��$�n��˜��9fy���=�miV�l����3���!i6��:#�`|F�qj0`�99N�B�Z2z���)4�W�{���qR��dR�&5�A)[/Δ�Z](Yx�N!�{���q�^��e&����q:��	��"�-��c�m��H���WU@�T��X+ӕϜ�sd���O���U��1U���"wAq	z�LԤ�ڶ��I��c�+K��2�"r�`1�h�A]�l�'��5!����0�Q��`�_5��t������TA!F������ J��yS�d`ɥ�@���VsWA�O3W������+��x��6ئt܎ДB��)��X�*�#�����>Fp��ϜZ�<ΐ�7�C-��1�U3������<���qR$v�NB���d�ˇ�+5��7k�6�<��%K��8'�]�P.�R'o��:~"ֵ��l�YY_�n�1u�;4ϯJ[�O&�����+B��;��9!e�1�h[��1�A�8A�NÄ��EəR](���Z���D�������ĳn/�w��q���6��#zwPCjV	�ʋ��}�]��%ߊ�AL�rh|���nY-(�9���%[D�n��)l$���<�yVy�ʝĈT���*�D�vp$C�B�C"���H,�܂���ڍ���ax=�E�,�;Rrx�]���Bm��R�_'�S��"�(@s0�L!OùE��j���vqJ��m�u���EX��_�ܣ�ϳ����Nl_A��ur���
�����J��\��}>�^��(߸�j�͋����,
������y�"��?̓X@�F�q�T&Y��K`�mf�A$�߯�I@)�`t*3B&��*?���L�Ħª9Z�tE�J�#��1������o���#�>]�1����u$��&<䒈P�=��-=��v�z�k,�`$�������yj��4� ���Pĭ^ʪ�R$]����Gmfk��M��g��b��"hͮy�o�i�:��}t#ы:�A��E1��X�HG��ћ0�_%�Pd�#8�.�e[s���4���ҵ�R=:q�ة��]��s|����\Wc�٤3	��Pb���hE�D}���L��TE��^i�4!��>`�|KM4z�9zG�`ݹ���{�@���rMp�J�iu�h;���UQ��Է��k��ϊ��J�U��v���2y0��� ��V��}t4��Ӧe���-n�>�uG�2'+��+X/�%W�p����)j���Ӧqq���}�BA�"Z�� ��1�@���Y
�*Ԅ��CN���n�:�|���������G*�+N���#&��������\��P�%�ˁ@±��ul�Τj��}�a�hC�����_�Ý��_ ��8T���v�"�Y%�����*Nxl������V5{z1�FO�Ū
��2_P�㣓���k����yi5C��4�0;7�gd�G�GtM3������#�ޗ]a����u� ��ǰ����9����g�&��e��q�/�t9�rG��cL�cr�~���Z;le�� :��8�#�}DyY+�4�"���Hl ���	���h��)I�����z�R/� �9����^������U���{Ӗ����q��.P�|i��|�}��`�"Ю������ފ�<�gݑ��
���'���g��=f=t�x���������:Tv�M+��U��,�l#��lwww�8���T��mfܩ�!��EO��s&����T>� a�D]L��C����	d--�Te�Z�(O���$A�#���&���n��~{	=8D5Z1Q?i 	3[x�UFAJ�
���(�"�o��<�M�>��%#��Fa5H������f�	�%���kݨ���9�47ec�x�|��o�չ�{ʁ�JY�L�("-}_���17y@�ki��FbRIN-� �s\yfŃzz��ݸ�DeXT:t���-*�`��m֯���m������)�9����ۗ�-��23��o������Ќ'"�|_��X(i��X�<*��R���E�k���,B�nUk��$*�ݦg��UI���W��I)�x��4�OK�_|пy�U�[�����J?��0����zƆ��7�W6g'��
Z�!!�[��Ck����rs}e-�kA]=�~��[�H%,C�ݗ��	B{hE�E)����F4�3U�Ї��v���lm��'���*�~�\�v\}�_�x����;�?N�����	�����v;}�����7S$��	Lj9�쐊Y��J>$�3üKdi�ʨ�昭���I�d8��Q�������鲨A��<�`YI�	��؟A�	]���n��a�Ę=Ctc�ww3/ ���
2f��#��ك�Ѱ�ܩSxk�� ��0*��@S�W�n��;���^/5�$Gej�$�`�]圏�ӊ4u�����bj?��DQ|̷㳓m8�_�44�O,��� �ף�N7�c�~�j=�u�J%��S�ҷR���ߪ/ƽ���;Fk�N���B(:�m�����\q;�|ʍ�g��w/7� �^S�S�U��#�%8����51��P��������"w��	�.xuu��Yј�P�|��v����ql��n3�G�75��c}4��>:�!]��w�+����^�Z
��a�(�7���=LD�H��7(������Dp�b\1+�4�Z�(qe��b8׾nu�O��I[�9�J"�*����Lj�g��z�S�eߋ�*k$�65L6X�Y9��{��ed8�T�#�I˵��ɦ߇��#N8�S�%�>ݼnPq�l*���ƒ`x�,�
�W�!��V:Ɩ�լy4�|���#��z�[K���J����#��Օ���h�����e4�U�W���_||�AO��^���ft�6�е��<���P�q��h��4�ǫfY7��Uf��B5�[n�3����o�[�X|����s*)����Ak��[��(���%�@0�\/��3}L]1~��(�$�����qM�Z�:������Z��+޷#¹�a�NO�|�Cv�_���J��࠲�Uz��8�UQ�����6Jc�%L�Ma�FqIĚ��=)3��^+l��j���%&1�6,,,�	���R-S��?��/us�#X�+ﺾ��V�Ө�����#�?��V6;F���6��o������(��q7C�ڨ�:ѹ��eFvo���(���M�A}]��p�*m������z�����<�^��l����AZo�����>�n�{�gP��] �����Z�D���~3�v��GE»@ZxIJ�R4+@�E�q��(�-d��h�!���&�mɞU��1<��A����1/�4�~{uD���gD�G;�.%�D�V_����a�Eer�%x#_ު/���A��C��^�I?�.z���{&y�[wssmӯ?K��^v���������c��l��(�����=_�a�]=�P �G���K(�!�M�_�Y,�o2ʐ�h\���-5��3����4F>����F5��`��ı#�sY���wcaƻ�). O?��B[�°Ն4��iQ���s����	>K�ɚt3�JF J�:ɧ�_�'1l�����IRZ���xA�- �^���`���W�=N#�Rn�r%����fJ&���1�,~w���lR�3T�C�v�P��@������"����=�B�0������i	+�[IB�~�*[��T	�*զy�ڼH�=&>��a�\5�f����^DD�䗼�G7"M�m�&����_g�I~��!���5K����Lp�E���푑��7�	 Zp|:�N�Y��uX&�"C�%�F���r�!���?|;����ܔm�l�Y�~�}��x'U��g\- ���GQa�!WIYD�h�=X�,>����M��Ǟz���@�g��|Trs�B�3��yh@�W�%�!��Ɗ��kjT=̂)�]�'�Q8T�}�߻�1J��'M3��fؚҋ�ܶq"n�V��vUը����/ �t��22:����H�O�X�-��Oװ����t�Fg<���Y���h���5�Mg*_6�T3���Jt������In6���!�]�h�X�.��2Y(vٺ���2�~�g�	K������Zq�/�ւ������h�\n�9%o�H	�η&6nU�g�O$.�~&߄��$V��/��b�=�䣬oAVo��jd�_��!���#DA��%UcR.�I+����� h]��/vC��;��gf�%�h|dQ��I�KZ���*2�M��b��6�%���ݏ��D�R�qR�8)1��Hg}��`4Gqp8���XCVo�!�'��mЉ�zw`ͥ	�q���E}��Mkh��`�)$�L6n�s,{����{�fGOO��W�����UM
zGH��Ȧ�Vb�P�ؿY����Xp;�c�.�-~�q�6F��Y�~�u ���}o�^׆��j�y��|�K��l��
�R{�{��M�i�������\�=�hҦ���.K}��������`0jG�7�)qu�����{�&��� ]1�O��b {};��r&,i�D�$��������+!؉� M>"�$;X�ӄ�I�7X�6X�R�xs�_�Ki6��N�p3�c]x����
#eDn��Y�T�H��W��ZT�UtH�Yg�I�m���a>��h�~^�:�!�õN��x)7��`�B����K"�H<��0!���5� WOBU�����<8[�khغKi`4����@�S3�y��\����p/�d�(���&��-}7��=��/�x��y,-��Ab��5�-"�V�������`��O(3:[���y�+:%L
E�@t��;bd�)1�\Zr<哩����y�X�ǨR���?e��ڄ�'{��܋�f]em2=�G����p!��ii�ja7��J^���]�pG�_v!+$i'ad�b��z�N�|�����S#5�)�������Y"�0M���c�j�9��Pf�3�,�	�,�!��#{�_��r��q��}z6a�P%��E��m�V@"~��R��+3eљ	*6�N4di��XV�9C��8�;C�/�����E��o�K����N	�Ōr$�F��1�h�&O��	t��;�C���:_(f:nw3�[
�� �)Z�B+�s��Dobܾ�]�����H.О'j
��I�~:۪��Z2��~���p��<��ѐ�E��%j:S��^|5�,��L:*O�R�4��N��S�q��7X��F���4!}F�μVUߓU��tr6�Q���$���鈨����f�Qz�X����&g�)��W;2F�P_��r�}T=�S�b)pb	�z�q���=��	��2+}b�eIP�ɢ�[��0��b.�W�I�/#���i���@B;��5p"����{��#����P�.�ν�"�eQ.aǳ��27q���0�}2�n����)p��?�w>�&�ZSg�#���1�e�p����'D��Fgn��O�h�
���h���b���o\]]w6��q�w>9J�����x*,��Gy��͹0��f��F��V���̽0O�p�����q�ܕ�B� �� [f���n�ot7���hH�ʧ����
Ps�5�7�w��BJv��?^��"N�R%��3lq��)��Z���S@��p��@�ؗO�����ׁt#,���t�2"׬�=0�yR��vNNb�`nU�9�(]��IBb	��h$�Z�Es,�3JY���_��F��^1D�&Bu���wT�Sٟ]�R��g�[LB����ţ�K��f0+%���t���[�yP~~�����S5�O�l�(�oc�7а�W��4�d�l���\Ϝ���菻���Zd���Wr��[S���b�6��v,�i�YT��WqN2 ��RVc&�������[���
�78��@$d����8�,���=�v�>�rg�{���?�/��E�C�#1�P>���|��֎�D��F/���I7�������.2 

��[h���(�g[��m��_D���EH�ரH��)�44%��0�P�v�_mk�����P�͹�p�)l(�7��]�ӧS�3����+�<�J�s�"e�w{�a����t-��o�Pl�?TAb���xT�|6��[��=��#�"�R�(�I���CVoooy���ɱ����n8*��>���q���s����N��x![���X��(���g�1�$���n���"K��9�Iq<h4��(�4��a��ײ˔�NR��oN;����h��e��;q�@^��P�Ne����������{� \u7�DQgJ�*{��4y��b�]tx���GC�?��(� c`I	3	"<��w=�e��a�P>��M�o�zU~N��}Z�cG.L�{,Q���6�7|7V��Ł��c�Ԩ8��B4��TkK���n��-fe��E�'����.N?�'�6��O��23Wg���b{�VT 1����tr&Od���[��x�k��ص����e �'���і�ss@ʋM�?�e"q�	J�7Cj�>������Ӽ<n�	2��a���/̿e�ڷ�?ٚeR?:o7�������"o?W��%Y�I)�׻����B�Iع�V4���x� ^+����,�NP��M�	���W׍�e���e�}���<���q��^ɰ�R��|9��c�Ͳ����x�in
kF��<1W77=}�/>N��i.���7�-���(h�L}<��'y������1)`Vg�uw#K)�N�U=��).I��*�W;=f�� ƥu�m�������!�%=7��W�L͝��X��,@��*�St�����o/ R
+�87w���K�L�����0��.�mϨX�5GE!���tFF]-�t�t���!M+��l����4&&&���Fšx�3Xjv�қ 8������Ƴ*r����4'��SH�\�2xQR΁�����$T��Lv�}��������%�Y&���-���뒤�5Z�(�`��h�`d�N�	�i/�?ڄ}�� �/���V*NV\�G�,K�TXǱ�ͥ�%�cfF���ƾ����L[�;� F���FtttR��E�b�g!��7�O(�a�i��N�Vo�/`���>���p����F?2O�����M��t��.�5,�^'G�r�u��q���\�ƀﶒh%�L����ټ���X��%�ʹ�-ZKp�N�6�2�(C>����tZX) T?��mޢ�;�}ؖ�>��na�n��!����nV�����E�� ����L��tӿ�*�r���~��4$9�Q͚7�H��*�r�����j��
%�{a�Gl�)�;�b��T0���e���ľ�-��K�7�C�<���)��8+.j��aTz�t��}�0fśkG>;;K:G������=����I��+�qb�@e 0y#�&O��[9��oSq���(s�ƤEV�{F�Y2�ԿGdWx��4�S؂�w׀Ͻ�����pu��]�,и��w"7�^x|�abs��+��!�n����9+f�U�7�;M�7�[�ag����]����:8܅��QK�/��K�{a���R�ت7|q��>�4`�9XK�����*�"�A�{G ��,�'T;��2��Z dk�fN��|�p����+ #�4��d02~�<�.�������F��N�h`�?��%�uՅ�j�Ҍ`O��"�z� (����Jn�8��u_��^�^�FܱrT�&�~Q��wZ��?!���XA����!��+0Ny
.9��ji���JH6T���B�S�?򏙇6'X��Ɂv�1K|�$b'H3��߄"'�(l�m��Ԑ��U�(��&5��Ҳgt\�W��g��63�"
� �(�b������_���}�t?r{�	�D����i.�'u��4�L
�n���
��}d�I����S�g����)u��IJ�T[S�1�J�icd�T�_�֥vPQ)����::ڟ�>j�2��~�4�"� XYp�ů9 Y,X� 
�Sƾ^}!�~� ?�A���[k��Tnp
,=��
�M���isSY�#�����;�����鴴�w)��j�R��h!�����N��fփ<1���Z�n���r���q�vt��r���C�����9o�\��Ġ�1�H&��\8�ۍEԳb^�M��� g]]�]�AQ<�nTa=+�\�*9�\1�R�s��yH�¹�梁�8>R�����D��cA.O��~�?�ז��cϊ�Õ��5Q�
ŏ� �����dj���S�o�}��/�yv�K뜍�@kg��&�G�^QLfΌ�e�C�̱�%!�P�+6�.]�V���)�hH�]SX�r`�DQ�=K���UZZ�#T3���XyQ8&��/��3�c��k����7s��������# ��	�����z����&x�*Z�\5-�5#�,'�11�\�M�{����5�'���j�f��n�G+�y�J3�֝7�y�f��xv^���T����������JR�W&a�0����u}�u�q��]�!��S�>Ǉ�+�;�mGX�6��^gn�qy<bkOǉ��_�5:;�NՆ���� �,����/�8
�s%Xf8U��4'M�3�f��%��4�G@>�sMz����YS�c5	����EiF<��Y>��b��K�S�=�_��t.�����W��x�@��.���G$��5*��%�Q��&��z6��7��R�D�o|*�dy�TJJJ\� ��h� ��3 �.2��d80�[\��]��03���@=��E�#�i�^O�[�����i�OŜ��=��4!a������B�9v���"Rb/T��� �]�c���Eч�z�����6�����VU,�bЖz0/��o��M20ּ�$R@��Xi���uE��<|v|����N��O,-����8%���F�T����<[�`��Ne�٧��o�[�Y�IsƖ��X�st�tX%��>�EN
�.�Һ���Z��?�@��("�"����θ7����YH0�%ԓ��%͙H]��{|P��7l�b���`���\=���w鉍�<�@��:������
��A���(_)vRB�[,,�+Cl/hs����gr\�5�ɷR"5QPzƳ�z�*����ן�7�c��Ф�"r�I�?f����}`e��W�U	:ï���E���[���ϔa���[�^O� ����K���5�pd#3�a��n��ID���`�߉�=b~���dymw��^��̑���^(s�go�ׄ�l�4Ң�7��(ķ2��]�8���.�����Zڊ���Bυ��n�X���5z-�7�8��Σp`/���(���yZ�N�θP����7W׷��~(đ��Ӎ#��S�k4�,�S�V0��붔�������jء��t�i�0�I��'!U���r9SL�[c!gb�s��DՎ���~L��=���/cmC�E>�,����?��ႈe�G^����&���'}�X�������Q�C4�O�ө(��N���(�#V�Ö��J �#@���d	=\��9Qh+t�2D%<��bh����"���9wK�I���Y�u.�n�,�-g,q�Wj<Z�*PRj���.nC���he���]�����/ӡ��Ҁ�=�~�Uo��)'il*~������B*C���J=[YoW��	�!W΃U���
@/�ϲ����b�:&�^�����W�J�Z�Dmܖ>����L+]��5��T�{Eo) �
�>�R�ܽC𕛄�䍝����r�~�@�Qƍ뢏h������hȎL��x!^���Kl	H,|FX.F<��z����N�qza�"�������(�J;I{��?�M|S���!Jգ�B_٧�ͅ�:���xȚ��2��D	�(����5�"}u6s�#�(}�W��>ϊ������i*"Q
w^����k}L�i{�y����S'�mL����v�k9+V�ZJ�U|�Zw9����)B-�O���5���5��ã#s�������";~���"B;+C�j������e� ��*Pf��J�s�F��xW��Gg�g�d'ͩ�$��5--#�L�����˻���s��Ju"�
����}�g�bi�f^wǱ4�=�U�9w����Rybn�;<��qS#s_�Ã��_�M����Pki�������f� N*�_��O�(]D|�B�L���+ׯ�~���R��8<
~odWW����Л��,e�~0��n�A����)
�'k�H�h�I�1m��b7�
ICV�J�Z8W ����],��H�Bb?kt�}�N}.寞]@7�����^��
袥���4�YsW��]H��mX���q��=+}=��:�ecbi�C�f%�2x��;���$�F$�w�����񯒯GV"�I�C���f9T�ٗĶ�r�c�t�=\���OM�2������֟�Ay��W�����[|f5��G-�_@������ͺ�rλ��s��M�ډ�1�蔃Q�o�J�L~>Y�H2���L���4��q�fL~b^�5e�1}��v�Nz�u��G)$x6��?�X���b��IG?��P�rrK�_�*<�ՙ���`�Ye73��I)���Զ��X�eg�9��G�o#���w�11�u"��q-0�uw���:Ȣǒd�͗:���Y3}�qu�B(lif�{���*�G�!���?�Blٺ�!�&ҭ6��$�9t8;�3�\���[ɜ�z/qڼrŕ+-/�x��}k�5��CZtT^��d,��Z
���E�P�>~u���6����Qs��Eѱ��A<�碚_�R�C��ԭ$�ǒ��)+���i�-�#8��z��.�j��|���B{۲�@���lr�>�}�O:���]ED̜;u�C��dy�lȓJ�}c���?;䓣c�miI� �/D4Y���G)�P�<%�v�x|e�"��#��]\�?���`Z��|�	��r���^Z�\l���:��sN�i��?��g�l-I�"W�:�"�����Jf�LTb���B����ge��^>Zn-='��%6���mZk���d@����+4Pk7��D�66���z�0+ќ��w������8d_9�{*�eTm����ޕj �L����ϧ��?	�r�Ҍ(��j�{�;��64ʵD�p'����v@�z�ne^�?PA���M(�j$�\���#�i�)j{{Ld�����,��QD���}2�Rͯ�G%��^���U3Ύ�7��/K6���+e�y�&���(g]�$)�pg��E�iԩ{  ��I����xִ*�.5�<OC���f���h��8L��|>H�VU�L�a�,��
RJ��n���������O��"ѣ�Sv��O��������qq5�C�r�X������,?�o��)^�"�̧�Ҋ2N*�U��ï��d�e�cJoޚl��ܟ��9�憫�e�d��K�Y/Bw�Ғ�L;�����B�{2Eܘ#"��"��F�i3�La��\�^���RId���^&l���*�Q�N�z�O�T."����:�A�)YU�o�Zo[<�Qh��Zj�pk1-P��\͛�2%D�b0�V�Tv���Z�+��aR��&G�-^d�F ���~�`i�P+�.�|��И�'�L������'�������&�������~[�:��a���< q���-����b����L���[��Ǉ�"""K-nY%%����;�!uI�9{�0�U?Ak)�#xRՆ�qB��8}S�v�*=�i�ی{�^jUOϨ��q��ŭ��V�Յ��L��������8���"o�$<�
�vR��kF�>˕�6)U��7g.��K�j3�s4��ͦ�`��d����#q�œ(�v�<�m��m0}�k�g��DA�.�Fp��_�o�0�Ϭx5����2D�M�QY>�n�����ݽ3�*������`�Q���k�2�.���I�b�=Os�@�68Sh,k�����gE�`��A���� (>�l���=wus�_��ZX�l�
�K�g�� s�����
T�"�x�Qd�$Ǹm�:&h�{�$(/�9��K�RӼ�����]\�X���H^Kn���Gm;tww#��ڝ5��͸S9��t�LQ�)*TKӿ;p��	c.�U��'�]Z�6���<hlL��-g)Zi�x�ơcGSb|��R�������ˀ��{I�g��<��x5�K��B��αQ�V��aDit]eI�o���R�k%�>�E
z4�k����6'[�gLT���<T\�-<�є��lJeI�F��#X�Y�F�۷���E�n&Yxć3�Idw���'S�_������urZ�h�9��c�]���	�����t�Ĭgax_v���ac�n�0b�I3�]���)/p	{~yYNq�`�	q�1JjF��!5��~W�&�~�E&���~�AG���RI�pML��a�66��Cd�,1�/�o���{[�<~����&Ny�}�AH�Æ�۠��p����[=_�[�7�Ot���>�5�1�����}9�#Eͭi��Ƅ/^S��nUK�.4����&Bs]P�^#<��2N3JM_�e���)A���"�`U[�����Mun����}/o&�T�z���wy�&��Ca���Ü��?������L��_�(�m0���
n���G�Gԯ;�&�ב8O;���wg~
�p;��1������h��C�s郙b>8P�g��l\������6R����Ҝ��a�ǔ�*Q��2���-{BB��x�2Gȴ� �ʇm�q�E�]�At�sS�3�Ԟ��*��� L�TP���Sd1��CL�N7阇�t[hV����O���'�i2��&%'sZ]_�m��n���WDr�n���Џ�g�&	��o��e� ���yA�Z��ؗ��1�/�����01⏙T3VG�?�
�q������A�p�	��|�fҨؘ%�QSdy*�%� �0��w,��}�����{�\�F�}�������h��a~_�c�b�#~�'�뿫!�ine��{%�s� ���z�A0���&��n�Kz��{���5=�����sR�nT4�Ǎ=���3�����+���gb�q#�޾z����,�S0���nD�����yŨy��
ܬ���H��2��L��3,K%�y�v��D"=��*�R�ofe��y�JJV>*�a��q��g ��segxJr*�#����tp� ����}�Vtn�x:9�U�~���=s�kAuM�� �VN�$�� ��ޚ����NҠDdZ\B����n�V��_R�����fV`�LV#�*���$�Y%�e5�v<������4��Υ��a�e��GZ�)hU�x�k��N��p�t$��Q�UqQw���)� )���!9ҝ�J	!-9� JJ+���!5t��Cw|������9�����}Ŋ�by���惭�������Œ���h��8o�a���?}A�Sr��v8ciJ�FT޾'#����fO����H�n�z�ѻu0��3:l����A���­�02��韇�'pYBb��������;��s]J<�7�7"^�uu�W�L^�s���VNB�f��~�3a,�/�H��tԨt��UG~)���*�3�?^�q���cr']�\�k�`T��Dm����v��I^�ܽ�˘C��7�*�%M2�PC2��L>0�Mଡ�����ԏ�oXd�q����R$�_���	:���=��sr>Dh�'w0K��b�[��kUϿC&��%0 ���b��e���}n�P��d����yr��m�y�1�T�OFU?�c����S8=�L�t^r�g_/_�
�j�q�-�իW/B��J쀿��]ɶ�G�6��vp���e�7�Pqj���-pbj$�0��UT�U)l�N��Q�u��"ck��<��55=�I��H���)�Tb��y���`�����H�����P�����SQw��VܘC�I�{��{j���8��Zn�E�+ņB�0��N\H"+v����VQ����g��=���=u`��Oh���*�;���t2���7	κ�ň?��3�C��Nе���Ӱqڣ{��;�)�|! 6��1�
�ͰN7�7[˺�2��<��֮���.�����&��UF��(Ƽ��:Àzcϰ(�����U�W�c+Ч9�i�z.�7��O|��8��x=c��#S�*�E�&˫��gV	�a<}���A�g]sOY���x�WF�������:��8�������ܾ�S�x��Ǎ��islE�Pr��*Ͼ��[�Rn����d��0��vk�+��w��uY��q�Py�� �_�6p�����������Z�\c���+�r�{ԽI׌���z�[�3�*r����)��L�Es����a����սl&�,s ����I�q��@�H����yy|��e��0V�a��E��Q���\��R����NseSӝ�yr�f��k=�W;�
8�kf;9Z�¡Ԑ����/9X[<p�n 䘄���-<�j���� ~O�NU���v�)��R@�u��{7� \�����=����W�b��n���Y�����֞g<�X��=	ѹ0�M��� ���r�$ېM|��qw!!���ˑ{A��& ��A��B塚�톶>m��p�'&��:}�t��t�I)5���%�Z2�H̱��پ�53�^M�BI!]�a��w�����r�t>����
轃/K����W��QZ)��+�a�����)�����]�X���
���:��Nu�n�d8��KN}��̬�mB��u�f�k?�-�o�b���3���.���x�Am_̎^��
���ј�é�A� %�KW�	\��[e-.-���`"(�cK	<O�t��G ���;}��R�Kh]�%4��+j 5
��,�s5������;ɖ�\>��*y2��)Tv���%�L
}G����I�*y��V� h$����87�r���PBp�x����Z�J�l~?�fNO5I����^p0Ӟg�O&V81=ۚ]�����_\�cI,�K����۞�"_��t�j�_Ƿ�>�a ��'o��1���U����kī�9�`�ް_�v��5���3�Q�����{��v���ধK��A>�]�`������cX��l�Uu��=�
	�`x�Yk�e.�ge&u���`���[��11����%MP���?�5�#��nU�<69��E�βb�Np�����GE(��^�$,�� ֘Z��)G�/�*���.�E�/�J�C�w��"H�m�k�\��q���nd�d��#u�DA�ZAZk ���k� FV����Y��u���0�I'(1S1��_�1�԰��4�m@@�U7{|.�G`��r�v烨s���~,�#~ܼwx���
�r��iE��c1o�-�_��ڑyC/Lt�<�2>(x�/����=������Vn�|�F;�үИ];�֜);pNW��dR��D���.{ͮ��������vvv�����b�5un{�5�s&w�TIa�'H�,��rEx�`�[�J8�r�Y%��c0}�ժ;�/��z���Mnh�(��z���#�%�]���7�����q�ۧ���
�~D����ޞn���*��M�����x�1��z0V�=~�(oA�5P�r���U��퉘��Hɨ����W�߾�l�@%YWbM�w�g��F�F���9��ҙF��X�fr�/G��\~῿ۿ<k�i_�Aq���u+W�B�|Cj[�6���i-���4��|�޳���v�^��s͠0�%��>�џGv��=�p���Z��)��(�94�໽��"�����=���@�?hY�f�0�#�r�Q2�񮝛>��.�E����Ք1O�;0GR�G����k�qfs�E|���1�w=d�����1�!�����`�`u�|�.�n�����pN6����d�U� �1-����*Y(:�!0r�D��m��
�6����+Λ���\#P���/�������n�Ue^���H�)'����9N�?��6��y���ș����\�o���}
�qV��߿������d��j�F�!�����,�S�t�J����n�`.�8j0+=5�?-������rRa���òG� ����ͳ�S�����M�����D�Շ{�u��׳Z�=��
J;b�<Fk2��1�p�E�'� t͘ꔉ���^Ve|��ʴ?���d�V�O$b۠�_�</�&T�*溒U�+� V���V�nA�1��Y+����Y�H��m��"0� ��׶e'rD�@W�S����s8�ڶ�8�ɦF���U��i'>2H�����U�L�9�dm�	*�(ē¼~�mM�t�����U���_<���u�/\�g��z�{@y�Uf	�u,M�WK?ĵ}�r��\�.�O�����GzӌI�f���T��� m�Ή?��7s���,\����n,�]ڗ��I�+G=�O��"��ի�	}���g��"T��\�����b��$��V����!b8��/��4�����d�*$�;:�eR�t�����~����	���7�	A��HB]�6/�]�y��z�8�3M�
T"hfSl��9��(C��#y^�h��b~�pK?���RFq����h��D<����S_<�
���4�)z? ��{5��`Ôޤ8�}"�t�T�8k����GHG�q����G����v�����1�m9��e�18%  0o���-F	�`/��Ui�D�E�N��+��[jI�[E۝�Ϝ��(���P�(d�}W��%a��ҞW��d�YJ��sE�/�B�(���P����-���Xv��W�E��uHk��ǝ�����$��V���������\�n4�#T[��V�}v9��o�_�Z���Ys��L�w�gN��q��+_�+o�}��4]\k���	�q��bM6�u	��
,%�&Vю��K�N�^�3�Y�VN�X��|��ŨE�B2� �%gs�3s$sd���DA�ޛL�FƹF�|&��l���x�ni�
)���ׯ��?���vEtk�&��AZ�.���l�`��HO��
�������1��yR�qn���
W��l1IϬ�ݹ������6�y_�"�y�p�ys�ռpu,m\}�5��`ʛ|�f���J]��ZY�g� ЮZ�+��ϯ��ɩh-ߊ����3c�����Dq�a#�%�K��ЗaI�x��0��Jɔc�5��]??�����9fR)�:%���U����U�5SJQ6�(��ڷ��6�n�.�z��}jN�yyT\ر���ȏ��3�ߧ]�\4+��M��K����wMo��U4�AK�i؝����$Y��:��S���4_Zhl֪X�X*P�7 �&��P��+k�#|Xs�h�~^������.c&X���^w�B<\�1�Dh���]t2�񩗟�_����n�c�B �[�>X����$_�҈;B?����������f��i�ԭ����;뮃�d��#�vY��	�p�������m���͂J�ng����C��e�q�gXUS�(�j�`n��RF<�A�/���Cz�})Dq)��CsM��%�D��[{�;�תŋ�w;��׹d*�cN�`�BȆ�(�=�x���lU���+S-@^�k�|���subxh�[�h��Pi�m}�k��igJ���߰�TUV���I(>+B)�?�p��^5
$�@��*�yp"V�V��0n��&jd�Ҡ�v�Qk���x�+-c������t3d }n��v��8���yii�HΌ8����[�=;Z��)�H�#وV-�p��%�/0�R�4�����Z�KT�9}9����R������-���b�q���T7w�^�rޫ�,�{?��`L�{���.�q�w�Q��zB�o\��yP�#�m
�J�g��!3Z(�����ʭ7�V'J�l��:1��i��i�މ.9"��Su𠟛ó��u~+"�-��\6$�Eb����C�t` �#�0� "Z0)S;�fCK���9x�J���V�)�4���%غ|�>��&�~tKw�X:P��[3�t�5$�
T��(���߬�S$J�*��4t\f}̉l9*����'���G�h�J_U2����_�71����ae���J0��}�\� {�t�k���
HIpb�V� Im5o���9�l��iH��M����|�3�I���*�ݬ�ua��q1�&�|?cY��pq{��. \-w�P��;��<���뼏1����;"�#N.���B&K�&��T����+�V�i[(�9='`�Zj�'�"�	󫄩��V��>��?ݝ�}ڮ�ya�n	��9�)_�f�Pc΀��h5ɬ�`^
�\!.˛�ˁ���x.��Gobp3����)Oj%�!�R�T�>H<�����򚲥���|o��{�~.�A�,��E�u�d������B���
~�= �Gmn���͎\�b����V%�cȲˤė���,���5V�&Cj�z�ؓ����*7`��B�ީ�w�@�K>n�r���G�B�Bdq��(���@�m��u���s���c�'�Myp4���K#��}��7fOcѮ�����MM�lS��Fn�L��`��]���Ū����ĩ�.!oݗ���,��,!�Z�J̈́�v�X?#rЬ��=*
;���������C�#�
�s�^���-����@��"����5R�y�U6�1�!����nz6D��;�~���J0U(�A:�<:r�i��L�s+�?�'��[��`S2ق�!�!�E�$q8�Xc|?񿋙aWF*��)y���y�v��%6���i�\��*��ð�����-P���o["�(�ʺJI�M�������=�)�C	�}Y!���v)�ΰб����%9:�ݳ��t:P�CD\��D���y����K��w�f3��~���������2�����,( �^�[�s�_f��vu%����l�[Yb��|�+ ���S�m��D���K���;�S`�v�6�L���f)D�G�޿�E
BM�̭ J�y���E�����9?
��~�Ɏ�[ �hb��p��4&#���#�f�� <�XOk[��a�����VFYO���C��WeR������k�$L��t7��ai����c��8�.s��`#h�K5�9�Aв�O�J�A���B��ۏI��2��!�l-��e��#OQ�!�h���p��mYܝM�P(�!R�g�Elή���[��6��O�3��'g�h5��s$EC��ʵ��������t}�����Rcd��"��VH��9p�}K�$ �\����,X[,	�8�U��ձ��vM۝{r�W��=$�5��R2}vQ�M��n��à����L{��Z���$�,�4Q�x�Z���B�nթ��mm�K���:�4b�!�q��S��/��zҏ7����%٠��f
�C�'�񜳪��[GW"(/��V�D�R��|=c�uW.�$�<E����,~#���F�l_w��i�/�@�����ΐ;/��mS9gL��u�
����/-��W�vx�LI�~��_�Ӓ�9��s�(��"�"�&b�ug}_ꮿ�$�촣�x�ԡ�4?/I��n4]�=Өf�r���*뒇��D@W������92�������^�n�����w�����5~`@�������Q��U�05	1���(r6�@~j:�gXT+y2>�n��Y���{G��l������1�-"=w��[��V<�������p}+��ҕO&a�Kb�5i�&��E��$K�aw���y�R�p�vJ�1G�|�H:C�#���V靆��0Ø���Ţ�{�`��ݽ�J_����<+����ف�����W։h،���`e�x�\Vp�1����c$sǴ�o�R�t(n۫t\F�������}Y��L��)˹ޕ������_�K�iCBˡ�
@�JrJ�KA729���PVW�����\_Ga���O6��=Wv�
���P�9��j�{%:�L1�D҇&���q����d�!Cb�%nw�!�S���\�#4��b�l&n���h{��%ߐkǫA�A��ƶJ�w�l�ӳk�G�枑e���C��a��r>ւ�Me~)��?9��]�,>D̐�[���{�<&fEfL
���-�>���زNU?�<���C��P��L����*�ԇ7�퉯v~֕|^&�e�����b#�.�=�R)�{��SX�@./����(�N�kQ�(��.�֞
L�{�|ew'�jW�~/(t���7�0xQ���U��"qA䅱?ʤ��2Z����P�\YJ��6����5`�+���O.�j��Y�=��mm�Z���U
iX`[ �wHMq~X|R�����x^�?�I���ٹ�Aa��q3V�o��z{����m�m��5��V�������*� �?�5u^��Bm�6o{�/��%���J�L�+DfF��VEs����Ȇ��5���6�X�2�����y���q����N,��5=�╩��ю���G�*��3���M���v<K�)����N]8�g�ô#�]��$�w��~�`6@�LX	�4�D�aqW<�̊�K*4���Ӣ?~�jS��@�]���Xl�91��覽�����Rk0��t�Mn�e��?+��?Gd�J�0f�w�� [~�EUU�
�3���(\ �U��8n=�q�~�r.�L�U��I�}
�<�����H�y5���k��l����m�ԃ���T�&�uc�#v�������qyuee�z��ʜ�$�v:_O��cV�ʜr:��|�և�PH�e"����uS��H�7^m�`���m��:�6Yw�l8���,1���Hބ�>�;���ި�'�
�ѳqh�y(��zβX�Wk���(ab�O�	�V�1�
�*f(����&�t���v�\?�G��ۦ���yDV�L �#�����w�0�����<�TI�	�)thF������t����X����!	�/JuwX.I6�}��r.���d ��Q�dd����_�k�b�����'������#Ni]ig����j<�F���?�!�}�9��	��Қ�]Ǭ�>���S�u��h�{+@���������A�E�=!b=(~��d�3kdN�A5�j���q�`��+������5JZ[��b�m��U�����o#����4���(�3�s:��n:$�>Muٰ�C>\�Z�xZb�x��W�l��>UAvZ�Uci�/�C�k�p�ih�d��
��]�}��6��@W�z����bW����?��IŻ>��Q�uNO����γINQ.964q�*�[fC�06�N�.|�O���l�+​1H�$���3_ƃ��yr�j����Jͳ+�'���#�H����?����h�}�rM*Z��)���=��o���[�.�S]__׆�O�W���'�W�(2�>�vt���?���G�!]4�<8��2��,��W��/�s}}��1T|�b�5�������aL�ݦD�~#𜝽�8�Xd���"y�`V�2�����N[� �k�au�E��ոr�u�`D� �
X����gN�jaS��^_n�����e�� d�+��ʆ��exÔ���e��}��K!ɞ����еYTc;�����c�Ou�儷a�������Oމ��)���E6}�2�&��[@�	�"JI�n�35�����Ď�VfJ�_�X7qy0jo�*d��^�=ӅaG�չ�d�,����K���sl�<�3,"��?���S	ʎ�)  ��BÉ
�����Y��\�\Sh�@�]}-,,\��,11Q�|,�A^f���|��U�p����^�ɗ��q��ms7��\9 -�vU��ׂ�$4$�������]�m>�7�l_=��*����|�o� S l�	����EE�H\��fS�=�F��B���;���{�5 �=O����ع��P-�;��I��S�/*�����-NK:���ళ)2����4��Ć���Lw<�\?�B>�ڏ/�t\��b�Q��Ԅe_�w8;XK!�`l�ɪ���}��95���\��"�sxsٿ1��Յ����������EK�;��~Is,q?r���O��Ĭ��Ά��yo5���J^>�w���W��$��D}ǟlث�z�%l|�\�}�<|��UN%�[HW�t@�%�Ƒ�����h�d�@�A���]�!�?��C�78�I�Ƿ���hSx%N����Vg`�%���Ϛx~rJS��(g��|Yr����L�x`ʘ+J-Y�bb{C�*�x���A!��ŧ�����Of4��⨡,뜞O����Y�Y�������s�\OUR�g�ih����]X�'T�-]�J�G%c��>Er *�I��U�p"<PJ$D�-MJ9���v����Rۧ¾����3f��8	�{�_�zn��w{���T�l�i��8NK�urrݣ��;iM�A�ۻ֩�W�E��a�1j�^�qLɟi��s5���^&mv��t&�;ړ���~�{M���<���z��NHu���V�m2湞~����o�m�wX��X�ET�Ob#�r5��i)^k)�)�Pee�P�'�;�J��M�V1��8��L�g����;�X�X�Fq�q�3��ECF�L�u��.��Q��ط�!�t(�#����'s�^�J������5W�1�g�rھ��p�+;z����\{!�;�UUAZ�߬��>�WSO�x�XB�H�^1��
kH�`>i�4��R�L�G�Z >%9�[��Xg$�O�#	��Y04n�A�AH�c('������oc�7⣎n�O�ϑ(S��qA��)���8�����`�qZZ--�О'�ɫt�1���m��u��ګ�O>7���T�~ycv&����T���˿l�7YJd�f�M�bZ�4�CGD��8b�A��j���r��KU��,�T�8-�{.�a��^h{q��v
�/�����;����� 3��ᣅ�[[� �g?��K�7z��~�0�$IG�PN����E�Tݯ�p 1������X�Ú!	$�蚬��%f��R�APq����k��NL����`i�O��!6���
O�(�N�t�=V ��s����Q����i���kg�Z������3��SXs����T���	��rH�s�q�ϰg(|�qhtq��xp9�C�{&+v�bG�]^�g�@��g��́I���pb�N��������I��͍��-��E�5xA����o}��66I11��55;�2�^�QcUaE���*�Pn�f�^�~D-�+�@*��4xd��Ա���&�rpĿ��8' �N>!���O����nl; 5pՅ1]�Cq=&{����7zz�V�G7Yo�~�C�[N{��Q��)��������w���S��D����|_j�B�UЎ�����]X���w�ި��oMj-s(Q�^^�o|������mh�6�y�x������=����I�B��0ol�+Q������^��qR:�^���qZ������ύ�&R.nv��S�o�v�>���ivw��=�7��!�bWH���w`C�pdU]a)&�����>� �X�J;�c �g������{[��,�h�[�6c����{=[�(++���������=�������.�7�ԍ^��9�$���F{ؙ�;��}L0�G��,3�oAh�[oZ��	�V6��i��N��'(��V��b�R��V1vĈ����I{=ID��*e�X��m�{qg�����Fy�o��0jc��'��#j��`~�q���@��C�����m�#gڗO_�>P���D��hO�������x��5,�)�������t)�
SP����*|>{��<=~�*�&�sO��l�6}4N�	���ZM}����t��1�0����Q"���s����̖q����3�����?ߵ>6��f�2�3��"�4��`4���O���6�~s��hWN�^	��o��VnY�#w+���OҚ/���������?'0JU�~���}�ʲ}���R��"�S�V�5n	׷�:��	�+	����X��O~�~0�����و�߬��X��>W!�-����Z���%|k{��H-�Y�j˒1y�Ă�"r�%���oU���3�o��M�����}����&�?8���d��\�ɞ��;G��Ӡ���U���r����"�[�â}uB|ꓡ[�P8��[�B��K�W�[.9��XV-�wV��bVw��ƍ���aƾ�)���x�a[+�cN#�>��Qc����h�h�zǙ�HI,=��g�<o�3���٢/�[S���.8T���i����:���Y��� ޕ�p�]6_�bJ���&��c��+8���"�ŐF!�l�����~����mL�f�������C/�������]IP������k����������'ULM�d
������x3����U�]U"H��RLo�������~�{ZΒ~|QU���n���b����+�HμKy)���I�q�>�^�aB�o����~�o٘z���#�e�/F�/Y֝lJ^u��k�!ɟ31]ٟo���Ӗ��(-�ryC�RI���(�l�2q�ݦr�H_�����?�OȒ��,�e����M�����j�-]"�Hwg�Y�ԕI`�h9�+���{�&��S�k����\}���g�z,�s|�9��uɣ!uN�O��A%�UAI<�Q���~B	�����u1d�}�Й4�
�1&��K���;e\߷��7]�=�⫘p��*Y�z�%�=�"�����t����b+�������.X����ސ��@8^�T�϶��C�9ͷ�P����6�tηSJE���!u}�w(�w���`�F�뜿�;iZ.�6*/�-�sk�I�3E�6� �[�6��t��m��6�χ* �\n�h���)�@�+�u>k&e��QU�.;�5e-������ �o,PyN5�[_�h䕤�k��8�Z�����le˘8^|2+��C%��j�˗7b�� �yF�n2�r�}�zw�{��f���#/9��C���M�����}�J'S�+����@��r0^��Ծ�+�1T���ѽJ͋E�X�y�!Ý9H��9T�YVF=p2ſ�=Nyb��pyz�~��_�5�\
?Fc+�	OBxHRKV��] ��8$����8�;���ƥ��� ����)���G� 7�2)�l���o��5�������A@�6�����	��	��-gv![��ܪ��=�s�-����m���>�^v��˔��[r������rv~NEG�RT��*qn��Z�p�@��q���'+V�|6��S�Z������N�&7�����N��II���g��Ț��C��g����9���-���RM�yi7x�ɰ��C��8y���-{74i#�0�M����y�>ø�@�l�M��?/��>��\�KŘEK��b���a%TfM�I�1nn
�
��}�M�.�Q$��u+>PYFk�%&Fy�t�x��<�yS$���>a
4��a*-8�a���E��{��ts��[�~K(r�<�t�?\^#E�Q����7H�R��L�ATo���#/$`P#V����lo�h�!�*���k�F��K�5k)��mz���Ӧ�8�V0!r	u߾�10�ug�r�m.�W󅎅�nCxF!��T,�^CCC4D㛺��~ďu����oS�d��C7���z�,t����g�B��h��ˣ� \|���K�M�͗�jt�w��!o�<v%�����V�aX�4�]Z3aƜ�Dr0{ru����_�|��w����w=��w&���3�{�����ՋO���Ӵ~�w��W3���;-��~B�D�G��a0�+�p����$3�]����րj�[K[��{��j�E`-b�ּv�� 
Q
9Ί?g�ۑ�@d�~�Y�)}k&�m��e�9�5��̈́���Nk���T����|n�V��C#g�+��}g���UmC��9dz�B�������|ݏ��B�y.@��^�?�蕙��"is��WQ]ݽR���	�gxI |�S�6���Ot��RW͵�U���'!��r�2X1��h�J��M� L�1"������Hd��M���馦����w�o(�(�*�kwF�eHqũDl;M�Dj�;� �;��g"�&NQ*�fy��k��h9���Q�Z�ޚ���1"�[��|��_�^�����-����
�����Ͻ�pJm�oOw�c���N.��_$S����t�!}��l�%<P�rj����Ēq��9)�L���"�>�Tk����B��U��Ԡ��Tǣ��F��S7��e�8,�GO8���d���i��y����gJ�I������5����v�o�^�Gi7�wQ��Y����O.��]'j���0�Vظ	��z��S7,.�	��&@i~��`�}TGd�S��d����p�rT���"���#���n�{ C�H�I-��x O<���x��R�Q�]�GCD%�m��N�W>�-�q6�/X��꾿j��ܤ����J���N�L����7�n��9������0Kn!dd-��U$Xd��@Iz�5X���}�~\Т�G��Zs��VH��Y�>���#ώ�T�����5�I�@"K���Ȁ��U�#�����K�?�D�ӯf�%S��wO]]Ѩ���H�����vM�N#�z渗���K�0^��R�����(�	|m���L������w��w"7�Ywdpz��<�ϯC��{��˒f`��H-R���oϊ2���TU�67m�_\|y��(�5�&��ةp��^ҧc�(������/fGę_?�o��+�h�Q��K|�1TѼ������>@���)���>��t{�Ć�t@��Ĵ['|�V�=��bM���Y���m-#�3��h����Ȃ�?�0<w`���y�?�I��F�9�wMM����dzF�ۧOH$A�җ�Ql�D�u�`w!����ٌʾ�c�=�Ao9+9�3]������ٜ{MWzHE�m�_9�ϳߌ��0�v3h������U�2~�WR�������=�ްÄ��DF���[����q���q��[z��E,>��yqb�f��?�����-L�؁���e��{ 7,�͗����r�4���e��-��J��|f|!�Zfk	|��A7:�M0�!�ӻ�*~iZ|��_�fT�������dQ�%n_�{���j�Ğ��$ ���K�1SlJ.�H��M�3f���G�^�����X��R�}���U���
�.5'��n�}��=�������Q/���P�i8�/�RJ��}����=&#bWj��`����^.�{!��tN�pw�:�� �6u��Rs�ȍ�_�o�ѥP���J���
'�^�K�q�<�Q���jf�1KHi�4��=Ň{8q���{o�l�\���|�ƹ:Q:[�[�=x ��������v��o�áxű۵������JwzF� m��5G�IQя�ToQ�bA���Rh2�ѱ�c+�j���dÑ���� �e7M�3�`��	da�}��ӾY3�ɺY��x���)2>���t�|D=�0!m�٪M����%��(M^�A7�-�~6���+�u�˹��i&���z��.7��i��������x䝻lZ��^C� ������k�9��4_jږ��P�]J��n�H��e�2um�G2��\L<h��%������� �[�&q3�C�������hQ1���X���������)&�Fi��Ȋ1y����dh_�{Q���?�	��"��A���]��N9P�Z��dq披��T�&�u���Qf}����o��2��&x���$�ц�Q�kF�M!����Z�h�w������+Eb�Q$��Ea#��7�*�lXTO��p��ny�4�條�-����eA�����ZQ>+F�/>�gu���I�w,o�2��~��g��v�}yQ?|F�CA�v튒�H��`��5]��=��Y� ȷ�Npy�<%xX������Z,��B�R0;H�P<�3�ͦ�q�2�/�yR,�e_��`
;6K��o[K�x���ˡ�z�H4m�N�rōQ����(�2����Cb}�>��9�K��:��d���x�Θ�l��J�n�l�8g6奊fJ\=�o�I�:��g��sk��;;��8#��M�86^�>'�oTu��ѱ�;&l�a�Kul���F�2
��^"mUd����p��C��`�6�:�U���?HSl��q����w���O���|m�ڗ������W7W�+����1�ic	E���SS�E;��I�V�6i�[�H�l�s����
�=V[����]r��j)�x��L���W�k�wr���%؊��9�fJ�P��H�B4~Uѥ�i�b�[��|�4G�"�ޤN��`ժ4�"�%|N�TWs޶UÏ�xP�𞫘��ŻYZH� ���
�� ��E:���G$8�4l):�;�����5�+W��'qq�)(�|Q'�;�1U|�] ��D���=�~d�*��f���."��<�\\nn.G�f�"�C1Q10������{�k���ZwN�ذ�'�|\�ɴ�c�;�ݏ~yC俸�O��֔�Y�I��95�������T�:��ߙ�tv���{�5x�F����V��e���K�җv�����E������ox�>��OW�v+��6�v�H��l{|4n�{X�1���s����7�E�!�x���p�r�w�@�fu���b�k��r��o/iN)S���߅M���q������~����1� �}WAzw �+�瓘�pZ'�K����H�p`o�۳S��$�F�y�c�K#<���nZv!x���fՂ���(}�׾��r�S��.�D�[	"��j�iFו�)� ������O !/9h�(�).�{�0d���p����ˈM-�-?�=��ǐd���?T:����T�s��ʄ������=�C��VVQ?=-8�̑i|	�3i�\P=̐��}tQ���S
~2z N��+����/�/�xA�	�l3�+����	�n�4N�,�w�}j9<$��Tc�(_X�����w~�{���U.֎�-�Ql��D���Q~'����-���OծD���@���O���R�:���G��^`VGnń@L��۠7���p��H�{��Pܐ�[�q��0
���_.���1g����q�)b$���]u�K�Ys�oKF/B�$(\�"����UM�o����R�qO��#�o}��-�i�����R���j~->�	k���\9���?��b%cb/?�u��ϴT<�E�Cc_E?6M���9߆/EH�B�<�Pag�`>x�9@�T=�z�b��S��*-.cE��|�9'ZΖy��ޘ�u�;55���y�mu^���H��̕�X
RtV� ��;�HP�Iq��Fñ�!�0`��<�(�4�u9���h=����7�=���p��1�ţ���{n��6���wG��}�.QI�Τ7�X�#6�|U���g� �L�f�*A�]_J���#]��\��lq��|�T�IL�t(L��S�p��wi�e4���>�w4��)�K-���< ��m@wB�;�HQv��Zm�qk���㝋y�F�ܬ�Aa$���Fv����X�e�L(S:� p���猤������ !��f���������g:��4�Ǳl��������L!��o�o�-_��
������z�V��X��Ձ����k/8JGrka��ڢ��B˷�h���"?Ψo���_��͡��!)|fG�;�+�_�o�ۃ%�V
������3�Բ�9]�<�/��&B��U���F\I�}��\}w4�[�"�� D'�=z/A"J����h��Nb�����k��F݈��A�r����{kY˚f�s�ޟ��~��d55��YQ_���1��y<��21~\zzQCmMD6x�wF����^Y{!Z�OB˱SIun�m��Ŝ��+�{��4e�a�O���_A	���y�P(Lt)���wuA��}ťh&@$i�w*6�o��]4�e�Yb}{;���z���K�e����5 �=z���3��b������ˁ������߿�uK��R7�䷏?1���R�;�n��UB�(�� Sh'-�g}\���j��Lr��O@����)�S���湡�}�hXv�3�x��*}�ظ
�!�W��@�6|�C9��i |���\�{lb~R(}�W�d�G�T��W �%^#��=$|g�0?t�M<����w���@��u�*((7����}������(	r�}\LR��+�Y
/Nn%\��8���xuhs2��F�}嗡�]M���(~��֣;�cgD����(y|~�~����8l]����,f?9��������6�T�G�Xϻ��X��̅*K�gZ�Y�oz� �;���@���$�������ۡުBl����Z��]�6>� �ϊ�eh*ߤ�A��}Y�o?�ϰQ�7���U���K����,��3M��S�h*�J`��#��Ŕ۟����.���9<F�$��j-L{��~�����>�t���W�СQa�L���j��lxaD�o�x�[�3�#x1Ϥ�2\1�
WT5h����(st��_����o�o��%�{t�9V�1n��'rT�9�����I��/��P��)�`�._��V�
��&ྮ�m	���J���N�g����\�&oJ��0��h(>�R�J�6��Zh��H\l�����Xj�|���X"$"$���^	�ɪ�k��$zD���F*��w���+u��(�׳װ�����{��n����gxC�M�ѯ������x�����O�~*q�3���k���{5S�`��|��~H(�uuTo����h��@�&�uY�}����2��TcW+ӹE��P'���ח�����GGd�%o#�(��,&D,�O��`�IT��	C�;P4EG�����J��	����S� ���J�V�ƛ���"�|�-��GYm�<Pp�iw�{K�doK!֫i�ʿ�i��)�YuGh�8�I�6g����RM����
�ݯ/P�2N����*���u��Q/��\I�yo��J3d����#�/�9�A��|��9�j�x�j˿�?��㏔���Í/5��L^����545����oD:1@E�ɑ]VǗ����h�i���]-��4ͻ���m,���q�4�&E�I^��&븢�������р���mh#��}�^G�$(�n�mܟA�>,�U�N��6=�q�B��z�0OX!hgg�!�k���N�B2�����r]�ov[~�f�q�Q0�����_�e&��6��Z�Ϗ�RV����כ�f[\?0��^���fд�9����F�2xz��$�G�5��u>�b~��o����`v��jۛ�P�|�K����N@����U<p2,kl��mg`
�ө�A6�@��<^q�$i8
�s����2M�k��4�mT����8����{(-2�����Խ�P���OsҮ���3DS���wN�JV�+�|;Moǣ�p������j�]��<��y �Tq� �V� ,�'�hгŢ� q֋�*�Q>X0��O5Y���H��z"���a<t0���z5wx0�~&�М�S����D�F�Vw������e�ua�b��f��߷_<����us����Rf��.v�8S�WS�'�q��$���>㋄����O$���jH��tZ���1� �d�%���pa��*D�e���w/k�E}Ѯ��vd�����K�Լ�j���E��-�N�#�dcӫ�������s��� SXM�]*L�ziL
��Rv��E��)~kJ�,i��f�aJ'��"wB(|:�z�(�8�s'�|gs����>�͸i�|���$�={ٌ��%�fS�t����F��\<���.�Q{4�?��ko�]&))r<��)&�k��}�Z铲�5��ګ<z)?�!0��V/��"9}Vhm��x���g���K��!>��bP�ެı"�1�">���l��7Uu�C���r�@�������k
���=o�)` %}�c�(yn���� m������L����X�D3�(���U�\K�.cq��r����HBx�(-j.���0����[C��ňf�Wg����������?|ȫd����̚f����PyO�1����[��*���1�LL�i�feg����������0��V�G"��|�p�L��A8��q��*Y��aլ�Ǔ%���,1�0�	� I��OoF餚�چl"W�߻v��]^ �{�xZV��@�V�Z��t&�^�-"���L����ւEݲ�oW��3b�UNg0 2X-��cs�)��3a@�Ƨ1��$��vk��!c8%'�Z}gb��L�C�%���_B�'�4s��h�; De�Q�S���憑zQ�{~�nnNo�}�c����M&�>[ ���.����QR2����P�C�HbEEۀ'B
[�@lE�J0�p�ܵR�@$�tO���!�D��{.� ����� ��B9�	[=Uߢ�9�J��cé�Mk���J���C�E8b��	!uQ�}��������j��%$���H%=K��x�M�K��-t@�=6d�g�����pMj9�%N����+3��L��[�����o�RI�#k��S5�,0��
�˸XV�6�O^��������.K�ԃ�^�nJZ�(�\�g374�̘%���<o���\��0.C���}�<2b��55"��Pٷw�6�mq��x�+XKð֡������\�@����"��j��Y��~x.���U�+F���aMF� $r��b�T��=�S�WZ�~Lxw��p� �&\���=�&�¢C�.�5�oҩ88ʖ�����]L�u[ԩ��Gy;ZQb��f�i/��y/d��/t����UX�j���@��;�����������A>Y�[�E4݌�z�`���6����b�)maP���lmug����c����+ph�R�4���]���Un��u:�v�߲��2Z�&���%�S�IŷE��1Ip0��7T�
hD�y3�x����h��*cƨf/F뵠$�# ��ՠ��W���eW'6�ۈ�ȡ����¼���a��<�B �Ha�ceռ�$��BY#�ެ]O��P*e�W�v��U�޻�Y��1"�i;��8IO���g$�m�à�h*�N���j�?�CB� K!ӟ���J�]V=dN7�X]QQ�7�T�	c�*.��-/a&���d/v&2��S�i��Bj��F@s'�*�N.z�T^�,k_����)L�2|٣c��؟��mk��<������k�w���kUZ�����d�=b�,����`l�0�Pl&~��}@sL\���(�X+���i�ت"
/��3��b���M�1[���}�3j����:�X�^��{�ane���Q��]u�/|�ٔ�)�uL���N�6���><�õ_"n�WӬ]���oL+fր�O62�6�{Z�����������<��6���rU\Q��A��&I��h����=�32�ը�R��-U /ƪ#p���Ik�q��j���JH!�ƞa�MF/臧�:��Uil�1w� ��8Y<��kJ��
( �� ��������q5�!�4�͘u�k*ڼ��{� � �}�ѧ(�1����~�����5�ǻ։��4��U�@S�>�:�J�����y�ڤ�CC�i�btx]����8�`i7޽�!{) ��;�|�L����E�E�j��߮����o������q�k����3�|������� �"rܘ��))\c���1Č�W$M���d
��z�k��D���!�ado�?�Ov���3a��G���N³���~��9�|2(Ō����N%`��tZ��ō|�L�# �A��m�I�4��v �US9,m�b�/z/DC���HXJ�m3�9��
�"F0������r5�ehYJllmK ���F�BS�sI����4��Rὑ�3~Qܦ�v� t�x�ǢLT��i~�5ӁY���U뷫��Q��a����H.t���:�qފ���]�˯�O��G�t]�tH��]�������V��9�.���{�vG ��b!�l�\�>�4��qϦ�����3)��7'�����ti 9����mյM,c���f��VՈw�g��xBs��.���0����a���wP� k8�#�}ԚaS��)(/�(oq}�Tׅ��=����ә��1�sq!F`����?����5�Z)�49T��s�� R�UE�\B(%-��")�oA�i/���Y��\|�1�#�`!����<+�\�a��?"p�����t�K��O��n]�RA�B�nn����u P��yE�@�p�d�'q�C-D%rV�7Qe�~F�M�\2+����Sa6�W��J+QM2UĒ
�O�_�فl��ӐD��1WrV	�a�z�����[�8�����GF
:�.�m��$�BSp+Ϥ��1�
C|��d�к��ݾ�VC�5��C@�i�s{H&뛍N�,#Z�p��x�5�sgk�\m��n�������x���<�j��V�U>պJ�����?Wd����+�ɷ���]����ȳt��w����266�o�媉=a�j���:�u�v���̚���y�����W�7L��7hs�oG�E���g����`�|�q��R;0[l��/#�q�$l[b0#׉+�����x7�߁��C9��h����΍����� �# ��]�4ԟ����Vb6�Ѹ��ԟ+�K߁ W��1#B]g���^v�]{�b�@�ŏ,�x?9��^�W��Ϧ��Mٽ.�ġ�����.r-�ׅ���AX��eܱ�<�*ݏ&�C��W�pQӘ�R��_�m{�ndf�FG�6�񗃫=�4Ο�����}���xIpJ��h�xrp� �N�B��0�b*}�b����/C��lt^Ů���3&?��}.A���94�0i v�u�l+~��,���z��i�y��w`���u<6K��ٷ��\�aI7q0w;T�D�D����C��m�mF�Ukþ*U�.��I؉GW� �F�ac����I��w�@j�(�[9�1{Hr���H��
[U�X{�[��D�m�M;]M	�$�-��E��2����?�g���l�?��l� �R�Z{��x������S6{,/�dۖ�� a]��N��."[D��=B�E���v� y��Z_��)��In�P�gԤi�*ϊ>�wg��T�`�ٽ6g��/�v��l��>�����1q�7�螤d1	��l.;6�X]��#ÌB���]
,���q����c����qnϠ�w�	�p~I!}�"P4Y:�m���r�~�&���H�k�K�F)���q���Y3(��Ϲ%��|&����̔��{���_>��9Y��>��
��K�|����ƫ��CrN���&�vB�pų���5CJp��l��o�{���8��@�Ԉ��=8�Ia5���J���ס�(�\�t���Ȋl/����Ϟ9-��١�J�=�dkE3��MA@��	XYR��B����ևS�3̃Gn��WBoU�-ڭ�=.MG�'�0��Yd��ƾ���*�'�k�Q-�}�Ӷq|�S7���һBw��:k2�����_�7x�Z.�����4D�M��7U�`��E�F�L������ߖz({�x�0�I���«�[}�5yQў���9!�@
Fh'(Fı�<�$R�nv�Y��ˉ���m�vm۞�T��R�З.�m��{p(��s� �C��8T�~F&�9�����#��!�Rݤ)�
�o+�1�.օ���4>��e,����
x9/�n��?A��Ěj�#?r�\z�]�J���x�5
_=�	���g����
���9�A3r�Q�wY���|�3�_���ۣ�6���,~oS�Ӹ�l��%���1x�Y�ptѲ��g	%d%���T�=(�ō�Q��i��g�g/��G��ĝś����f�
R���<��	V9U���M?�E���9�1jh�g����RIV�$�x۶��j� -N�T��,g*ܒN	�)#�������o�b���K�����T֫ �.F���~n�?��T�Mv*���x����m.�I�yx�7]Qc����v�p�͈����P��ʷ~9$����7���̃oùsgZ���aaπD��T	��w �3�����u�' gyrrq�9��G��S�M���F�;b���=�2�rTi���C��O��,��>BN8O�M�b�Ɲ�7�vὛ|ڏA1�!�G�TLw��T"�J{J.��Ҳ'��E���*8*v7+��?~�o�Wݶ��8-s��>�G'�ߊ�07PI�ٴ���=̊n�.	�@*X:
l~Ӂד	^��d:)$pO.��L| �����6((7�[��=���>�
�8ެ;�������̎��<�i��WLV���ю������)�Nw⼈��S�*��;�x��� �-5��g>����H�E��:r-~�'CK�ia�m��C����e�v����s���N����5�6�2t���a��ibl�;@]8���W������ͪ�О^����E�8&7!=4�Ҹw@�ӟ������ y��R%�s��V���[穝j����y�gKpDgyZ�N��+K�|���֎�v)��a�q��D3S�ő�]�(2fx�7���ʔش��-"�˃�P>��L'�)(�%i$��)��"��l�:��pI������ԭ�rrB��`�&boݵ�/zna��5[�2���)�ò��E@Bb`:(�Q��������J_?��n0_�b��)޶���P�����3�,b*�SU�.�2��H8�$r���W+�ǭ������zn��i�9�BSU�I��z�2�z�a�(��;-yʯ�%��=~�0�֟��4ASt��=��� )�}a��{��*��!���AC��[�zvY�|��YfD�{��,$0( ���z��'UZ���I�P��Ef�)N׫��a�Fsk�c��aqȓo�;�?��K����lO0A��#�cj�Q�U���z2�2Ӈ�є~�y+&i��'����@���l9��_P'*?�A��(��(����32}@H�:PL�LI��q��b�3� 陘P�s�q"�%5����KUo�й��>�7zײ]���~U!I@�*��l�D�T8�ھ�yچ��a	%6K�\���Y2R����~[���cج�: Mcf�쳥/���mD�\���6\LM���].�:����H�?�H}qO����&:l��h �}�ީ"w�6��f��UNG��D����V���/&�hB�lX|��(�Е�o|��3��tORi�K���%�'}�M�
� �lL?�R�{N�s&ꚺy9��[�	��!���_[i�x�Ni��z��)������?"&q�{��T�oK����T�	������������yڹ����<M��K(Gm��F幈�X��Ǽ%��� ׁ�v�m݁ǝC�ȴ��WR�W#T�@X\�wL:����b��%6%�rةF�$�0�=y{Zj���󙪗n����:� 0�Q�ϟ�Y�)#�h�U�ʈ��߾�����C�T[�@��(�����k�?��"W�A���0ׯ�����ր���:�ju�ۨ��{�R���%�N;�/� ��Z-+��f�L��LW�޳��_�+'���:�`�I�|�s�_3G�_�zb�n��0�pO>�̞��r�f��񸗞�^K�֩�O�� ��ut�:yW����r�r:���e�N���/o��x���s�$��+�����*.�1�;R�}2_;S�I4�O1��f���,���`��qm��'#���.H{���%w������œ�����N�?GB'ҥ(�'����v�3��O�a���z�7�� �l�-T������C��-%���a��(7��uԏ�����a6J����±굖vm,k�KeA΀� #)�����i8��CGj[�BKj�~���#�P������RW�''��
�<�V:[�k-���`s��t;la�t��R���y�ũ�����:-���!�[���Ssx�|���{�z$_J�9�\��{Y�*���)�]�p��qqw����6_'[o��wQg�L���`��4��Pf-�FK�02�awxTU��Q����$����[�Ax�ڶ��`���D���-�R��&�.ې��+��;.C���$����\W�z�n�ĭ6�O�r$�er��ܚx1#��;:�1xW�_ZG �a*����:Hݍcv���n���|l��lFn10Et9 �Qq��b�R y�$����tХ��5�A��,����?-�DN<��Os�;���/t!�X]҉�a~�D�>I��l��w����n�sI���B}��������Ŏ{��-���^�[�>��S!�&ZD�/>��X\��bj�Qfw��^r���u�D>媢�*>�Z%��;+��0kMzJ�\E�0#�[�\�G0�xֲ�s��b�������	�4�|W��zXO���s��G���w������+S�������n����C�f� ���qy���=����t�JsE�o��zi�˥_�X?5}į���i��z���-ն.Z�� d�q�\ e�m��-�C��7��i?�t���c�̈-�[�}�ר��\Mv��\0���p��"������>;�±��K��u k��$�v�>�]Z�3���ߔ�x�Yo�d�|��ޣPM�k�]׃�fQ;����ԽUƴ�b/g�݄1#���tT��a�@|[SU{�<��B�*._�����#q���p�1O���ms�s��B$?��0����X�3���[yT&�������}Ox���������������I�zIH��U��@*O���{��X�H��e���{��l?���م�rY4E��!�WZ'�}�n�t���$��圖�p��p^�"���Gdh'�4�9(���]������j9�y0x'=�K��gl�WK>捗�֤��C^�����v��s���3J��1�nX���'�!�Uqgò���t�Z����ͪ�Jo����n_g�gZvX�����M?M��@�������MN�x����P��F�:��3y<�<A��yVȂ�(B��M�����w�V��|ـ�m�;�s�7�-u�&Q���N���*%����YN (%#�����xv��w5M����8�fvW	s-�K1I?�S	3uٚ���)�v*ϰE��
)��fm�˼��{W7���ՆM]�5c�k�[okGV�D��A�I�|��g�_�Y�?�o��n�;8�^*?��n�������:-�ԡ�[O�J���S�b��5j�,c^��	��w�:e[P���t��^O��0���&׷�}�]Br����/9E����;���P���v��Q�t�&mr��������/Q�������y��c|��P����~e�!�⣵��5f���/�����nO1q��P�j�~KUg��5J%�ۿ�j��c�˹]p�idDgP�����������?���3��&a�EU�$z�Z�)V����hЗ� 5G�R�Ҡ-��\O�H~|��#c�0�dqM�%�;���w�*�J:�W\�v�c��^1��ذ���B��g����Q���?��:�����(�Զ�<ŋ1��W{��k:ϕ������Q1�6�?~���KCȈ�d�5���$��ަ�*086��y����[���!��C�=FjT0W	{]��׃i3��]��mAח��<�]iI��@��p�a>q'��/�_�P��m�t���ژ̴o�b�L�2�bQ�$�2Z�>���������G�����EE�}���7F�8�y���ϵgҸ@��?�wcK�d$,2��J�+䏣����1�"U�*�\�]���A#/u0R���+YK� U���rJ��!���J��&4p2���P�w��~�BPVV���1٭+X�W�V,�[�!ڪ�ih��-P���_�F)���Y۽�W:9�e�զ�/ejj&�ck� <�Z�-?b|�\N/��Y�}{��w��\��Zz"����8�X�<�&ޕ솞e@r���2���^�n�F\S-P���-�����X�吁3(�dN�鴾��
`d%��y�� *���4Y�τ-+<}dm3/�Y��;1~��Bn�>�����ׅ=ұ ��Y��j�ٳ/ ��dv�;֥��mc.�NA\Q�i�6n\A�Z��n"����-�X����\1�<n�kl-���8���A�7����7�������l/��4S�it������XBٯ���	j�m\җ��u4%:���3y�-H�Ld}���[e7o��Q��g�V�T�r��W�)����N��E|�m�57�-����tHp�y��s��a�3G��E*�W��qT{i*JA�	fѼ%oұ�1"�@O��;0�d }��
^K�.H �:=��3�����z^���u�G��'N>b?�R�	�A����;��H���u�x���~����BB�������ms�-�z���������˽v�q�j���/s��4�g��Ǫ����L���N]jO&�IR֮$���w��YV�	�QYQG}�Msbً��^�LLJ���in����JG��*4��s��L)�b�/��?�]@]y�s�{��IA@UtĴ\��q��~��@�v���6t#���&��R,��DcϞ��W��tꨂ��4V\l�i]$(�|n��/�������K(��Wl�9���r�r7��L�9c֜?i�����X� ��WU9N[y+���?�<��6�D�绀�mf?��g\�]V����7��h�"j�fH����m�:������l���&I�ޞ��w)���-�cc����E4Le���#���
��n�H�W�>^�������b����6���<����r~��բ!��:�����b{�	t��e~!�}Vu�}��1lM�:=���S�]����:���*˹���e��t5<2�K)�`Yj�%W�YC�Wg�d_�'dAK�S��U��~��xnnW�4�a�%�ݰ"�gw���70M�(�O��"�b���p�*euV��<r<���-0��ܜO��������럙�]7[�M��o3>���"A�w�:��C�`S��_�d�����,�{C�N�h��~7�1µ�$���L6�O�46�iۋ�mE2ƆQ���'�F_4��ՙ�N��y���eS�Ϸ�����l�#��Ҳ��$nє���P�ٕ:p��٢��[�;@SW��i|`n7H�"|��<�z���zUaԡVp:�E�x�0�0��s<=b93���$@�?S�����F��p/L�}ow��zduu����l���V�Wbssy�Ϗ��nÈ
�(뗻�.>�����R�Ǝ5g(U����Tm�*����6&�F�b�A�V�T��~R����8h���>Ͼ�eW�9Yߔ�>�1`�C�Y�a2&�ʱ�X5�u�q�"�	�>7z��i��{��a/���$�k+�9O����CV��o���TB�+��;��C/c�T�Mڡ��J��H��_��s��k�/ÜK�	<��:
��z={��_\Н�/S��-�1�!�Uu!�m8��A �"����'���*�.{^/�,ӼU�	MU������*h�k��G.�/s�
�3�D�Y|�I�
 �%�X�c�����Mf-���lR��u�ԭ�6�&�b�+`�a�u�ey2�0�>m��
�X*���I����5��O� J��G$
D��0K=z:-Ã��7�=������s��Î!C�o���kJ�](Qx��sc˺��^��,�(S�WP�j�E�.��4���[���_O��[��-_�.<?_O���+RI���A�cbbQ��m��Pi-^y@Ɂw�#~��,���i�\u�)5'.]I��hi(l�k���y�!�����h��p�҈0�Gp�e���;��y8�!	�p��4_�\#r������QЂ���S�͟$��Iϔi�Hj8��k�� �k�qznٶ_�T�+�uZ	���(��򨆗��6|]Zm�޿�k��|-f̿R���kA�v��eR](��_��`�9T6���PRS�]���C� ��Ko4G�?=����mdg���[^��ɭr��N��[�i)e�s��2�23|��l�]�.�{e���d+K^�7�h[$�DY
r�j'@��P�E(�л��.8��7u_�u�����;���P�o���ȫN�BӜ�~ɖ��~b��;J�jߘ���||�/Z�3��p�&1�\0EqN��i�ab�;?�#�-B�b��k��v�m�큔����x��w�`�ʮ��BWE�ըCE9+��r��`E\�S�߶��]�F���y���B��������L���(eE��D��f��>S��T��:��&��89�P��4n�!� A��q���R�0W�;U8� @V��U�[�_5��K^�,��܌C�ۘd�SP5#���i�}��{2��a�~�^�����!����E̼�+�D��xb����#;hŞ4Ѵ#���n��1���o?�����{n�#qvC�vc�5`�f�
ciCʫT:뼬ˤ17����g����_U��Ή�&���y���'*�i�2�������G��R�Ǒ��v��^�l�����G�:A\���6|ˮ�
ExC�wc(R����TRw$����(sxnc��j�'����Eg�����%����0p�~�`Y�<�pR�(��� �h����a�r8*��N�e*�xkN�B
F�x����i\R._j��r��.`B�R�!���ɩrs�Z}�� �vsQt��[R��]z}F�^d�J�����.�גLo���R�v��d^�Q\3������Ŵ��@%B0뤣v�ACp�]\\�����i}s��@��һ5�øG��l���ܜ�?�ƎTh��^P�����#Ԟ�.���	1�����=)Q됀*�/�#0j[��m����2>��pP��R���@Z��kF�Y�gVo���=8!�vO�ڽ�����H��fM}?�V�:�~�q���|��Y44�II�/,H�{�:ˡ9��Iq
��Ռ�JL×J���l���݌wpS_����0�ILDG#�ʅ��;����jV/��+e>�����ں:������1b_�Y8�]HH>b<����Y�e���b��8kw��� ���X�O۷���]Z��f�j�J�Z�Wx%��I�5,�+l%ʃ����v�����`�������6����.��[�q�n[�d�z3�s3��W�Ϲ;�"xk
Ҕ���V�02�J`�qZ�8+�Փ��8�H��[۬�:Sm��9�Y9� Iy��\��O"�B�^�5�N���7�߆��Nm�L�/ĵ�-#�.�:,>"�逊)�Vj����wZ)��6��B����|��������`^��E�ÉXI�^�P��H����"4
�s�p���2���`�Jh�ьl��b���b�V�"?JHd#>J�����]����k�\����x�J���Qql��c��}��u�i����`+:�0�T��=���ɀ
)�����������^Σ$�'x��k7����V/w:��A��ooԳu�<(юj���
v��o�jl�TLg1�w3:�4���lY4$�0���J�[�(R��;wG��_%����.�14���_"k���������/˷�@z;O�h�� Z�|#_���#��e�7�|&������k��̽���O�b���!`�ꨒF$(I��_��ƕ!۸^uL�;0}��z��f������t"��v�d}�[i�s+WBl�j�����?�q)n��fUն	��Wp��C�/�v()�
�-s��݈z���e�1�@3�~б�~ZE�_��5x����n���V�YNr�(ޡ(�瞄����4�P6Ǻ����]e:�kll����z��U�f����[�Ӽ�x`��I-��2J����B�y^��� 'h�U{I}.n��ei{#��zoJ˵�m蝟٣�h���)V��6���|cO֞[�N�i�Jg!a�I�*�O�Ȯ��֕��Y�<p*}!�$�#��H\&VA�jG�Q��!��c��N`������Ӝ�`?�s��4{ݵ�90-*ލ���_Q�D��T��-�� �Q�&\n�WZP�Q^�w�/'�ӗ��G~v57���_\�2#�~���f�H٣�t&�ւo������K}�[U�h�]v�2�H��h��
��snpLhszC" �"�,�/g��	�/�Gv�6/j�� �����ewI�Kl�[��sI�yMZ��7G�8-�V	{�Ŝ�#>5M����'7<d�O-En D���s1�7��!'۸M�y䪯���X~2B>�v&"�����y��om�̳�OOLL�<!���
�|��I!�[�JCQ��p4&�8��v�pm	d���0+�̣�~6E=�.����@Y��k=�X��;	Z��l�Y+��w�>�R�T�

PM$���?|�x���mn*��@�]�v�V��Q����P	M,: �q��R�|pX���ώ�1����M�y�J��]���M�zv�_���~�H�\�t���0� �Ux�a�^��;ش�[�4$�������@t�9��E�g�������Y��8�:?���^��'7���{����铓:P(t�m;��(�U&�;��KJ�1N{@6�c����I4V{#5���X�;�㴉�@mUoS�b�OI/���c_&�)�'+ N=�����M����_~z���z	�,	��p�Bl*�̰iECY5�iV�����x� ��h�%L�D��,B�Hz}���v�}do����R+����6_b��@G�I���2W�9i,�t*�w��ERx[������if>"�bF�C~�m�r��L��Lu��÷�J\F�����[�Ⱦn���a�{�9���j�d=���ZB���oF�Y�h�/^�IBkE�a-Uȡ��O�8���Ө�ʑHs�_GR�
PP���ɵ���c��C�ݠ`�k/����6��͂=�n@��%:�Uf���I�&4�h?v��^��Y�bH-4B��mg�����@Ǧ�h�fF��w�`����U7�m����M�m�zig�a$��eU�H��6�G]__w���/S�n�0@���n}{���x�F_������x;Z25o��:d}`�T��b�I+���H���4-=֯ycj�q�l��K�^!_c}TR�XZ�_�ʕ�?plD}��V&pi�a�'KI5QF���D�W�M^�I�J�xG�p��e�މU�:�1�mQ�f�f��7̮D�>�w��6׹�-�yWj+_Ҩ#�f�0Yc-�v�R�4Dg�%F��̕*g������g渵��8����ңn��]��W�*�RV�n){U<n{::Z�,iOP��(ۼz���`)is�ծ2{ު6����g��X��᛹vO�(7�����J���:�R[��)r��|��j]U����U���n�Q?4����Ҁ/�����g,RD<�~TB�lp�wp')4�e!K,�� :�ˈ5�)�a}q+ H�(���Z7���~�t������t ���~s/P��2כ���FW�{6A�����%����]�!�#A6�� HRQQ`I\�+Q���q0��2T�t�g%g_j����i,�3��{E�f���*.UO'+�Ɖ�����j�ɍ��4'��%��
R�U8����)`m,Պ0�1/q��c�R��Ĝ�Wmp)/��X<��ߧ���H��'�V,�Jj������G,5zT��ij0��m��Xk;�*����?*���N�Ws]�}�[�3cw�t\28���B��䐆/'Y_�Dܘb]���7!�3���ͱ��%��B�[ڻR�]X�m����}iߒ���=8@_�b���$����7�[,�壝���{��H_hV�_���yZ}O�J����pT�n�٧�{�Խk��U�)D�b�B���Ȃ�������\bvNߍvvVí���@xfx,o1n���PV(��
��(��P�n�ߠ�Y�Z$�f���]*H�7M��
���g׸��+��2�#֪�N������f}��q�ՏH���ג[��]��h,����}[���P�g8�i�\�;��a�Sc�s���O~���љ��[$'�:+�D@yք�]�3SB�h!_yJ"=�=�}ju�g���}�i�9��0����7���Pۓ�0�G<\�*�p���^U-�#1]%�AdgG����e�NB��T�'�dv>h?w�T݆��]!���F��>=�{H�Mw�����; ����X�;,7��N�"��G⿽ l�f�C���{�I�5�퇹'�[�P3J����eH^�����r�]��Xda��q]sb���gFqe/=.6�R�#��t}/O8dU�	�6��\�#���.�e-�X"	I�m셲S�}��wƘ,Y"*�d��%1������Y�>c_>��9��?|�?�>�{_�}_�}?�����5���g�Y��w_H����r+A����\���4iJq����OY?1T�s^�cο���^�g��>?;'��2~7�H�}y�o�[~c�%�E��Nը�)>?ޙ��nn�9z�O��¶�@��(�@ϭ�B�C�Fj����e�����dC��u�>���C oN]��!��-��Z1oL{��.~P��_w٦wϬ����Uk?���ai!<~Ăp^��9�3�tɒ���>�vnH/�����NS��,����.Di*�27����Ъ`y%��A��5��):M�\@�7
z֜~���s�W
n\=�����:x�c_�m�?[��Cá�@��yb3�M��{��2�%e�v؞�GQR3�X�l���Ii�n��S��b�#L�A����BR+q��`u��Z�ߊ�W1r�]�w�k��f���ߕ�'���{���(A z������.t3�#����<\�{�	:��)F�Waf�}�ӹ�;�����4Yv���t1˾yu��7��Z��6�����Y�eK<�_�ځѓu�\������n���_znm�<�0�(&s�}Xz����gC�i3�^mA�xL�V��{n���06i���-�������J[d����a���r}�[q̢4�L�����~���~V)8�g}����^�J�@<;��|�I"��_��E������u�� 7�`����1,�
hu܈���O6EB2+��� ���,�+ސ��xۚX�9^�_"�ŀ��[.f��Xn������zr�2��T���6XrZ�
�)���l\�kիo�3l�iM�@n_���"Śi��J�����>90l3�{���f7���{B{�g'00='١0�칳����~���qP��&�\����i2$�o7�-]�=S��5礼i�����A���X�2�fG	��z�S2��V�J�aRs���#C~�AM�'&�7�5�wj�;Ws��?l�g`T��ݏ}��%��h�F�Y��}q�"�Q�ߠN�T�ݔmHTۻf�cD��x��+�/>ݧ��!�mr��90�*�T�,�O�g�~u]։j9�e`�6���*	�G���;z,��k�0�1z!�`�uS�/���,��]]y�_�4:�p9o��^��~q�����d���%o����\�r`����
����볒���t؟̇���T��B��I6�.����Z�"���ֿ��j���?_zY�"Z��#OW��m~�
P�	+��,��ϡ�Yp��4St�ڻAv4)��EEv�ė��p�����BER�B~p/��)7����U�#�a������4o�Y>�?a��vF�hXЦ��_��r(u�&��G*'�}��on������� ;2�4$�O����pQ�V@e�>]?��}V�Q�a����vƧ�=���π�	��>�����g��4���Z��.6-Q�YǮ���u���<��]��C��4�;,�^ea1�>�x���1T��G������튾MQ��+Efs�C�������H1����˻i��)���(����;�����ѱ1��4��[V[��Ip�/*��T/ѐ5��n��@$W����$�R)
ǃ�_*G�kz�8.������M]��Q�煴�iQ��2���"��U�@f�]��"9�Ir�>�Cܶy¡8�-���Q��~�X�`�����z.����|s�9��I�)�"J j��J�L��]|R�pUz��ʨ�s��y-��W��	�o�
����S-Hw���M�I,v1���o�yVJs;;�C���2�83���tqҮ�1������П�)�c�P��>� Me�+Ԙ�e��~ǫ�!J��@���Yz%@�u9Wd'�:*vp?v^l&��{� �N]��JH�Ș�q�=�eJP�E�����d!�ŧ�A<���8:d�L`��#�����C��'H�,u�+�v�� NX�;�Fӝӧ��IzJ'���.�GkԻ�����V��/�f%W�Y�y�B��3�� bm.�{��_&ʇ�$��l6ݩ5���mSf�����/o=z"�ӏK�M底���`�$�26�"C�!�M4ߛ�_�9XIep��!;r�x����@0��/(��^�
��^���x�Q	��px��;�� FM�0ă0clb2����B#롛j��-�ni�@�[�]n���̓A�w1LVA[d����
H)o7׌�m@֏�f��2���qN���Yz�s�q.���Ń;qbQ�H��"���Z�L���$G��-���YO/]]]�ܺ�>�-��M�m���=]�怰=&�Lk�^Mk{��3�\���?��Eet�"��KS۫�N0�5l�U�O/R���3����'J�Ս>F	�p�����[���F���u��ԋ������>�]�Ui�A�D�)�T��!ެ?I�=�"s�G�wwX��Z!V@99���׉<6��l?�\��v�NQ>��g�ə����xR����!҃f���Em3�F�GI=7+��,��[��
G��<W>S���XjITTJ���lPr�K�_5*� �]0�S��]���pS��?H���ś_9!��ѷ�<`���C��>%�/�R�(�jQ��%��鸗b�1)�ksu�V�h��a��W�[��3�e����2���_�u�О���8Su�<�� ��J��Q��Ds�C� �)�>E0(��p~���ƀ��86faT�R��j���KZ"%�8}�h��z��Fܦc��?���-�?�A�ӿ�O=�����1뽲�����Bt�-�6�\Wn9R��6��yRQ[U�v���O>��r�mOnv��$s�D���Z�5��M�ߕｑok�����ʻ�+41��'�:��pH?6��Fm_x@XGu�C-�ȷEX�s�X�&��hރa׹��B��Զ�L�6T���r�v��}��J%�}�#�W�KX�q=�81��;���������Μ^W��敉�	gW������}$����zU�!�m�I��s'�7���Nۻ#Uͣ���ZTkùB���^��"Mҧ�Fj4�ݻq�|���~�<�hu���E'e!�j�ez���-��N�����|[�bڸ�K����4Ú��� %7~:7�Gb&�"�5`|�ӑ3G*E�3�}���d]/Q�f�8X-�6�;.�>��(�"��m������u{��w�]&~
�=�y���BK�VX�TK?�R�A�N����>��7�9�t0��ΊH!�<|ΐ�F�dl�����7[O#j�.i����8�Q�\�(��6�h���8�l��va�c�SL
=�lW�(���Hp�9�U'��W_�EJ�)��O"3Ty�E��65��^o�6�v��#�xU��7��.�0`���s��S�]���e[
��n5�8GWU�����f�1�+]H�J<�lc}.b�P+�&�p,E����z���(wX.�F4�%��3{H�3w'�|���;�AM�ZN���#���O��~0�;��~gl����lF>^_��Vz�<(�~t���\d���ƴ?�����e6Y�-��ǝr�iў���~}a���q���sI}}7
En|��Վ�b$�(k������c����(Bv����hw%���)~��͎�y�\ǽ��Δwi����"4����*s��L;�����[�����P��VF�x�Y�O�xCy�lk��3n#�q3Y��E���BB%�cmo��Q?�J�]a�{�"���D��-[���#�b��OX��2>t�DFF�]&����f�]]�K~� �����Y-�
+�/��]�_�h��LU���׷��gd�@�tT*>{�y(�̱=�@�K�OL��F���<����X)A��4�g�&���u,���2<�s��ּ�@�,]�d6ߩ�oYQ�
�Ξ���-�lF��3\��uM�y��������qJ�*t�oe!fҲ��hV]S_�����[��<���r���9۲��+��4����q���A�ߗ螽�+�>���a�+�(��YA'eڟ��O�uP	4������h[,x0�b|k�jf^�H�i{�,����4*F��x՚���MQ<
psp/5��p{��Z�4�-��[������K�K����z�?�6�C}_�Q�MZV̼�T����hzp������^=衟��WZ$=��8�ї��~�6����c�Uv��jS����[��"=��F�;�L�GbQ�7�)�"�o����<H��f8�Y�qd��:�q�,b��N���؍C���~����06�4�Q���Y�p�*�O���ُF��,o���=�֜�-)+��ܘF�#�g����o��q�J��m(-����*��8a���z+`�2P�o��>�t��կ@�Q�m��:��īc�m��*�2�TEC݃�P����f�_�-pӰ/���s���
��@�6�hێ>q\޵�7�� ê+��U)u
�U:2d���l��~V!MP�����Rf��8���z͡h]�ȶa�����l�h���<@�U0�I�4GY�ɻ���c�X\�PF&��.*��ޞ�E<�Vg�2g��]�U�ֵ�կŴ�/j&�b��[��51�ji�1O
T���P���OW�b��У	�Hz��j�{�|� 7�k^�>EU�̐H=���Ȣ������� ��W��i1b�W,M��8Q��u��+!���G�����һ��������ǰES�fffA�ޘOeXf�����<�Ʊ�?�)�&|����ݫ>�w�G�5|�ZhrQGe�7�'/��Z-�%��.Nz 1��p��:��`�,�X�P�0�CE��Ye1c�5�9�GeFsu�JG���'��Q/���R�Ͻx�D�%hGB<�\���78�*{��4<��犵]�@(!u�|2�ם�D��0����X_�.[�ښ�W	�5�/> �8�uTZ�r����Sb�KR�Lż�I���6�*�d�6���Ɯwruk��1EX�o�W�P�?��q�ͤ��d�۪�hs��.0|����R�+~�%N�K\�ZQDGޙP��fr�9R×i����6�
(�����c��Xl�Pc���_��������������g�yk.�hM_Bq0�0�����D�"�y]E�OZ�5Q��q��u�:�WW�e\�B0C
p��3�6�]YUu�..��^��|(�㛂�Ei��~�W2[���ǫ�s�/1������ i��8�[��yE���+B{A�"�`Ý����91��9��_B&R�y�0:�Q:�����p0��5�K_!��ЀPfYu@S�,���f@+s9h�{畁氯�F�0�7��_�YϩO��2��.r�.h��_���ȕ�W.���ᝯa]���x�.ڂ=�|V�����`�4O��h4�sXL(�C)����L�u�[���J|@��M��fO���$p���hz3U?�h1�v������]��e%��mP�8f�t��\��zk���V�[�k.��K�^��zn�>��W��Sz���̈́�e�*��*N(,:n(�g&�&Fwo+��q�4(�������%1�i�G.�)��䡰"_%a�0�_��]d:�)�`�LTV�+����*���Ԑ�e�^h��T	���	���D�'���b��i��HY��������=W,��W|�_��@����|5��JG�8O�����B��ԩ��������Y=�0��<�������݃�F��������7��h�j����SH2����� \GG�]5#��3�j�7��M��&�Q���;)��I��Q����l}b�Qq1��8Ƌ����ΙXX,,��V�N-�r��A�����(�jc�J�<�T�p�,�.��ԫ�o����T��6����KCb�����PH3��&�i�ّ���b���2u�Q������:SD�M]C� 5�5�=��ޗk�Y���`��Il�iR��۞_��)d�9a;��G�v��<m/w|bG�E^���~<�1lk�v)���S̸����S3�TU��f��{�gp$�j4�C��-X�A�Z8���O���]W�)�<��ܪa0I�M�H)?�i�wj��nc$���� �ͨ��ǚ�$��.�bO?/xs�b5�G�k���ݹ�Z�I2>>d�����LE�w@x?����A��j�	0q��
��ىھ�Ăvt�= Шy��Ul8�Q5 �22�R��J�e�A��dC�}�j�I���v�i��r�=̙�	[��Y�Xhv��q"���l*t6=���%�^e�L{:�kfm}UIw�[s��b���+��8N�g�xَ�|~^��m�85
B�����w�H��YV�0��-y��ʱ�;4��H>M~'ͩ���8C#cɠGc��k,0�2�8������cT� *�__���]����h#�h&E�G��`�ax}�ʩ.v�۰8ݟ>g���T��&tp����suq�����1L�ܾʓ�#�ō����'�w���幛�����^���i��V}�8�u�@L�P`��:����y�;��0�kU�C�f�oq>�&#�*u`ؒ���!	�Ӹ�6J������^���c+���{h�7[�O<p
\56JS3a|�}f����&gd��J��|�����j2=�;�����:��1d�5��Qv��g*g�����*�e��m�E�Ã�_���iV9�O�7y�͘�h��w���?�|p��1�O�S����5����,�!7���%��v��߫/\��u��G�d��}t�:��׶o�庎�QΓY���4�X��#%졘NXY-�M7!ZT[(p(�r`��I����?Pd��zP!�5~�y:=����Y12����e�G�#"��"�|���z�*� � I��_�s�}S���^ ��;�.�ه�� �Hm�zη0��U�o=�o%ʥ�J��D�����9ق&f�~u"Y��Z5�vq�_��y��|_�}�/��nA=�~�q
C�8�6&���b��ň�/���wק�<��~@��'�R�:z�EZ��=~ؚ>�0��㺖�8��l�j1Mx{J�0'�tp�>w/g>0R�8efD
���/�1�ϖѿ\nc�̭J�}��VBq���Ǩm	z�K��Y,<�މm�.�c[��F|K_Yx^�ݜ&|+'�Û0���^	''�]:�Q9����E�}� �܆;ی��?�愞���[��G�X��VSlǄ�����Y���,�9!=�&���浉)9�Zb&r����F�QD]�����ꞻ�c�[�d ���� j��\?빊�O��&��=�O#A脈����PEwW�5m�۲NSa����mxz�0�E��E�R)��e�G�r��h�~� '��G��m���<BePO�fs��u���0��lı����1rh��c�ٳH��s��ꨨx���Ƶ9Ѷ��M������DL���뒪�L�X�82 G��_�����û��.����^(�0��N��#�n��x޸����,��l1&���x��
O��0��r]��o�����#ɢj�݅�q�7s+�DǍ�j�}S�B�\Ɩ��,�>Ω���]�y��-TO�wCڻ�NN��G~N�R+�*���O	��f��`I%L�#E�&E��S�tF��/���)�H��z�C5H�����y�e��`�%��<���T�֢)P�U�P<6�ْ�S�df���v�kO3�kr��[�ƙ@$�ƶ4�Ym 
޹�3v#�]��#eWM�"܉�6�Їh�2GE��p�q�O8��D�R)�v_�s�8�2���㽹/�8��!�W�U.�Ėl�ls�Ӱ}�ǚ��-�ʺ��zV��XF�й�N�d�M!�j��P�L."�����5���j�'>%%������ϼ}�����5�`PG�3h��0��$3{֖��/8�YT)��+�����޻�"Q�:7.0�&�F����V������::���>�:eꃬ�z�*`~ETF$��v��ۤ&hI]K`d7�U�6��fFQ'�>R��eu���'����=�8%0ҁ���K�A�%���\�9g�p�u�˾��|�`�1VTu�Eh�Q,0��?R&���F1���]�A��/�kU.�0P�Rf\��Z�8	tqy{2%�>�U���Z���㵳��Ɍ��)S��*�j��̀jS�7&:O�s��uˈ�C�?<ҾX�4'���a$[��)Ζ"��I�Mـ(���Ȳ�����-�D#��^��Y�ʁ��m�79����M
+��V2$�$����zWkN�r|��D�mF���� �%~�'�#�K7���&��UyB��w��]q�	j�!���ߙ���)��ޑ���t��ww�lcmz�iRS��p�F50q@�B��TK�j�;Ο��f�����\ʝ�ʔ�u�*��ם�s$�}{��^Z���ĺ�#�WȢ�7����w����>�o��W�J�C乘�e�L��}��<V㑫nwSb��I]TC�i��� z��>��j/��@�ƒ��І	Ծ�5��A1d�l͟S�F=�w�J��d��؂�;��N����dG�Έ�E�;}�3\�]�S��JQՌ&�B��[�o ��Br(ykDs-�FyΆ����U;smP��N����>��d�����ڑb*�J��66<��;>)�������K���%s4n�'I;�9aFX��Y.ω\ �t�>��(A%t7������ተ1'~��8=(NpH�oǈ_"��1����e���&6���{^���3�-�[��Pq��
+7�]n�Ś��|b��d/�Y�綷��ͥ-�T���E΁(�N�����Nڢ�y�9��J��i��i[;,|��E���#K�G8�f����K�����$���Af��J�r01�RX��ƱJ��⤧�
,�l�
�	���vp>��'%��s��I1r]_��޶%�ƸVȣ���^J�z����)��io�䂢����ڍ�z������]į*U�K���{��9����(��y����έJ$d�
:� �dR�P�u�87�vT�O�j�#��HS{1��zi�s���K�+�y%m	��f��W�x�ZƯ-��N̓��g��Ȕ�b�ùl��]2��;o��
���ܸM����i��0 ���*2�j�)W�g����Ю�\_w��߭����@�u�o.��|G�ܥtR��8P8�t��C?�����&�6+�a_��51;ݘ�����o���]�ͦz��eQ5ښ�~{"Ӂ���[�Gla)�I���sB߃ţ�͋=Aw �NuA�,��⨡����/��*A����N�o����f��l��{��$���66��)(���K��_���h���L�x���~'��`i�H�,��O���e�H�)���b*��{u~�
�d/h����G��ͯ�"�]_����է,1W{M"���o�M~�*J��ܸ�H9L��.��(^<)w��8%�_�[����!���x��n\j�2���l�Nh�
bϘ�Y���������1�����q��D�o�M����#�^��O�"bFZ��� 854��nLLU�'���V�d�o� ��Hq����*�z�r5(̢Pq��-�C(�i�ʌS��X���i�v�嚜KOp_�WE�e�P�M�	o�t�.�zĻ
2G��,�S�I?q��F�V�_�a��;{S�U�����E�E�\��R�+g'7ˍ�|KV��g�G�}��eu��Jy%H�E�~\�㚥�,�6 �����K{�]&0�1����UC���k�'�ڟ�e��b�+���Jgggw��ɮ�e	R�S؂K,�	��S�}�ّר��s�l'˗�`]�~����q-��>ị�G$`�FZ|��?˰>yD���s��Ds�!GC�A��k^K(�\�}����T�o5��\��lf�g}�|[W�עѸ`��W{p;�@�/^���/�<��|�|�1}�΢�b�<&O J:�1�v�+��c%�"T�>j���Od���r*�%M<{a�I�:��&mn��-�E�7��)��� ¯=Eh�@򉪝�:	c��
���Om�}U���7:D��OI�i����]`C]���Z<ҠX�֟���K8J�����Ô �YWJ�8S{݄�.I��ϥ,�d?�	.)Cבo�@�d�����#�[(��[����S���v�Es��4;DƐ�}u�Kp�w+�\��<� ��xR����B�4���m{:=�1D�{Um�Q��q��<�2��8N��n뱦��"%��de�B�������������!2��%Iz�}
���ޓ9r����1J����`6���7'��$�J�%v0"��}6����.�]En)ڼkn:2�?��&��Z�O���wR�����S8��`0 �X����G�����Ղ����=r�7�e����~������P��l�3�Ɋ:XsY��3"�h�1E{�D1�p��zY��T���Ӹ��ge�
�Izdg�Y<����UUUk�;6�ay�Ŗ��S����Y&�0���u�+�%����Gs�t�jS��O�D����<,&�߾k.�W,��U$o$�7y��ز^]ת�(������uz��״ݬA��ra���6�K�rF�D�E�K�-"�����N{ؽcDx���g�!��{[|�3y��A���O����aǷ�ǻ�P��Õ���ӧ�-��St@�� �Jasj`�}[��1�f��:�Gp02P�f��j�.�ynɜvA3��|����TzqW�&�l�w��
���O���7|Ezg(�nF=�fj�F�F�E������ۖ���?z#��G޹r�m]�##�[�LQd`�dgbc�W�{�����Ƃmq�?(k��
�!�^��z�>[X�^����?rzi�,��"���M ��^JF�sVЫv4�AZ����{������,����BDL�X��?zfAd�\dhв�����m���2��7�Q���*�S=KG�)�F!�=^U�����2����:��#��������Iӹq�bdd$�d�q1��:;�����?-��gux���V���1ϳSH��t��U�a�f��t;&z�Ya�~C�B����`�hˊ''�S�8i�i~5����9��vm!��&���<rB.���fV��zE����Ӿd�E	�l�*DmP�
#=:]�|����9�Ұc�v)���p��Մ�:��4*��hc�r6�4c����������L9�':VE�������kTB���+�V�U���U��R�^' A]����dE�@�.L-�+Pъ}@��������v�A]�������� ɀ��V|������p��9�y0A�0p�3<��G���}�Y�z�b����3��0����kX+� ��[����4olV5�n�Y^fV���Қ�I�F��
��	�{B� nt���=�8k��؂�/!���[-��N�3��;�wo�Sz���N�[)8�΃��y�\�n��U�Y�Jv��s����8�io�*���ϓ^
plt|�n����n�2u�c+�yk�{J�	D%��>
�vvq��cv��"��}���/&�N�c�=�Q��v�į��-6s$���7刲�m��iu0�=�yl ���z���y6����c�?�{{餵�{��E���-X����H���{gt���_�xU�d�^�0,��[��׹˛��6V�������x�H��:w��Rv�@i�����^"����p%�?I����q�q��:���d�]2Q&��_�41]e�H�����!���I��a�l��r7��Un�>̽���#����p �.O>ZnM��ݑܜhz8,/��y��it��^�ʛ�h.S\�	�,W��n�*����w2'�)�� w{�l^���|QJ�Z����Tr7C�ICE���W���)$m��J�OX1�,})������YAQc�X���"��ڊR�*�p�S������>A�ytzz��m�?/��m`y����v��~�~b���֫6-4w��d�V�^22B����y�8�"{jmL��=��U���������]8~��q��y�E]�/	5gv�!��h<
��@���2��gW0L���0��]��jV��j�5�ф�mokLi�ޘ�*>���2Lj�����[i���WN����X��6�j�u�:K�������ܦ�P+��℩Ac���M�7�ӏs��H�ѴaOBG-���D��LW�O�a��i�Oi����dY���%ִd�v�?�' ���X�8��>*�j���V������r�_�["ε����J.� �=Ip��X�=�iT�6}����s`Or#ir���9^�f`��*R'$IIU@��i.�:��)?aJk����H�䒁r�6gK��./���ݸ�9��N��N6��%���� �Z������8̡4m(iG-���.L�/I	��QA��Z��S�ϯ��J1�>�{���bd�{hf��V�rOjW���)Oٷ�bnK��i�T	��R$�9�/�:��?^O��ǧ6�͍)	�)�^ޣ?�F�x(��79K��x���5��5q~TzloE���틜!��K+��9<��s�M���@z5q��	����	ǎ�G�$��O*r��&�7���7H�P䈠5ǎΏw^iwt\���Z{���n<�X����<��ڡ.�/.����J�I�6�>1'�y��j�c�Swj��e�9?B��f�c= ��Aa��ǜQ9�7��]�v���,�4�b�sΟ]�F�r\&�Alu��]oFR���-�K����)��̕dv�*D�K�`h�p���|�ؼ�깡�,�t� 3�M�?ٱIA8��3�e�g��W���_�yk��q=��i��X��-nؾ�s�v�E`�x�Ύ��'�A		�9��^ �R'�m��Q�\���oS�S��2��U�8��:�����c�~mF@d�q�$e��ī�I�¤Ē�s�_�M#o˶3�P�����b#iveQ�N3�A��Ԋ��|�ꃪ���UY��1�ӏ�}*����L-9�����N"�Q��~�_*��A����	�Fs��xFD,Kz�C	���Y:�6����hg�K��G+��/�-w��ٹ3]�_�l� �p��1���|��H��+,�]�u*����G�����Q�۷>�kn�I����O;�cb$2xYaA�\x�k�L8�����r^Ih�t�n��p�2!Spߏ#�����wH����t��b��cL,�{κ#��[A�UQ�@+kdi�N}zϘ��e�C�^�=�Lh����H�j�"s�_����j��U{����;,���w1�9|��q�z���}���³t��=�VR�����ӄ$l�j�s]��T�xZ�pm8���ۇ�#j%��w"��mx�5��8!�"Y�#�[�R�<��[���w��z����Nz�/+�"7�A�Έ���I˝(�˹�5|Ď�S�skG�.��R�ãF�-��wꦃ��/���ŧj��2����(���H���W��5�M��%��Lk�����w7���{��Z�>5[�ʵ������]:( �$��x��TF!�e ,���l	3Z_�b�k�-�;j�{�Fj +Kd�G�Mv)�.ҭ5���b�V����v:\~���.�{H6���e��Cc���W����ok���@c]� 8�v��
������Udbأa�J�F��b�2Ҝ��%ډ(�+s��sd/�:��gK�y����Y��O��*	����f&��̢Ք��R�S'
�8=�����������OS �%��w��p�nu T�G�]�O;�u�(V*|�HE`}���`2���)�AF��I{ū/���9�
+%tT܃T8��\��\�o�b���:��*fWr��9a�Chl�����?
�@`�vv��<}@S�Ѻ�d��.����NRq�֕w]j�Xz��ǒ�c����7�@r*�W�-z���$��B�N~�Ӷ0gU6t/�U*�]��^�9W�f��`�7���w�����gS�A۝z'��G��(�ט~2���Ӣ瀎��.�;�_�Nɵ^t8v�A�3��T
��B�s�cWK����zqK���a!�v�D��v˟�*���S���ؤedϟ���'�ױ����U��<5�n$�ۈٰ3�+��c[�߇:VH�O�`�Pq&4/�v?��ZvˮZ�#G^��٭0������߄�d
��2�zU����hׇ:8��\���ܝc@#t5���q��γ��K������̓��p�/��'�?b�;��w��
+�]Blg�<3"��)N�PY��v�$��J�}S^t��f�����P���;!HA�v�v�pBB#ZW�֗��w?�~w[����f_3��,9[{���hqN]�>���dG!�VA�}ϫGe�v5eJ��1o��쾻�d��G�>��4�`;"��A`�ې����e�.�w�,��[�<ˍ����7��>ݯxgYۛ!f�n�&�X�ĵ�� �O)<�n�G�����^��H�7~B)�*w�~O�̍�I���GJ�N�:��}�=�Fɋ�Ds9��y����G1�CJ�r���oNLǫ^��^���6�*c�כ��޾v4�9�~�x`��*�XG�l +��<S2-������`�O:��e�d�%>P,!$�23L�~���i���C��r�rjS�fL󶼧,�1 �"h�%��s����zU2��K���6��1gã�l	1X��JI�`�۷��H>�+8e��E������fi�v-(�#������t�q��&8ͪ��=oBW�^�B�_4��o�l&e�4��c2�"lmD�"�����d6�;7q�ˬ���D鴚i>���.����d��;�
�kg<�>T���q������eJ@a2��Tn�&qrY�U�=9R{�Q�����%�Uh��I-�k{ٛK�t��=]ܒ�&��g*��n�\��ٷ��M���%7�|]�j����!�%�v�t����A������tq�l����e���E!�Γ�<�+��JS��4�Y��u=.>^&xi�Ox�j���G;o�ta>"��g����ژ��F�,��p����k���2�Z6�0�{M�S8�ѱ1;;;��WW�B����[k?�����zz��d�8���n�y�Z#�}V'��ζa��_I���1��^�~O��`g��ڞ)�UV6�b�\pF�
�$ ���
Q�T�5d��h�t\m���ߓ���i|]� n<���H��K������߮R$0�!S{�#��#L��-��Ly^�Nm^�O�v_�i�;�h:�<>yo�̌��b�#�.��[��K��^7֍����Ň�[4��A7�U�r�ͱvb��D�%�#��T�|��E,��\�<���zӤe�2����YrI���O���U
(�.k� kE�x���8�K5�OP�u-�,�d�"�/r��GO���[�j�w��Fm��*M$���"�L�#U7/�docjn7c�P[����yhu����Jx%��s��H�����4�v���@6�VL�E��+nw�;<4&���^�E��J�=C�m�Q?�>6:jm畐���o�l3��Ƞ��/�m/U��n��W��o�
�������Ue%����>=�+7�'�Fm���v���y�?��q�v�����#5�Ƀ�q�
AU�O�~���6���ކ�Aa��c[[s���
�xA�&���΢�$:�����"�N{09'0LcsL6�;@�o��_�k_D�W����j%
b��:�2�Ӹ�T��^���_�}�����Ӷ_��N�i3�����/�l8a���u#���M�����\�o!�ixfy�B=CZd�lj� "�FUA�_�ͱ/e KL����k\�0�}� m1dug��C�}�^Z�d�9�NWS<(��]���w�VaR~0�F7,�>b�l��/��F,�3ȷ�=���OK�0q��.�'���-�\���NhO������;��FoN����X�.ˍֿB%��ܸp�4�)[��PK   �I�U�Ra�  }     jsons/user_defined.json��[k�0��ʢg[X7[�[��҇�����R�W�JvK��5��.���GIg�9�9;4n�hJ6�2v�5�@O6&<<T��nҤ�4�����p�>�ګ�M4];�M�[Р ~[��
�(���p�JRYr�M�U�J˵�B+mT�l�X��d��/m�ƃ�w[7���ǃ�@����_��!?=.]�v�=��?D��rP�?݆���1km��,&��L`�_��1:��в $�}^�n�� \6XpF2¥��j���[m�����4��B��>}`�^��6��"�yW16��u�yc]�g�5��������c��T���Ɩ@楔mSr�L+���_����l�3��O�A9V������NJ�
RK\7������m|۟�"�:r��?9�q�<?*�Ǽ_�_ PK
   �I�U�G^!  �]                  cirkitFile.jsonPK
   1�_U���R�$  �/  /             �!  images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   �H�U�T�S� a� /             �F  images/dd298255-0ede-4bb4-88a7-459da88d83a5.pngPK
   �I�U�Ra�  }               ( jsons/user_defined.jsonPK      <  �   