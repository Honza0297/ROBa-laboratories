PK   �PrU!/�#  y    cirkitFile.json�_��ʑſJ� �44��f���Mv/6�ds�dl��D�Zع#�Fs���w�.rl�DqF=u��1p�Xd�T,Ydw��ž���mֻ}����ﶻ�ŵ�W�w���}���Z���6�]��}�nq�A��~{�g�}�v�]�iօ�U��٦]�k��u!Y^���kW�ºq�[\�~{�r1+�F�V��f��k
3�U�5��`UpMif�*�&��
���V��f��k�f�B�Q�������}���\�y��i���o��naLx��H���+��_׻���n��C����*]��]2_�E���e斮�æ���n�`��=k�=m�%"�=q�%"�=u�%"�=y�%"�=}�%"�=��%"�=��%�=�5��r�m��1�����s�Y"R n��y8��a�D���a�D�(MWUo�l{��9�,)�9�,)�9�,)�9�,kd��D���]�D���]�D� <����w���~�k�pZ�)칳��N�D���N�D���N��k�=w�%"�=w�%"�=w�%"�=w�%"࡯=wz{�4KD
{�4KD
{�4KD
{�4KD
{�4K����N�D���N�D���N�D���N�D���N�D� �2���Ҟ;��;��;��;��	��i����i����9�H�}�.����Q��D���~�LL�N� ��H�;(�`�\�c}��ҽ��S@��L�������P:�����;���N�t����;(�`��M�w�;(�`�\Sa}Wa}�,�kj��j��t��s��%�wP:��M�V>��{�PO��\�`�t$)��A6��\���h	 `>��\���E
�O�|:v�?p���0��z�\�`�̧���,X>��Hs���E�O�|:F�?p��0����\�`��w<� �l{ro)�r[9$��'g~��]��%�/X>��������O�|:q�?p���0�N��\�`�̧�����/X>��T%�����O�|:�
�?p���0�N�\�`�̧����/X>��<���,���t2!����'`>�	�����	�O'p������?
p�Q��,���t�,����'`>�������	�O'*���?�|��)�`���,���tr8����'`>�֎���X>��|�����O�|�J �?p���0�6A �\`�̧���C�3AO4�\xp���0��� �\`�̧�>���X>�i������O�|�`�?p���0�������X>�iS�����O�|ڎ�?p���0�6�\`�̧-����X>�i�&���s�ѓ���G	�?Jp���0�6��\`�̧�����X>�i�2�����O�|�^� �?�|���p`���,���������'��%v;�k�h~ڐ0����`�B!6s�{j	�'VTK$9�}�h~ڴ4����h��i��D�����h�`cOVpK�7�dմT{c�MV*K�7F�du�T{c�MV�J���Pc�M֜J�7��d��T{c�M�GJ�7��dM��k�1�&� ��[����+���/Z��������������?Y�&�����`R��?Y�%��zk̾�Kқ��<�e,(�P�,�jo������P�,��jo��2���P�,��jo���r�����,q�jo��ɲ�������"�����1�*c�U�����W�2�_e}�d����1�jc�������W�6�_=�(�2��ޕ���fm�^f�ڻ媗.��'�D_d>�}�\�m.�l��&�K��]I���Z���o��|���N:�U�u�6�>y�\e�_�֕a���z
������"���� �y���>������.O��l\YO���̇��q�o�f�����,%u$Z��W/����!	9�H�ib�@BN�/a�@BN�3a�@BN_]a�@BN߆a�@BN_�a�@BN��a�@Bâ	Q�� )��qi��eȷ��v��`�[`���ת &X�X�F)���/�	����QJnxMb�eq��q����yP������sXG)��?�	��sXG)�ax�	���!�n6 &X�ay�䆡 &X�ay��!$ &X/`QPJn�b�����QJn�b�����QJn�b�����QJndb�����QJnb��q��(%7�1���q�����p��q�ay���8J��@L�<�ay��Q{ &X��<�Rr��BЫX/ay��Q� &X/ay��њ &��M��MX/ay�䆑� &X/ay��� &X�<�Rr��_,�X�S2�>��ڤ:�G��V�*��5��	�@�2X��z47��������{��*gY�8�W�+�U(��������V���� �_O��a<�`
k�G����;�V����_\�W�PX]s���
�+�U(��9��W���*VL)��Sq��E�"}K*�HU����]�)��Q��V8�:֜�[N�E�������S�Qh�C�c�9��TaZ����o9��V8�:��[N5F���)���S�Qh�C�sc8��TeZ���΋�s����.;Kp�.�9u�V8�:��[N]F������S�Qh�C�s�8���eZ���\>�o9u�V8�:'��[N]F��έ���S�Qh�C�sD9���eZ���\W�o9u�V8�:g�30��B+Z�{��-�.��
�V�Ps|˩�(�¡չ�ߒF+��+r겂S����B+Z����-�.��
�V{p|˩�(�¡�^	�r�2
�ph��Ƿ���B+Z�]��-�.��
�V{pP|�9u�V8��K��[N]F���D���S�Qh�C��]8���eZ��j��oI3�HS�8u���e�S�Qh�C�=�8���eZ��j�#�o9u�V8��É�[N]F�������S�Qh�C�=�(�-9u�V8����[N]F���8���S�Qh�C���8���eZ��j�9�o9u�V8��;��[R�R�N]Vr겒S�Qh�C��9���eZ��jOF�o9u�V8��[��[N]F���Ȥ�6p�2
�ph��'Ƿ���B+Z�Y��-�.���e��K��t�MT��M��2�M6Qe��w���y{�)Qe�Wv��Lw�D��~ԩK�CTfz>�F(x1�;��k�&~�VM��D����2��[&4U�s�q�ʀr0&��V�L��D��Z��2�(�[q1U�s��^u1Q<�z`��V��z�EMSe0Q<.^7]�<U�sKĥ�`�xn!�TL�-w�*�#���u�Rer�i�TL�-��*���e�Re0Q<��S�&��TJ��D���E�2�(�[(U�s���`�xn��TLL��	LLLLW�(�0Q\a���Dq���
��1&�+LW�(�1Q\c���Dq������Q��*��Y�]�y	m�V�e���[�z�B�|�y�E*�'�\�m.�l��&�K��]I���Z���y��T�e�;��W]֭�h[�>[�r�u~ZW�����=�E*�g��"�g��/��2�Y_����o�:/�{�ʷ�qe]<T��� �v�ݡ=��_d�+T�����oo�Ur�o����O"��bBr��<H��!D !7�g������Br��OH��R!D !7��ŤH\�ƥmX�X�F)���3�	����QJn|1�a��o�%p��_�c�`9\`I����&X�ay���a&��7���sXG)�q4�	��sXG)�q�	�	��sXG)�q�	��sXG)�ql������QJn5�a�=I�=J�����QJn�a�����QJn��a�����QJnP�a��q��(%7u�0���q���a�p��q�ay���8Jɍc1L�<�ay���Q�&X��<�Rr��L̫X/ay��Ƒ�&X/ay���1�&��M��MX/ay��ơ�&X/ay���A�&X�<�Rr�pg,�X�SJ��?�,�V'�T��*V�L�J�U�~e�
��5��hU�_�Bauͤ�Z�W�PXc�E����V���� �_'�� `�
�5ޣP�:i�� �U(���t�C���`
�k&�Ъ@�2X���I7?�*ЯV���`Na���(�¡ձ�ߒ�.R�ũ��Sx	���
�Vǚs|˩�(�¡�1��r*0
�phu�?Ƿ�*�B+Z����-���
�V�bp|˩�(�¡�9%�r*2
�phunǷ���B+Z���y����(�¡չJ�r�2
�phu�Ƿ�7b�Wb��,��e9�.��
�V��q|˩�(�¡չ|�r�2
�phuN"Ƿ���B+Z�[��-�.��
�V�r|˩�(�¡չ��r�2
�phu�.g`�.��
�V�s|˩�(�¡�9��r�2
�phu.8Ƿ�ъ�ኜ����e�.��
�V��s|˩�(�¡��r�2
�ph�WǷ���B+Z����-�.��
�V{Wp|˩�(�¡��zN]F������S�Qh�C�=Q8���eZ��jo�o9u�V8�ڣ��[�L2�T2N]�9u���eZ��j� �o9u�V8�����[N]F���p���S�Qh�C���8���eZ��jO-�oKN]F������S�Qh�C�=�8���eZ��j�6�o9u�V8��s��[N]F�����������S�������eZ��j/C�o9u�V8�ړ��[N]F�������S�Qh�C�=2)����B+Z����-�.��
�V{�r|˩�(�rm�:�3�nUfz�&��t�MT��㝨2�y;Qe�Wv��Lw�D��~ԉ*3�Ufz>�F(x1�;��k�&~�VM��D����2��[&4U�s�q�ʀr0&��V�L��D��Z��2�(�[q1U�s��^u1Q<�z`��V�s���`�xn�TL�-�*��⹅�Re0Q<��Y���s뀥�`�xn��TLϭi�Zu`�xn�TLϭϔ**�0Q<�pQ�&��J��D��"<�2�(�[�&U���|����&�+LW�(�0Q\a���Dqz̆��
�&�kLט(�1Q\c���Dq�l���ʸ{�{Wf^B���z��k^�P.���ʳ��-�y��&�����҇�nW��.���*��y��"�gY�N:�U�u�6�־�V�\e�_�֕a��/x�q�
����H���� �y���>������.�^��l\Y���"��~�x�﯇f����m��⺸Z����w���v�w�����~��~���T�p�2�y�x{�ڤ�l��ק���|��?B1����	��g'!Q`�K_(M�����y
�z:���s*Grc��O��p��9]���G�o�~�&���v?ǋR{۝�>���q���Ͽ���_�&��+�½�@�G}�w��ۺ�;=p���1���eg��{���\}Ճvz;��}4��f}���*��pc�8�K<	�+t�E8�/)´�_x���5w���/�?�{�ٌ��a��o����>�l,w�b�pÓR#�Y�O��f	7<�6R�%�0��Ha�p�L#�Y�3�f	7�T0R�%�0��Ha�p�L	#�Y3-��ӓ%�X�l
H��ԏ��F,@~@��k�q.���c�d�n�c� �Y$Z����X9 �V �֮��A'�0ޭ�mȶv7NQ�r �kH�v7N��r ��0��$l��ms@��k�qڗ��ms@��k�q♕�m������Y9 � �W��'�Y9 � �W����Y9 �� �S��' Z9 �� �S���@Z9 ���]Í�0��|��Ԯ��i�V��V�W@>��|j�p�LV+ �z@>�k�q.���O= ��5�8���j �OK@>�k�q>���OK@>�k�qF����
�OK@>�k�qR���OK@>�k�qZ���O ��5�81��ȧ�O��z�G�ơ9���&\���� |G#|���ߋ�0��@?��&�;O�[l?�+S\�ϟ���Ӄ�#�O�|��o�T���b���>���,�`��X>�Ż��&K/�O�|���n�Ӄ��'`>�LV0��A���0�k&��� ���	�o:����6}��5�@��Mt��Q�E
�J9�p��]��	u�,ڇ��L(hB��!�@
�P�'�}�.R���&ԡ�h�0��	uX8ڇ�bL(hBҎ�!�`
�P��}�.Z���&<��y�=���������e
l� �l��e�PЄ:��Ct�&4�N?A�]��	M�Sg�>D�-`BA���e�PЄ:G	�Ct�&4�ίB�]��	M�s��>D�-`BA�6��e�PЄ:'=\�zL(hB�O��!�N
�P�B�}��S���&�y�h��~���]��:L(hB�?��!�N
�P���}��S���&�y�h��0��	u�5ڇ�:L(hB�/��!�N
�P纃}��u
�PЄ:O�Ct�&4��@�]��	M���>D�)`BAjo���T�U�u�G�)]��	M�=5�>D�)`BAj?��u
�PЄ���Ct�&4��aA�]��	M�=d�>,�u
�PЄ���Ct�&4���A�]��	M�}��>D�)`BAj�$��u
�PЄ��	�C��z��zt�R��]��	M�}��>D�)`BAj�0��u
�PЄ���Ct�&4��f�0��0��	��ڇ�:L(hB퉇�!�N�s���;N�#&�O�&�O��.Ni��~�O�/L���EM���3M���!M���M����L's<Zr��[��5$�+��
X�p�fY��5����
X#q�W��95Z#q�fU��5��B�
X#q�S��5�K�^⬑8]l(U�|��Fbq�:�,z���yj%�T=k�NW�I���t-�Tk�NW_I0�NZ3�t��T�3�)=k`N��H��tQ�Tk`N��H��t�Tk`N�jH�F�tq�Tk$N�#H�F�t�Tk$k$s�m��`��`��`�����5+k$V�H���XY#�2?�Fbe�����5kk$��H���X[#�~"CQVe�1˽+3/���j���w�U/](�O=����c��˼�e�m|�d~�CV�+�||[KB�<���?��y'���˺u�j�g+_��ίB�ʰ^�O>�����O��E�OD`_	eȳ�^�Ѿ�du^v1���oe�ʺx��_d?���W�/vۮ9�(x�����$�ׯZ�k��O�E�����:����_�[�>Î��订���,�������Z�j��j��E��Z�j��E��ZjQ�E1�E��ZjQ�E��Zx��j����@-�Zx��j��«E��Z�jQ�E9�h�(բT�R-J�j�"�EP��a�Z�jԢR�J-*��ԢR�J-���jQ�E��Z�jQ�E��Z�D�V������`F�K��#�K�~.��h}�M1b��@���Mܨ��Ϛ����գ��>���2{���Z�	.��NޏN�#�gt�z#�	O�$��VB�[֘y�����CsӮ�=�'������!�3hؔO7��&�n*6�M�a��n*6�z�lon�G��nv����.��}��A���}�*��~s.8��&�U$�9yٗY���l�/۪(�y�:ퟜ7ߵ7w}�����o�M��\�ܿף��}��F����C�>}�߽���m?�5���V�� ��;췷?��z����֭W��ۛ{�׿*�p廿�F�E�w�v�����Qwq�џ7����oﶫ���g�����[\"f<D?����'����)�ǻ="�w����$���o{��^g�«�/���WuQ�*�;��O�l���M(��}_d�2�l�i��Ȳ^����'ޖ�����%7gW��~�W;�,bdģ�ݯo��#�:���Uy���۫�W�z���A��̆j�"�Y�9�b�BN,�Ӗ�dC�iC��l(�,��E>g!��Ö�У�U���wm)>�3��������˓�?�I\5�!��(N,§��JaY���q�v�|���ϧ�?�:o����z���χ-�x�0���0{�0̇�P����LΜ��x99�>m(�̆j΢���݌E.sŜ�'A�iC��0�|HN��:��:Г�f~~���d��"-w��^��W3����������2��;�U�߿�f�/g��3��3�����l=I=��t�sGv�׹#;�˝'y8��ϫ�����~f�bf��ߝ����N?�f�/g��3��3�����Ⱦ�I�g{��p�mw��w�튼�W.�~[o3����>+����׾���~�v����4���˽f}�~�/��˫�w�u�U�t�^�*7Y/�X�z�m6���[�|�I��:/z�t�]g9�)�ܯ�G	���,�m}I؜�,^s��g~��iWe�^��������b���/�%��3߯�l�tE���*/W�XV�S�]���c���]���#>���D?������?��tY��?��7p���_��w�\��O�<� ����<j��?:&�N���%�l}o��<�7}�nSUe�Y-��Ӡ��Q�Eŝ��_�ҟ9���=����]����yQ�r�O�pUV�U)�:�J�xу���\�ŏ��B�Oev���p�v1
E�po�d8������/���N����g����t�P���zj�ۑ���i�����}����������w�l�Ûx�nv�7��7���A��fq�&�{������Oݰ��d|�o�3r�O��}����ew��,~~9g#����~��=|��b޼y��'s�|�~rܝ~z�Z�W/�_RM���M��puf�x������������=��/�8�֗����]m����gͲvg���n��8z4r�~!?��^���|����ef�o��a�qv75��A̓����n��nE]�d7wY�� |^�>A.)�W��f��t>9q��2�$.yQ\p�z�WhH����! �8��S�E!p�ۥ�|���!��E��M��/�l�b�,�~�ns��*���R]t����毛���~���~,�b����������޷7����C�ӝ���PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   �PrU�]7;8  n     jsons/user_defined.json�MO�0��
ʹ��6eko�]vBNhBM�K]R������qVƄ�Ip�1��'�?v�Z`��75jP,`�`M�8�#N�K/u�x����.�%��4U���؁4셀7�o�*`�H��R*!Ґ�j
�*�y�� �L2�K��Ǜ9��������bۍ�N���#>j���Z�s]V��73tmS�������H�N�������I�LF�8�^�GO�\=u�NC����\`C�8�b:	xe"���NW��R�ͦ���l�'��dq	]����^�?��ߢ�1�)dM��Î��*��9W��z��8{��PK
   �PrU!/�#  y                  cirkitFile.jsonPK
   1�_U���R�$  �/  /             �#  images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   �PrU�]7;8  n               �H  jsons/user_defined.jsonPK      �   PJ    