PK   t�>V����V  &�     cirkitFile.json՝Ks�8ǿ��j��7����0��I�l�b���c�ZE�R�dfS�3�ć�߲�>ı��h? 4LN���z�(�m���nw��&��*�P�էb���*�_m�v�K[�Hn>��i��}��ۏ��M����Y��K�&/S��.��ҦB.+�tN�,�ywu����%��0u��L��)e!�*[��T�M)R�s�ڬ�U�y���'@�s�c�9HJ,�� � ��V��
��	?�'A�$:e��I�?	�'A�$ȟ�� �O��)�?��� 
�O��)�?�@�ȟ���{$�h]�ƛ �DW��j]��At���N�g@����3 �π��?�gA�,ȟ�� �q��Y�?�gA�ȟ�s �ρ�9�?��@�ȟ�� �σ�y�?�������*lV���:�Yդyi�4+3YU�TV�g�gG�n&����L�u-�/�"�UY�K�"�*�A5��ҙ{f��=���9Jy~�E�Ϗ��-��s�����LՑ� 5k�f�����5�x�jvH�Pgy�й�(���4nd�#�Grq��h�����#��8�>���-��mfo���+���V$��bE�X1,V,��bųX�y�c���^�����W� ,x<�Ă�b�C�d��y(�<K�%Œ�b�C��X�P�x(V<+�P��b�C��X�P�x(V<+�5ź�8���=b��b��P�y(�<k�5Ś�b�C�ᙋņ�bô����Plx(6<�-Ŗ�b�C����Pl��'x(�<[�-Ŏ�b�C����P�x(v<;�c6�Ŏ�b�C����P�y(�<���f�����4�Vb3��w��=��͂�/u�CPF�x��&���S���T��֍M;3��Ivc3�ǩ��
3�rr����rP�/���љ\3'g��.���1Dt����s�w�]�&{7�C�k0ً[�,V��bŰX�,V��b%硎	^z���_���!X� ,x<�%Œi�X�P,y(�<K�%Œ�b�C��X�P��B	�Ŋ�b�C��X�P�x(�<k�5Ś)"�X�P�y(�<k�5ņ�b�C����Pl�6v<�ņ�b�C����Ply(�<[�-��Ŗ�b�C����P�x(v<;�Ŏ�b�t��C����P�y(�<{�=Ş�b���d/n�d?E'{q+'}�N��Vx|9�ot��r��d/n����ŭ��~����1��C��<G|��������^3��
���{���Ū�-��U�i�ֻ���(�j��,�mU���{���<��~�۴-V����-E��辶��gSV��t��V/�ʳ�߮�v���n�_����=1��4�)]���\�Zz�B�i��|YW�v��!O��sE���gWCWps�o��o��L���\��=B��:2�Z��qKb��u�k�/�	6��e��"]J���,�m�1�X@�y����@���0�j�T��U�J�)����M����0 �̛,�J��B}U�e�:����uT�o��]�E��:�h>_r�ɷ
̵J�TJ�J�F�x8��.�ԑ*Y���YfB@'�O�dne��$�
�c�$�jl����,��0�˱��8n��2k�L�|\Y��E�SWٲ�*���q��(W�!tlO����E�Q�\f�{+9�c��_|��6����in���g�~�k��trX�Ԍ<��4Ru����qP�����բ�TS��A��߿���K?����o�78a>���~��m�#���	���c����6-6��\�q�ϝ"�=BC���I� ��;o 6�	��:�6���ݯ���=@��q�4 ���'�u�?6^�``a�xb>x�D ��E�WI�����I����F�p���%�w<~����eߦ}`��!:����o`���7'��[��/�i�z����dt�}�.wz�e�.j��)���x�?]�Ͻ�p����K`�]tW�:�<��Ew�����X�u6��������ʷ�(�{�|_�H|��p��=&�!���7��э�[�����$ٽ�K�_l�y�.�#�����z]�y7��t̻��_g��"���XF�!��p�2�����q�1�x�˝��O����\H��zXm��K���i��K�V���0l�/A}�kP߀��l��s�;��Q�`Q J�@�(����d �P� 
�D��(�%Q�$J�D��(Q%J�DI�(�
%Q�$*x�FIT(�
%Q�$*�D���P5Jb�.�A��P05?�`jL���Q05
�F�4(��"J�AI4�V%Ѡ$�D��hP-J�EI�(�%Ѣ$ZxW��hQ-J�EIt(�%ѡ$:�D���PJ�CIt(�%ѣ$z�D���Q=J�?Bb�ˬ��\�9���s3��_o=0� s�i�D��ѯ�F�e��)�m�q���k��>z����Ȍ~vܸ�~����!2a�Q���ǿ�2pdn��5d�H�������YqUQ~0X�Q�0f�In�'#�MC�&�4�PZ���tɀ�l��$I
$+HX�� qA�iHҐ�mҐ�!IC��$I�4$i(�P��zwHC��"E�4i(�Ф�'_�����' M�M��tפaHÐ�!C�h�0�aHÐ�!K�4,iXҰ�a�v"K�4,i8�p��HÑ�#G�oZ�p��HÓ�'O�4<i�0��*�Y��;3(�,�
1���r ~x�vSw��"T�͘7o����j0�̫��k��Π��μ���!	��Ұq� �^.yd�-�u���4�ƃ,�G���:b�|_$�E�k���Ej\���q��Zdhu+��Ų��j�-Zz�Y�]�W���3�w��Z��?ۇ:|S�u�t�ƨ{�*{�T��,R�_��Fыv�ˇ��{�ǻ��y�ע��s�ѻv{_�ݪ����F��~׵��/��M�~�ҫ��b�@?�~V}جBI�����ӏ����MS�wu(���ϫ�j���>k��<�ںJn��L�i?���(����"7_��س�WE�>��?���H��1xܺ��V�j��v��*����*�yv-C����-L��,$�J�YSWaY�J���,����)U��� �+6�N�By�l�n��ѱ�� Z���ک�v׆��������z*s��μ�3�yE���������j���nw�5�kq��0�a	�E�&T B=�[�+�k�"�K�25�5��6O�:�c\a2�,M��[�D��=���%����-5!'�@Α�wC9���C�~f_ '�XNN�ec{��>��\�Ӈ.���Q��ȧ��N��%$��N=�d�M	
5�#�81�L���ʱ�|����уL��q;��ă!�_�`���yM�k�	����:+�҄حv���L�ˠ�Vڻ84yX��c6j�1fS�%M[.���a˾��Y����{���_����x�}�K��Gx�k���s�X�:o��6�
��!�)�BWWB�>�KQ��:b�ߌ�f;Ch����e�@�Jfj�P�|�P����D���J�_h�X�)T�4�@��f�|�?R�;R�9�'�|����7�~�h�R�=�:�w�����_��DZQ��v�����C�g�s���#������)A=Ŕ�$!S��N	�@����y�ᰚ�Y���t��l���t���EJ�C����44�En޾��R�:z��"�k;�t���㪕q��j��z�2JL���8	�S�z1�GY��B��"g��ZkZN�89i/��'�8{�Eڳ��t�=iOD��;��^1�@�b����3r#~��� ���ϔ���3<#8�xFpL���i�	�g� ��I��<#8fyFp����	�S{?:�>l�~��m�)I�v�il�̇���?�����dB�`êG~��}�Mbͳ�oC���Sn�(?�՟��fߵu������/��t���6��6�mrs�|������m�m�n�����N ���Mu�T\�7��~�t-���w��զ{Wtz[�ooo:
��yG?��}z��=��,¤��3	\MH����I*��r����Y��w���r�|	�]"Q\��"��{!D��@4�2��s�;�������R�[�yΚ��3�Ǚ`�̲r&��,r6Mƀ1=	�!��r�R����Rv(6͙,�F{N�Tgq��9S�����rvxV9;��,j��I;�ک�)�O����9����LKN�4j�S�fE�)m����Ρ���^��'��7G�M3�[_Ԭӕ��57D�5��gQ$���L4�j:2g��>�ne��1���j����{���X��!���X����^l������;z��/ɗ�PK   ]�'V�cŌ ~ �� /   images/40a6b5df-e714-4004-b865-d48720df955d.png�eP]��.
�����-�-�������݂��w�.��!�%�����{������=�V1�{�7z|�Cz-��dD�ap`@@@��ń@@@{�|� >z<�F�A@p;ݕ��]l�m��,��l��\͌A@\W�������k�u���S�+\��.�=�Xn���" C�lBC���{�Z��*v��KY(�?~J����>z�1i��9xx~U�:Q|rz؅�!ß=����~������tww7��?�=���!��M%6���wz�O����=v=���K:~���������wv��I���y��r0A��E��"����+��������E��bOj������Ъ�4�����]��ד�E��"]�o�/g't��b|���k>#�ի�������]�ޛ,�ĪE���s��&���0��\�*^�6�Hg�X|�U:��c��*5H������<U��Cx1sT�-����&vƯ���Ik��#w�Y�/��K�.M�]���5ݪo�1�m�-�rP=_Z����e���С,�ҷ.�u�K��`0~�H���$_ғ�UO�!b��a�Y�|�ܙ�	�\�!F:��INV���3�S�X�c�O�j<�/ާ�m�Dq[��4!�W1�����Ȁ}��/'MQ07+Ĥ�/J�(ml�R��m<�0kl\Ho�V��]ѼX�]c
=C�R��V`?��A�e�d����Դ\���4;IUݩq>��vW�mɩy��̮77I�wonV��y�p�ڞm��ĪY�mWt�s�wqv�|�r�#U!b�W����NDd!ra�|���iҜ�|�}�a�2���l��I��MT"�o�k�.��0�Е��*[$��i�'9P�oV�e�ܷ�Y�L��?��%���E.��jh��:vu^�~}O@LԤ�.�8Q�T18-G?��jF�>�����b;]�о9׀$ݞ]<�q�P,�>�j�&E��<*���=����Ӹ.������n?�vYJ���F �
u[s�e#�pR�}�z�I��O#����њ>=B����%��8 ~R�p+�-��Q��^������[��m�l?��w$銜�<���.͝��a����U��݄fxG�ި��|�F�A�������b n��Nt��S[��&񍣉5y1�Hk�w�U�V��]��j9�g �-[|Ԃ~��n�<}��C��a���u��jz��r�3x�ЗA?z\�~Sc��%@�������E�=��R�������@�ѹ8_#Y��W�ʁ&���U��f-ƗXJ���bv;�bi� 8��"�����(�$��a�Ndk�,��q�Nv�7[���L_�%����75?��l���wq��D�(2�;t��d+�#�|��^x�6��q9k��(�;3h�Y���82_¡�c��c��t���0��3a�ih�y��w�����"�v�Wݚ�9�.@����{L���OHgp��E�o;k8�2�Ԩ�y;�΅����S���r�i�4˃.0��mՂ����g�Z�I��rU�C2�n'n����:�_Pkk�-����H0�t�猾���KpS�� ���S�\؆s���E1���L��� ��Ær[�����&#�j�GS	K�l��}��fV�§��F��T�,2^�[�,�����������_x�h�น��N,��rm������!�H���98Q��~��&913j ]*�*NG���2V 1����?5���
���(�M"QX��?D�2�zXkS!H��%�-zl1-\��D�(M��*��i#Df[q��qK˪TRD��JA�1鏗�H��ll�!�Q�R�؁�*okC�p��-�A�98C�CQ��>	ί�0��}-k��x��Ϝ$�Yѹ��Ð<���̓�-d���+`���(��P9�o�[b���+�P��%���1F	�cEZ.��g3G9��v�Ce+����3tx��y!/`c/�;_3��B���`w
>5�%0��zj���"���9�o����Z��m4�2���/��� 0�7�R��u������I�x8�!��4K�f4D�1����<�j(s�%���05�%`IŢ
�]��%ǁ�+t�P��:������S>t�pUȼĘ&i� ��o�X����W���[	���uS��F�e�i�K��kCB��^�jZ�6�|_vl^��v�QU-�f����Dp���F���4�5(�\��POc^Ƒ0�4�����o>d��Ӡ	�C�����̩Ϛ_���&�f��|�����@�E{�*��1�N�'�#8�}&�mf�ݛ�()��0·������#��¼ U�X��$�kK��~�L�����&�h0 ��D�\ ���� �̨";/����Ӑ��bj9�-����T�}b�3%�&��~b����8G��F�P��W2ҭ�T�6B�C,Ra=�/H�8��3�t�C�����V�c�T����p�>��ف��K'<��)��#P�"hzg��ψеvO&��	9c���D��OpI��\���^>D#�oYߧ�q��_��4f.�{^�N8����
ϸH;A���z�@F�n�� G�y��� �w��!*��rU��zpgic�Kn���ᗏ>�E���x������,t��Mey�U]���B�i	N#K���K�Ks;Sc�x��1�Cy�ÖR�߳4~:'6ts
d6e��HL��5��P!�Gs�2���JгtsP��A/2�C��'�k��`��]�ځ�9[�6�\�[:t.A�$�:ظ�$�fQ.��V ��B�2�)z��L�
�:���mx� ,�]��`�'	���q)�g�qZ�2�������c����XW��/=C>foo�t�o��C�#�Z}�
r��q=�_y\l������5���po��4��8h ���4@����]�6s���T����R��>�V�K<v}ފmI�,f=�3L��1��ب@��h���]�������}\jM0��T"�)p�cuIw-y �m0��n�f�=�6�6J�C���HeQp����&[T� �.H�}5Xe��EW��9���,���>B+ș����%_�7�E�)�+/�@�� w�(1�fs��Lߎo=:#"4�=�����tv^f�M�>J��T�4��ەya�����h�0(��ӡv�8 � �.wi1H���0#=q�d66O��BȎ�Dl����W�Fo6}�!�w"��3��23�oJ}ˢ*�:<��Em�'����t��q}^(�ٹ�P~�����f"�N����q�ݘT?e]S� �e���6	�>�\H�_[&M�"r����$z�y|C��
��VA��ۿ*|�<BcGr]�R�SQD�A�E���.-����Y��!wf�}K�L�ҽE�Td�܈���(a��!��������������W��mT�$���\a�v>�PY���ˢ}p_�mv	��m�߰#!�SX�=jǣ/F��!�
Wb��g��@��D!�UNn�2�2�@�`��T3گ�)�Q��
���fn3.����}t���vcS�*א���q^9��"�#�2��J���q_fd�Jg����COz�*t��Z��T�O ��K:��ǻ�~��&D�Ƅ�ߝ��B7`)�u�"[��R�`7O�Q�~}FN0Z��S��
V�K�p��D&��+'FŠ�?��L?�7?UQ�{�[h#n"z�i�ᗞ9'�_��j����~�XTph��0|̋2��	�]ƈ��y��
;�E�#�����_Y
RJ" 3[�2��h�� 5�(u��=1���JD^�Q��!��[мQ+LLC�_�U��SY��s�,��#Bww�M�״e����<~r�0�a7�ўѥ���n�k=r_u��-+��؍oG\����+˔#2����@����M����Q7��d��0���r�O�n�tV�w�9ݠ=~堂6瘲���(o�!���V�Û�s�/�Ԉ��MG����h�8�������$yw��Q�����D�������yBU�+���
���Mh0w�1�PĿ��V��Q��at�ңp�����c��#D�axݪ�!�<r �{\�y�G}us|w�5M�k�H��(��v,�_�ʾ�R�%�̆Ɗ�Gl��
ZXhD��	 %����\/�W�P���O��HLN&Ks�R���@��̍H�������Z�S�+�Y��'�� a!l��s�CzR��'zt	o?E�FE ��iH*���s��=�RY$a+U�38-�짌>@}�8[�P�4��v�Qy����2�1yeMkT��[yױ2t�D����ρ1�`�_��|銣( pv��I�?ӆ�'T6*"��6�#�@Сq~B���V����9G��e<�:=�^��?�]����!??�|�Q�����堓n:�+k����6<�<�
hG�a�m���ՂC�&- n�q�����ɉ5�@FR�T�K�#�`���j�{�D&^?�iz����b�r�]�!� e���bY�sU���A�B�b��?194
��&�Џ�q���}eIp��H\ڗ{��!C�NK�֩j'���	a�����U�g����ΒH#/#��%�lj��H��Q�-}��$.9#绉��m3�AX�F�ݒ���S
R8P�sᯎ/e�])�/"�~�c8��5��A7���YvGz=���S"���~V*�����A�G��Zz6��fb1;{����a�J/��� ����'ɑ��J
/ٮ�0O)4*vuu��N��U���&�=���!-C�ϼ��B�+��$��������Z�_A�vZ�7�7�H����USkK���*�(�ۢ��.x糑�P�p#�*�xN���9aTu6����X2'���j�1�e��ƒ-Qx��s65�i��W�C�5(�5�/g�WW8�x��4��K��u��B�CP\�_d�`%6ֽ�M{�W�y���$��_���ʮ��)�C؛�t������]L��ۢh�Y�Qv!��W�z����A`ꡦE ���#g�48Ƶ�W��s��^O����DK��I��Q����ԟ�l'a�%A	������*Fx�����������8�G�QCm�&aQ��0���٣�����|/��sFKK�P^����XY�^��}��g�D��/d̂'	�%�Q��ZP�1�Jiu3(� !d��m�YZ�o�����xK �����,����ɭ�maE���l�q�H��3z�v'��&�t-��:Js`}bx�t	2a�G����q�L��|ھ�:ό��
ħ"u6���cw�=H��mW���Y��C�H���5��A%���%�bV�;��:�>ꁤZz٪Q�$�}�K�(|�G1{�UD����rK��L����c�����JF�a�`4�&U� `����Z5��C�у2��H,f�zQq�9�N�k��1�``�H\Asb�!L,����T�m�~U.E��|��5m'�)�R�1�w�{�:��տ0H'���gXQH��2��`j���}���]g��F-!�`@���!ވ��9g�u�O�.����{T3h=����5�7��Ie<ԿBZiu��cC��DF�2Y�54Q����h��Q?T���L$��KPG��J)�������9j_Z{��T�L�5>��^e��`��$)���ņ��[%25�:l��?Dk���$�D�f�\dT��$�hOEmB��}>��h�tn'����J8Ka"���gL|"��p�^�'�"x;b/�0~�&�7(W�[Ìh
*�aj1�U�OMܽ��?t�"t����|,����s����~��KM�Ɓ�,)�-��Y��N�q�P�B������[`�s��ؙ���DT,�;u�
�1�cx�R��N�#;�.��|�R��a@��Ť���n�NN�z�1'�cv=�o��Pv�ع��߭��('!��ǈaW�oJLU�
���8�#��(�#Qī���bo�k�bpf|,�L�%��+4W��!�R�������R>��.�ା��LƜ�A���?n�."�JmE+e�ȍ2��x�N �����
D����q�~�$ŶӠ�v^�X[/��3�Z�vKYPZ�7��
������e���*����IN�̓���	�RjM�H�?�`u{�ZE�A.6n6�,����;;��!A��-�m�h�������!�&���;� !�t�
I�Ps��3-88��y�T�=iթ)�~%�����̌������_o�������]eRw�-?��0|п�\�$uu�3j���j�K��g�琧�:�x������*�x��b%� �}�㢑[��u�`k�M"�]H�u���E�|V7h͈[E�JН/_��fe��ѥG�)ś���{��E[-ҝ4�s�һ��1��8�Q�BOY�֙-Z_�"����ɛ��?y)���a?�X/���:s"-��?�|8_i��#_�3J����[��`p4��	H�"�jޥtLv5h��m53�]պ�#�8��")>�kY�bF�C%����"H����cj�����.'�*���mD��0褵p7
�p��'�(x�֒R�y�ć]$@���:~�i9���zl}���&t��ߢ�����Ɣ8r�q	"c�(Ĳ,�j�l: --Bԁ��=�@� �a"������'�*�E�*�g��w��[J�����>���2G����A4ɡ��*ޙ!Hբܶbq��=���C@�~���Q�@9ɗ�	T���;zS�J�{�7��e�YH�/��,���؞��� ��� �}gcW@0+(+>e�Q(ge��9	ؓ�V��ψ���K�1�x�	��4F�O�i�Flݠ*���V
�16��y[�~��P?�A�I��j�� $��W��D��:Z�*C_l�Q����	Y�~ ����(
��Ŕ����k4���K�J��s�����U�S쩙BdL_ۘ���[8M���]�p�Q:���:��Z3ru�P�YFg��7�D;"���Q��b
�{�m�(�P�� ��V�C�J�+�|��:l����`�{������msJء.���=�3|2S������f��,Ӈw�;�%?$=��7�7>���};�@�o��Ŀ}��_�@@\3��x���Ђd���B�Kd0���HÅk�V`*9S�oӘI(��-zz��"���	?���n��i��n_�N�\o��N�0�<Na^gU��W������!���n�</M?�4yzxU�2�0��'���� MZ�@x�@Q�P]q\��c�x�jݹ�=���0���@ժ����̅���z�Ԏ�Eԫ��.�<���y��tʂ�Q������:]�`@(|�tG>R['�Y)W��u��K����HF��!b�3,W;G�%�8d��c�%a�\�w�p�����=ऩx�;�E�p$Vz9ɿ!Pԕ/�f4���"-E���?�N�����΃������}��3(V�}�^��'xg3%5G5i)N����������-ȟ����Vha�H``dbf�Ct��ED`f�C��"� m����L���H�]F	�n�0$���v�� �2r�'p���v�t�!����������ை�����7{#f:f:ZaW3gF"^n{CcN!�B|�x�Lm9��]\\�\��l�M���􌌴�n֎����� ��!d� �7�u4��&���7�qr�!"�'���Y�JK�7���?Y����Uߖ@�@oeE��3����3��l���l��F��F֎��
a����N���1�YY}�:|` �M����ܿQ`bfe�w����M�������?#�����l�_�q
� ��,O\���~NC��!��Wc��>�!�!;�-3�-�#- �����J���Q�h�꣇��ǀ���d�J��Чefef��ggf���g 0�22������ǩԷ��U��2��b34b�`bg�56be�e2��| 32q�0�L�����"6�V��if�obDokm�w��r�<D�t��#g��h�1��̬m\�gH���H�Q�� V6& ������������T��>��T �ߑ?�ǜ#�����N�o�F��6�J66�<D ����a��2�w��w4� e`d�d p2�)889YX��4�E�������K���p��f13��n���S�Fv�h��ii���_�����}g#C���[�}���7�� �33-�1#;-3;-�>+-;����>�ǿ�8�;���	�|����ǩ���?�����]L���A-��H`'������j-7�����K������>"!��������%�Q�%�Q�%�Q�%�W)���˔��G��qU���5�q͂0��{�y������VL����4����Q\Z� �3�U�� D\H@�u�ã�D������paw�����|�44�U"?X����Y7(�5D��494!by*3�S��(+zj��[bj�B�MM��A�0X�@i��$+��65�=3�cȩ��O6V�i{nS�Q��Q՗yo�xx� ��������DB����������K%����(0u���B+D�(��T�(H�(�3=�T)W~[���q}#OR���u)��-�O�������^�.==������S����뚻x�كЈA.UѸg�Ӯ�X�>��T�徊j�DSs�ܦ8T_�����p��eռ�8Y�Z��}������M��W�ŧ����+"LzC���F�|�ݫ��`qc�	.�H����J��o�V>�I/e%�ſ�	�ݲd׫P*}�8�T�'oJ_��*�%b��*P���Wm�54�8E�N�6t�9�%)k��ީ�}$�>S�aFW�d�m�����³;ܷ{�=1Y��8͐.,,,���J��$�u%)�>�A�H�܄��A�W�߈Յ��TO�7��n�rc�B�'b_�e��]�~/��S��l�������i��HDV�W (�'"��>�(><�b%��D��;�I��_�����x]�� @�A=��O���+�HbfuyY�[����"ʵ���i~��C���8����^ռ��$�(S��D�@��3�*����*�_K�a�o�$!B@��7 e����U�2hZ��^�ۀ�43��p��Z+��Q���H����p�zu�H*�F'���8��rZ(�������
������z�D:�M
Uw�� ]�0v�I&u�m���[�u7�AdET\���#4װ�z%ZVRޯ�|#����>�H�nur1)�U3M$�>[ �ȴr�&�{r�.�{2��!�*v�D&���q<��`k/L��${im�m������������A<ސL� �pǂ�R��v�ް�ੴgw�0�R�4�QB�@�Zti�d�0&��r\�����Y�pA�{HM�Ji
^�iX��&箼�c���D�֐�_���R�vG�z��z6�~�,����ﾓt�(�z�lVU����455=��|���^�����CHsp���,�ϗ!s��{$#�{>@���� �$����z8S��Oe����i�����>P� ˂:�7JHY�M1�����M'^/���ʍ�.;�}V�8�'-ù|�51/���%5����V���n@�y &}U]�s,&ݕf� " Y�Q�$��gI�#xĔm4ը�Ք���o�%SX;d��F�Mݱ��97B�ݚ4��x�C��x��^���.�b-��R���wa^�g�&�D��a�J��)��:\~͘ϠP��])��\����a�uvN��������]��rqq��7�W����0^���Ea���=/�!�>7�@�Vw<��Ѥ��2�����o��ڦ�t9D�u�ՠ�~�v����jG��������+��祡�΄Q�����m�i�/�#&v@�oצܴ���o�&ѠU����q_��Πf^l����g�6�(���~R~&-�Q�B�@��í�����....b�K��5��=o��x�tC��n�+��c��Q��(?hb�	~T��V4��hd�	��g�mlo�G7�,�Ud!X��Ő�� �8�&��rLZ|�~�uO�2����h�O��D���o���E���"�扃꼅=�gCL��EGJm�>Rf����.?���O�_7���<@.7mr	ѡ�>K�N������(9x*��L���z�ֻT9��e�]�������zm��A����#Kh�����9�����I*S]Eh׿�9�1;<V�.�����<�$���3��ۢs������c�M�]�DX���]��~���kR7B��!�����x��=}��)�� y2�}�`���]��VV�r�"�Y�'��VG_Ҙӑ��A�ՙtP��I��ZN��QVw�(JW��*I��Qn��,h!��n����4���;ƹ<��/,��(��.��l���A���L �}�)�9������I(ؘ]-ᾠQ����m�;��$��;�����77j٠F���t�zn6�Z.��P��a͟�*4��0��*�x�Kr|q1�x���6C�����6`g�PV�����d���@��N��E�Hy'����εo��Qj�6Iu��\�����;��%�������5�-� M�ȕ�`�wf9�x���L�T����Q)�@�~�i�����s��Q��3�)w^�k�88�ڽb-��j��0�Y�-�u8���HH�I�O��}��ӦEs�UY3D�
�a���IH��Ҏϔ]�Ϗ^���X�TӏA⳩E�:�+ŪgL���e>N;��\c���^��?�r{f���K/���(�ŋ�����奥nϯOâ���(c����l�����E�U���c�̔-ZQ��;���?�gܬ@����ʐRa��W1��3S!�H;8�X:鞯f#p�"wٱ�>� z�ۇ� X��#�:���������9s|�OF�n�e-�=G�B���0)+c�h�s7�T���HZ�U5
q�&������R̳�-M�;U����_�Lk����Xt�K�3�	����@&y|F�x<�?��,���n��A,����T�������v�P6�����j��Tx?	e_�g�D@z?�ڃ����C�׭F�<D��M�Z
C��cQ�Cǥ�G�ti
U��7y�"���Ib�@?�OU��fv�lޟ��&���{)>O)���F����g�k2��/V��NF�ej^>,&�1��FXd�Z�t�<Cc+hU�n:7]E�����W6�☄e7�Z�UI9���ݽ=�f*�7s1= (��;�`�[VTV~�t؇��{���_���~��
�KC̡��B��,E���of�����e�X�aȝ�����>ym�:]d�>���1��4���z��&�ψuZ	ߗ�R�]��^�t	ӂ*�=���1a;R����>R�k��������IS��=8]���E	�Ɂ�!	Ӆ��V����s��tA0v-B�S�:��rRx`��l�e�����m޾ڱ��\/�Q=u��9o|o� P�䘬���HO��du����%��O�����#�����}մu�U?���Ər������o�vؕ�>xr�ɶ�ze�9�R�=1��-4-�Y�VП!P�Ѽ��Y�c� ��v�����U�+�o����ޅWHۑ�	:A��Q�Q�V�-C���Ion�������r\j�_H�X䪘8)�ٸ�@�[�T���;�Ϝg0aYL90>6�[k啇6p��u���"W	��-�~��RM*^�����t^ܞ���#��#n$����������N�h�w]o���!F����(�b͍��-O���;o���9�����"X`�p0A��bB�υI{���`�H*�'P5(P{�l��M(��`*i<��:F�OEGn^�Nӿ��+�_ۺ�w%ȆS e�������V��<���X��=��a�)�e�wv��I6��o��&\�o�b�3��ż��C|��=/�ݬLUY�v׸�,��z�ɏ�������siF�i�JD�<����� a�F9hX��i	��2/��Zs&!�	)-��<&�dy��MB��ԑ�zE��ڽ31�
�
J�i�����2���%�P�6���׻��[�z5��;'w������%2|�����bZ��ܣ��R�Jw��4��@%���xI��zO��4���O0��B,�'׾�a���A�������G�����;�|C)F��`!��Ե<�hd�(dA���5�h�@~�+��'䢒A4� ZA9�U�hX�5��ޙh�#nbK�.*����D[�X�X
�^��r� ��&�� ��MJpH�6�g<��KeZZ��,����b(������L��+��0�%~T~%Є���E���1�d��Cf�;�QY�]�f�Z�ˎ�ӎy��/��̻FA�yS$CaM	�Я��kgyݫ;;;/--m=�\ b�%�T��SM�>��@�B�8�V�&!n�Iǵ/�d�*�B��@�fz:g�������p~P�d�Ί��,bh̆kP(��QG�.W��W�����d���x6��K��a}�o�Ih�;_-����rަc��f�ҡ"3�ʑ�-�0>�nk���M~]��J�vf�@�R�Q8��|@9J�{�r�ډ�f;@��hR�y�P�L�x8�|F���?���NG��7��������������6D��V;���} RQC��(��/�3#����tY$ֵH�B��,���J{��5��cq��yq��Dj�u�������o�L+��%1cO\��Ĕ[WhV�����,��(C7�Z1�0Z���M�r?�2Y�;��B�E�)�WSSU�9�R���Ԉ�V���=�ak�;M�l��7皘�h�П|�������ks����R��]y�G�M">��+��?&�X��.�
���ǥҰ2��&��k�3�Zۿ�zz�������s�q�����}�8��K�f]�h<XnF�NFT�¸��iZ�oSC�,��Z����L�<����2ѝ7"̺X�����I]�@���)�Lѵ�<w�$@�������L�Mf3�����#���ﹺ�>"J;�����3f�;� &����3q���vB{>Q�6�H`�$?2c��[�̤�Ծ�癒!*�[���ެ��b�6tC�4fB�Qi�D��8͗v�̇HE���k�?w1WنMR�9C7�4�=� �۾i7�U�]\
�R"�ʬ��;H(�؎�(Fl���Qθ۵d-<~;��{�vT��t��g�:&Lt5�,vm�/@���ml~K�E�`�z���������� M��
��61{���_\��߷�*�����fљ@Q�5�EQ��/�I�Ҍ�k����x5?o�����o}}�d1:�i�@uzm7	^�Q���r�p�|aY=������`s6F���P�q��g]��/�l3��3���F�k�b>��D����M�Ƿ!n���/�Hw�9]����5Ry���^�9��V�Qdժ��8N$��=ߝ|�؋w���A��ߦ��[���_�)���(�)�ЦMHb5�z�g=�r�q3��3
w��׻O�eW,�����Y���V�:� ���.�����_=���4	L+�����$���M����z�� }�5p�df���U�lZ�Fٜ�� m�Qz5�?%��X���GWnM�p��];<�":
���Z��^;�F05�o�e���A�ey�ғ骗r�
ٲ���e��w��L�r{��<�\ABp�oK�ic+c	�1��ܣduғ���7:����ל�ő"����IHF��k�̦��2��GR��[Peu�g�]��-��<	����hP?NO0�N�q���NMR+�J�
ɏa���u6�賨���h�\�~0ϯ�φ�g)�^<����P�����1����?C��zSڄ�*i.���[2������I�	̺���Z�4���3#j�[��]N0lOYD��,p������۲��Ĝ�#I�H�	�\�nV�)Y�a3�g��%�D��݂gh0!��H�!���Md�
]U��٣�+1�4hg����a�"��d4����cO��j��l�L+�2 K���q��в�Xe"�*3F�+N����Վ��_E6��]L�K��*И�I}��d [��_��Ebv�H�QY��(W�>��fH� y���Ջ���4|��V=f:GLhx�[M�@�HѮK���k���*�4o�J���Ob��\eb'�^	�V��S/V`����p���e�It�%J���L-=�QE� �Jײ�����^Å��нI\f,���ز���l��A4K���1Cb��T""U�?s�(����2�õ�t#�{�Ȃ`c`����*�5X�5+� 5`��X�����D�HGXՈ��k��6�*�k�j�\z��B��T�
�Jyf���	_���t�8�Y�������D۴�3o����;��b8!,��LAN��m��N���,����9ʖ%F�
7���ܶ���lE�~��X�j�x
�\�04B��U�IR9FA��;J��Qd��$r5m\(� �yb8���L)�vf&�+�n�Z��:�B!5,<�0�$*�M��c�4 �V��S����a�U�얽�fZ����#��ǻ6?�(�(O��}q8�Læڕ{���v�����ݥ�`4�v�1|��^I	���x|����#gf^j���3��qX�b�t�AY��	i��3ʉF3��K�&$�D�L�mޚ��"��@"L��+\J��Ue��0z�i�NG�T�9�@�m����y���ET�*���$�+NI_Q�������/�(bᇠ���Mr��1?��>ke��W�m�셸"9d��Y{ �)��$X�*����Eʰ\	��+�p�M|���A�@��B^�Aj%Ҋ��ѯR��_���ú˳��o���ERB	����+Y�%p��U�&[A���F�e�$�IV���E�J3@1Qv�A#b�G���u�sA�yU���Cͽ�������o0]/s<� #ǥ�W�T�t��rNK�|q+/*Q����$7#�)���m�2�&�v�e�r��0{&��-�'S"�s\� )n6���� T�)�
J~0|�T�yu ճH��g�*"Mgy.�b�W_�Ms�z��,B���F�%ع�`�G"P���E�M�^���|i�Gjgc�q%b?}��QҍS�T�h���pj��0|�����^T�&�Ð�ٌ,���'6c�"oh@U�~{��Sr��Qa�Mڕ�w Q���(�ZHiEr�%k�����dhu��SL�.�&?n�i�T�k�-%�z��2cuR����]���_�	i -���n�0���:.L�R�_dүß!�=�;ѫ�~�3�8�c=m^15oKoܧcd������_B^�p ��V4������1~����p�&�tX9c�G�ml�^�_�N1��]�khP��=?��ێ�)��߶NWu2��~���EЩ�\z\�Ќ���c�,�;ĭ5�n-PdWS��nY_a�ll��G~K�&�cЫ��V۽	z�s<o����xӐ�g�m�L����-��}"/e��+���3����Uϐ�Wꯤ��F�f�Fr����%G�(���:��Re�����,-����}�ÇfS�lĎ?E��"|�9��p���1hɁ���]ͫ�&H��&�Ky*8�]��BU�E9�$��M3���7w������Q�C�eNl�ӵK��~�(%��M�H�}(w�/f������K��kO�P��_*F�g��H($UFt��]��"��o�_|?2`��ynsi���z�<��\8������O<I���EL���3ŉ�b��[o�7bŠ��fʄX��r���������`x,��������0�����Un�{4��˙�R�r��Ap7����ps�4۴aG�ּq����}v/�9���߂��m04�J����N�C>\>0R�.��|����wu�!6�<�9?XD׼��
�+�G�һ�M���j��\�2�ǚ����y�JAN��07����m�.һK�f��~ل��\K�^�[�9��U�s[  �GO�=�-����Ц)��6udǛ��d��R�;/�R�h�0Mc��J�P)Q��	*� ��_���\��r{��Z6z�{�M�D\=���
v��,M������[@�K#L���+N *b�I�+]�`�ަ#v�e���AԞ��[����M�g��)
g���t���]�� ��.2mb��8���`�Q,��3G�o7n�F'9%e�Ie?�1,�'~oψ��T������N����swsKS�{9<�QC�b��f���|a��ʼ�NGK!oV-qP�`1�_,Ku\�L��viY��2��(w���vjJ�kg��)@l�̅���kP у<*�#fٷ�]�g��N]�����)����0,�țۤ�?�w��D$C�^Ǝ�z�<f�7>���������y�0	 ��\>/h�st�,������������qu��O�$���h��l0acO�ƶ�hb۶�4��ƞ��;������9��g�uc��Q��5�Kw��=���p<�j�W����5�\�&x�^QQ�}ve������p�]���A���M�c	��w���Ў�,!/�.��+��p�&LTJ�K�E-���<`��3�@F���ڿ�`�a5�*��#o��h���v�H
.�\�hMS?&*ϒ}��B�hX�T�<����^�}�� �.�E5�J.����q���ə�X�@�/�2$�nXF��#a�Z~$[:���Ю#_Ǵ����@�l����T;'���/珜��ʣ��8L�U�wS����O?�x��,;uE��=���DK�W
�JĬ�DBBB���;ħb~/�b��i��p4wK^�K������Fnn-:M/� ����Ƒ*r�x�ɰ����h�O;�r��`RY@z�M<�.�	������g�R?��N�E����a��K�?���8�UmR����*u�a�~�����%�xP!w}��t�\E�E�g"�6�dp���{����75!;d��T��mL6�N���ճ�D
��x�hb�!��[�i���b-�y�&�cl��딧��d
�{�h�ܟ�J��R�|և��K�n�z��&T�&3��-�4��w��	�fB����-I�����+*D�Z[��LeC/l�VVv������hx���df/�#f�����:k��e��-���~O6�6�It�Q2ohlTTD��^�4���1 I&߃�Y�l��!��c�'ss�lx�q�ݛ���˳D9%:�������Vl\bĵ[�5җ7�),M_�����TrC$�͔٢�r�A�8aO4���t(A99)�̵�j8*
%�����%Te���M8�3�V��7��𛳴P�^�Y�܆��[�N�ǻ�cW��A wO��8���Ѽ�e�޿Ƨ��^C^�����+�	b���~4�	���_��>�����?ϥ��ؖ�J�7�����vjֶ��ܱ1h��5�~:-s���F���Yg�ϻ�>^o2y�~AF�����gt rz}t���5����v��~�I#��:�UZ���S�ΪU+ރO~��R|����ƚ(��h��<*�Pmc� ���
�3a�-ؙGSD#����]���w�&�`m���=���1��,��.�����V���c����h;N��?;����-R�������Ţ �D���yuu��y>�/��b�H���=o�o��U���#��Wj�������Ii���P�y�Uv�!�1r���	���Ǒ�����r}}}��������������$�Ͱ���������t�夝o�X(�U�[g��S���b�/�����?����kk{��b��Ḡn�nҗ�?�n�b��ݺo�:���G%9	9�To�9 �A	?��o>�w�����1��+��!����	�4�B�����nW{�W2�d����u}����D[:>�,��'�^�x��c��8���c�ᑦm�������n��}�I3�i����&�OI�Z�V�e�k��O�U멉� ��@�]�5���� B�qa�Ә7.�`��K�{Qtm���66W�	;\t=@�;�>����w�]��<�QR��Ѥ��-'�7E!�<�T�ZC��?���n����9����a�����8�F�y�gc�xѲ��A�eU�J�eu����3@���\������뤚ZHqo��~K��/��]ڶ�C�B�l�B$�[PC�l\ ���uG�K��H�+����{[����B�&�}� ��d��Cm�Y�v�0�nׅ�̫�Fs^��%��]o<t���LC�8�mZ����f K��q7���+ƭ�%TI�
���49���%�'�p�;4���o����l�9o�����l��9�V|���'Ҿy�7� $��*1[��ȅ���������W���ϳt�(Ix��ֆ�lQ���9Y5��`]�_hO׸�p�!�����bkV��4@R��|��6F�7�q�I�TO~ש�k������%Sfxg �|z���6Offf������K*v=m>�n�������RD&����<;/|.��{��-���m[ƽ��!)�o�Ї�p�.�66/��帓�w!���E��P�o;�O�7߄�Gh�*z���YUˆL<��%)]��$��D���%�&H�?�����伷��wf%I�!�!��(�v3���v�A�E|���������~9߅��mÃ�m�޳�(L���TQS��C�s�3��J7��G�玮ܵd�NMb����Q����h��@&�FA��HV�+"/�2��|���ĥ�2������l�&�b|@*%��E&������|l��z�䤜�m{��ypb�-�O]�t�bx�����n������6ZJv.�Uw�ߍ�;���ɿ ^���/��vݩ��%-�C�
$A�Y��s���a/�r���7�o(����뛝�HF&&�M��Yۖ�p7�*i�}}����|��X��Jr��W�,S)yܘ���O���B��G�e��fIއ?�U���o��v��q*�txܲ3��2�Ѯ��I?�6��U^�(s�(59�k�3c���ٳ���<�?9][^���v��vF4���O�9��w��wK��ЗOܺ��F���?| �6S��9A�-(j�n�wI�5�|���p�{
�?ޒ�J����"Z╎�OT�������p��]�㐴+��Ь���B	;���WG���?�3|lj�돣<��>��lx]�k+(y�xd�T}"��FKNOOU6nX>����`��\c}Ҟ秙R�{Msw�n)��� r�6�)�Ъ8!�Tb�������ق$*��5<??���'�-��Ǹ�k$sq=>/�L�S��H��)��~9���t��d,��m4�T�\x��ᣆ�&<O(�.(8�уY�r��KH_��&�3~W��y�������>��a���g���X�{��%��!0����U:9P����cP�&w]w�s����A������C6oxmq�vF�o..�1u�k��p�h��u^M���V���1�++i#���z]� ��"aإ�=\,e����x��v^S��W	��m�&T��-=�5oϒ�_.�,�B�f,���������]f��N~�7٤�ͫv4���DZ�b�ƽV��p��N�${n�>o'�9)h���'I�}�M��_�dB-�@ځ=�?�o4ؚ�+k����Gؿ)|�SߊRQ�7��U�����5�@�n6f�����M�-������O��[f����/�rY��K��]B1]�|6�^�vH�~��8(����gx��Z:G�:������7n
.z��Ȓ��;�a���nP�� �S���㒰�T�� �'pN��	y��kReU�ͤ�Od(�/>��t���[��ϱJ�}S�~օ7͙�"��m"W��m; =���Z%q�)�/JC0'�0���C3�T�zi:��h�E�m�j,uE6F?.�ٲ}%� �M(���ꍹm��f�qĻ�+jhū����B��@� �q���Mt���o�~�n�4/)=I�ta�YCd�� 5�����)\�d{_ۍ#*oޞg70�܄�=J��t����[��_�8k��K���g���vZ%nq:����~�&������I�]--4����	#}0V�����Q�*}H-��d��m��tД��1�E��0�X�����*��:,����5���<<�������mѫ��{�2z����|��o-|_Z�2�%ޠ��UN��_\�;Gd}vn�4I+Ǫ55�;�����d!B��0PX����Y�9�7&y�F>�bVH�;�5xf����	,���9�?~�`���֑��g� OO�!����-*Y�1���f|��kq)t2�!i�jN�zIJ�2� FR~G�׍�8<�jL@�
ۯV?��4�2�xE@ȸ睧N����ܺ.�)[̩l�k7ѕ�:�2��W��ysl�(~�Pn0U�*��R`z��my:MՆ�d��ȵc��o�K�Ƽq:�o���G4��JY$d�DY9���=���ܖ74�؅�H��l��u�j!nhj�_�e��c�-vz��`�k�*����ֲ�������a%bH-k y'�ф��k��*5�rJ�G���.@)�#��ɻ��e�ʶ��3���4B���#��!�ʿ6��6J��T_2��JW N��=�F�{�7�J���@�Rf*�΄J��������D���K��df��Փ6yNC�J_�_�D�c�tA$���aȠym_�G�1�4�
/\�q���Q�q���+jP�o��u
��>޻TגKͤC�&�_��Jؼ5�3%�T�}���q���ݿK��b�����kf�bO��BxZ9�D8dc��,`	Ef�\�vD8"�	o�a{��ܿ�Bܱ���`�;�F��[q^����խ�ԢZZ�h�XrF�b9_���'1�7_0g ���<������~�T��f�0lڈ���X)�a��.��ɰ�ӕxqj���h�'Z������Z{_d_������lCvW`1��b�2_�4�`\��)�O�~��`�����7��#��'�M�aMII	WS�sg�S5	�W���vk �O"����U� D*>��I"�5���z�K���r�ku�P�d�=�~r?���<[�;�<�HḾ��k#]��>�D�C>�EA-�n��g��*���б������#؟�a�E4���DT݃WLhDW���ӣ�����9�*�qm�+GÍ�kV�R��Eḋ���F�ek�
Vm�F���5�U���^>�*�w�����Ge�	����N(�����2�6e����l[dmkƾ�#+�`@L�K�na���z��W�mv��g�ު+>+If���x�:���޶��f*_����g�9�!ꭠU�<����~0u�T#��s�_{�D��4�# �	������XE!��y(�J� a���j�躇9PŎ�ܘ�UЊ�S���i��Y�S�))�ϜQ�ϺO�ȆS"�=� \Q�|��6k E�?�N��G��H������ cXr{�[�ò�-Ċ�/1QR��\�Es��rcs�Z�|)��{=����-v�v`����g�ĕ����Rk����r*U��q���ex��g: �_-�$-a�g=�h	���ȥ��T�[�(5��15��"��M���ؗ�7�(0�Z7�+�hŵ�yG�prB��z\H
NB����ԩZ5���u-l��)�6�.���c���l�ߨ�m��Z$��+�T����Ň�bb�h�ʖ�����P�0�u?U"�Frڊ&�fe$����B�h�n�N�%��N)-	y �8eZX>��R�s��`�36��C6sB@k+T�P+U��d'�݃�m�Z$�N�"��`��!�(T1�$'�]�* �I@M��$f�Nm��[��&��|�Ă��n_���7/R

_����c����	8Ӻ����P0н�G��̼���񬿡�8YNr*R!Ɯw��Г=j�$�� ��x @����&�Y�/Bվ��������I���>b4���7��D�%���m���+�"O���L6j�X����7Ԫ����t�^!�2�$�ǎoa[�I����'L�L%o��M�X�rX���}��`Q�A�"'��u���+`:��Y%vrρ����Xr�+�2f��iG`tE��aUNG��|�U%�Ac�z+����h{�"YN�z����'y�Q�V�1���)�NU�_����ZDࠑ��;���e�j���s�a���Q �`@&NQ!㸹[���
�X%�Z����Q5� X�T��a�!�d��o���*�͚"3��#����76���WTP�����G��d�W4�7���Ц���2������6..�Y_�����j���=wf��.�5mf��)84�b��}��"������l�B�G�*��yv��͂��zo�wBv� .[GQ��QY���͵�䦽#��0#�Ot���	�ߕN��ftN�z�r�~�ID��}u\mJ�����r�}�6��2,9�a���|�e��V�l�'C�Q6�;r2=4�#���y���Tx*wUm��ٕ���\FFD�f$�tt�����0f�x>�w�0-������V�+�rw_��n��n�8e�BCc�
����o^ۻ���c�G�!Y(
��)���F9��nQ�?�3W��VǓE	K��v��H�=���$"�,P��iMBUO�o�o�qMB����Aq���2w �%N�` �tFg��b�����1�s�� ��<j�t�][�7������:��6��P�,f��ö���%�~j)�57Rh$R!�k���MY���Ed����g���
ӎ�䩠��5�3�ly��kB��Q���m������Č�d}_��O�p��]�s�7%r��&�"Ȉ�3��0����p�h�I����z6��� �p����.�6'cXU�2��e�1G�Db�Y�	UE�}e��Yd�����$�,;WV{�� %� Ǎ!�=�0�'4%�sl�2L��Ʀ�P��}���o���{�^�U6��-���g�Ѱ��.{�0&oR�R�4�8f�j�h6����d�5H�׶��B̺��6H��9�?"�*=߲e�2�.p���";�b�U�����g���#���x: �Ɔ��*���^˨��Rs�e ��ԭ�t�Y+�2��j�B�Ƃ��n�٤篹���Ks�bG ��YCJ���A��@��ˏ�ӓ�� !J�-J/MEŎK�@[�(ΐֽ�U=�����B�^o�C��~���h<�Q�#�:��h�vTg�u�M�}lDÑ�Y{��;_���K3���#�3=ޝ	�'n2���q	���N�4��`6V��CnkL�@�ɌQ��k߾��]��X�Q�
�q�Y�  �	�� 9	J  �+O=�:{�&oܒ�ڳ�SD�5�g2Y�ޙo9��^�>�ok�]z��Z������*�� �\6qQCD�y|7"�9DP�ޠoc����zD[ޮ{�_}[�)J<2���ݴ��-���2�%`�zƶ�;;I̺���h�0���܀�+ ���{�つc�O�w=����V3P>���'K�G�2��NyF���11)	Ƕm?9�us��Z�v�*�]��e��ٝ?W+����w��FA�\����u�TQ��YX�"��G��Qw�o�ńz���(19����	>K@����W�O|ƥM"�A�1�5LCDv�-��,0ԓ(�5ñ��D�cE�6�0m�B�C�4���B��[���S����匑�֧��t˘|ǵ�}��#���\��36Ә7�l&��s[���id��]Gʘ;����4X���h������SӍ���(��q�mn���^s0����jjn-�=29{���/x�T�.]8��e�/�|^���zX���\�2 �:G�n���ח~_���_�4a���G��o3+g��'�gC�?�y�Ki������'��c�3pL*�6�E�	�/>-8b�����4��֫;T��j���nPHg�^����I���D��e1Ѭ���\m��.K�d ����ŲS�P�&B�[�]�:��L�>�0�4�
�Ho�փz愘Di�?����w��|�%�}��OaHSz%|�g��R~�w���jLu��� *��y0���o�`s����c����*�H��D���P��Gw�Ƞ�u[��In��+��͹*=��P�<�$�4�HQ��+�ݸ��h��@��C�-����k�z�\�9牮��������Md86��'dRU)���z��������}37mt���~����ꦵ��S�э����F��*u�����ֲ*DrJ_�;�	�@�H�t�N�6f_�J�C'߇��� ���SP|��^��d�y�$>�TK5و�455��9e�a����<$J:F̭���,u�8��s���7Í$
`�a���J$��[���f�"մ�.���55r�M`����߷D�i>�?���w��-h��l��ځR�_s��
#���)A�{��1��R��Zqn��;e�j��屃�DM�8u\
�Ҵl�#sw�C���o�9wUr;<?9��Ifы��g��U;�z?�Ę`�S�̦I l#$�U����L|��|�:W���ۢ���4�*��+{bޮ=%�(�B�pq�ੵ4���.n�>���=��i�16RK߃J|3��FeK#$� _>���X{��C����F��)\���v ��H�Q�@�Hb�X�r2-�t�h�Ec����S�-���>,KD�?������1��]�3�=�p*�t��躆�1G�4qQa�O�xP�q|�q%�sC*A�$��!Q���"��A��+W��/	��{�_Y���a��3�{i���~���C�y(�A�d6�&I%��u��ԱŊ�)o�§M��傴���i�Q���`��X���J�8R�:��Ƴ9|�X��i%�i��[�2	�?ܦ�Z���&�޾����J�zO�l����6D2��Fw���H�Q���9zئ8EA2tf%1�C>ؓ"�]YҺ���8|�b���Ҫ���L�]E�mn�S3C�E���#��Z+�b�-�SiT
�IB�ۥà�,���`�Q����Â�s�L�j�0Q;�O�#�M�{����+���Y�M�[���Cf��y��dQ`�U%H�@��}~����1��O2j��ڱ���p�ɘjH��5��+�u�����_(��u1�M�,^��y�;�(���
!�V\�=,�<.��Q������<�B4I	C4��ӒͶ����^�rFJ��Ey_�� 5kڍ���x/��~Cox��oϽ�A�S		���9̶e���$���G��� *ܧ�%�U��N��5������M���+O˦/��T<U}j[��������Z||%I?�T�.�!�L����Z��S�I�CO�$�.ya�ԗ��v����RMG���S ���p�6��\�W\k�Arە��ޗ �B��SunΒ�����Y��#��R��R*pﻸR��!w��F��y]ck�,�l[�H��R�yE�EQ�|��T�O�}֎�tq���s4^��F ���2�Zd�B� 1��V�|�]nn]v���{p:�B��u4��6���C �y9U5�@ �Oh�Yo^�k퓚ͺ3Ĩ��6���?+�e|�Ev��]W>�b�vs�q�.j	�J*���#���Ƶ55<<�Uړ��y� �SVޜ&�"��-�6���a����KJ'[��?Tv�q�N|�r�,���apQ#}|,ۄ��x�?Ih7�W��u� G&�$7)�x�d�PC�u�n�@s��(3�F����|Pxƕ�!��P�1���]4ȏo�c��#ƾ���B�s���Mwf*9��ҺJA@���_G�[��s`�c]���H�y�ں����;@̍�h>�����*��|�����l�����t�㣺�l��*�U'8��[t�}�	�7�	X1�.�%K�K�i�ӕ��\�ur�S�8P�'iA��l�G�N9����tGd�;AJ�����{nK���J)��f��/٠?�0�|�q�plQYF]]}̾��&��T����j1�����V`�6'*
�כ�s���1��ЋKYxA���+)\g�yJ�G�V�П0�j�F;��~U�p"r[s}K�E3�`ZL��B�� �s+�khƍ�5��A����4L�m�NY$�1���)��`��c鹥��Y~�ŵ524�aƸ�8qvs��꼿�3s���\mW�)�~�9XG9�x�,9Eڞ$&c\��5���2x|��_8>���t., ��>��6�Qۜ1T,u���%g%��������n��T m��1K���bAd,G3����x���Z��ܻ�b]���R�eӠ3��Ed�O�2_��� ���M�<\����2܂_$�P.��_p���$R�2���b����M�0������~���U&ˇ'�>s-�dL��,L�X�V�<�#���K�{��"<��L�D��q��H(�_��`J�\f��E)�X��Q0��R?���~�I�3;�Ș�w�YI�LP��(�hX����>A继��0�FB#��9L�q�om7�=~����*y��`Qog��F5k��c!�y:�}�Ԛ�������U�`���q����}z�6��^��yx�M����h��D�w���E�9{���
�.�|���5�U:�e�|� �R�Wx����B�	��n��-�
�ay'�#O*�U�[�:{����85����ig]-���s�m�4�4��e�()���ꑑ�׫�+���,�F��CK~ez���u��3�َT:@�X���F�2j"(1�A���|�mr��lq����x5��I��(�y�΋j���@����D`�b�w'\�jM��<��sN�tGww��b]�$Q�)�Ά��/�����+�1�+���\e#��;J����f+ڽ��q�[~��"�����o�A<��_E�������F�A�C?ѲI��[As�m��� &������Q���
>�Ns�/���'M44�N������࿐i���T�ZY�/�Ǳ�}컽��Hz~w.äbm Q,j������K�gѵ�Q�����ݻ����?���/Mu�|�,ݡ�_��)����ڠ��g�T欔KPBD�~2��G��̙S�QRͥ�����\
���������,������`�`b9�]��=��|�y�9���mO]�L�{��`�����]��s�vmYL�A�z�0p6`Gx_�� �!~�/��o���p�e�}>����O
�%J������0�U٪MU�V�{@����͵�߹%�.����|8�K�����q���,3C���`��C0��'"3-��/���"����Ԍc�&���hRx�T������w��,�L��(G�����BT (e�Nϯ��'�#e�G�lLq��wR\�Fԛ����g*.�SI�Z�/6w�g�,�����C��g��X��S���z�<�WI�v84n�h/χ��㈠P���n�v�[V�����3g���nr]~ˇ��I���B2�k�úqls	2� �V/!Pɩ��������^W�g,d�nۇ���o�1� �x&�SY��rY_�8��� kH�T��w�¶ӱk�za|��3�>͓��w\�.s\`ܛ}x�(�,�=v:��������ՎR��jIg�HiSPk��U[O�K�܏�D쐝N���]�z��0$�w�]��Ԍ�&�NeNy�-�-�|�����`�.��0�S���Z;70��+��}��^xp��[7&�#��Z!\�,���V$^<Z )��f)B��wf\���L�����@n���Xi�U�y��ێ�`�0�z� Bj�s1(�ǡ`��V�.��(�/V�Q�s���(�����4�e-�6;����v7�hF��')�\�	��Ϛ�e0���FU[�3���x�$�t����ꪣV�e��B=ޞ�lT
��֠���V�u�o���*loW�Ĳ�N��5(�tҜ��/m�˚��|�D9�����t�����^��R��"#�5��������>�_�*	ѷ,�_]��Ɖ��1�q	'�@s�����,�Tԃ�5Mh�P0�i$���	-D0=r�@�u�"˜sſ���g�n	Y�"ou���Z�pl0�V��ʼ�:���>V����O�����0԰Z�X�B+�R�J��	�͜M6��U��*AKr��Yn����
�2�-�*�,	XH�9����Ĥɗ�A<��D����i����Z�bOy�D�BQ��.��Z\��U�o���Smٸ�N�ȥ��������Y&t�ᢡN�2OJ%3�5ʶ�_���QK<�%��u�(q�����#��1� )R�W����o�c����ɬ4aL�<�*6����@���+�v���A��M ۯz�I��pL�f��d��e��Q����8lB�gЮ�g8�ľl4o�<򲸈�"�����1�<���ji	�X7T�)b2��:��Xz����]!
9ݬ�<=V|��ǝH�?�]ps�[�J&k�_�L��*�e���D��d��4�N��7/�ȡd���M>(��`��;:����G���~�OV|t ���.����$X-l�TD�q.�$-�wL�3I��_P?e����@I�sz�@�)8��dY�F����:B�U���I�Ʉ���}O7iE���3M'9.�w�\>�W�QQ��	W�c�����P -G��\��~�nޟ�2Ƿ0���;���'e�����ː%QM�I��Lڭ��y��������N5����N�p��ے&�Ś���P0H��|��l�~|z=����O�k���Pn#�i\p	Gs���c��iB�O��%�^6g�P����w�rx�����B��|'l_/�Y�kA��p��ƃ�?"��ǡ�DIA�U�5�dp�a��_&��%����qۈH�6�!Kɜ ,��	}g�����%&H��}�lI!I71k]G^rƠ�f�#\t�&r9�������|Ʋ���.�V̪-Ǿ�͙H*��\��R���W�ל�ѐt���egBG��1���q�\�Y��y������%����!$�Ԕd�ĈQq�
L�|;�������zFdѽ��� ��ܮB���oi��j^@'�L���+0D�2��3'��{^z-� 6p;�јhX� ���e���;H�ZQp��C}�V�߫����
%��6rZZcs�0��5(2�4��V��\Y~z�A��M�?~:�UnE��}��ڈd��"��۶D�x7#T�Zwu�?�Ed�
��L�}�F�Vg�U�52ʒ{�罸R��2������zo�9��R����G�A����)�ȁ�m>���kԍ��/�*���E����I$�E��v�Ϫ�������oGͶY+�6�kQ� k�${>���M��M>O����Ң�*CES<aJ�<�r!b0�
e!TmE +am���	���GP,��4��&��#n�#s�tv!�/�*ܳ��~�o'���+e�(b�ۄ���睩�<����GC<Y���yT�!��o�k�����AdDa�p��o���MǋT�NW<]�G�������e�V�.����U�<NMR���X��k�ݑ\�o�<��*.r�m�,���BLJ��j�vb�Q\�������^K�o����Y��|��A��q�MS-�;�X��aP�w�j-����Úײ�n�p-��񽇍8{�'�1|l����roq�s����P�hE��dZ@�@��h�pG��
���B}��԰I|*����	b�Z��&�H�g���ĮՏ���$$�+��*�����2ۊ�G��LJ��(*�U	7r
o
���S+5V*�p��L�w�P�����d�UT�ڶ�bb0�c.��R�Ғ�H}]�/�#�E̓X`Bp^rn���%�{������Y��n~<�=m3��ݙm��S�&ۧ/>5qz_�5����挈~�_�����g]�gv���D�Փ��M4���=r��=N���8��/�����������ꗝ�ŧ�9�ҧ��ʿ�B�ڗrM>cΦ=��t�Rҁ΂��Op'�-��o�mSQ��'�95�%�Y��y�$�QI�Ͳ\��'����](�8����?2GD=r��K ���Fv�a�In����Q�X�DB�Ŋ�a>�\�ȒȢ��E���?�S6X���Vqf[��rHm�F��FU�e~]9)������YQ}֩�K�@� ˣFP�����Y��j��;1�D���;$pm��������b*)��N�ie;7>ƶQ�PY-4Xx x$!!���+���kXT��&��_�O"� �t�1d\�d�%�.�˧���������u�[>fƧ[;˲��H������C��(�B�9�h�d��6뼹����{:�|8_IP��{�Pâ�޷ݼq���DMs��������ǲL���J�LTz�d㒋�P�N�x�[��!/-�w2F5���r��]I��'�;�(��*���ɑ�אm�,�,���릐d��Y>��W���3қP_��oTg�g��m7sr�g}�켿�w��zH���P={��%�t�8ьɓBG`�=�̰�=~�z��]<�)R4��`�=��uZ�N)��ن'$ɰ](D��Ȼ#�D�0�aN���RM�Z2�'� <~d�H���=�=�Hi�[&��;�gQ��@��P�ƕ;�~"بw�y��*�	TZs��h� ��JL��T���'��\G�T���DF����^�tv�3������	u��"o��Zgݰ����s�R�t�;;��VSMτ��������a��s<>c�_F��������d���:�\u�d��+��׼�&�(spŁ��f�("(���y���ݺ�ݘ+�e]�_|�i�x��	��t�t���8m�eŊ�f;j-ܗ�n�
��9~����g�<�2�AC7N�W�dyςܗvߖ����n(����6u5����]��=�E�,OP�����.q������Ă*@�v�m�\� �^<!�s�Ã��>XD؈--�иY:��^y��WK>{Fc�$l𵹪�w��
�����Ǜ�y��Z%�d��)naW��̟��R	uUa��[d7d��9&��0��"@]W���;u5uߝ	�K�����b�)ѭ's�E�.^��U�f�z�z�������ѫY�H4�����C�}y���=C�ӎ���&�����l�_:��h,}�������t���(2��|39�Xp��)��~!o/���K+�Y�sr��=�ދ��~���5ˤ絻����C�`7:�9�,)X�V��{oǌ2&"�R"�]z�|:���D�M����;�c�'(�o֕��_��������Љp��t,Ӫ�r��B��(�����ZQ�(]���J]j�=De�ލ��(nvp���v�ƿ7�X�����R�{��D۲�ZMF!�Z��G�L�9���I6���1��&4��G�$�csu%=�rO�D���>�$\&�7)�dZ�LP#��ciyC/�ތ�
�w�J�^MX_-���->N$ G��W*��pk��;*a��~��V��&@;�a�:�«�hxM-PY��M�	�#�<�p�v�j��2͛=��/��Nd���~�D��hL�؆�����.>JY�����j�{��%G�o��yꉛ�a�U�W�ܯ&B+���xu����{�����[AV��d�i��/�����[ Gm���Q�m~�����/�jҧ��;�wK+;<�m�_[�>�ي����7fu�d����]zs�<�����U�����n�V������.�i��s4���D��V�����W�p>m*FJ��Ƙ�Z[q��D�tC�୙� N8�OR��'�qg��ej&�M��݋D�{.���SU�J.�I��x�(�]e�d�swN�MK��^]tM�O�Șox������������	�?�Rx��_ߦ}%�GF���/��.��AGw0�Q�L1��E����q.��z��jI
�~�XQ�\"�:�W{N�u��Bl���t+�rn�v*���/E�;�u�ZR��F�����).Z�j�WWl��n�������t��AI���6�6~~���\�ᬷ����E��4"n`��B��*K�چ��5�h�y#N�F�f�G��(p���Z4�tb���@����(�}j�]4��%�ee�	�X0"���&\�8���',����^�
�����u5�x9�0��"Jl�i��'�Ւ�Ҟ����.�S��S�hO n��^����T���(���I����!--�_��[b���v[Zx(��7U&Z���ߖФ ��p���G��JW�e�"��2�n:Yen5}
�� կΑ���<m�%(�j0E�x�
���o/l�5��F��a�'� �\(aO������3lY0əh���%9���BKN�(��9�.aPI�;�(��^7��>o�·�������#��pt >
�D��ׂH'��懕���[�~ʼ*�N�Y7�-��#�4���AK>���Q\OK}YD��{��%��ߧ�i����MmVU�T�pvq'U�e6c1��$IDqw�F*�{��N^�
�%�9��Lj���F������V�G/9��ɬ .ek�hp��O1������;�[�)�sV��\�<�.�����a[��a������W_���:�U�J�C��l��ο�I�N�*��9�r]��y���b��O�-	�.*�I�t�a^nL���P���3=A�\�E��?vSs�$�K�,�lAoW����p�ț�Ef?���G�6Q���/U��L�r���5�p�hy� ~��;��r>m!�@e#-\^�8�~�fR�����'o����mԄ��;�
�����j���0N��.���J���!�k)�R������
ww(w�/<���e֚�L��}���9s��S�Y^X���y��K�%��A���Mye��42�P+�F�9�x�_y�Ys�<����w�rt�@bXq^�#����I��AI.X {�9��셊��?Ǡ��r�b�('�ζ��U�N��x{w땱VV�屳��'9��z`ۅ]�n���$�h��^�ܼ�K<+�p��r塼i��n��t�-0/���ѵ�>`�}Sy"D*�o�i�r:/�Eͼm��0.���������g�v/���b�a�`�D���w��^�_�ŕ�	V���Ӽ1���.�U��^���S_��j�8W9eL���@/Y 2C@-�����u�c%�^z����0��4��$3�$�B
M�ܹ��XxM@�ӪP����T䔢�x�O��^�"c&���"��Z������2+no��v�}�n��hLӪ=OI�uQ&|Ji�k��HNlz������g~�s=�sj�w�lp��t���#��r�g�B���J��i�_0�+tG4����vj�Z�@�A<��R�T�ϨH�_Jٔ����Z'7��J�=�%��<��j�p����?�r���_>����v���A�}~�����*�<��#p�y�0���A%�����2����t�Ϧ�)�����?6@�d���bI��,��y�g����w�ۯI���������EKm8����+o��C�Pu+���C�HK�ྲྀ�>��T��8V��_�F��)�^��������
��P�5Yp
��Kxt����]��v~Fp"q�d)`7��^�5����ʒ�_3��r���-),�M��o��%��va�[t����4��A`�րѤ��9�	�-a|���5�.R:
������!�9��1���#���mpND�:A��t�_b{E������!����v�ͨ��V8�0a��S�#]�����*��]Obj-���!�{h�:PY[�t��H�Md%���[�f��堮��y�߉,Ք��b�Vb���\�6��`�]5�.��-��@*u�Cd��l0�j�w*�L���0��U/
�+��R�Y����×ฏ�S�1�h�m�8��,���f4���*R��n8Ӂ��s��L�z���jGMP03��f!�[	��������u{@>'�Y�Ι�-ڄ�ȧG�	�v�[2�=�5���E���)�l$!mb�[��.��->��tn�h��43U�i0�Ed�|K�/�U� ��F��7��ЙO��z�V��Sr�r1M�Xu�"dv]�ܱ��h<�\�l���R[!�ܚS�ψ>#]�&����[t���G�
��D�q��đSm��p���C�e��@=�������I	17�*�)4b����{�����\�$V�]�L���9��U�~�p.��7ĿT�2p>�I������'w��K��1=[�&e(s����D�gv��8����LP��}�H���������9{�$�V,����ݡ=�]�����.�r���y��m.�����t?��_�u������{{�p�ؖm�\h��X��D6&�� �`C����l�Wd�n�WV�)�S b��mn��]�2�y�
��#9@�9"��^?1�)���a"���S�ȥ(�綂+��@�Ƅ��vC���g|j�	���̓t�&�c��P>Y��Rk�+������+#5��B�cMnT�yI�i]��5�C��/z��Uq��XT�R;*��8��-�-9E߈��_�-3��DOG�������:�+����%X�_���D�A�R�\�G2Q5i�����p�о=5�4�_� ��61��ة�%�%�����-�r%y�h阍�O�ݫA�fޚ�˒���k���8,�77�u�\�)G�/�d��k8��<�_$1��Q�Y���żC*�8�H�#s�Pa�6�Zf���ġ���K��$\�?ϷW� 6WmK�k�d�yR��A�g��o�w�C�/�s�a��*��Elh��95?~�gw�1��$J�5��l������d$�(��a��U�~[-��Ec���c�Tp�~$눯:�(�O⿐~@�8��gr��D8$��pMe ,�
�,=���R�l{f%&g�����4�8�&�E��.WyRZ���D�̲������a�2N�����t��ȯ%�����z�ݸކ�T<�h-ˢ�-������f�����h������غ��吂VZ�]"��"�������N..��(����T�#
��_/w�@��f�O�*+�[A���E�|��_��<���B gA�!P�v����I-E�@��x�7%���؅S'�b��ܫ����gk�O|���F�D��k">A�;��?xo�f	'�'#�Ef� ,B��'���GaZ�o�E7�>�g�+L�sӃ�e�7�I��r"	.WQ9!����PH5�%]�P��r2C��y��ޏ�q��
T,�$s�;�*\3I�p���F\�b��H�qO���|=m�q	�z�僝e�`n^�Nc�$j��n�
��ڮ0r��T��9mo�&�V�j�$x�}���x	t�1�g>}kq�TvdpVRQ�m-ޮ�:��������y�K�GvP-`��HC2J�
���h�L�SW��Zb�Cv<
r߁���:6s�����ǧha����RGg!�!���W�/�>��;���A>������i褣һ�g�m{�����zk��2�#��k|v5�ol�J0o�L�:�J	�ŀ��d$M�N(�O+��t��4vRm����+������qim$�}�iFs�t*��qI�t�>��LUc�}wX6�m�p�0z�Q3��I�1��`f�D����a�Q��@?�}���_lk���CY/6���<�����B��Y���'� z�Yp�;�l|�E����v"���:��J�X
إB�}$mqX�=����C*�:�~
��.Dv� $+q�bح�������=�RHw|u	�'�"%26�s�+Q������j-�<�NSE�XS۳���H�Gng���ݷ�'��ˊ���X��zB�
"o�+���(�Ja�i	�)�z�Z<=G���餑�(Znݠ����YU�Y/|%���(��Ħ^ᒩ<b ��S��G�]1	�i�����B.@�8+5
����wY���A�B.�q�5���#�s��3A���[�
������?��_��M�m�u��+?�l����O�V��0���Tuw��np������NI�7�+� =Ã�b�3|�ݖ�ǐ�H�$�!8��FN�3%SVm,0?jp<5(��̙K��>@s��j������h�ܰ.�����ӅB�7<��PDT��<r���OY�{�1�i������q�[�㮯ۃ"�a��2���*�W"���\$w��%�[����M s���6n �F�J�q�z�R�ʷ� <�����,�IO��cJ�@#9w�N�6����|�|��0��KHk]��
kw�yw�X&�jN�R��~�.g}�A�������?������hp���4��Z�\�:]�r�Pm�E�a��)��l�a��$<\ƠG��m����#���|�B����)�.]Y��26�a����ϱ�g���o	:L�zڄ�拻0�<��Z� �"�aFڐ�X���6�!r{ɨ�,E-3�
�˶-RN�o���9��A�
LI&0D�i��]h��u�#�+8��j&��2�N������c���P�*l�m���e-ն111AkG�`ˆ1�:#v�����|��߳FS�y�j9}�+�3��M��&��o�ͲOx��/]Xv�g�,^Rb�3}�{`)�_r!��:xu����u���$��i���MA��e�	��4��+
t���?��k>��SU��n�=ھ��u�O i�Ჳ��AJU䥿�a�[O%,5��A����i��1��T�,������m��綟���&JѴ�we��h)/L������=4B,{TAQ�O�kFCdVd��K���]�[���9ڑ㣵Z���?����h3�3N��+E�\x��8�n%I�M�?���Dl44��1��B�����]݃���\� ��������+�MQ�81����AP�,%8'~�x����wM��V}W>�	lP�"�
�	ώ[���MPx�>��� ����U�����HkK`�aP�ނq���t�)��0���������y�0pQN@_9��l�(�( �c����a٫VYN�Ȟ��C�������̇ҋU;��2
�j���m�ȸf���Ɏ��i�D�ز@P����6?�L�qE���T�q�w6c���*?�s��^}��a[4��=,�$B���C��WJ�Zvʋ4g�F�,uozZYL��31+�<n{>�q�/���|�ebI�]E���h�@��J2t�M7�s�I��-�9���aƴ Ç��t�ﳩ3Ժ&�<΄�>�at@_@=`�#�.����G_�>������MM��!�wG3۬�9����2�+��?�r�^vZ6@���a�F5|J%l�g����J1E��3SZ��oƈ�U�弝��#Q��|�L,?Q4�d�tBQ$���j+��p��n��:��H�F)�ϭ��l"_yҭf[bL�AӘ�O�or��7Px�S�<*55���&����C�.��S�]�ԴM�K�<l³��^X'Ҕ�`�d�I��a-�l�ޏ/��a��l�%U?y�$aN�vx֒���ϳU0/��&qHv�n�j��^���5�>����F+X�S�&~��K�����)
F0��إ�
�5Y�~v?�jo��	��LZ6":���e2�O�i�Gl�r��NHѕ����7�4A͞��̛��2�]�
rw�+�dl
;���>Q�A(�[���i��5��i5����E?>�ꢉ�~9��D-WW������`ܝm�ݻ�>���C{��݌�y�+��W������F�_�@/I���"�����EZ0�B�d�X����Mш������K���i��쓖�L��h��i��f�3��U�ؕԞ��s9r</�� q}�Y[��5�\%	<�;�v�'V�T�����̽v��:D�b���tFe�c�Eh?�����8�����(\�7ؠSPsS����:j�/�c"
j����B|�@i�v?�M�P�]������n��Z�W2���j�wt���I�YZZ2f'�@�7몐Q5X��\5�҂�B&��{j
3r)���t6��^Z�/T^�:��cZ�l�G�!gy�W����[[7J4�'�S��A��������Z�\j	�3e��hx���cVz�G��R�����'�+�&��(ء��]Bۻ��^疇���(��crl��7Zۅ��_�8#bE��k:�bEHH;'*�6��8��Oڥ(P�L��8�C9RT�BJD ��&��-nT}e��Q/���g�vt�0I{= ,���pdo��7!�eG	�;5���{˿��9��s�	�f�-?#����t��r�̩��{���'I(QTj܅����߶����f۫�Z<�W������#��g�މ�����������H��%5m�ó�9�s�9��T�.����50��a,ޥ/"�ۥjl����9�@���5ZfE5Pb��q���0��3�߳��eGr����WC�����[�.lI�ee?�����0�y�ݰ�LW��8��q&�cB�~F����k5;������l����p��g��ɱc����:�2)�Lr�N�Ғ�����]�����,���O��a�W�KL���b�Cэ�8e���)�1;	')�6Uky�1΀MUӥ��\����(\�������bعS^�e��
�y�ߡVr��YƲ���q�2Y�m��3��I0a�A��:g�X�����~s?��S�W�_�����︓@�����2b!p��V��"���)47^��"Y �
}OY�f>�Q��Q�,���A�c1�c��
'��^�J�.,z �w�ާ�x3�z-丘����]�t�./;�/��.j��Xn�ё���s	/�W��:{���wH�Ѕ����mwH]����͘P��ϕ"~�-���Ow�����<�Og�W�o��X�4ѽ!��*�!e��ĳ�^?P�M|�N��������Nmy䋎�Y{J�7�9TIzXz(V���P�șф���U���'�$k��l,����*}�[���g"Ĭ���j��/9�{�#��tم�~��,�^�����wr�{��������o�7�	���1�wb%����B\��v�2
�0^��E��Q{�&���5*	����j/UR�� 3A�dPB�/z��u�h��%��9��!�2ס�
��GVW � Y��N�J��4K�w�Y���/Ep�f�W��;?���ȿ��`s|/��G�W]Hr����ѝ'���Ar�'mzh��}zJ������.���F)B��sD��ء�v�I�dU�ݪ��C�����|V"����깿�3V��f��o��h���/��SV��͹��^��}� �s��X��=Uh�Q��=V���F�6Vp����jr�-���0E�⺒��"��^ �>�d:wq>��������.Z�[ς;[-EǠ�o=�9��~P[E)s�}4�v�T�A~xL�](3U�q�oQ�9�鶏���x�0�2r��=�!'OK����B|��Q��ȵYO瑯�gΔ�-�^$ðnT�j����Ya�=9|/��d��_�K����������`Ff&uTf�iU2����'0zd�2h-+c�lM�wC��:�%�����KkT������>
�6��)+8��3w$�/�2?��U���eIP.m��}�,����7])$�8n!o�<�rK�XW��1*�"p�����A���QmV��������!�_�V$(NDaXAK��r�=Mqt]*�gb1d�3~�pU$���F�S.�"���XųO]xbH&E��[�� ���$���py���"ܫ�%tl�Z�1����?q|��#�2��E����x=��(iΝCfb� S)~w�lu��MV���s�>�B�����|���O|��<�)E_�*�M��+���L�kCS|�Z-�':/x
���nۛwG:h?�t�ZLΛ��r�(�1����֌7ӝ�N�(Y��y{��̫�c��©��[��뫰8�a�C!����?�%��B��q��P��۶��M{wM����˨N��n��7�L>.�6�:�
8�c��F����>E�kX8$�ŭ���/��i�o���'JL���#%�ri�����y
�����ihuϘڠٵ�,�UVD���=��Y�E�8�j����ֹ�_�s�q&SDu�-���&�z�(������T�A�ncbm��CuU��d⳧���>��I8��9cͬ�₂H0�8 ��K���b��Q�����Yq�f�k��$�D}r��B�l�i~[�=�Dי�JF��WUmw��߱<�3n�mG5��6A�tʤK>�g#��7yzQ
J�e��M)��8�Y�#�~z���@�<� 6��CU1w��7
�$^���"��5�ٜ3�|���G���q�
*Nz�N�"LD	^yn�	1�Vv��έďث���l1�j�p��aќ�>�o�
�\�صѕ�Y��f��u;��면��{]�q���lYR��1C?�j���Ӹ�=�c�Q�V4랛v,�-�}8�d�<eK�X�4�n<Q�-$�Y�Qh���������7+V��sn���m ��MQH�O���F[~4hK�{�t�C��n?~��m��1^ļ�1I��1��sW�A�/� ��1x%t{{�*އ�ݡ���V����Q�G�P�X�ђ�b<1n���J1���&���-1��?~s���{���O�cf(�+u$����l'v������*��U)��ާ*�G
���G��3�]2���O̥���{��Q`w4n��k�k����E*9T�[��к��R������%gz�9a���W
H�������|����t�]�|(`����5j� ���(�V.�b��B�D�X����W��XiK��<!t&�N����kk�m���eW��)b_v�iMM|�H;��Yc�k���cSS8�k�Aʣ�����M��B�S-ox�!\��C5ZޑpAf���ٵ�����As��k+�.�'��+)��"�Ս���-�4�U0d�4y��L?	��i��xY%��s��bPFV��x���s�1ypo��h+2@8o���D�y�?��R�?�h�z���yr(�K��<���t�@���(f�\,��#�c2�������`̯J�o��[�����>��Ixwn׸��
�;Eu����ƽ(�X�I&�L-S����X�bנp���{��F9��|�6sۉ�Ơ��
�ګ������)d<��m�P����V�����*҇�܋h����.q��3�s�Cv{�b�`���R_Vq�A�'v�1]b%�m�vd�)������ݫꕒ�y=oұ�h�����%�_���W!I���a���J��9\��3�Q�k�W��s2�K%�ȡ_U��JĄ���W�OO�#MJ��Z�TЄ��\3˘���e���Nq���_�<���������(n�Ȧ Q��B�
��亶�����Z�;�6��
x�����|+�&i<4���@���݋�1�~F1�C������#�
�)��HHL���ihR��I1��R"�k�(o���$�I��ڢ�̙!���ۚ�8�9�z�i��*��GI%���h�q�1�4���z�^jj&����=QLa
���,��!%�P�>"�ջᒓn���8��=Mg,Ͳ�I$jg�k�#iCZ��?�~�]Y�.�/��yG��}�I�G����>���l�=a�hJ�+G��Y"i)�l�V�������3���ʢ^6n���m)E�5���fse+^|[�?���&y&`n����x�����zC�VI�IE�x�҇�����2^�l������/}ǔ���_�e�o��E%��b�Y�
���TO΄蠈f�	NH�\9y��܇$�J��;w5+oM�z�|ȓ6�>y*����	8�ĉJ/t����^FO_O��+6ΰ�)��o440C��g��\ND�pWb� T6�:MU�6�^b�{��5�������3�F"`� 	"D$�$����G~��	��<%�P���n9��oE�9��������p��Z"l��1��#�8>��f�qAcK����U�`�b�b�I1�v�T� ��ו�o:��k���o�P�&zէ��T��uG�	�%>��%e�覘��7��^*b���?u�X��:Tb-ӊc�+��g�(M0� ��^��Q̲��!��$����˥�~�������p���&�6CZܓ$�i�'S";�ְ2���İK�7Ǖ�um��Q�w�|~��!�^@/�j���P'Z<Q�ߟP�R3�6[)�;�:�yt��ws�dމ�̲ S�w�%|g���[��Q�ٿ9<JK���sWpK�{�.��^��|��&��T+W*��\냾qG�5`Q`Q���I@0O��i�s;@.�OxK*�O�'�86�z�>�a�it���Ƌk\#��%���?�Ab��M��U<���?X�N��HB2:ZI��5�Bg�0'���A�c����v��]���O��T�
�gƴ#BG��m�5��]a��I�-:�.GO���ö'�Q����1n��͙:����9����]e���Hֺ���vT���f��FGʆ�3;H�9*���-c7���y���N�A�ka�9՚�3x�����D�oV���jE�K�&b��NY�s��=���OUMc��K�!��}��r2��BT&͇��Q\����v��'ܴ�����|�Aú�k���C�vvv:)�F��%k��n�|�Ai�!�J[�A Jrڴ�B#@!��C�@/�T3�R��HB���p]�{�������kବOar#tedj�K�{��M�������xL��YY��}b�ȵ�ܼc*>�r�������� �i����(n���zHf��kVF�
`3�|��x3�?D�W�g�./e�9��z���3�h�O��F>�+|��Sݪ��M[����5�3���]̀��v��a%�r�\��E͂���Y�(�g��i�B�0���.��4l}�h� я�����xz
d���rT�m�(�>�����M#U�ѱ��i���\�X�RF,��t֑������f���׳mܾ��w�9aff����7�0�ٹ&�TY�w,���8���--�3�N�4��JR)d�X�F������f���)��j���0�g�|$yk��e��U�mѪ��@H�>b�Ie�W��R~�R@OQ �4u6��#�W����=M��8�I���sr%���[OM�����0m�w�:�����g��u5W�\�J�����:�å{z��0���_�p�k�T[�	G�p�녷���Ɔ-+V�*Ga�o��]2{�e��1��2�ܔN��}suu���q�zu][i�*�)��+�g]��X�_vܣ���o�0�b෶���3}�9sA��Yi��?��T��>wO5�j���� ;�Y���}�[���	p�}y�E�ȵ�Օ��> ���Q)SJ�+�۔�ⴤ����R �`�|�o=0�%����9�,E��.�߰?�d��)��(���Grt7�QG��8�����R��o�����E=��emD���M�{���L-ط����Z,��l�� <RkZ��Ɉ��]Cܶ���p�'�\ۡY��y�9���q|�ڤq���[���\��RDu:��u��2Y�y���
�:�H��H�3��HR�ͤR!�W��2�Ψ�D͕f�d
�7���^����I����d�K%�UI��R�񈕕Ih4�"F}Zi�%�/��=2ӑ"���h��C6���R-��/�V����X���t� Pm����#|yQ0���C-Y~.U��!,�f���q��r��˪�(�v*h��R��J�`��,�hp�h�X���f&�_u��կЊ��eE�P�|@�ui(7��`g4;-���b�����uA{^`���J��pc�ܡ�8!e�(]F�.��J�hi�/��@����	��֋""mdi�����|s�����")�"\�[����]41&�[pb"�L��'N�rѽ�r>Vm1���W@P��s(D�8ED�*�`t����k�*���H��ElwT�Ŀ�߄:c�R�8��2��GP:T;�������b������ %�� �@��e&�+6�6.R攐�-�JG��@�ܴȥ�pO���+�����NR�c�0��S�,Z;;�m���q�3��
��e t��|�����-]�:9A��z�������_We��֯�����R�^;mD�@o�n�t8Wy-��� �l/I�)��Q��.����7zZ�u�'�/uy�'޲d�l��η��ZVې�K����5��2|��y�u�"�9�q�	�>�l4��]H�"�Z���C�ʫ8�x����o'3������V����B�%�A�2Ú��RĦ~m�Y��N���5�����I>MmۏTp0Y[�9���爊 �a(�5�Ղ_������4�����ʕ���šHGT����"��I�X�>\�z:�v���đU�Y�%�_3~!2Kr�@w=A������i�V������X.uqi��XT�k��0:1�V��1��"g��LFbqpu�G�����?l�,����\ʏ��-s����NJ�ʹ�����t.���a|��S���.�����\����ެw��u���^k����4ѳX��P��g3�ESt9)�����f4).I ����$�K"+��K]"��W�%��Ve�Sڣ3���fn�ԛ�[VuEN���`�s�������3�øs{:������!��H����ju�M�[��8}@%��	���C~��3`����i���Z:y����>��l����r�,m�,9��+*�?}fR�	4:���o��Pm����`go/P+�ZO]��u�#ӣ�v���^�%�m�`I,��u#K���������f+�Y�C�e��5��[d�*H�ZY���b�v�ȧI��6��:K�<+RP�#l�'�ro�L��_�s�ޅ�������V�y��s�e[��G٥]l.	��F��� �YV�l��*�HL��ԁp8>�b�sm�S�y�� qUMM��Hj�����*�9{n"_��gw0��8����/;� ���I��m�Vp�X��Ń�|T|�Y
�������-���OI�����~ooS���H�qDP���!����Ե����MZK�R���133�%�@�>bqm��&�I􍙭��	|�$� m-��`��U����-ˀIW]m"����\���f���Nd�a�msc��k��7J^�2�S�������F9�$Z��%�Q�@�����7���6��*��1ɺdʱ��y�*�b���������Ԋ:��Tc��>���L��E�'n�H߶��{e��~��Ltd@�3�n����{��t����@E��>c�
!���y���G���Ҩ�����_�v��|1X����)J5�����[�����ˉ��d�䐀�����G�?ߺIv��`�a�y]��:���+�\9<P�s�4�b�\4Wa�pڞhֺVSjґ)��1��츨�ƕ//Zъ���� 2��M��3��J��4����>`4WL(��!��Q�#��?��@A�VKK���;���ZM�a#j�D����d������5�7��~ߺ]��U��c�L���&�8g.������ѲT��)��ɽE�r.�-��{�N�Ã'/��S��7D�}ϼ�Ѕ��e�s>� �������:�<��	�{&4����e͍����������1��S��]䑑�����U����w[э�Sw�wFbǎ���щ���?;��gۧ�g{Ct��ޝ����ޣ�nͷ�[W�I�ݢ�5�s<�S�����4��Vk�<_7R�@��qOA�cL�K���N	�2]-� �E9)���cP7��o������ub����v���(��0��	���M��pQڠȅ+��;l��v�bY����U�uD��l�*��ug�S�ϣ=f�80ㆿ�+�1�����Rh���W+fwc��] e�UO^�3F��D�Q3j�HW=澩?|�-���I����W�KL?ȇ��\����wkKHz�;`�Fm_�puMv�~Z�y{�@���>�r|�s��L@z��v8�U�������)�g]�_I=�W��[[[{��tA��a�χ���<�O�I���3�v�Ž��k����G�����8���u�Y�h�����{�����!<rzK�0��r�q5���wg�r3�����������ӎ'�[77�-��L=/ �˹������S��j}W�U����:��{`����/��x��@-�LI�l�T�&ٔb�L��SԾ8ex�4qƊ�5���Xƍs���Ȱ��޳���)n-_�+M�`�Z�⨹���{��N��y��y�j�K����W�`+�:2 �C�4eį��OP��^�����/�)j[~��̣�B�~,�K���V��́��2c��MB�q��}Q�W8n"���5��U�ۺ؋w����!��_��o���?N�ݯ��oW�\�.es6�h�]2�mYR�-��H�qb?�j��\����u?(8��4`߼;2�i�l��ޭ���t\��r��*��w6��i���	_ �z_�%u�?_	=�Kz��y�f��z�E�;���/�o�o�s5���}ӗ�LLL��W>g�;/g�"�"���lf1﹁o�S�o��	�w��!t���q=-�slJ�c�vcX�Y��������(!SYY	9P��KKO�����o� ���������e��>����Xq����s뻟����i���0 zzG�	_�|V�&���6m����~<N��x���&2��.o�rg�[�hs;!�}���m�]� 8�~-�2�q���k�xa��H�F�t>�|mHSx%�<�*�ࠋ<�w��u�#C������ݪ6~�������*s�_��c)Jm���C�z�n);m�����=�0�-�g����,��~ݽ�K���.�aQgC�mMG�Ү9�㺙�u�f��@4q�ۋH��e����;/��d�_]�R��;M�[��|��S ���W������O���힬����y�x�>��4����=��i6�����o��;���}5��_I�꾊�?�Z>�������'�	ݓ��p��[��>k���|lY7��������=|ErD��n$�K�ԑ�Ә��QH2�ɟ���Y��	j7D<��N�Bǻ���7��#��$L��O��~IYu�?hs�@+?�I4��4���$*	A��k���t��L/��P G�ɉ��~�k1_��軣(�9C�bo�2W�A��U��2RF3J"���s�}�1K粆�s���߻k]m��	��R��j`���'�~]�T�J	ǧ���ˉ*`�T��.$.���l�0�^��2�|N�^����^�����	��.����B��Umg�B����G�����g!%��5�T��������Y5��|t_ ̈́�3H����3ܻ�=������� 8����}�T���ԹQ8sP[_����n*������v�*���!G*i:=:�a��Ќ��\� nO4�����:��\�
���,Ξw�Z�.Tt0�7�{Z�=��G��u��;�c�����O�B4�o� 4�^�a๋��e���y���un;�ZZ5�hc�s�9{����=��I>�v���ܝ�1b��CcG�ؑԚ���h��$��{���H��х��}�r�t�����:����=�&����T֋��c;G��m&�F��?l����Mt�]�hl��v�M���pg(t�V>�nܣ�v�����hS�u]s�H�^�}�6<��v���{��t�?	6y%J�7�D��>:���7CÇ��w�`cusg۟�\���F5kź����5o�*8���k�3d>i�]��c
�Ն�S�����wK��׉�!G�Sg�v�h��D�1ND�5��Ll��h�����g�=�?7�8o�P�����l`밐����s�HE�÷w�w�	�e�sK��hU�(�����Q�`��3u�fݲ��I9�i�~���d؃��[;��!�ÿ5��o81e$|���_ ]���H�6�;Ʒ�n���w���� 
�kcc$�ڻ ��6�#<Sꤜ��M'�s|7�xO^Ƿ[W�L��4*.-��E>�6�Vl_1�?A {؟0�٭L���d[-Ísd۽X�40�N�41j�r���7�O4�vS�>�-.���S�~[����4m��n\���s��G�}���u$[��&���~�@z��Q�7��r�o�;��.�[5Y ;A�>�����ng�@��st9���LQ(�||����)c,�>k����8��F�U�E�F�����Q���K�AU&ӭ{;0�ctl���]o?�7Sa��d� C�I���ۻ=���FG�/�:OӢ��3�����_|�R���ZFҹ,��t^>�&P��1F-�);�O��X%NgY_\�l}b�'�ǚ�p���:M��n����}��'{[x�Ҥ"��_оP<_�R��p�eh��S�jZ�Oc=�9�.�b��՝9Kg��f���h�R�w���{��O<���)S�� :�J�B#O���f4��?9�Wd�K�X�����^:�xQI��r��֦��y��=�e��e �7ƨ8�"�)�m,�d��/iQ/5���n
1p?dD���>����O-�}�B�J�:9���)�Et]"����� Z��$�d��1��.���ܪiř#��@���L)���� ���#��d���!X\_7���U�#�Dq���ײ������5Z��1я�ɵ��3���mm���X���_9 @���}n��3�~?+T#��p�md�>���� u2�OA�m��5;��+хO�<��E��⮽�"*40C�x��2!-x0��Y�}[#t�{�Vi��� �Iu�ݽ�<Ê,�t������EB�x��{`����%dH��\*�>���YU��[j��pm��=�N���,�W�4;��Lv]�?]�wSA��igqQ�2�t�I_OP����W�(!�%�����+�i�Z��#e�0���%�p4.��!��%�"�����]��:���X�f�=\�̛��h���{�M��W��sל�D
`�����Cbׯ�gЌ�W4%� 0	�MQ�qnr(sk�[}<N[z�v,�f\�������Jf�*"�׉���ޔA} �!\��^��9_7�K5=M��-��\�w���B��a��!11��>-G����@������M>HI�5�3*�� ~o��B�H(pa^���q9�íb��TVT����hJH�?��2(����n�Kp��%��www�����Np������W�?��t��K�W�)V�����yq��&Q7��b� Cm��A쫹v��2�Rs�kU�c��W+و�~n����A
�	���.�k�o���j���*�`a�e fw�A��q�hhP��0N�m�?jo=��L�ݑx]�IE�1�)U���ڐ,6��I�r���S�i`��4���柞B�DL��ؿ�JZƗ;v}}=S�S3UP+��W�M:�=����DJ|�PJ��4�K�M�qr��Tu��;��$l<��$�oPb��i�����|��S��u6.	��H���XK�M�$�~8���(Rq�ڠ;�{����9K -�b/�V<
HMMGW7�a�e�yu��J���5�a�G55��!�6�2T8�ճ�
2i�mv���?�ۚ��i�u�aw�
���B�c�l�}74+����[�b_�lEnQ�������<K�a�Z
	n-� �Z�Ml�h���{v��x=� :�sW�%�&wb���F�����LU4�_�+Ϊ����r��N��o�'?3����#��W�c\�Bݞ�P����x;��v%�M/~[���$Q
`����cMA��r"jˁe1@'B�8�l��,����2_HorƱqB=��iV�zN�6��ˇ	���d�������Ȝ��T�X��Ԧ�)��̉�&2��A���cT��_8R��� ���I�'�UU��E��c�(��{b��B?Å����yz�����vvlU�C�Х�ۋP"���#,�0���DB
H@K��>x:�T!��ǤK٫o�����{#?�߇_>�`�J*��pe���G�
��p0bzX@d}@��Z(�%g��	��d��3�A�{��T(��J���_�.�K_U~�r���y�	�qv�xЕ�֍�/��"�Vo8��>.o^cQ��,�ni_��T!��Fú�A�찑ҁF�}��cF��y%A*�q��2������(d���3҈R��H�c���x��z��ch
U՘��>�:��_0��,#���x����tR�3}��`�J����ΊEwS���\X� ��h97�<�u��V�!���Ab��Cu��T��a5�����+x�{!���Ԫd P�����Ϊ���E�A�6�ER��a�H���Z���r�"��?�}�j�>���6�Y�i��).�1J�5����e_D��$R)(L�&X�mo'�	�)zL��O��i3����
��r�� |�C�Q"H��>p�nDgc*3��3�g/���,�9�r h��6?e��ڈ~'Q$=��^�L�C�Z0��@�#��=�u��C�Ze�)@#E���9��뀈�Ė>J�L���U��� �\�)� �n�a%�d���*�~6��MX)z����-�!���a��U�io��>(��^$0�i�����^�o+��v���4ݼ�6��	O
�<�Όr�B$��KG1]�i�u�]K�R�V���d��P�$�_D�����]�@ƆGŖ�K���ff��t���r�O30�][���0�_n����i�>rR>?�P ��rk�º�"��Q�n��N���K���H�p�a/�eh%���)!���#�4�ap%H0�{�ctp-2B�����l9��r��L�Gb];�!����eY�n?;������,�A��W̩�@U��kJ� �LWCy�*kS.8i�ng�1d�g28GE�S�������2�&�O�k���7��':�\y�Q�z�H�_!u�[�т�g����g*����c��q������@vøRW��w|��[^�3���8&�,,��K�i�&�7������E=�LZ<�?z�H��%>V��9�S9��S�|�pW���خE6����JNvu䓳̻5(����o�(\4�Č��H4�8"����<R0�jc�=�����t,���z�����)��9���iC��fվA�xi�ML265�K��G7�>��i�f�'�������7�|�BN��PE�����ʊ�1��L��+�Lm�K�i����]��|̓��l�nM����Ru�fNH�/pd��Hsߌz��1Ĉ��d�%o5��A��4�ˊn)�K�(/�����K�b�>N�7sR#Ir���o��\l�V�N��}4�ph���?ɑu����y�V��a�jzq�Z��S�HxP�ȡ���kQ�\)i@�+I�·8��}�=���>�5F�^�9j��˕˞�N	>:��x��Z�boY�~��C$dT`h�#�t׺��"r��o}��Ӎg����<�(7�����{�a�,�5�N��2us;:��enǴLsy�G����|w�T���Hq�M���5[�-|�k	<2��G��U�Y���k���w��AƣZ�<D�nA�u����c�rRk5���K̓�F��
�zu]��6�|��2|t��<�1&h�TH � ���� =�9�L^4���-|!F����4w<1�{����Bp���!'&`J����gӼޓ�/㦏���K�� �.9�@��*���9��q}�vٍ�����ł�׽z�Ͷ�7��cz��.�H,r<Õ-�7j�-Ny��;�b�v���n��J��nh�PM��pJ����OUd� ��ɽ/���L�n����r�n3���+�W��P�s+�V�J���L�"~SR|X������L&*�9���c��C8AZ?�.B��ԭ���z�NWn+~�l~~��c��8�*�Q�Hڒ��2��zIqrJ�Q�zC����z��2�PY��ٵagP4�|Oz����"!�?%n���/z�ۂx;sF�6ѐ���\l6r<H���"�����%�_
TƸ�y�%�Ӡ�K�!K�����Cy�ʨ�b��2�ˡ[tT��k\���E���~�?[�grU"LrM���A��J
��U罾��]G�c,�\��T�}�I�'�V�0"��gFp~�'
ݦ����vK�ֳ���Ͼ������Φ�P�}I{쥀��v?f��|�uH��b}�&��#$�>����`].�Do壩)�K�R� �Ӏ�y�{C��6i��� ��0���{O���Z�aM���L�)��@��f�]����TM���C�c�b<(ž$��!y���&�EO����NL$d(ؠ.�86�EG��T Fʂ_�gI֭3:/#��z����i��0�ב�b�k�.}��p�����zg������E���OOW�VW��c������&x��u+ˀ�����}_���#��]ߔBzN<�U�u��Hi���#X]�٤�h�<�绺Z�8	~ػ�V�Ⱦ:`�<�Q��#��n a��卩p�wi sX��ټ�K����a���o�%c�/srS��#`�[�o��r���Eҋ==sv>���1J��Ds��#>���m������a���e.{'A��i�&u���ff7�A�x�w�ܾnZ������d=,�^[և_�e����ipAw�'v��ټ��ד�)a��i�xqV\�EJ���P���H�I��#7k-�CT����9�o�4xq��_V��C��]}�C��G�` ��hX��&# %�r<oʓ�P�4�����B�b��=����	�l��//�h�ULI"�x�gs�W~k�0��=5�-R���uN����wUk��^t�u,��BҏfǷ~�A�/�KDM���Mj}��r���*i�B�ͺ�Aq�4s�D�6R����-��Bz���N�6�u�V4�4���)�I�J�B>���3�B���0U���S�MA�9vs_	�]����2��"0��k����%e�?.�S)�E'z��.�H�;5멞^4�@9�v��OQO+��$��aS7���E=���^�`�):��F���}��L"`V}��O� �7�٭���뀺(��2]���~7w�b���i4�����ͪ�����;d��G<�p��O��iǎ�O�ݵ���|���giU8�����<zڭ3�ύ�=|�M�]��<
1�	�Dy�WML��Z3O�夨��/����w�:�-j�6�&l�j�d�+�����7�
)
X��C^2{h���x�D�ܔ����3�#���p��e�g�S�R�S�A0�K7Tӟ��]���ۢ "�0ctKp��q��exͮ��z1��L2�z�ݐu�aF!��]����ګ���eMR��d%��n�����B����~Ӎ���B��N�.��Dc+
�	���'��6H9�\�&�/�@�C.m�%^N;k�>dQ��~���U��srr2a�?=;�I��D�寞Cin��QD*�%�5a[`�/SA`�Q�ͦ��7���lB`�AԱJ��B�����oQ�G�@e�{8��?@L�s��3p[_���#��#�˅��lj!��M'�$�(oX���.����f������)xZ�@���WaJ�c�g���|'��P��j���#�+L3:q����U�V�B�B(y.�������B�/��bu��rE}G4v� �������q�R�GS'��sfj�@������G��誮;h/�K�h����$����O�@�2�(䡝s{���fe�w�����k�hpR��=�S���y4"R�X
� m�i���4��TQh��R�9R�G�������9�E��0uE�r��ͱ%s��,*�|�u|}��c+x��[�W�� 3��t���>���[����v������0�E5|��������}�sAKS�-b"�W����Y�_P����?pqyY��=-2���Ӥa���ٻ�{�)�jI<o}�eu6ge�.�?��>#lI��N��ɸ�o���a�fHB��_�P��vww���B��=gv+6.	_ ��-�A��G�����S{�y�\��`G�Uϖ���4;%0�$ns|�v��m����3��X��=���y��ƍ���~�b�8��(1_�q^��J�`e='���#��²���ŷ:(�`��'�r��Q�Jq �
���2Q��G�<��#.61��}H�:��$zDd
?q6L�p�ݦ��y&��t�3���fgA���x.F���+��]��h�Z;_[S����ɵ��Δ9�n��n��F��)��C�&���@O���yh��������4��ӞnQ�Nܚyx�5���+(Dppp����7���U���#�{z������wN� u�̧l���-�����oJD:�U�K
��GUd]�9���4�f��(n%k.���!�{��y����,-e�ώ�q��+�7W(�����_pW�5e/h�㈃K�G�t�7�S1�Z�^yWVVꛚ �-"�����p��"�*P����h��?z�����'j�8eC�;b����Q ��J��|����̜}����U�>���YY�eݡ=7Wvzz�����,V����d�$]6�q����[��J��Y i��z������G@�#���I�hrg�=^QG���
B-��zJ��kjq.uI6�W�.Ob��� t���(*�SbѪ��v�����ʪu0�l�(niii��w��������~[��'�>宎�%��S�}^kU?=[�o@�l�X������h��O\��n`F(�glJI�T�H����{Y�~;�|
��o�Q���uҝ�<�<���g^��ӊAq�� ��.��6� MC��J�Z�p�4���&猌���V�X�Ҁ�d��ĉ��Ή�e����IFL����ڸ���/���Op^U��11�����˨�[�H}���A�W 閮���};A���V���m��}?�2[�H\ �_�뛟���ȉ��C���#�O������8xM��Μ£f����j���q��hz�q��%i1��1�|f�QM���r"����R1�x�
������*�V����]����_d������KaK�ZZ�2��?ݞXTX�W-4�V�����r�*F�`K�dUc����u#�v\7mL�^��i�����ed�{N}�nl�)r<9E�td6� ��#�Ȃ�`�Qy}��A�ݻ}�yVVV����Xc��m;�de�+)��66֐>P�mR��:�����W�hnN\�W��(�߮E��b��@/�Ѷ�.h�N�!��f�����i(I�[��V���=��-���Ĵ�8(7��4���k|�6�K~�k�P�7�7�$����j����j@�������ڲd1:>UK���j%���{��7v���|�����+�C��&�.����"s�M���z�����hΤ����Ҿ��p��w~9�z�ŝ�8�#yc����������D�|�m�����@䦚v� ��R�XqryxK��|UKy%}[WC�ls�DC5��C�ʿ�׾s΀��gw�8�V���H>��'�S�z�����m�{a�6���M��8�h�t���mA�`�&�H]'	l>;����0z1U�V�����D0���%	����G����ok��!Љ;���OO���pT�´FFF�`C��0߲/�]�c��w��z��;O?N�~ȦdR���$���m~0�)��_�Rgn��o�D�f�V��_�TӅ����#c���	�9xK��L�qZ���?��	<#��������B$
�$JJN/��lY��3�*U�fO��V��D���|ʐ9H�� 欽�4P��a�wW�y�c�4a�9>���~�C)�T��ג�N���Ykkͼ�������g\T��f8����i���2h�t��oφ�ρ.m�Y[��Cr��DF�3�4����������j�G����h�����{�2��@���ނƀ��;b�U�����l2��&��p��g��R�����?l�ӻup����Q5��9�2���즥|�'��c��p�T2��l^�@O�¤���#�	��C�"��t�:�c]uu��4ҭ[�Y��O�ϳϔ߿&�6��=p�J�� �*0;%�rY
����8ԑ����FU�8����5M��#d�b9�h�<V6y��)��������N��U��޽�$��K�^�		���ʰk�4f�"11�ɔ1?�B��)/����q!䫖ն�G����s����׍��D�B��M�+�u ����!�Vy♳ �R����Jb�0�����&%����Ώ.r�&��$��֭o,;fz\3��L{���2
ď��L	����b��)'�'?�\2u`��ЦU�mU����]=�,����G*>�A��������Q�!�JK���69�9����������`#U����AA��b��^���W}�y�U(����,����%���&86A�c��ƪj����\�B��iŪQ�m �a)@'�@٠�]58�F��y#�	�P,b�+�qm�Y���F��>�oҲ����@�Yvm�f(�Dg��,��e-w�|��VJ�Z��텪z�$�����3��k,X����B���ؔ��%�!;��lY��W���1���� ==��f*�!��)�g���8����H.�C�^�S�A��S��sC�L0h��f�Y�4�C7��*�]�@|8�'��a:.f�������j��5͐E郧t�6�j2�%����H��ϰ�Z�:����H|p��hz$H���xl�����wq�W���JR�삃�?r��c�!�;?� P�@H��qZ���z8&��z�ᱺ�X�/����aln��u��^N0�^����y�|��5���6i�������މ;�΃o��Z�}1VM��o�C���&n7��ΏBnM+kV�Do\�r���&��]�1���ڈ�������R��m_f`g��UKz�K��|����y]�}����e��3k+Z���:'�#�4ҫn�R_�}�4ӭsf�	��4���Ϛ6��ަv.{&��Ih������G���:�EM5^����M�	�����z��W�o��|؉�9�/�yU��ֱ����l ���e�&>M᭯w+���ۃy�6ʖS�Wh�?�KN4Mz�C�<����~�#�ʃ�3��U��ʿ}3;�!��|/M��]�����iu��)Nt����=�ץ�����E�%t�>���z�0:N������'��o���p��ү���W��8������:2u?�`��m��?�:�"�p�[*�~�\BGW�:6��S���e2�q�����/(���� �.G��r� ��
���L:�s���ن��+^\��_5Dw>._5̸Q�DU�ٱ[�Bd�����n�������w֊Gx$PPX�/��o����r�|��~-�Hʧ���������>#n��L��`���`	�*���e�<�M4>.;��P�)jڹsf
%�k֒��C�����h���.�Q�#�%ԣZڣqM9���#T�ǵa .b0�r�/Z�e%HCc�x��������{�
[0ӎ�V��n.�~�U�2H)vlӲZU�9w?L��lK�q����7�p�9�+�g	b3��)`��Z����Ǖ�uC}}�#+�XJں�q亸��o���S�XV��=	�A�;�|$d��F�{��^���~g�X���2�3+����bH�����q{��z�	�P10����9�p�"=�[�.�|�_2��FmKヺ����]jb��5�a���u��F����Ť��� LY*���n��Z5�qN�s
>��7[���q6��Q0�N�ĸ<���f��|ΐ�nh���@�L��ѡ�健����J�UK!N#�]�������rf�b٤е�H{na�PŇ�z֡ոД��Q�ߒ�10 � J�^+�M��"��3�/��vN�vE�e�YX����� ��J��7^�$�3�I�OEC�����Ҹ�9#�2]��r&<�B��YJ4;=�j�hS~�鸺�&^g�4(���D+z}��xG�>a���.���,R��>;�0Ce�A��r�r�j��1X.Lts��7٣���hI��I��/z��su�����:�BHث���wh�'�>�酡OWj��&��w/������p@�u�����=s:��1��pCY��0ut#��i�/p�5o�W�f[�¥�Ӊ�C�Mwbcn��/̟�
%�W��~���zE��[^���K��l�ֿ�5� ��58�b�4�ڪ9p�� ����`�
P~��GA��� �!���(��+���F � C���P�Y@���FbO�lw��0����m����3?~���+��mG�2����n�h��;O�Hl]��O*"Ӌ�	H���##x���	�Ygg�Ɵ�C��3s���R�/>���2��#c�"ɐ��������VD,��o�O+�/*wP��Wӧ;� ��L[�����r�C���d����,D��F �mn��*�[��㣢���e��Y�D�YAL=�0��b�;�eܲ�[��zAl_����[[7��\�ł'�"���Ơ;�y��5�Y�1KK .Z�g�ā�J���P ��ÑUp78O�M�W�����.�$��R"���gg��M��`��q1	u���i\-n�t�/['�A+B� 'ggx3c�f���q���ꕏ�yk�H}��m~&G�g߫��|�U�cv|T���-�Om�5N4|�y��+�"{Rw���ʊ��Mq������P��B��l���I4��Ý�X�u���K��އ���2�o��|6��2�L�ih�[YE�����N&�~�����\gsrqI�;�u��рi�:-�ooaˬ�:�º�s�s�E*|ߕ{r1�\r������9� &�	�!,N�N�5J�e�C����}������8 s�F�`��|{d�kiq5m�PWח�8��n�o�SJ*�A�W��"G=���4 :��g���� C!��B�hu,B�1�"��YXay�����+g�\��06a�c����4���u�w�o�---�C���0f��]U�"���d��/����A>�Ѩw�y�������x�l��zE��Rл�GV�UZ�����Tp��< �&�X�����/��Y�+'X�*l��ک�<�։��U��)����X5��˥���$&%�"***r����*``���*��c��f�> ��;��j#B/�qΑU$�_���1�����֯�\�q<�9
&9�|L��g��3�r=:�-�'K�J��㔄���?ُ���0-i�F[b�esp�����3r��n��3�\H%�Cd��uP�(��N)`��kL�ē��S�J��vt��W�7� ��3U�љd`�@E�Ka��S�4�|�)�������&���9SN�C
�@�9f
�V��b.��	�W#�)�r{EB�5�X��q�oY1P�"�I��n@�s[��߽-����v��^#W=��ex�u���A��b�9U"�en~��z·B� ��e �k7��5���q����^��݁�]6_mL�[c�����Ѐ|�ԣ;�Ó<m�nc�v������*z��R���YK��c՟?�.XG�T&�y>n$͙%}�	|߰��$�Iٗ�L�\c���[��f���_a�1)�;;�R����)C��r�t[�g6�"��������_�NbI�G6��f����,P̙9b�Q*�Y�T�ߣ���v�9�ѥ����]���D�lL-����\=�F��_�`àK�Y<26:g;�u�����`���5��H��
GmP�P�P�Ymעe3>-C��a�}փy�p�;@��i*+����јUӉ#¡oyEEMc�~��녔_�Lĥ�9?�On�$\����^U�Z?$���T<�<��q%1�(��n�CZ1^Q9�Rq�ݘ��S�o�l /�]v	�.�+bY��j�̾���sδ�-��z����<Ҕ�?|�9r�H���'�ݜp����3/�3�����R^v��cyE��W�����y�H�@]>0�^�h���c>֐vΌ;Z��J�^u�0��%y��&�/�e�/Z�U�����T�`xt~��Z�̕��n�W�۶�qyH8�ǅi�]]��0��~����%_9sB��� �Z�*���S�f�1j�����˹L��o�: _��
z��83��}�Fн�A\�
��%c�aht~�t� ��+�R�%[l'gE	��Z�z(N���BuhjҀ�<�"0����)@Z�u$f�B����X�B� �h);�%-�ƺ0��a��v��]�r�"-/�#/ 	u�%�� �ݕ�H�X�ї���jOS�n�f782Ji%���#񳢕
�����c��;e�.�IH.�ӻ�Ÿ�h%}��D�u�N���w#�R��rrqLl�i,3�lT��FD?
?a�)��>*A+�F���F�QN|f]��pU�xurڰ~�5���`�F���}��F8�����>$""�k��B����N�.����I�,V��wjۉ�:�nn���~����}��,�ଇ�,]5.��_/�����5;�`u1r�Z�02��\�}����O�l>Ŕ���?m�=&�U:��J��tP��`�X�C�Ĭ�dxY2>w���Kf��������U�ژ�9�۪��5	ز)��O#.mb�/@��>�q}��'�q'K�h���a �E�����Qx�+x�h�)�j�eL�QǑ�=��eײ�2���-��X�EǢZ��؎���`+�(^8qk�*�='~�#��0�#����nj
����z�$�����>����F6�ߢ�錨�{��F!���!U	�Zq�8=\��#ɓ]���b)|�O@,��f������k~��6���աY{s�Y�v�An<��欜�ɪp(��&���a(e���l� ��S��'���J#a:zƚ.�A�O5R�o�U��7�R��u-FT�tc�E�XR ���"�a�D�g��<�J�Ǝ������	R�q1Z.��b�BcqmM; �WmIp0�5x��5��β��z��v��8w=ky�
����O��M��V������#�)%��h���ORW�����J���
��O)�cFB+�qKm>찀��I�هEWMsAt�P"qO|�N�`Y���5���Z�*U�`�����i �S��P� ��[�Ǐ���өZ#���w6㔜o��G�+�j�U��6e"m(����+��F���Jq�I̯tjKC}~|]~�ܺ���&띁���4.kr E�@�f�˧�{�/[�}.~BuĨ�=��}}r|y���q��ɾ�����fag(�෈��,^�i��'s̔���ܭ���H�����T(�mbb"3!�����f���G
�� E������߆%Y����ϮRmɰA�4����Q0�sb2����~������z�z~˧�c�iI��a�9���{���Yq�+�_*;:��dҁhr�p��g��.{	?7�Ѧ��篈q�RNut|���f��>��>�؅����%3�!K�)H��Ϭ�tt�J+37�cn~�d��ʩ��J��V�LI��$"���!�G{�odT� -&�y���|�4���.���EW�D��AazM ��cRH���%:�%+C��ȼ�#��ճ��o4���J<�N����VI�x�ܙ�[�se	�ΖZz�f�zN/�>��8����r�O��G�{LPZC4h�=���@��/\V"�#�g��U�r�գ}��c"���?�xg���h"xI�t���ލ|�%	�A�C��k���{p3�r��a]e��1`mVˀ�K[U�~���W��+��&�$ZQ��ؕ�Љ�(B⋲�d�`�|�<+$j�fk-�ҙ es��Jৈ��H���1�!��A\���������Q5uu�$o��GEY�<j��5$�%E��WǼ��q���3��+«+��_��"���%}�8�_�Bw�U4�?��]�E��	�����sN��~��oai���M��Ƿ	�2K5ad�^��[2�Q,���#1pV{��Oke�c��,Bмv��<WD�2�3Q�:_m��-8�����CcX�P	;�&�+�ǚI
8�Ê��HTcR�E�<0�a��b,G����? �_X�\�x����?;��O��:����[����h(��rx�������0����jZZOǩ�WF���X��hV-���]m�4a6g��JY����O�Ǒ8�=���do�ڃM���OJY��w�j���)аVU�r�8��.��׫�֍(R�J@i�>뷳�����t]�պ��e_�)n�#��������b������O�O��!����"[�<w��u���E�M���'<"�M�p i�B�w�>�+5,Z��\@`�UUPu�Õ��ˬ-w�l�]�E@������Ac!Λ9"Em�/�tC?���E׻@.i�Z[��ύ74�>b!
�&������� \�S�V@���㑕p�/����~T�O���P��&���)���(��G@2�"L�P��rfQ�(�2�ǆ0��h)�~�?��SG1��`��nn������q�o�U;�7�<=��#��QPQV��3:#�����ߧ��{�#�4���$��`|���K��A�!Ń����f�-�� ÐX�%�}���\U��-ǋ�������Ut����\�����U�,�����3�E�f��h�.��V����	e?zk(��^�SQ���
�"���]�DnۣiJ���ˌ�'�K����xWΌ
�}%l��s�{3�+��˥��ㄸ)�?im���4����,zja	)�]67e�� -��Y>C2��Y�X;� ���j{����� ������˩��'�>P(�~~Xhd�1$��?��(��e��uu�e%�`�t �qx��E�ᓵt���� (�K��Zʧ䳋��@\
a者�f�(᫑ʓVn�7�R���!(���*��*�����S&��l>Ex�,-<�[���i<��{�D{�����*m�M�&s�y��"��`��4*'֍�<`�Jӥ���L�jPS�~�sH��:&|n���$���v-�;�vw�����*��j�k#�:�2e���@1(�0�(Ʈ��>�9�º=��L�>����p�+Pjc��C�#9�R��Wp(�t�!��θ�Ȗ�r�#�<�C(���i��V����ĭ�G@3O�ų�����1�ԣ���f�#��8�ޕ��M�nM�G�L�# E�����%4ǣ$2�	��Dӻ]�'H����d��x�\*���J��ib�_����d���|!�	��35J�{?:p�������i������ΤW���G�tQ�G�'l�0\�"6��'݂����b�����������"�I�S���i"�x0ƓL�r�X�hvx�3��ㆪc��0n�V�q2S�),1�FL��c%�q�ǻ��:Hon���o�����	���sk<7_�K���z��ݙ:�
���6��#X���yE�l����X�K�$�����zE���ɢ�"��w[mtF�9��0����O��X��z��rЋRA@ŏ�Be�4�9�_�V p���sI��b��dP��T�F��S@�=Bo��<�RS-�h>�]��qo��P*�Z|��	ų�gt(<���yVo\�.� z��u_��2P����;
�� .+������m���q�1�/���d%��1�m�3Ӌ�OB>eg�����Pn����@C0S�jb1+�*�<1���Z�r�?K���aF1�����l����'`Q�6=[�eH��Eχ��ؑ��m���{�j��q�KD����F!��(K���2������W���M �O[�ݝ ,���H�� r��'�m�Xȶ�o�ZH�?"f���$��n�Ϳ���"E��ф@��D
�l�+���f���-��k��,�j
os�Y�1������x�93�(l�O����T�}2Xy[�BɅ��Ц�=�Z`�X��#��ی�)N'P�-���ܓ���v�� ���Ϲb��YT��/�(C�2!=�ԠOd0pd��G��^~mmw�,�X1���=�/�Y�oN"l�emP���63R1����R>���EXi,�N%<��m\|4z���(E?����@�o^�հ5�>N�5<���u���I����ι����B��$���E~��Dtw;��\�mkp�|m!;�m�DC]GG���}B��:���ֲ�.�4R�`��*QE�o��M1D\~yi�g}�X��x�q`��I�J�#4���D1�q��w;��/�a��k�ƈ(F2�ɺj���fX�%�������k}LE��)������{��vY�����,�h=-�4��.5�Ū�⇷n���"]+	a���|LLf�)�����5���'���Hh�rR?_�H�5cjj*%'S��.U>䖛�]�MH�7���h�%�|'S���K����d׃�S���m���E������-!�ȶ{ӭ���jzDV["g��Ȱ�yn,,}.nz��}|7r��+�d�
;��wul��;м�JXt��Y�
U��q�+ӥҖJ���X[��M�C�e�k��Ț����>I�L~:y^d�G㌏�8���f#�X����^<gVm��3a���;��h�F�. D8�ޒ��z]�mMn����\LNF 
�4���V���<�;I���������i׀��� X{*��8�k`@�K����T,��'6��W����7 T��aGE5�6C���\+c�He��Ke̲�Ir���zB���
`(�bÏ�yW���=]��|�i�����ŕ��J���������t�!3�^Sl�ӕ%0�vkƦ7�Ȫ��rE�Fu<��v��>�h-�"�޼��P��x�d�*��%�=>JY9�&[er�?��dn�,--?��c�谢��B���eUD�������1���}�%<T!4 m�$wY�b
iGa*z�+� �8R�뇑�^4��{��n�_Hm�\k��������=>̜�\ٜ�ij�x�yѺ}�j��s����u�)�pG�{��b�1b��\��D!�J�D	t��	�(��0jzzzx&N��;X�nƯ_�Y�6�k�[�F1`��{����姆-�ڋ��t'CJ2�!B
}��%X���jT��U�)�%���O��	�YC���?h��m�q�R-�q2�㭬�P�?�`>���:���a���ub����M�.�c������ ��� ��l����� �$\&ٯQ���ҖM��tK�GGv��Q��}�8D�k����tt	a�_��/��GUn�H�ܒu��~}��!�QֳXm������'O�x���yDT?�:��Z�� ��sr0��,p�'f��a���D/p7�����#C`�9_�qɤ~�~nv� >��U����CuKK(�I���|E�������4�5�o�5��FX��F��q�7g��]����l�lYߔ�&)���d�i|#��R<�j�6���Fklj���B�HEU�Z����-����I؎��*/����,��vm�=A�!�f3i{�?e�������aP��➛Aa�;D�TA."b��5S&h|l��7� ���u�t/w�[n����7�DK�2�~H6b�f�������0u��+E+}��eV?�Gcy����X�A�궶p����RB��eG�j����jq�����Q�⮭�M'"g��� ��h�ʰ(��kb��Ap�!��A@�A:��Ni����F�[@�A��ޙ��y��e�k���}�Zk��ظ���a�a��ӫ�Gt������h���?�;�?d�?���j|�{{ ��}g� �L�����>J�Y�;���RSGgng�J����F���_M��a�yl6��l���������?~-�Li<�L�{����-���8<��Y���h>�*G��Ij�H*6|"�|a����\��y��Q���A�D���U����/�����_\]{��fg�-/V�ܶ��~&����۵`�5|�s�`�������n̿~�ᠣ����J��h��B����̅�V���t=}����+��^�Xq���;B~�=�y�Swr�#5�sd�kAUL.y����~��B,�Ŋ�UT�� �K5�y�����U�Q��/$Ϥo�F@�P�nVs���
�EDD�7O޿`��Jh��aJQ$srF|��w������ׯ[k�=({���p%��]�!ja�����Ua�z"�b�qi�xzdL�"&!1�"�+`�%���=���搛5_
��UQ��"�_~����M��~���3�q�B���O�l8W��GG��sSz�;�x����̒��`&���������0-�SG:�Ҡϧ?���5�A[���l�@��O�o>z��ڕ�L��D1j;���c���m8CS��U����W��M�[:��h����ǝ܍
�)q�h������J�ھKqe�br'M�S�/[to��(p�[6iGcap��^Y��P_+����w��9��j�j�h�vF_�V���������*22�-�w����am�#��*v, �0xP',�~\�[<=K�:@x� F��:�P s�v���xrRì|/($��F,~�̴s�@��Wa��$/�����p�ˮrIH.a`1�:�}���E��/����������� )C�r�[�����F�M�Yߝh�ÿ*����>5t�����9�eN��j��Wy��DD@��-1X��j�r��RLD�Ӳ�O��-�5CS[[�h�h��Q$��%���������P�@&���e*�[1��e�dɅ����(��#�*� ���6�2�T�?�a��E��A_\�u��W/���XaSvt)�'e!�c��;�������ϙ�tʝ���>k�"ng��\��nY���U̊�[C� .B��'��璊��Bk⧝�2%Fp�������ݧQ��G�-���Y*%}P)@��4��gTġ��C&�nֻJ@릊��yG6ԚCc^��y��]+�
�%��=*d31�� �N�������}���E�t�*���]���t�45qW��~��T�l�sc���������BjԦ��o�=i%�x���\1�3��?8��̱�T��3|Ok���Z0��Z��Gnbb⺆ځ��SX@^��_�NN6H����Xf3�}u�
��B$�&�eQ�DZ��	=S�P#M$zQ� �j��!�Hn�p�\�V����(<7�Beq���i��0��/������7�U=�X"�-����{86L	v��^�]�3����n�'*�~�w�˯�����ј�,���|ԕ�J��ܑ��4��|wa������oKw4��y$?���Z3g�r�����o�пB���'}A����~%<%�j���}m�6�S�W�&뛻8�u�e����~O�i��og�>(�EI�mj�P�4D�R�>�'e��sRSr �(ӌ�7�duH�le}�" �� ?��׷/��S�����S��L��ZF�x�Rj�J���Lh>p����$RPN+�2�uUUi�eɓ	?�3�n���ꢥCJ��6�jAU�W��j�!��d42�"q���;�A���w���5œ#���E�
��
k;"�zs��s�Tr��A�~b�0QUF�����ϵ��Ͻ>W&���K
 ����M��vo��ޥ�v^�{�C�����/S'�k)�F9��P�8����l��\@h���<�O[_����£� I�b�ލІ�鴺�X�b�L�yI"��	$P��ֶO��L��#>o��j ߤ�J��Đ��-���Z?�4��I;N"/a䪤�t������h�pUZCo��b�<ʛ����@�yc����2�� �"�B|͆g��� ��=^	�����c��1�y�Wwΐ�$,�mR��o٩3�W{ЋO�+£�J��NNU���̈̆��w�������T�A���I��}/�M=�W�%[{�}w��{�q{d!�=uGC`������q홮�<�~�g�3�H���@RJ�Ĥ�1�b_m��/�|j�� Z>W�7�I���G�^�J7q(f�d�L�v��v�`|9�= ��+&
	���<�:�M�P=�S6�-�YewP�'�.�ˇ0��Y�Gcy�Z���|S��*ϩd���g��P��F��"�$d#2j�K��<6�M��PŲȒ�r���C�վ�S�ٟ�v��F$>C,wM�bG�Hw��>5��~sd�S�k��0����ť�[�6t�A�D�Fp�lmqso��!�����#x�o�x�"�D���amw���;Z��X8�I�6�M�ɢ(q��:p��?�B]SS�'.\�Xr�i�h�'�&��D>�x?��{ �p�俯gm�Wq8ҟ��6<�X��"m[Ic�N��5G�"�nX�!1G���u�vMpί�]Z����?�J�S���5s��rCv��MGH?B������j�Me+`(�Vٝ�!��:�Ok�8�^h�DJ��	�e�;ѫ\��e6��*��"L*��ϝdl�DZ%'?��vNW �ݶpᏎq��
�ψ"���]}�^�Q4X.HSН���f�B�Լop{��%1�R6@f�19xI�N����}��bl�[p��NKՑn{�_ή�Qn�٘Un����F����jO-���	����3oJ����L���Re@y��-�,Sm��>��n8�ZeX�)�k&�Ҩy���|�@��j��G��m�ܾ!۟���"K.2�ƧU�	�#�g�N_������%�[�
����*߲8Q�h�s�K#�F�;@�k���8�i�s�%��e�.�ǌ�h��g����b��+cI"�g�}4Q��"㶱?-h�{MGV�8ϒ�)��hM��W"綾|e���cD2�{�Q8��241A5x����U5,�p��p<�.6��a�@�vX݂H�a������ق�����Xs�mLf�G� �ʣg�ش��	MV�5	���{�2p�
�T��I ��&���-�f�&4�����c���A!&���L�ݵ8�F�ni�� �C�
|SW�p�\�6;^[�]]{�a�����lӯBL�	����C(�fl�D�,����:����#���>fKi�$�����K�1��!���1&��7u]]1mO��r��u/�6Yv��4#�@��>��n�9l�
8� �w�K/��]�����V�c2���քe�� M�[��N��P�3���"�G�Q�Z�튕Me�G*��H�R����+t!�6��g�qP���9BL�����D0����[ ���'�yk��!�����Z.�l�&y�&;D� Y���G�g:���+�� ��*�]T�����?�㝅A��QV��f�4jϯ�⚹�vDS*zP	[c�������|�����J�ì��I�$[�B��PIX$<��1|	���M�JC�1&U55��9���;��?��|Oo�>v���5�����#O�>�Q̩G���u��8d�����۪y ���>:��wW��j=�������]t�Yjpd��<N	#����t�sI�^/�[=��qi-�S�o�H�d� �	�r������D`P�y�K�[��H<���.>�,i��98��%�" l�}���[��hT" �'�����K�ð�q?!��U$6r\�^q���OM\r�.zAFa�ٯ�*>o�z_�m �濑����9	vL�������zA� ��t��B\�P���hʴ�
�=K
�x��X�`P&��Pi����з�˕��L[�ͽZ?��-l<���㶉	g������j�$��>�v�]h�E�J5���^�eu��w^&��U���E���{��88p���po���:})������"�m/����nsNh�#�t��&�����w�(FZ�k�7��4Ƒ�+�
?(C� 9{�	 e�|��D���O��Mث�VT�%�}�_3\��'}�c"iΌ�Q�X���o��/�
A)��fys��m��U�5�A>��bX�}�Z�S�����C�R�W%���(�o���=n��"w����#���t��K��P��m�Xe�a� �r���a�YѼ�19��]�u�ba5�{�f[[[yBS�9�,Ӽ�4���?Sc���EVI�0�7!�5EVX�iVt���%UH_����q�V7�/����5_��p���k�[fV�Oq���)��?F�$��J�K���_�{g4c Y��}]�fi�����>lF�����U*���7A^�D,PJp��.Q��S�`tm�U���.�"����O��Bu��v����?WV��.�L���f�u+�D_Ȧ�f[�$�}�-��h�DKϨ��~1�,r�:�q�.1+Ǯ��gHg���[�>�_on���d����]!�h_�q��.,.#�m�9>��׼�f�� )#�����O�X��WNo6�u��mW�N�3��+���;U�_P&�	�֡ ��<�*;���ս��g����Q'F?}ɱU�7����`�z얕�pM��a�b@�,��)���.�C�Ȕ��(��Gu��<�LMP��	Hր��vq_x�d_���b���"vz�vfI4��t5����Sq�;�Di=cJѼw�c��e����E�%����G
T�'�8�d�6Y(��
-d)`��N~����)�j�?~i�HAV�X �vnB<�[��
˲҇eͮ�J�z���!�����9���Ff�ҹ^�6��g[�SK�9�]��][ԧ���< i�\�/���o8�1��:E�Z�Φv���sP3/�J�����şU~�c!���N���F����3�e�����X��\��XC�w�n�!������`��@��n�-�,㳗[��|2�ZD����	��Q��Fm� ���
]��.m��a��v-"��5[�\d}�A�\�N�r���p� fi�3�-�=�ttt�.�-f�Z�އZ����l��/�\�Сisc��i��� ��4_��E Qb�W�Nk�I�C?7$4��&lZ:�8��,�DK��]���]�a�#��^?���FX���%��(���Pl�]zn�ؒ�<�(�)��;C49�,�!�"[v�hl,�wφ�o&q��A�1���� �=}��ɂg���Ƒ8�|-Dz#5KČ� ��w9O�W��]F��ؙJ��*OF5z{v�������%C���$)��;�*�&�|uabIU�Λ�[e��%�|9���8%�]���Ϧq�LSڏ��>l�=�����B�6\�M4��U�R�l�S�=4RȎ<�R�) �N��\pVQd����{e��B׮��/�e
Cq�*�]{�mՈ�����ܙ=��>��t��@,0(T/m�� �$��{�����I$f�D]nN���w��A�}�R �(m
9NQ�C62\�J��j���� Q�#��7�V�S-�~�-;���p�(t�i��p��^[z���ǆ��C���ѱ1�o�äI͏9W����o�����P�$žɗ-����n����t���7��a��Gc�u��S:yOo{�¥C��F�������}�G�g�뽓�['���jFjh�g�<e��RsD5�T@�l���YV�%uu��a8m�5��J�k�7�
�p����\E��G&�Ȍ���n�k�:f鑈��R�������+K�=����k���m9��X�aɟ�Ã.F�Wx�n��+5�geY��C<��/5��-�P�0S��5Ny�q�r�@$���^p0Z���7h"��z��bix�����{~Y�@���^�(X�NG˶|�ܮ�r�c̖T(��̣ٵ�km�����uT��$���v�������7=�T���S��V	���_p��;S��cT��������Q�S�>���9�D�|r"��h�	���l3*��G���l�����Ut(�x��L����W�|�O�f��M6O�AFr{��|�����fIĞ��Z�eq�ж���	��o��\DH�����YX�¶:�F��z��EO���;d8���)rA g��[c[@��:yb	�����b��+�0���zr��e��B�r�y#f"�
�0���H7B�՗7�lAWV����X�"��^��sY�}䓞-��3k:p��N��ϩG��_���"mD�M'��_�ӣ名D�2�����O�C#>��n,B�o�H@dR(�R�P遀�8�p�f\��&bJ��?ifL#jT��!?��sh����l�{3�C=j��X'$,m�+���;���!L���[tg���!c�"y�7��e��g��'��C��lG����!���D��I�l]�L���
��-Ġd �כ��0.za(N����Լ9��7���(�$q�Y��S���C�C�="q��3�6�<[��bq��4�����%��sv���s��{��^W3�̶jN�P�T��s�� ڡ����@��1�M,���Z�z�C40�g�'>0��S��~���%�c�3顖�(���.����S�_���c쵼�*P?����\���R'z�j}�9��h��p�4�k���;��e\�]݇/�ri�������\����W�̻��e����:0�a�JD���R`ځaN
ۿ����L�>�/�O�RA���MCͥ8�pB�s���?w�֏�G�HH����[ɩ#	��}��'�{"��6�.m�=�U��R*�*T��77N0*�3gi]�4�)���p��~�5I��Yƌ��?�f)�U��^�R��$#������?������G5�����Q�R���zMoTi%0ee��?���{pp�?T'Q�>�mkJ�$��"?�,X��ȶFJk
�k��V��>��8"CQ)�,�3i�%oD��c(ItK�*ȵR�.8(���*Jj�-��x���s}+}Ye2F�z�l %=~U���	~Z�A�ce1������2J~���u����-��k�15��0��#[u�/�l*>��q鮽��Ѥ3{G�%�Kz�=��'S�-'t,�u����>�T("�E�f��H��B�1��g���/�k|R���؞��py9�p3�B%�rL��Z-�����^VB�Bk�u���J��1I?���� ��i���{ޚ�hl���=r����Q�Y��|�8A�i%�"�����3�&ҍ�ih�+�v�ݭ����������֫�D�0�6��BcW�ԥR�:��S�
.:�D��͖��{N�P }��27��OV`�*f��҄����ǘ���I.x7����{�z�a!�� x������B���uR�3V�Ea�0릊�X����Λߞ`MK�?d���"�}8�Gd�;;�}�c���Y�z�]oy��ɥ��[�(�A�v�D�f�T͍�`�J���c!�ɉ�^�x��1�^��g�i`)&�����d�2�6<к�;���Z��4P�ŏfT�^�e��x�� �-/H��m��ݮ�>pCk'���zZʳva�a]evM�F\�S��QٙP��x���+�F�\����^Ȉk"�X���������?�*˥�y ��]^8�K���W4�J���/�����5�I|���+B��[m�<����H	��BjH����A�<򆫎\7B��A��h�*�s���MBfmE�Tq~9+�_xP�Z����������vȤ"���/V�I�3C���KۿnL�%��5�=A DNrp}�^����|�t���}X�џ!���>���{�n�n�X�����t�Jx]w?��^<_r�%kք*o�Q��ya��{9�UE0���DMե�"M��Kb�B�"�1[\f�ũ���K�p�
W�->a:-v��ݑpD�a@7��v����H/9�uw�jW����q�a�h����(_�C����mUAQB�G�
�ٰL��g�Xc~˪���0�׺�}g��E�r�D.A Y�h��u������"�4��kX��wh�6���g��w�t��?&���Щ��^)�
`�g2
�w!�P� 	�^��d���R��������~�c}@���ScF��l��lC�9a� ��)�t�SU������֐�����+�4>�6ˡ���'M=}�W�J���`�H�~��D���J�!���r�W��?��8�=e}X�������-�Z������T 6��T��3�

��B7EH ���$:2�����!O��x2W�5=�E�r]�N�AՑ�<�Y��w�ֿ��M�Ʊ��|���~6d�4�d��u,d�W��q�m<�c�e��7�ec���[��w>�ϷB� UPOPT����^�V�JlIt9v�9.4NgJ�^\-�Q^�2��ITM�Q�&�:��V)�����d�:�v�i/�0L�=��u�`!�8�R��"ݞ:�j��m��H��H*Y�#W~` R�i�́O�?�f������&VZ)>���Jϊ	8�`�?:��Fc�-rL�*��U�����%W�i�-���'� H_D:@�Y��i��a޲%T���	(ʃ�R�q��Z�S��_,�=O?�I�a�-@j�d˧i��7�%"���CFg�M�ଊ�/�h����t!�_=v�FH�[ʿ�L�
������s�|]�efeUL���'
nl�Yc������H$<���^�A����֚���+��_�3������X�E=ޏͲSg�Bc��j?�͞,gS+��7���2&ER�(,0���0�l^ŲZ�5�k�w�|�ѯ�յ����f�L��e$������R&������OL74�j�j��Ot�6gJ��	:�0*4Z�s�E��h���߾�z�����G���
T�,M�_LO��Y��y�zް���5Nm:��C�:�t�1A�B�v�su�Cŗw��=���^�:�J��Q�Wz�AI�_��=���c4�xh�~`�G�G==�i;���9xa�z\3���`�>����'_ K�U󾛲� ��3&t�3���X��>7$Pb�5x���a��`�tl7$�������xH[YV����������d�$� %�\�Io��������r�@��I[|L?$��ʨ��\��JLL�T�z��HB*���κ����1A��g~�~�7b����lllz�pt[�ّt	�خ�׵ t����V	���j=1��F�c�MUm�X�R��Z)J:KI����I���O��b&_y��ӓ ϻw��x�Hؑ�e�+�àl�ε�m�p�ҷ�9E�q1)�Ԩ�sJ p���� ���sI��"���A�*n&(�P��`�k�����ڋ1��P9���3��v;B�N~!"�9��7��LLu���D������>��sU�9$O�D�v%��6�,�9�*U+2�I��Md�M�x2�e�aR�O��1P�p����y����$ʠ���Mw��--";�{�X^�5����긅f�N��#Z� n�9FR&�0mK9�NF� Ȳ��NV�� Շ�����d0�J@��� tKn�:�@RBIh����9h�|��m�qn��d9��d}KK��.���RWH$�d��l�c��$�8�!A�2�P�< I�p�1��g������MK�mܟeF��#£N5�[.��:O��o���c�" �����R�Hv��N�P�N#� P[
	cVdT٠�V�!T$�_���ݚ��$n��k�Ӈ����n}B��v6vX0�b��uА�'�$�K�PK0�F< w��M�6,�����8[3`O���Z(k���/�o��/���Q��IFU�� ;����蓘(.��o��R��=��y0.A<�dX�>����D��Bz;��KG]�k�ر��:��ꍝ~8C��ŗ\���0'��vX��<��*����#1�A����<��T�B��:^�2F����Ğ墭Jݹ���Q��+TE"	{F%r>5e�eaF���i�wD��r�另4ܤ�1�eH.�H����`�R� ���|�c��̛�p��N+����+�}V�J�=��:��%�7�bi��������h��ذSYu%�Ѐ�����|/{?&0�7�5>���~�럋�� ��)�rPW�D����o۲� ��*�@�P_�u��v������
'Oq�X|���i����ŹN��A��f{�U��v�z��L�Q�k#ŵ}�G<c�겂(q���8�U۱o/.Ȓ{�F슬2@H�}h?ݟ����p$7b��~�T劥��%+����4ƧU�J7�^�l�4@*W�!�8�ǅ��]������	��R�3?��?�WGg9�W�G��@l��~��5R��sɵ�D�;��vF-�Mp���>/˝�%��r�)r���C�Y������љs]��|y1d�bdhff&��2����}�(z���n3�%|J7:Fr<;�~:�]ν���2/Q� �0�S�/�ׁ\��0��\�=�� &J���,��@9�����ӌH��Niג��_�p0�\�D1���B�ɜ�`���IW��x�;c݄ha �|�s,�!���J% �%�,R!�7��s�6}�;;*YӬCҏf��
�H$"�]�c�<�릐y%y*͘�C`���@X҂��� ��`�H�dpc�GFOǔ-��6sr��h@d�l�waOD����B�E�� �ˇ�м�;�W�
V��a(lӢ�'�.9��ڃ�F�&2����v\wܦ��B����E���! ��[�����M�P����h���z�`r�RiҽjZ_�F�F
��/
t{�(�;��O�x3�B3��H����_�ގg��#��/�}y�`�9�p$�G��N�(i�S����Z�t��t�������+�~0�����D����7y�˫8�8�"�	�A�m�E� (�,(�l�&=�y�Ɍ�<�\�cR,N`�4��5:��mȆ�_�5�|��G)�N	��ɝ�^���_�B�k�����9�0�L8Yb���sD-j��@R�� Su_�|�V�r^&^l��G[���F>F�˧�pr��Xq�:B>�Az`>0"Ic��*!V�S9v��>�����,�n0�g�_��$�ˉT����BbS~4%$Rڽk@*�j�n`\ɼ\<E���y���ś��Zr#^e�)F~O+��D6�4��.��xI�M9s��u�.T�D�"�`5��7��8Wj��������F�\Q��Ѓ�y4;ʤ�H�ֶ��{�{��z�p����h�<�5��l��ևS
��W47*T8"���/j��m��A��,{{|���g��Ɲ2��"�?����#�Dh6C����	��=���ZTF9�X�xGȊ�Ñ���l@z3$K�Ĥ�B(�j�m2N�L�����#+��jH��	胆X�*S=,[���}!�"
�����R4H�l�[�,r����,��$
�=��di>�72�������t^� ��Γ��.M�G~YBA殠�E��i�H��6:�� �6H�{yQEr�>&Ф�����(����H����֛6�b�-�K�������7�/T?t1�!�ư����ͦѡ�����,��]O-)�5�JA[m����\�O�	�E�S�'η�kwپm_(���26욅����e��Ĺ�9�����AQ�Q�r�/�O��ER��(L����$���20����Xc��и���N���pP�a3��3t�S��Gw���SwtSd�������paP0ŁiV�VIuEm��!G#!���Q-+�<�)��7�p%l`����T�|��,��!l4������T�bQiH��5�25�`ҁ�{jKZ�f�z���s�L�O� ��5�����!�����Ͽ|}�}�F�T\s��m��0S��w�������k�ш�b`�Ե�ŹdV�Z`�6���`���dܥ�A@QJ������L��7H��\�#�X�Q;de��£_l��%b�麿�0�P��a0˛����a�����!f��ؘU�p�Hg�z>C΢�e8������Ȓj�SC����dp���*�>���NّE�L�+SaLaq�x6Vp����xU�n�������gx�i����~�QF��_|�����<���sN�K�|���E�h{;7jZ��y�'9���t����D2V6	0e�U�a6tg�aJ�,��!�J�{��P�KE�4�=U��wC6�D�2�
��R�p���o8QȢJ��U�O�l�r��PYΞ8�H�J��� $B���<")�$�x�+��;:����QF���E<� -�����u��Y��4� �����=-0q������3���+���m��/[T�����(����F�M�ا�6a�������i?���D\��p���v��HJ�;D84���>�!%ped�y�Xu~mz��-��[6SCo4�a  r��#�s����n�Q����/��愵	���1�Ž�?��HX��|[	c��^�-Xb)�(_��}2�^���Sv��~������L�^�a`��2 a���+Ӵ���$fS�^�b>�i�.�WPs�3c�^��w�`�n�J��B�	{C��D�E��±�FKP^���<K�*�����$?2z��D��Ð�cR�%���Wҥr�_ p�˙�
K��^v'v\a�z���M�=%@xwJ
���/��'��Q�%��i���D��nc�楧�*�><u~�3]�ۻ��k�<�٠W�v���Ʊ�6,��5�a��_�@7�5i���,�1�	�E-�%E�7^�ɾu��N��8-��\�r��|:�y�a��Df�9<��[�-}ϳK�����#���Aր�ě�#父�����|���Ur���w�ǻ�)g?�}�Cϩ��"$DA�Vq�No�>-�:9>��rZL��|���;XR�jJ��~&՝�a:m���70�ñ˿��w�0��Jn�pnk�=�k����Q/��.�q�3�;kcG�čq�ASt[��L!3�Zߤ��d��σ�8��;[�_a����05��HieG9Q��P���2zoE��w�2�l�"$�w����7`� k�w4��s뎿c��^����'�?�,�֤A۴�IrU���G�B��M���t���V��l�m�3-�w��J���&x�˾�o����$��" А��7-mmc.���2����w'���L���>c �
l�I����;C��l8��J
>�}��t�j�E/ECcZ�e\��Dn#_�����SIzѡBDD4HG��s�!��Y�D�-q�݇������*"��7Lv������GU+�AZ����%���%đ'�?0��zfV=�&��(k���F%iU׹/�K�/����X�u�t���(afe%1rԩ]bx����S�Ūe�c��vC�gG��c[	-@MU��<�"	�5���:��
Ax�4�������f�� �V?��A7��K���绀���t4�oa�s�i9~��Ey��%_��ϡ%l��Zs�ؒxN��t�z.ݷJ	w��:7�j�f���;�屁����~Ֆ*���}F<'���0�c�mDX�$�|V�b��w/�i�,r�K��SV�}��5�C��g�[V�g,AC�[�i�:��Vj�dB}�=DU��%:�L�q	��Sr�J=5��� 5�㽖+������S�ے!�;m�ۂg)��P�v��Okv�o�������ݿe���X��,�Q��.�����GF���(�߯�1��s�nC��-�.�!��I1��V+��@v��Έ�;���_r,a!Q�j�fز�Т;�`��$�m%�}����=�\����f3�͔���cy9��\o�Z/�S��K�O����Q��P!�5{�bbh�^�qJ,`D%qV&�*�;�2o� ��x����S���#5�Pb��[��`��j��߲��Ś�m�~@���nT�%�}5�����N��(b��7ƺJ����wC"��g��}=o��2H�%�Ӓ��$�I]՛�ī ��N�ɤ%��>9��Y��$��91qLi��Q�f�Vڊ��*����5��a�&��G��yfN���tW�P��c�p�B�Y��a�իWg��l�w�Ok��"���i}�U���+���ׯ̲��Ro��[kt�0��;l3Jc6�Dҥ/��+8M�^0Ѝ�j�_$k��U�"V��/�)	˪�9�k�5��4���L	8i�t�X[���y�'����\��|/}4����h_\�\��4���}b�@���"��Z@Z�R&��F�a�Y����"YŕK�/�Ě7e��P�Zs��u���2tq�t�Aq.�I���b[�g��O�Sl�	��^Y��|u�a��GV��~�z��5�I��!���2����tk	p��n�0 i�e~��Pj��E@w�7�%����P�"*�U���y*}*o�p�����I�z�0jX�G�ߘ��5LjL�)3�DU��/���i�Iy�ы�OgBZ���Z4�{V4���F��K���K�b;Ҳ�&�})0�8�&����\b�S��L;`�,�	˳ȋ0i��I�`�Ֆ����u��5�+�������D����2u]01��Y�f��7d Ҝ��?I^���87MWxɨ#������i�4w���W([c��,�l�%��^	� �#k�E�j����
 )T��f��=��5
����z�'���Zwl[Ύ'��=���	yr���m���L��VgR�Cr����YQ�
W�o���VZ]�4S��d�l3��ڴ4M&2ט�ᾬ��!)��t�s�U��s��4�=-	WO����T���dXJ���f>���3�4������kA	Pf�b���y��Y͗���ɟ����9 ɜ�+�kV��/�K�hD�D>���j�s���ǧG�Sj�Z↫C!���F����Q���� 3�p�vQ���bۚ�ko�N�Ǵ��Z=R����~�r�z����ޯ/��ʗ�fҌ�k(,�t���8d#�����~�ɖ�y^_��tJ���{?W�g�V\�/
+���Տ�^Ta*Ǵ�1��T�4�%O�ײ3�`����5���fABй�e0�n�48qY=�-�.S�e�#s�1�\,��u���ڞE=lgٲ�V�
�Me9�X{�xx�z����?\�������p+?����g[s�|O�l����u$�&�4Q"�����|M,l���\�_�4�P��Bb�X*K~S�z%�$uH?%��җ5�wK�����u�)�3F��Ke�3��)݁b�GEC����MHݣ�tR�q�56�v���7ɗrK`�q�?��K͆qE�#	� �4�ʨoa��z��$�v�ٲonc�~h��NA5�U�l��A���
�L=M���U���32B��Ȳ�ۗ�	�'�/�K%&<⢬݈��M�דa�ZԒ]��6�=.3�*�ҧ;����2��=y$E�n��bd�������0fޡX�
G�׎a1aפ�f�f���$����|�֒�"2T���NxolAɱ�}���>5�2TAeS��'�K
&&�7�ԏ<m��N<��7����H� �F�ԏ�����{����I1�Ѝ��~�1F��%ܴ��Q�8�R&�Ǩ~Ȉ@b��ǐ>`�o*1��X:�i��\�����%��	L���7d�8H�hY5���wG�&+)�3�s�eY}�׾X-��3�#�� sVn�^2=��`\��h�a��d�A�8�ӮN�_e�,[����i�)�=�~W�t�b�&����N�GA��ϖ�sFf.�^q�n�-��笂�_g�Z
~��n�%]�q��/&K��s��(��u�FYB�m�ی�-4a�̲�w+��erϟ�·�<:}.�Ov�&��%V`п-rV:���
�^�O�Hg&���,�A�:8��U�W�55��6��`6]�����Z�φ\y��]H��4��&�a[��+WR��
r��\������'�-akC�(��9`�/�����o�W�����?o��l����垃�G����� DE��u��@	CF�����\޷32\���B���\{���a�A�OŪ̷��tQ��[���U+���@J�l��V>K�QMg�N�h��tI��H͆8����p#^���_�ֽ��E��5Dl��MD�,$(�)�wy\3�*do.�>.�=�������'\��c����hMO+�.bŻ�؇H��|z�I��y��o��'<fa��9$�:D�������Ly����C�%_c�4��^r���C��ɕ3I�����$�K����~����������fξ��+T*��
��I�'3���2r��>1��H��JtC,J��(��3���~�_ D�����S�}��n���L!�_�ޞ��Ͻ������t��$��z+���:�~U�4ޣK��np�Yt�p�~����4��Ճ�&�}��p����k
��o'���⋐@�1�ec������Qm�K��R�b�)N�R�
hq).�Hqww/^�ݡ���5���]_������ˏd嬬�s����{����T��3��t�2y.�Yi��Usz�)�(�uas�?BlU�Z v�ِ��볁2�α��Ǩˏ�M���� �U��D� �_����t�S:7��|l�6�/�M�~�cFy{�  �SF�d���'�l{ 1��f=3�7'?����	YQ��״��T��S�D�ZՋ�{��闔����N��¯����AR��HZt�Wl�]/�@$�=�^�~PI�UX]�xi�+��)�	Z�U�Fn�����=Ϋc�ȇ�\�3�j�x�hy,�2w4��uE-�$J������3m��5c&��Gx�6��&�ჶ^{:79��9G+��e[�����ݘǿ��eU+ᨀC!�����:E��`n��${�_J9VO�Ncg��"glY{.�}h.���r�(����������e�z�l���*�B��k��.b�4F|0O�������sе��:p�О:r$����_��RCx@u^/���@�A��&oO�i��Pۄ��h��k���R�쉨i�(�W�I������m�ṡ�������RVL��";~��!=a�V���M|�T�]����h����v���X}�]R&A��F�:�L�Z�q#�d�좂�����_�ydҖ�,�*����357��$�54�Ե��͑y��;9�U�S�b�౺���_w�mS��Q��%��0>�I��d��/���X:Nd4Q;T<�TLBd��L!��I��c�@bys-Y�e�6��ɗs�����ޫ�m�٘�ɢcRc���jV�'�Y�7�#f	�[ք�y)T�Ʉ�
GEz�Nw8�.�=�;���!��䪛R7�P)� U�Z����1�-nOq�H���mb2�.ծP�"Spro��~�7w;��ps^$*նT8�;�i2���IWT��������W���ձv�i��΍۩��r"ï_;��̐���8-���fAdSvtآ���y��Jx�[��_��,8m�ǆ�ɥ�r9G�#`��^��i�S�(��j�����{T~��ό!#N�7�lԥ#���������|���/7����)|�47U ���V�k���£�Vh����r��2�+TE�yS�����)W���6�x~"��X���\��.{`��L�Wb)��ڴ�JhT���|�<^���Xn�!+s�G���F������p�P�����9����q���rv���p�2/����rZKF+eH�D)��$2�ٞ��#Rr]ZA��{?\�r��^���-usa�������!����=%�q'{���z���}�� ��K��1y+��@�`���e3����9Ww��*�Ԟ�6��o0�<�����P�ޅیP����!��2*�5���i��,�j��F$���"���"�$�F�u�};��\�p��9�m��2�8���˜�r�u�	��m�ttJ������2}����`��Li����]T�jъ^��&��|���Y�e,n�֫�!4����Y���hN�� ����ԛ��ESk���D�E��_���Tשa
��%\T�@���������P�?�Y���"���3��\�g��A=�b��	p2y���w)��h)o ��ϖ(�{!����?��c2E�?p~�⤥����aM.�`F�ם�ķK�+��W���H��+��"9A��s&W�nY����w�斢gX��,l�t�H�Hğ�){��<���u�:�`z�1�2fTo�yd-5�Ť;:��]�/�c�}������rJ
�� ��v9�����+u��Zt�vu�.�~�[��9&7��Mrlr� �R2#�����t�T�,��ī������aJ1��U-�0�r�?�L��(p�����~Im��B��g>#xK
P�9��5����|���2�
�'N�3�hk������軼D}��]G��?]V�M%��y����d/��l�%�FH�_�Eo�(@W}<��3(W��
�5�E7�;g�c�sf�'�}�7>aT��38���Nc�7`hH>�'��i���KOM�O��jԟJ�{AXWғɦ�Y�Ȇ��ؙ��U���`��kyr ���A���٘ыQ��.�<)7�%АW��7����R��C\y$]:�d<b��!ʔE+7Ih��ޒ�����<{cp�1�Dq�,��s��5��t�E��_H&�6*�]1�U ?!P��.O��3Mh�KX�bD.�ݷ	�loQ;ny����i�O8����z�����$�DSnͮaS��7;oj	.�y�����D��.���!nSM>B�NacO�T����T�I?�| '��p�U`/E
�G��Sn����݉��n@��O�б��"�$���(w�*sm0IA�l��&���鴭#e�ۅ�Y��F�Ut�M�D5��1�T�`d�3C�C0#������3G��u�*�BE8��e�뷣12@H�4mv��5�Dو�o,r�����Aeb�����D�v2y~%�.��kс�{�G��p6�7����:�;<��yy�$�R*�ǂ� �[���^�zEm��t�8#���uLz�������(�n焸��<���f��U�9�D�./v]����9:	��
O�"R;�����b���y=�cm�4R����R?[����cۙ����Q�>�t/�G�c�ow��]��������9�z�Ü����4�ޢ�V��j���t��9�ϓXS&{��T� ����Y�������֡��4�ܰ���M"K`n��^��P�_�\V���R��5i�i�v��aF����_�]��ݿ�L�1�:d]����E�0�2X�Z9�@X�D�h��&Ǐ��� ���z&�A|*�_�3���C����I?���S̱��%tV�V���3+�ZΔi�=��=\���#�Q��U/��slջ������L=�9L�vn�ȓq�(3	ۀ�.,��B�_R�K<ޏ=e(q7���O�]pT76(����9,��{�<\Tz���)Z���WpA��'bm�x�8�n�3�Β7���:�����.vxn1�I<�Ā�����;�L�rD�F�*t�aƍME���{�p�qT�+0��5�����	����"�fV'G���{b�O�ﻥ�Up˚9�t�햰HF�Y6aIĕ���/�����2-����F��t�{�g�^��l@Z.�+���mX!@HΌ'0x����ws(e��n�}����# ��� �N(����z�t5��$&_�o5����i.���,�I��^(��Yr���� �:pY�:ZM��Kc:��ٺI1p��9�j����{vBf褭�k�wy���}.�-�@��+%:��W�(�y�R�(6�H��|4,�[%\P�� �z��{���{s�'Ɯ}���p�x��.5�7�+.6इ��"��-���઻������:����.=���E��y��)��������'��(�D��M~��2�P�����yt�FvMq�iC�af�	t�mm�#c�)?���6VWWo>�گ�;��r:l�S@�Pl��_�v$��Gt�<�h;{����	��TY�Y��#�!���X�eݳW-�{���C�s cw�O�����I�nd9��m��E��kwd;�:��t�7]٫����Dgɵ�Q�
Ĉ��O�SS�3ڪ��3�2��ŷtYE2�t��p��U�fP�t��#������-���=�`,�4Y-�T�g�/ϸ3�	����C]<�>.[�7��f9�Ϣs�b��{��3c,�)[�Q/�O�6�40�#��Cv�������%��i5��֞!o�^CJ�����1��L����W�
k���e�w�K�u�[�	��Bh����4l9��dv�l��&vn��(eH�{޻U��5G��.�70{K�Ns%Bnp�B����yG��&�G���{#�kQ�/F��G�����:[���
3D}��;N�~�E�nl=&R��:jy�p~��3��/�ܶ�*���T��}1�X6�f�+�H�y�ߕ������*���;�mz@����K�SˏM��5_�����X�\�
|�š~��:��u�pD�Ԅ��|CYs�ЎZ����$F�+O�J��w�ϣV�
� �ܚ6o�p��^��w�^$� 2{G�̯kyh��B��{������w�kg7c�ц�]9�2��Ug_\RN�z߷GdE[�T���u����Mļ�l�5�{IG���/ �����q#�����^�M���������ݑ����̓�K��2�|`,h]:#=�xO�j�Y�R��y;���s�;ʱs�� ��]�E���)W�zD{�H�~�|<ݹ�Hrr�YyEuA��7YW��¡A��s��8
z��TCRثkjT�����7���5�It<{N=&�*`>ΔJ���A��"�����AfN�S�����=�z*�����Ʌ­��f�n��;?�p�W�L�'��>�7��}K
�2)u��E�C�In~{��)
z���P�%��|��$z�&گ�ط�B�\���xM�y������a��Q6��l�,�t���7�*O��m���&Trj��Xr�a�$�T�0�D��jdí��?�z���GE�Ӿ�O����T	���|�i�b�?$��A��A}82�(<���J�m����
mmm$Ƴ�榦AN|P؎S۾���0�zm6:r�unڠe�55P	'��+�A@�F%<����SG5�6{�y��"�BB�?6߱�4g���sϩT"ݽP��&|ul<�5d^fԺ��l�����K2uOa�=;w�Ŧ���h� sv�3ϑs`�vt�of�oP]mgBxĮ��f@צ|��T��y��ٵ���Y�Hw��_���~	�KXI�gHK�(�23 -�bz�gR<�2@��>2�G�?����ux�i�+�ND[�N�zȕ��!S�B��)++������B\�� J��lX�"������1kv���i�I���L{�-D�u$wvv���s�b�4�y"o_�5�A�g�^m7PS�0���$F�ĞT�U� �v���VQ�v� �y�(�;��P��bW�\E���~���}6|*X^�5K^�N���Z��ɵ�A�I=z-m���8C;�ު��@r��9�����ag�;�5hWX����r`!�^/�e]�r�����,�ٯ�r-�n��`ka����>E-�E�b�5b��x�r��oS5ft8R0D*�M�l:�nT"�o�+�`{P��������|���}#?�����Km	�E(�.�`���F)�B�߿��[�����g��ʵA�
e����B}H>�޸^	�S�*z���/�����.�&���2!�T+f���_������%�����`�"e���a�\�g�ů��U�����	���燑⋓ ˬ��`z���	&h�{۽�b�i�;/�k��sJNI���2PP�'�Fl�9�G)}�)�ב�\|��g;��L���ݖ���F��/e����R{|V���GVHA}.�\���n�Z���4��i.����������q��92����Uk�0 �,(ms�H�R_����*����e�T�+�ʕ%_�����(����Efm[[�z8`�f�"��s��#a�1*	-F���e+�ꪼ�Uc��a<�4�O�`��K�}O�h��:��,4,��FP�Uy��%6_�Xq�����x�s(�����L*x3i��Cb���D�𑮢���Q�g��Kؑ����j�T��ݤ82T���WPP�m�twԙ}�q��Q�lJ�����9���o�\Й
gShMPͲC�k�-�	R�~t��20^�\��VU���������C��X�L%RL��|�9 �@܉&�3��D_�Z�m�'�=��)������\�o���e�m������`M��<���Ƚ��^���+�X	�s�n?ا��3UQc�f)�i1�K�NSЃ���s�^#��.�X�S����� -��<�6�FQ�?�{�0��wk��D ���V����g�_�2c�X��UAQ��I��M��f�Cc����y67�b���a,����b�G�ߩ���P��ll�@-m����3ϡ&O�·�N��#�ۍ���#|5�k�u|���d|�d��"j
�`���"fo-��xx�A%#��`���a��es��R���2�y�Q.c�������8��;�B-�rP��u��2���� �pc��&�� ��U�2����x�Rk9�sEH�b�i7I����J/Ў$J:2Xb�8�]�u8�FnM4:o~��B̀5\��zy��9�Wb]��\~{�1H�@��:ʇ2�ʈﴅ�:g�@��"��*"��FM�c�eH2E��K� q �ԕ�7���� E#�U���B�8A�!U��[�4�-k�KL�ЗS��i�L�'�V̅��Y�_��K�}D���\�oWDmO&�Օd0dh�F?�ɱ!"$��k:M���~���Gpg4�v Ty�R&���v��C�A ��ȹqY�.��'D���?ƛʾ'�Z�z�q����y�q��R���މk_ʒ����"T]�jf\�0
]BgHm�y��G�����msv~>wΚ�,*�k�Ry�Bg��Ik�ܨ�Β�9�o�Dor9����=.����@o_O�H��R��[�bY�0���FZ6�+2�T�8��ጎ��#�T	���.�sF	Si�[qAc���[��!Ž�"3�(>_�f���E��2j�����s��{��o s���_O�f��:uyh�xaE~l�e�$sB}�,�e#`�,�/�N$11�:%5]��1ᾂ!b��=]v�1�����=R�I�c'�r�6��C~r�w�I�A{�=�12�X�`!���=�;2\tn$P>�T$l�;��~���n��ֿ_'�K̅U�\�7���D��jFI�c��0U�(d����~�=��C��������Iw�|�(h7_w��P�%>�c�B(|2��}z��1�<�(O�:c������a?���G��p�X�e|���2���D�0�P~|\W�2-�.�D���x�u��+��Ϙ�B����y{4׆��z�N�����'�~�E��?ډd#H���i:�R*}���sٛ�#��nc�(~ʶ�2a(k��z)C)�����{�$���:6HO�s�OQj���E��� �+ݿ�|�E� �mͤQ��i�H��]I"���5�Q�5+Ѽ��u!�4Ht�Z�Nz)�h�#	ï=]�=Ⲇv��,-v7�5�g�ʪ���4N����*��`�1���>�E@��#ط��,_���<�~ё�9�I���K�b���9z�뷄rbPc�6g�Bb�r�YtsZ�O�M�3��,��c�-��(ݥc�|�" ٜ��Xۇ<f��8,d���j�Ny7ɼ��
��fVܾxwH�qTW�Hm����HV}՗�3Mf, "��B����.Q��d�ȊBZ�"I���M�*��G�A>�l�R�&�4�)�1������s��B2^�������"�UO���N��'��¥1�A�4o
����2��l;��`���t���S�I4\� v+��CpV:��xC�,��J�fDv��i91�������T�'o�x�* �L´�L�MJ+�f�]O����B%�2�
)X۠|ň>6��6g
�M[�Z5���+�M�X�-Lcj��OCh���:����d��ö��3�\�\���E]���1���W��?`KM'>���Ǝ=���#�?[|�,�x�� ����!�ʊ��� ��9��D��;�K��/� �d�>�x�]F������竹(�V9q��Z��Uy4cԠQ���A���JJ��7��
�W���x��ox(�����wд2zt?z��������{v��hEP��q�(1�B%i��䤝,�-UP��u˄?�DP���o�:�}�S���:�S�g���lW��������X��_˫5Y��)�2�����)�Sr�3S	�gK�.oy�S�������^:�xw���_0#nm��tB,�b��o���Á��=�J�ʙ��?I,�S�JdQ�v'@C��2�4U\+��Sz�w/S��Y��"C� �rF!=Ã�\
,lX���v<�-��X*�%Mɳ���dЏ!��zԀ�
4���i��ڨLK�"L�O��bD�L�i��叽(�Q�W��xz���NNS~7#XZ�ś'_!�B*M�ߧi8�T�4���F�����~��Q�MGa����gn���Ȧй�/pSm����Q���~C�&s"� �|�M��~�r-���L������!���~��hЮ'S�OdecC�nA��&�pR��ՠ�./oEv]��l�QS�l].��Wgk�	6	a�r���r���(�&��#��ɇm�R�ţ��	��4�Dv��v���%�0'��J�e/�$�m3i���pm��B�bg<�8Xn�D�p�_�N\e y ໬b�1݀/r�A�4;��8�tKċ���,�?o��u���/����	���iOT]t�?<�2 _�̈́<j��R���F�u������(�����M��,3��2XF��r�f~�N-��B��]�ת�C���x����a���{Aw��P~�.��*��76&Sd�������Dẏ�X�7�t�"%�����9��wd��[����	�?�����n�1<�ɥ�K\�ҢH(�v�l�l 
���onӜ9���\VF�E���d�s�$�~���.j k�	�+~>������	w)=�B{9��o�Y�*����w̟4u/hi����p���.�b`E�)c@H�7�j���C/��5����&Mn-S�:�02��
K�"g���y<�=SC�7����q=q����a�ԡ�v��`sv��[JQ���u�=/ܑ�t��
,��H���',�mi}*�p�6�wX������=�k���o����!��п�Z���y塩��:��܉ k�9�{�lP#���Z�{�z�T�\����Zϫ�,�!�u�*���)�#�t�_v��h�>�#V��'0�%�I"9���M����S�����KZB��}Mm��˸�w���W"@�c�����c"�t���/�C�A�T�P�����n͹"�蘁X�(c�I��4�X�Ȳ�H=��M���_�<�\4����=s�Lh�������]����KF}������;A�5:o������B"Q�<>�!�2"M�O��WɓO(9/������}	�"3��F�_a�ʺX�󪼼�a�}~	�`Iye3Z��<�},<���Z4- E�Nj��`{G��� ��D/�G
g>���@f?x�LYt��T*zq�fg����G3�*]������{����[c�uä����<�k�X�/������Uq��2��y��������u���
r�n7"�y�E�D7��I��I:�6 s�(����2��:o�3��Lʱ����_�sˤ\Jr:���$&�}{+x�	r�hz,�_��'폘2G��`�a�k��c��{H�mR�rZa��(�hoo@�3��GqZ�� ��~ސ��EW�V�e�O7����'�E�=��ڷjݶ9\��w�2)6T��k��*}���d�!׻U�V��8�+8H"Cs��r�+�_uo>���2��<����p0]< � ���=�1	"r)�
(*�ms�r�
�/��x�	���ڜN���5i-i�w0�͍mC��goI��ُtM�I΃Y����SE�n_����g:V���z��PU����Z��������/)��E��e}��$�E"k@�"n�F���T�R�1z6P�����E�]��5�=#�g�Пȟ$�[/�1���8�{D�qr�MCo����a"U3V�u��qu]�U $j/̖-&�t�[~#����|���/f`�i!$f܊mjg|���<:C/�˿��KP^YɅA��zM3Ju(� n���
+�A��R�nW1�vdk6������]q�� ߙ��J�F6��;�4�w���y�"��ѓ0e/�
^��h�"up����L%܂/�v���֠Mկy��:Hb��I��(���os��˫�л9�b�����	5�2�� �!;A]o�%��]�Z��3�p��#�t�$���6�����;����U��;)�a�+.�ٱ��/�8��f>���nQuR8��o�0���㌊#-q��!�ӟ�|#Fnn-�r�7#UA���}�A/
��t�cؚڗ<) GMC�AW��5����F�s���2�!ɤ;�X�����H���ENU����I�����%O�[Z(L����c��O0������P�<���(�����7�[7p�9K��ﻺ��+�/��PL�R��69�S�DUœs���ē5�K�'��m���b9}G�_�`x��ƒ@��o챓%	F� ������T�����������9b�빴��(�qW��5�Lz�XV������W��
m�[��0��$�\Cw�\x��"N4�Y%r�&��h,��O��e��W��ڌ#m,���������ʙ����n�ad����nb�'�7�6��qHG�����	���P7v2S+�i8u��eD������78��%����ԛ�ޏ�+�����ǐ��E�II��')��y�"�.�.�+�!���[.V=�J�Z�a!��~�WiB�+�s�y��S��M]8�����j �������FgsǗ������EKw�]h�e+����3��\��zʝ���Up:QL�ͽ-7�dʼ�w	0�!����������q�Q�[��-rj�6����.m��(����U/��Ϊ�f�"9𥡻�H�7���KԸ�|�᳜�-�Gc��qk�5��������F���il�H�H� ��@?d&,f9���O��fO�n�m�V.ṲW�iE��mvl$���)!��<4�Q������t-q�i�-2�(���G˗|�'����T�1i��>w���G>{yO+\J4�ccV���1��HLA�B�������X�T�?�uP�o����&�T�L]��F�-��ĉZFǩ�~�y�4���k�Z���U�J$u�MJ�J����̀fI�7�ߠ�gE��'B�y��uWz�ڇ���o�F�*�0+�
Q�ޒ@�{��J����{Fi�@��`25��|������ǈ;��(P(����Lb������$UЛ�d�f�YvM��w �mg��=��h���&O��!
&�������'J�1�3�v��sI�A$�M��۞��� v#�����+t�d�!��3�G������{x�&qVs�TlR��T�<�z�j�}8�\!݆�^*�ؓ�i�S����2�D|3lR��Ta� �7O���k����c�_���c�,`lS�ʛ��W����R�M ������l�@)Iɴ���s��6�d9|kp��8U7Τy��9�g�Z�� �G����'�J]C08�������̚DV����gz^�֪���o�~@��'6�)N�ߝ&�-c
��)X�p��v�m�YLG�Q��:T�J洨A$�K��"õ�?�[�͌� ���?Y�l������W�K���gE8Ѕ��"Q�&-�@����Lj����8z�U����70ҳ"��i�27�7��zL�_1IN��#i�~M$�
9f�𘤎�P�h$�E#���߰G�̗��0�N|w	�.��l Җ��*8��������Ѿ[V��+<_��'�m4C������G����C{��X:��� ��!5�||�_Ϫ	��*�]~�#+��f�����+�fY4���ٽ �������wp�Ete�;��Wb�b��.Y��*|"3aVZJ�*��o�&��4u�9���* �
�ܿ�z����4WF����6�9	Pc����v����Y.������ø������ę�#�稐$���A{`������L7O�4xR�#f�k�|2-�K h|�!ϻ�A���U�[��U�?�÷l�ly�$��bA�	� y�ɟ ��$mQt�>����L�d�XT
%�ZB�3�	����AլRq"�5N\x�3S�\~� �T�6���]ib,M-�z߲��Zy
-�f)�
}7^H函r(I��o��ՠ���#��yA	�iq��R�X��x�AKL+Ib�+��q��ꎭkLL0ǉ���D���!-���W	�H$�WuA��9LJ�L8HG>5tm�_�]�,�}��<_߾�*r��	�Fn\+�p�E!�S�g�*���/N��qz&��_j���x��.��;��-Ú��3�����?M��Et`(�լ\3a�R���zT�����LU^c��723 �Q�X.s��~�>m���!_�H��Isܽ`��LǬ���z�1��1��0�'�n	��u)oD2��A�P�RV�`�����ۺ�ޮ����u�Vfx�\��'�뗓�}��Nk۝�=���w�=ݱ�t�b  �_ۘ��i��\Vqϓ�W����+���G���2xޝE����~�����*�>k4p��?��i��ٛCOfƬT?�-��0���6�3o� �+���6�ƛ�r ?ǃ�곸�G�z�s�Ԉ־���(n���1&r��󉹴���͘�u#�﹑�ا��H~�D욝$Ith.I�*�eX���1ɽN�4��d`LR-�Q�HG�����̏(8�8v�0�����	�0X�Wr=�%:��i�ps4?��R�	�I��GZ��ʬj�d��3�vK@���@=���S�������rv�w��]Nz��8��<�L��>�?Qc�ճ�ߦ�,2�p�Ma�$�k[0��r�Є����Y�Y���$m�F1G��1Nt��w�b���9�/9��N;��Zw����������bz{�Y:8UGp s�$)�+ی^9�hDH{Ӄ����	�^rj�<��Zt��!���>��E�An4��Mo�=�=��g�0�ǜ��*�M�:Ͷ�;O+����%�_x�LK��b���2�r�������Y�J%�����QE�Y%�8��x+R�f��nG#��]=X�V5睾��7��ڛIb��G�;#N�Zc��݁x�Wcu�κ�7/l/Ƭ���k�uU4���-�)��p��p���2�^཭w��v�,$qr��5o��j�62��o�(Y���}�M��z�f՞��W����KӞ�"·��f^��(��L��
~|���g����8~� �q��D��99���4U�Vq=o��U��И�⒇��ф�Ĕ��Y���hX�Q�zo�/��I�k`���[�4����*��[k���u��!�Ɠ��������  �_e�g�z�Y@��k��3������H�1�>����4Y&'��������wC�$�έk��}ى"B5� 1�\�}yh��x�ǸG��Q��(.eV���!di<ӷ�c��f�6���}v����	h��Pg����W�Kv8��������crZj�oٽ��_夔$+ſ��PK   �>VS'49߈/ q�/ /   images/a09c37b2-5d65-4269-9e69-57a504bc5c33.png ~@���PNG

   IHDR  �  �   <rc�   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���wI���5O3��OWU&5�֚ZKh-B�@Bkh��&�	j��T���YY���ݫ�>����� dUߞ�~˗��m�#�ͷ}a��_���6ȿ�헿�������~���o����~x���_|���/^�����yr��ӫ�\���/��x~���7�yqS��7�n|��&@�׾|v����\|��G�����G�ϯ~���/�}����on~���w���������?�����W�_>:����/�����o^?���o�<����/�-�{z���Ë�_>����@� }���[ ſ~u��רAỷ�G�^ރ'�j -߿��w��J��eAd�xvM�y|�������_x�������o�E�?}��?���e���O���z�>|���_��>���ի�߾����~��䧯�����=����?��_=����|e/^~z����gޜ�wm������	fܘ{tkayi�ŃKp�G{�_�]�:�<�9������>\|���O.}����+_=������;s˷f�ܘz|} ���􃫉Wc��Dɽ�r{1 �\"��Z|�v�����ٍ��n�w�7�ۧ���C@]zr�;�-�����W�^?�/�>[�z|+��z�Υ�ҕȣ�ɧw20>�7�����{W�p`��|�_��FlQY��On�^ޙzq{r�F�������'�Ⱦ�?�ţ��̿^�A����+����.���z�w/�pt<L�ҥ��	�;��o$a�:繾0~����	:�,>��Ӏ�_,M�{|�ó����K�`�v����ҥ���>��yn��yԣ���k���s���{'^	=�yr=
� ��y��^��0^_�\]p_�w]�s$���\?�}x�I��հ�����K���Y���Lld>i8?i�0m�2���Lt�Ҕa1=t6�Χ�B�o6ҝ?����
v̄���uN�����xW����:O�l'����3z`�p���T�u������jq��x��|��~�>�t�q8d?����G�k��m��s�[� n���`�yD��Qvܸ��� P
F�p8���T���N��ٿ�pӿ���]U��jso����>��n�Gw'<8��`�|t�|�p1c�4i"qy�
�L�T�8�p��tzz+��[�� ��;$p�H����<x[���$�3�,M>�7�|�ك��0j����^>�G���yt'X���7'ޚzt{���٧Ks����_x���N0���{u�ۗ�w\H ����?���riC
G����i\��FN�sv�ǈ�'��C~�d��ӳo���| ����oepE�uwW��{� ���� �<Ұ`/�>��}p)�A [؅�02p���?���ԋ{��K��;�'��o�݈޽4�t9p�J������X`��/�r������gQ��<�:�<k��Dۖ��o^^��ե�^_���+ �_\�����[�d0�ܻ��l���c�݋8������'���W0v)`��&lQ#�%���8<�xx-�4@YY9�bAeD�s]��]���Ō�O�ϥL >����N�1�c>1|65z>c�0e�8mH,N/�X��Y�ǭE��ޛ��H�K�YH��,��$`�.���n7ι ���\G�����ʜ�M#M���aDh��N���#���A�F�Y�� ��?A�L��$���@7���C'�U�[Gm(��D��c`�v�o=�7��L���# �<v
�1�aX�H�Yaƀe���P�s���WG�����H��L��@�����W��ut��:���@�-� 	da��w��7�m�F���փ	ۡ�a,�c/|����-�ml�7ֆ^�3��jcG���||��o؍�Q����ؤ��L�}>Ё���]�wU�#� M�Q?���v�GZǇ�����Z[W���
Y⃛��3��Ũ��iv79��}��6PO��u��WKF;*�H{9>SD7����=G�;�l?�۵�8���m=����-�9��_�����y�̾]��ޝ�p��4}v�e��֭'ڶ��?�8�:�������$��7G�m;N�����>^�y���pٙC������u��ÝMc=�ƾ����t�giػ®ޘw �J�q��ϦpU:'����f�/�����a�O�f�橰LGLsq+,Z�,�\�S�K��+�l�>���r~҆��'җ���"}q�qc���z����i���.&-�fp.n:3.D ��x�b�=	_*0�fBC ��19�O���zgbc`6n�K瓦���l��J�l��ru���0A��>�>~۩���:�(�>���Rh��C���H�\����0��'C�%��焕��^�q��AS����Fd��zRt� �"��!�'<F~J恽 �qz�pV����f�<��T-OԌs؆ ��>�b�q���D5`w���ZGUzF;���-����&�4,��VK�n`�nCZ���i�t&p���!�����}�1����ۇ8�:G��a�4����>K�^@7ွ�e���1��O��JO�Ǎ���7��1G�LS�+�nX��y/,�Χ��R��I�B��@F|ԩ�P:2��DGf��������M�^���^��;W#H��]�zi�'~"|AT�}��ߙA������`�w�Jܾ�.�n^�޸j�8�����9�a��/ߛ�w=��O�=8����O�*,�z�����g��y����^����|�d��g��x�j������o^,�}����3����/^� ��o^�o_~x����=_�]_��7O����c���'_�|���ˏ�={�?�ŋei�'ٴR�?��Uj~���_<�����f����^������/��>_���*a��3/�`�:><9���ů�/ $�||���iLw�"�H��)+fH`�)�_������߽��-f�0b֊I<^K��{���K�]�j��7��|����On|�����W�>�����w/�����ֹ�g��>�}?<�����?������1 ��<���{߾�Ԇ���@F���E�߽\BU��O_��?~��?����_������)jC���@���ETP��Jp �2�@������O�|����o�����?���7?,_����ŗK�^�;��ۇ��G����ë�K�w��ޥ�w/$�_N?�����ק�����˧W��WϮ��7.<�1�]7��ֹ������;g�K�/E�^K<��~ug���i$��']��[����8�9�s�{{�sk�nιn�:��8���s�Jً-Ұܻ�w9Ʈ4-�����L#�H�o��a���v��������E�.�o��<�|t5�|3�[�'ף�/�.����<����s~���?v!X��w3o�&_b��D����KA��|4���_<�}v#�n�p�N���i;�G��H`ץ�y1a ���|`�2i=�	�/D��FG���.�Lb/>%�aA�3����/D�Ň������ȥ����bڀĕ)3�<iB���.e�.O�R#�C��G��Ez19��ڜ�Ҥ�l|x*Г�	ۏO��M��C�=����0t���9Sm쪷�6��[�m>����h�q"�:5����������h{����S�'��h{����=��C��5�����{{���8���ޭ]����(%C'ˆO����k�2tT���y`��=[FΔ�*�;������C�z���?��vQ9��șb�5�Qj�*7�TZz��+`�E{��yp�}��(�jO����EpCHcW�������8nh�����ͭP�w�����K���.@�iꪵ�7���ZŜ��	�锧33�=��HL�zp�������׽E?N]�Ϸ1�����9�����b>��<��|� ��H�4����c��	�����0���q��%��#�fU$�4UHd��La���Ɵ\�?�H`�H��V[&8���7�����3��r�����������W�(�ܹ�G��C�ܿbW�g0o��zi�f�Vda���K�2"-�\ �`�0��z�',�s��8��EPv���'�q\�Q\�
���\��\�6]�1_��ܜ��Z��9�{޵��2��:,;��W���(��>���x���&:3�v��0&=�R^X`�L�w$=gbΓ�q�3����`�t��Τ��>q�)7-8�.Am�C^�c���#؅�P	4����h�o��V���~)�#a�1$|� ��*������f潘�����11X�E�]�MثL�G���^��*���]��4}�������
�Ȣ~�B=ޱV�@��^��$7dQ*�(�?^�w, 1|��5�u�h��U�8nh���'�Tw�6zb�H�褡�b���ҨF��ZdN�,¨t�h��]hN�J=��G>�9������ӻF;
��Ŗ�2k� Yso)0����K"�ְ�90�����b;1Z������_9>T�,bֶ�coڵ?�ؗ��i랔e7H�� ��ƍ-1C3@B	�a!��}��3<� �@��m��$�{H��
"����u����h#[DǦ���P'��	[	���C���z01TP�0��#����)��q�a�-hkX[����on�����k����)�6xFqZ�t�I��_(�4�ٛ��"�ۓ����=(�����q��wm��3t�d�t�����]c���؉�k�X;�
H�O:X{�@F�4,�7�)�9R
z����m�Y�l�o�;�K�[ػ��/8�{�����Z�o�u�-��ޢ���G*��U�A��pE�����%���nǚw��z�nˁ�ϱ=ڴ��9t���}�JQ��`9�7�Ԟ]pVZ<Ѷ�X�6lO��	��>\�-8�'�����W�u���`qϡp�m'8�{>
����G=�
G7t
�K�XG����n�kH #�^2r���p>�E#�8Q	�Ib�O�D+h�0>O�:P�����{��A�(�@��
���C{]����J�5?�6�js��ő�S�E��JP�84������<X�" 	4�c��j�n���������do�E���iD<"ds2x�r�XE���#e���;Sg�h����>Y#z�bKO�BY��AZ�9UC:���	�"��BTn�lt��΁=����}���ޑ`|� �{�=-�G��@7�+�x<�,h�]Mp@����ř����;�� $������j�<S��hW��������n�Y�zM�=�C����&lǱ71����[���#��n�t�L�wǽ=QwW��r�+¥�٘� �,w�g��SA���D�}&>ޙ	��ƆϥL���7��7�/�f�<8����/�\z�|����'7�=�����o�~��o_}x����Ϟ,=z���o_-�{������ݫ�oU��b��WυX���S�}E�y�am�F�4@�i�<��Ų�L�|��ë�@8������K-�/����?� �/?�����o��������������������ݷϮ>������ީ��\ܬ��S�K��k���.L��+��Y[N.f�҆s�����l�Q`�	L�WfLw/�^�?�6�����\�5_���X��:縳�&Ꮾ�]I<��|r-��zz�F<�9��rF$^ޙyuw��=���̳���7��\� $^ޙ{�����/��;��۳��ٷ��a�����Y&`�'�*||5��Rbi1z�|�ι��[A�,�/�^N>��B�pFVEP	+�v@�O�V��鸓~~;�|3��z�����+��C��&_ߛzs��wڥI�<��|z#��7<Wg3�Ŕ���<��[��\�@��EQ!<�.��v>i����E�b�g�c�����,�� ��s�[󞳑��P�l�{�ב��N8O��Ǣ����ǑH���F�G���1Ǒ��h�sb&б��6m�>c�9g��`�s�vkނ���ȅ�"[�ut�Bڌv�E�E��E=���Kz���3�)eم�Tr�d�{"�>u;����a�{�$��ꆐ�V�G[CM��k=���a�߼/h;����{|c��G�<�-�f�`� ^鮱!:�w4]p ��nF �YEX�ш��PW5��G�Ӿ����q/�A��S����Ԣ~������C~Ckм'`��i��՘:�m�Ֆ�JC{���b��0��3�u��Zl�F�P�FXF���G;K����6X�k��N�.n/�*���_�]��WL�� v������;@߉<�R�e��*{�����U8֞7|j����Ƕ`;xb������e��7v;�\C��!��#�~��	�`������]Cծ�J=�᪜�u9	�'L~c��X�w����9X!�	�<#Հ��i�ᠭ��S���(+�z�kO0wU�`�厝)��<r�d�D���0z�l�vU�<^�����.�v�,����i�.�����.��P'�d#�#����q�����E{�%�C2����؍����;��[�l��L����Ϲ������'��3��S����)\ڣ�^�4�~sޱ��m;:���_H��K)Õ����br�)_Wң\�zp��84�p3/j�kW4�������X/�		�q�q/.C=��1�:��#�i���^�>�E���7�?�q�_�z0dُ+w��f��8�q��R��kS����yE��9U4t�`�x����������Epz�6�X.
֣�� C�^>z�e9A��#OĶ?l݇FY	�L��,�>Z����h���ı����� ZA�aǧ��;%\���#�cʅ�'hi�%��K{��(.m^� �x��D렭V\��
qi���b���6�} .��T���̲H�~=�pP�Y��:��4�Hǜ�#�Vd��I��s��:�A����Ɛ�D�q{SҦ��7�- �l�e��6��=��=�ޓ�y�9����ig@Y�i�w�,�IsC��4�h�]��gڳQ�<�h�)k�x%p�9I{v�ݭ����a���d�Z?a�X�`�g���oS{:�N�~��r��<g��Y�C���Ի�� ��A��5��j{?�˛��[l}�̢�AE=4v+�uVre��2��>�wz�֣-�9��o�Z{j�ʢ�S{v�ܽ���y�:��x�u�����2����� gxv*�>\ְ��mGC'�|~b�gh�H�C� Fpf��vu]R��]�^���Ÿu+�M��H~��<�C��*�6�Nā=���:@������փCM삛����[�{�P���[�ag=\`���Mc��Q��D� ƕ��Z`8�9Į��ᎆxwy��Z�,�� �^D�����_"0�Ԉ��� ����z���%>�0���������F{�2�ko�k�[���SK�0 �@�}�PY� g�	(�z8����Ϋ'�HsR��k@Z;�@��J"�C&�k�i�τ������W� ��n~���O��*�?Q�{���h>.����C�qn�H���8����n��7so=��5�Y���J�9��n���Yg��-���Y���ƾ��y����_�{���嫏^x��ҳ��߾���'/��}����g�^,/�����GO�^~���yVIy��)���^������<}��񃗏�c�v��/�}��ٳ7�?�����O�}������/����_�y��/����7����.���z���O޿x����7���'��}�\�r^>A�F�ŬO��2�V����{X�����~A�����/_|�f��Ӌw�&/͌�K;SCAg{b��g9�Z��m�"��u�9A��t�t�v�pa�T"6�XI�����x�ߩ)��i�(&��/�����s�p1i,��`��|p�R�|!n<]��ѱ�	�������y��9@b�������Ǘ.���w�O�]����I��i��׭Y7^I[QZ!������j�(�-ҋ1� ��9A��Ӿ�IoO�ӝvw�-��2
�N�����F�EY�G�����G�x�w�[�����F[O�����>�V���(#,��_b�{�J5���]�讱wU�u�\���(3��jHx�\8z�=�uށ����P��)8֚��t�Y�E�{	�q�~�����c?�>�ܧz�,{�N��L��GB���,�#�G(�9�vb�@F�7N0��3
1�@�l�*�E����K��9�׺�<�?7�F����c- G��Ʊ;��\�5��@��U	h��K�І-,��v��:+�@% 	d���Sy��"W_��.hh��L#1>T���13`h�V��\��ξ
�,ޡ���Z��~�0Z?1�Y�'-~c#B:� ��
��r׸�".D��83L90hE�w��:5����[{� j@AuB��z�\0���j�G�܃���R{o��� ��+�v�P�w�>�#��':�>���'� �Cs��$���"9��V���I�� ���	C-{�� �M@7�j�?�v8h��a��EaK#�B%j�~)8|�U�x�=e��RkW��W9�<�N��)����ϔ�:�'���1��i�)4��<�m^؅����SG�X�-|�?|�WY�Q\q�C'��$ �	cG%,�z��h8h���=1��C���U��u��o�����Ycn��e�tL�H��期*���#���3�9QT�\�Ac[Ĳ7j݇-���q�{Q�P}8p�3G�Oz�M�O:�L��Ɩ��	Wk`�W(/^��U9X�˖�� 7�'��\���J���+kpu䂭�E!lE*\�EC\��,�EOD��*��K�X��$�#� WC����m����$ao��#�z=q{S���6 6ׅL�AcH8��
� �a$��	�j�`A���!��Ζ��-�jH�aP��k �#�ѮȢ��xv�Q�'�{�֦'���9')OA:�jqg#H��*GӤ�L�Z �Z˴�u��6�n�w��gς{7s�V��0j�Z�s޽�NZ2��)k㬣ve�g��7�@N�͛"ek�	�W"�h�'�*j���갍9��ِ� ��2�3�TxO�n+9�݄wL��E:'��(����6T��s@bS8�J�����Y	BE�Q�amŻn(������9�[�,p��;�H!�w����*Iߑ|!�`KK���w~fϖ�}����@AG:�0�?��Mw��lH��;CD�N�.I���ة"��៽��Z�wq�Qn��T���])l��cv�i�z�Oޏ���"�����emإnQA����:�c��q�!lQ*�{�R�ʲ8�*Z��A	���(�x�D͢r:�Wz�7'�M|2Hh���-��.�U~VY�N�[�:�>����(E�`���#�=db�9'�&�����> ��X�@sL4�}��Y���]�޵�G����#p�����1⃅NcF���-�H �BY|��F�δ6$�g��5��t��zkQ�;ڠ��KT<z��0���|l�J�t�����~���k��/?{�����'��=������w_>����K^?z����K_�|�������_��W_|���/�)Ј� ��q�>{�嫇_�| @�}����gKH��	@�7�w_?���"�޿xL�,?@m�]q��>k*5��G*5B�?���\P;�~���o��}vw�l���L�I��p�qb�r0`��
�p6�	S�Z���>C@٠�-jݓp�XZ1Q�$�3I�I8o�E��h���n�H�����`�| d��#����p�|(0��7��;�
ƇPj7�a�A2�٘�H�v�?���&[W����t�
 ��o��`��?��cI��E����[ ��^�	���v�= ;r�6:z�[W�9���sG�n$BA��AF'n��}���܁P��n�nE����ʭ7ݞ*��y�d���<�B�|���B{G�����U
l�E"�-�p���L�����]]���[��/���e:��pb0��	��U�~�H��(��9ZG�LM�]��D,��c�ޱj��tW8���e@�"��{�D%@H�R~b��QDPk�����aj�	��!����u^3�DM\�����Z��iGF.�f�����7P=�_�P-U��<gw��@qp�"j�IX듶��阹6b�H ��7���,� ��Q`���6����2U	���C�:���;V�-�DQ��1�#X�����z�" h�K��jT�4�ҍ�*cV�As5bS������LU����A�賶�d����ȪbG+�@�9a��'l�H�N��Z-��Zg�,���)���3��!L�Q�ߎ��x��C���Ҟ��yv�T�i�4���t��V��4��s��p�*�����Ԏ++ib��%��_�M�fsG�P�`GkW	���֍pΈh����sG���+{�0�.:����V���c��o<�u��lG��=���C� ��Q��B$�"���:���d�چ�	\��T���@x9�[NP	�S1�nܰ��=�բ!�8X <S��i���Æ:1�GM13��椭K��c�ޚv��i�>0��;�ړq��n�b���L{����$6���?��2�`��K�ٌ-�X8.��,k����_�V�,v�*�Fq�d\� �l��o��0�i���s�Q�z�h����쬯mο{~b� Y ��l[8�-k�m����.�"+����yޖ�x��)+��e���M
�ƌ�~�Q?�l Ӯ����4�iFZ�s�0�n^p�����u�0�-��&�=�mH #�HL[�����n����aO���zxDz�����sГv֧�	W}܉A�Fs���T��U����Q��	�`���-����"�Z���V*�GU�����g��M��/��2@��?���e>��i�?�(qT_9��2sw���h�� :
�t����S��:�M]���-=��n��!�k��ή��w��wt���]�g
��@Y̉�������ZD��g���qT�c����S�FN���]��"�1%�#H����Ҹe�x7�����%lk!kkľ;�ڗp��셛��(��]�EO:KD{���EPʢ9�z`����*ԏڸ�{�E��V��ʱ�Ĝ{�P�M����^��((��H���?�S[��؞�o`e��-��k!��,+����L0��[A���֓��IZw#�i�^�BAdQgH�*ad�� ��3��v#�@����N���G!7�"(H�0�U�`m�I�,� Ix�Q�4i�~nph��3M[&�������P�{FyIܴ�ڢw�z��R������^_�޿>͗�>�q<�u��;/�~�d����z����O��o���������͛���=����ۧ�
����^�������-d�<���������E�Ʒϖ^=�^?]z������x���W�?�~�4,o��	T�G�"�9�SC�F�4����J�_��?��;l���������'7SS���T�ە�t��Ǔ�S����P�\�}>xf.prv�����I¹;�h��ZH�ފlұ{ʻ1(BO�� ���2��)�K%���<\�	���`B��Ҵn8kc���Xsp��?���uwWOOpvVGGa��UEO�mg�,�J ��r�T��_?�W��Q�����K�������dE%��Z���W�*f�C� 0\�}��E;���S��-�^�=4���:�%��(b�(��ɷ�γ�8��Q����N`W�ȟ�T�����5�Ѻ�X}�А06z�K�{J}�e��r�,�����bq`�tb�d���ݕ<��Ύ��Ѿ[d}}E���0���
�-��~�yb�&b���6�a�#c�ET([P��s�kwʽ w�Fm�!sC�PU�9bn�s�&�i����幚������@����A:ij�[|V��CF7�줭-miA�tFv�ޒ��g�j �2HYk��긩2f� H ��*z�Us�v0��L�s!�+f�Ť+d���j5"|d�h1%cMM�Lx�HЌO^��'�
���"l�BC��U 4V	#�$8Z�,��Ai
O<�Q�A��M�	j�	���,$�}@�űH�g~)�xt�	�=�-v	�5	s���y³��u�O'����9�	?��8iqGk�C���Q׀�X����p���<'9�EP��������Q"�\��f1�`x����.����X�Ƿ��2����{� 1z�s��m�3�Sy�;��=]%�sj��J+9�����O�\���CFZ�}�)6�n#-D��V�EX
� ?�>a�M���ֆ��q��<�l�q�*k�mH ;io�.8�,��s������f�a)�]6�
՚[8�� �6l9� �?��Ώ�JZ�q�i�~�)�A�u��>�H�da{��Mp�G�+��'�-	����`mz�Y�nm�Ȟ�]������C�����N$P��Vց��c=�[gUzf������x��6Oy�Ȥ�����n�:�|R�Ђ]L�Y����fl�s�F���Ԉv������JZ�����X�K�k��V��Y� �L������G�J��?J�31\�*Ŗ����h	�a��p]�����!��3�q��%`|�������r�d��%���
�@5kw!�t�;�My��]��]d�*4w`k�-q��bk�)� �e;H���1p����N�4u��O7�	��JM���{�U��E��2o�� '{_� -��J�� Öƈ�)foA��p�!�-�J��؋�vĖ��	[��F�,��FO�	���5r�	�e��ղ�ܸ��J���{�����hH����	�f����>�a��������c��A;�X[s2e��#7!Zk#,%�20���$-�u�hK��O5�]��JD=ye��D ĠHjp�QQ�MuB3��F��u���k�����{F;���>��t��\z��]yy����߿����;_?����k/��?�u���/�_{~����էw�`����_?���˗o"��ٽ/��z�i!�<{xP�y���Y*80�y���;��.Q�y��!��4,����@)Fe����]F 	4����:�����/?��?���?|x����K��@��>���Ǖ���F��E�φO-�N·����M�#99����������D���7�݃�&!��pɟ�&��y��9����=�������-���cF�9��qe�H#���e�Ն3	�%By�H�I�8��CĉH$p����Q	g⌤�r�r1�A�7�{[����}O�=�B)�P7e�7V2���S%n�1Lȭ5#%��R���{�o������"+Ֆ�բBX�0>XX�ݗ<��ށZ���B��$<RA���VFǪb�긱[d�#eQCy�T�@�������B*
#+�Rb@6<���1�oآ{�&�l�,�p�Q�XХ�����$f�!s	[*��Q�X2U�������ZLD�Hq*<a�,�X�_}�#p�ф��L�ea>� b�%�T��0��� �)��9��Q?�p��Ӯ�IGu�^ER֊��<a.��J�v�0R�6�j@l��{~b7�"#F͕��Ҡ����%Q[y�Y�r�d�uH�����-�@�E�� 0�*�Eb�P1eOT|�Zĉ��'$�)���#Zl���z��V�gΦ�YGp��O֣u�����ԌR8�qb��������`i����EG	���M\��] �5'08��+㌊6���"� F-e�pi@A�
�ՁK�b&�q��/WO��#�rf�͈���EYWW����q&�rb���6`=���^ ����~:�vj�z�K��U��i�M�Ȏb�e/^��'vQG�o4�jN��C�pA��f����)��^:���!mW��_ 13�|3[������,��7�����vN��u@QA���#�q���@rpt�H��5�>?ޘ���f�o iT+�#v�gš1'���)g�v����3@�0+�q7��E�FhY�`/-H {n�m1�[����B��{9�'[�� !��l��
DA�E�9�����b���<��4L��3.�M�&]�������xgǛȜ���bD��ƵX�4I�8�j�s�-@�z���q�d�Mh[��zp�"�M�6��l�$l��a��m�Y���r�Ӹ���[� �!���v!
bx��&�����1tD8 ����}�dY�R�H��p�w��3X�(r�8z�k'�u���a���c��}�����Uh�,���[��/���Sl�]�#��]��+�V�����.��a����AO�u�v�4v�������ǅc�}�7$����b�Z����	Gc�ٔr5#�,@{�O삅Yl��%�i��,�����!�BX?>��Óa-p@��ig�ؕv�p�֎�(EO�Yi�Y!"g}O����D��	�����31V��0�g�@�
����>��1c$ϸ�a��Y � ���Fab�4��ELC�D����r"�C`�!��6�B��P�\M�&��/̝1�����FeYW��c�ޱF�g�5��)�����<>zpz��r�~{~�ѥ�Ë�Ǘ3o��~q�Ë%��魗�>[�^ܿ����׏��zxF�4�=�������w�<��E4_�~�����~�i ��'7�=������˪�3�w��$^?�����oh^|�,��ˆ�'�R���2�����������H���������/ߜ�����{������h��Oye��h���sѓ���φ�-��>8�DN�G�����)MƳ ~U�Wg㌧e��
��8�R����6 v�8�j���$�����ӹqx�MY��l�V�R�Ȟ$��)�4V�Ɩ	;��'���-�G+"��(&� Ɩ
��g���g�m���0�
�U�N�W��<��AĀ>�G��QSYwtKE�Z	������Ɗ	���G�Y�Y�2Q�W�%�!���	���h	����*���F���K@h�D��b#剱ʤ�*e����Xy�X�2U�f��E�Blc�%�bo�R�6Wbot�84XS:�#�a$�e�=G�z�D<�,1{� �K{�3��0*j���p� ��!C��������NO�K�#���2|Qce�\p�ꙴ7L����������q��H���w뼫e��<co�
�c �6WO٫����r�4�vT�8����1iQN~�� q&�����T���E1kI�V��1G�����ĝ�D���Ff#撤�&i�U�Xj ?L���Y�!����'!�L��,�*�E4�?"� 1S����h}p��8�1�YeG���G����'�7��z�.=�?8��%>Z���"���!�&���?O{� |�}�Z0t���C�^��1c]�T��4��YYEK�֌Dp���[��*pv�c��)���wz:���y �ޒ@_)���"og�����hM�P�2"XY���1�.�&��z���	#|��MY8�7=�J�[�J(�Ѝv8�v&�t7)�I�Yg=�T`��VO�j��ÁT-�8q�|U�Y��_ˢ��"��j�=�Y���Cʬ�g�뉾��| �d�]��E$X�>Z7��`A�����9�2Q׃��*?dd���s��h�g�^|\9��EYE� �������<���a-��� ͂,��\�gV�R�ž��37㊼��Z�6� ��E�Q2�]D��Ux�H�N�n�#��2:`��\jO�Pg�#DBr#W]�Y�9��1�ު��H.�bL�FK1�r�����c}����?X�@E��a-@|�@wb��K���6���0�(F U���<���W��/�޳�ֽ `$�:z �@>���֝o�����W�(q�;z�&��R�h��X�o�iX� ����;T��jAǈ���>�@!>C�����(?ҬD�,�����D,�L�½p���Oa��iiw�t��jA�J�`[l�aGZA�ѓ�@��9�j����	�� �O	�*��
����3��r�"�i�ƪr">	�YVKc��&N`��(H7KI�J�ŀ�a���a�	"7�g��D�1�WkCYFq��� �P�&����>NO�|3��(�F�٠]���O�YV�5d��S�&D�	sHY[���(�۶��y�P���v����,9^ܹg���nb�`��q!b���_K9�,�.MOܾ�y���ׯ��{��Ww�-�x����o�yr����O�{tk<�{~yi����K��ܻ�����7^>��G�����m�޿�슛'���Ƿ$^<R^N���u��/�٨RCF�/?�^�5B�!�S����WX�>[zx=ss�3=ї�v-DgC=��3���]�b�.�O��ѣ
����r������HL{[�e���&�Ȃ��r�_�c����:����[�Ci[e�R�,ҶԦ�u�c#6e.M�'L�Is@ט2�)C�ʔ��4�j�r4�,ѱ
���Je��#�L#�Aز���@�K����)[Y�^N2�
�t�Z����LEiX��#����iw���
L:+E�np��H ��((��ީ0��0�%�r(��GJ��� �l� �c��������.�Ӧ��H~|�  ��������Bp\��Hx�����RA�^&�æ�(j)H 4"r���]qk%�)G��S���a�Y�lvJ��!�J����K�]�^�2ݚ4W���2m� )C�0J���)K5�E���DY��31V�6g,ES��i{錣l�YDBbƉK �G,X�gn.E:i�H�+ӎ*��	k�$�	Gq�^�F�K~؜2�QK�Y"#J� �i��t�U�Xl�����1�����OWS�
�����D�P1�XҰh�k*5lE���E*.���Agaa	da����T���EH������->����0c����)6\L�#�8EQ
$� ��C%�S1�b���k �؊�	 Yր�1cYd�$4R*����w���'��C%�b��
�� c&Ұ���/�t�rvl���b9����＝;�U|]���y=���)��FKb�8���5^�ʣ�R=������č���ݼ�(?��w�S��@�v��E;��dU�����SV�H�i��@����̡����Ӷ�{5��w�YO@B��p/@",k!<����O��s�59C͜�b�]I��jfiAV���~�WK��C��eiA(K�>���Jd�n��'&�
�9o#`�����H�`%H�8,�JX�Y�=?�$܀h�5���T� ���g�lN��,��k��Y=�J��Tr�3Y����<Ɂ�Ԉ� �焃�� $�X��.b/.j%�^�z�p��	�Q~r� ���+�h60H�R1b<W��HG��[�z��.���lN�W�,�lN��o ����[ �^�b/���yvy�w��v8{�9��a!H���w��9{v:�w�z�?>X�(�qb�D}V�tsA�X�#�^v�d|� �у�%2>����C��o��E�?!aiX�����K���$Av.�RN���B�%#Lz��v�,��{E+�!m��a�#ʝ�6
O��
/ �E�Ch��DLe�HF@�����Q�hW�1=a|/��^Q����pŉ�� �9ᵩGԂp(eR~ �4�Q�HceHП�?~lE%®�����]LF��A��WEH�����
F��D�!�+GdH��>�7�>�5��k"��k)o����M����*go���z�h��ъ'��hʳ��ٻ��k�#�oL=�;�|����.- d��޹{7�>�x�����^��ɽ�Ⱦ|r�x|��w��M�\|p�xx��;��,]yz����k�	�4D5^�����ǟd�����O���������������?��3,��ˏ��������Q:qg~���Blt��;�	vN�N�G�����������y�j&���z�i��(���k��� �kq�U���h�XMM�F��N��R�
ؑ�z��dל��#���C�BG��[�v!,P��cW�\+��r� g����R��84�����i���~$��� �F�\!�BmB���b5RI�6<��B���vC�Y�J��( %M�qCat4?4�38�#0�}�@����H���
��0�v������B��0�P������c�Tj���]��������t�^�m�XL�[����3�*v�=D����c�3�p����$fUtaA٘�z��� ��� ��G�1�*+}4B��%�\i3f�YĘ�Q���
>@x�"J!�Ws�U��ÜsVϻ�)ʹ�:l��uV�8*&��`�V&@6��*�D��(2B���F�MXKc�"����05iW�^����0l* !c>�Y�i�6n+I:��|)V�	�����)a0�h"�B����1S>�ʪsiª��*Y���R��D��*8��k|>:�F�JY��<�W�Fۥ 8R��+D�+�T�ҌY�/K�6�˪�;N$^�<���R3T���D|�46Z)V�c9�H���L�b�٥p�1ch��J���c߅�QN��Q�.�A"2T�/
�ҘR#�i��v������9ѓ�� ��@Q��0�W�mt�/�#;陶�N�j���)\e�,-���I�EjY�"2"��`/| raUT�Xom�3\�1�.��W��p��6v�f�ud�Q�e�ِ������99,�4PD=B(��?F�i{9Fl1�`:���p�]��
	�1RU������@#KziV>�R�-=B�����P��oY�5#K!>.|h��>؊� ��	I��r	�A9Fk@7���$XJ��f��
;���g�Y�DM�����x���;�m��8�)� Fk8���k�Y=�^pM�J�X�Ĕ`ODz�F�{*��B�'�P��9KHn1�Q#*5 i��8�ǖ��`:0�p.���K(Ӭ(,Y�|�w���7PgQ�5P��e��~4�,��8�|�kT�}P�ھ��qe}J��w��g��{���m����ٵO��|��/���<>zO!&8V�4��Ξ�|[�p1}DA j7z\�;ѐ ���ѡw;5�4Tj(� �L#���@q��k>�̷�倖�����Ki��8X�;��&((�Y�4v	9C��hw	O��L��i�=�k�+��;�dʎ�3j��Q	�e�`sz��hW �l]O_J.Dm���'Y�ڽ�=�Q���s=j<�x�QDS�)�1De�`�\�,���D�7Ue,]j�E:a@xV�-�S�:��is5,�g� ��n@xҁ���~=�Ĥ��9��`�#f@�y@ȗ^��r8���s�.qP�44�-ѱ��Xͤ�e�ٖ�4b���t8����N��(�T[nV��Z�7�����G���H�v2���\��]�?�}y7���ܗO><=����_������߽_��Ã￼��ۥ/_�|�|����.��w�>�1s����Kp�B���4�K�gܚt�쓥�O�->�������W�?R�<yp�ѽk�^��J�=���_����~��~�5�����矾��ţK�o���
&��)ߙ��������Б�С�Ё�о� 9 �W��88�?���g�������::$��i���B�i>�Oď��O(�x����Q%n�ʉT�@}�c=�'t�)"���	d1��S�2=1U�����$j*"Z�����<@%%4�#ؿ��$`إ���_��hQN��9	���R�IKS�kV�r}��Ne9�EV�x��⸡8a,I�JZiK9�H $��[t�02R � ��"	k�X+&m�S�IUH���<m*����g(��	��i,���=��&��ғu�G�j�:���3��I�*��d̨��-i*N��6�/=	kiN�r��E-� b.	��A�X��vE#�*?��kV�������D��pQ�U�w�✄F
@x�DƊ4�D��ւd"�V2X�]���*j��;����r��2JQޛS��
ꇰB1��0�L��cE�7Z�G
��R=)��OF��qP84fp8�G�]�=D|��ƭ > ����h9�����p�"묜�8�y2��<�����"��)�Hv8�� �Z`ʢ,����W��P9���	�����!<P@	D��ME��W"��4�p���XGb�^O�Q�:�8���(/+u5f���sB7=b�d05�t	
@Hp��<��Z�!3����1&l��yw��T��(��E9��U�`���y�,�k�]5�p����@�#A�B�Ӷ**,<@�P��g52͢���X	�"9aA!�Ј"�9�
��d@�[�3��/EUg��D�V�a-���X3���ٜ�ya��VY{��o�0;�R�9�T��՗�)gͤ+��@��t �H��Ȫv��9��H?W5\r��ʋ�$Ҷʜ�9-b9���(?�bbD�A�fAp� ��|=>j
��?X8�/k�R@��V|��R����������
���`b�(0X�lN�W(5k��p+dW�g�vg�G��UsA7�mߴ������E����m�%�]�-@�'N��H� 8\C�+	�����#6|�������9���TDm�@Yr�>��p��H;�v���O�)�V�� ���$d.ˉT�$lU�9��[	��z1mL�
�r\z�nH���;��vW@������I�@��
BÈ�q� c�I��c��"�l�T�56�)�{�c�Qe�
�IsM�Z7��6�B���B�	m-{c��W�-����j1Uj.|��O�������\�K����+xV^	�}+���Č���{w���X:�,��kg1Ҧ3���c'w��(4w֎��<^�w�l�X���:kO�kp�{�o�h�|&j�ٻ@�՛��'�ݓ}��+���|����_�ܻ�r~�����k���ξxz�ٓ;��?�w���7O�P���NB�!�R�_���?�����?���_����������?����x����s������xg�w*=qb*xl6rl6|x6|p>�,�����᳁#`a�0P���TjV�-R�i&ݍ`�keW^�(!i4��4����AR'��U=R���D�RM��2��3U*5�|U��C!E	!=Hh�
-��u6�F��C��|ȋ��
���� 	X v�h�-��h�-Z��"X��q�GJ�"�B���:5�dH��HS�^�J���҉(g�X��������B� �r�+����.�e+�{�4�~�K;� �B�ɢN�7� =��GV~!�T�_0 �P�����?�(�u��@�T2U+�{�&���>c�35��E�Ś�X�F���-��Rc�@���Wd�&�-�ʏo&^��%��iu@yo�*� ����p!b&E����l���i�Qj�Ǹ�ɩ� �X�2)Z�!� �Z�)ѡ��!+�Z�'�v\��"��2�#����]�J1T�^z��V%F��Õ 6T,'���P�صb�`� /v��S]��W.��Ui����꙱���,���?�0ko s��yg@Ш�A=%��Hw(2�j�T���$�ōE�J[����EQ5"��ѓ��q��CB��.V�S�n�.IT. �z�W58�fXD����tB7"*�V�/���P�vQ-�B�� �"��j̭��K�)�0��z���2u$�7����]=���`�[��tW����J�E?F�_�Ԭ�	aR���� ��G�nr#U+���J� �Z2��1<�%x���X�ߨ��`b���TjւJ��5�FC6��L���h%���"oOV����:�� i�b�ӽ��v�:w�5Z�e}$AG ,R��+�v �?<(�m����b*2B�!�!�-��NAgE����o�/��K�?M)�n��S���A�V�U�6��C�C�T�P��FPɕ�_���2���J#"*2�rڃ��G�Jp� �	$�,��嘗�q���$�#��������h5C#$�Mk2I5�:�nSf�АMX�OY��������@g�m��Qe5��Ǒ�4#�*5	�Y�|#�z��{��*
7qc���s�������BW�.��� oOҰ;�w��l���stWX:*����ʌ��m]u�����=Ξf��^�����C�ჾ��N�4u�Y������6�h+��X�Z����@:f97X�u������?yx�œ�?x��!��5���h��~��?������_~�����?���?���7o���9{mޗ	Ƽ��)����љ��5����0��Fk|m�Kj��?����;�V���ݪk��k+ B"���Z�e#PL�#U+��G��Rq`""&�Tj�Y�A�Vv�BUB���A�L��F�4�_��Hn1㴐�����~ BM�#%�k���Lt�V�-��q֪��!˹+{x80���_���le5u�! 
�,�Ӈ6�>�5�	� ,���F=��C�uc�*UeĔ� �Q>aͲU*5�F⪚�,d����n�cM������*+8�W����	��f�X#�3�e5�H]�#��BE��R��~{j4*�<�o�T���f)g��h�A�P�x"0Z���ң�sG=��(���kV��i&�@,VQN`���<8[p��<�	���c(S"W�^���F�jG���hE|��ǆ�zYt�+��	��W*5�<� q,/\ʵ�<<��/�S��4�p�2�+k(P�!�FCg=Ts$f�:���7,$�Ʃ.���غe��*�b1c'KIN���ȣG����@u`���k�s��.1�q�5Z��蛣��<I k�Er"i44�!��k ?Q'j7>~���Sc�k�Z����RB�ղ|���W���)����$�v�g��␵�XG��4�*�}Ђ�)��9\�50�+�W��Et5gb���F[V�<mj͞0�$�����S!�U�.r�{�q��^�"��<�����)o�ɽ\E�}�B��ݓ5����>�hXJ�#�ݵS�4Ύ���\S�_VC�F�V�,"i7��+kjԎ�ΰ�j���5��mb0��V��Pp`T~U�/L\����ȁ��ߑ���j}���D���{	}��S��_BT(!P��Q�3_�V u[ :��V�ZZˮU[��\4H��@r˒Ujr�@H"��k�RA�P�5���@6iP��*��Ԣ E�	�7+�]2f�7�\у>�3����� �c�]�|�*��V��Ѭ�Y�p�[�SQ̊�l�+�r��X�X�'Tc�ǡؕE+:�����_��u��8{�\}���&�p�����8>�������os��:�[�MA����@м?`��3����نZL�c�-6�a��L40v�|�K��<��٣{/�{����z�&��������O?�����~ ���O���o�>[��pun<=1��'�'��c��#ӡ#k)5�@shE�!�R�w	��7�� ��R+W���!�"p�a��GH$�&��R��{�^!�"��D�(���F��l!��%���Y1T$��6��p�Grh'`B�+K	�5�DyZ�Hǫ<Ĵ���)�vʪXF�ݽ�������,gNJ��4�?˲8�l�Hnh&��n�"�����4����ʢ�"�	�M�Ġ��=U��T*�hL�L3a�*'Ʋ����M
z���Dk��q�HbP�s	��P���K��VԄ5@��i�Ϟ�hA�����+�U�W�!�����BgH(���L#�h��! �549�I�	�P�:�!O�0��\8��J��ʻ�$��$���LD4ꌖM+5�L�sv���Ek䵰�RC��&c�ύ���PوFC�#1eS�e�Ȩ�E�	E�q(OWI������AҦ�3��hF�5i���r=sv������{1L�9�I����$�	�I  ��~"���K�0Y�� Ki���m�L�M�5��	�Y�,'�"$�FH-t�#i44�r
4����i[Y�Q�v����h������Rj�9KL٫�Rj(��X�-B�Ѣ��YC��՜EH6HӓJ�n��\}���q��F�i�P�h�)$iF�oP�r"ԙ�x���P$���,��@�Y(m|j i�2B>j4�۲tn�we��X���=�L˲����3��8(:�y��w�x�N_�.|�?�� r�ʘD#�(�D��$�5�4�o׃���F�_eV$��V�B�`v�hJ�"���5둊Es\yA���$�3?Rs���#b\��i-��Z$>�-��.7��E�e�A�:��GOV
YmQDڤR�LO��L#jH����F�C��"=�OD�UIb�䫃������P��t��C		�5��?�YK�aV��_Dh�4<R��H��|{�0G�}�վ�:�h��XS��4�e1�	��E-Aа�?�� 2Y������^�~�a��|x�~�ck�G7���ymq���g�����zͧ���X�￥R���Tj�y������Yo��q��{�'Ə���'������g�{�\�������h����{ʨ/�W�J�I��3n�otĳ�Z2+��־�H�iuc:�����H�
��L �gZ��	7a�Ζ�p��Y8��$��0��ʳND�4�_��p��G*���"L(sQuY醑P��`y�<dm�b֧��d��h��bW���/b}X`gq%JS���E�#ն�u��4_M�o�,�-z²R�"�,���[Ht���H��@r#�z%��Z�gE�P�(��s+5|�ܯ�X.dTD���	��X#�Z�b�@�����(=D �-,%�2T��*��U��J01\51\)��k�ר/�Q^kG9&0V�!O� v��;�g${D�(�4���)�Ʒ��ڷ�0ͷ�(�H�ǋN{�l�9w��Hq`Hy+Ap���'�9Q�v^-�P���j�7�԰�ڞ��_��x�D����c������-0��T5�j�ɉ(�er��b��N�渪F��úz���G4��o����(+�h� {NT�&�Z��Y�As����ѾG�VCr�E�d�Q%�E�웰0����	ߪ�������sV�!����qE1ɉ^�aV�5=ki4h>j4j:c-M��EϤ�d�:dS�R2����h�g"1eW��IJ��=�>hIX�A�Z"���h�G�V�}���.:��+�Eu7;��k�V��Îy"�q�8痘XYA#n�ˤ�Jʁ�\Y�QP��Of|`��/��D�J�^�p�d��q���DX�Ҍ@h4�3[���[�6{W�F�7-��2��j����he��=�������!�!��#e@��	Fڃʝ�~u9p.���ݨ����3Pt���4�T%���e��òz$7���i,i&,����\��K�	�jW�^q���Zˎ��_����$����MC6�� Q5�Y
%L��TN�,�A����ѕ?)&��&��ht"=�r2�P~��9�߸���7�-���͢�zR�W�lJ��r4�U�?�D�CA��l.f�	�BƆ��)ji�Yۢ�ֈ�E�Ԗ��K;g\GR�#I�a�D`lOа7h��������փщ������L��_�޼:����.�^�w�b�&������U5�i��_~����~x���͹�3���/�<u�{��|�2''�ON읞�f�d��7����ɩ�d�Ը�']��sB�Fį"��Z�W�3=���!IB�V �^��4�*$`aq�R��&��G��4�>�r'ww�E���V�٬R��k�� gb�ay�]�Nh9���*�Ae�m�3R1��[d��h�/�Y�F��V��V��v�m�w��{�x�϶`�N�Z����X�mƋ�<P(�����VPdu��.h�F^�gW+Ө?%)�L؜��'�Uξ�Oq�[I�X}���5)Ľ!:�.�#�HX빔&4VM�fb��?T�R�Q����e�ђl��J�)�F#�4�����]>.-��*��U�͝2E*2Tj(���<<�h�Eq*
*J�mL B-���l�{�i�@#�5J���
$;���KN$���$��^$�F������?j�2�$�U��JWas�z�IRF�z��G�0i��=�S��~���z�[�q0�G���5�δ��n@���p�q-D%,.��z�� w	�"+���VF��<�&$	z���%+ʬ�hW��W���h�4�#)��n�M1i[%�+�q)!: !�f?��H�
�}���np���T��%8�Y+��?ꍀ�	����w;�^#���9޷)�<���A�bE;���A��ٱ�P��C�C�����`=���c�^�ھi�݀����9et�Y�V�5�ӳS(5Zu�ш�R��*`��s�5+�bT�7Fg%��]��0�hD��	�>,Hύòz$��2�(�T<�i�ֵ�>h�	&>(�O9����A�����lسD��������h���GjQ��L�� !Eh;����H�8Y|�:�b�h�"=��	Jes�4�ʋĤ��tC��@�ZA�R����>jm��c�f�(�M�P��&{Ӯ�)��v�t��h��+L��L�N�}'�Q��������c9p�/�En_?{��w�=]��R�S��XS��?|��������_��?����}�|���K���x/����pr�`� �ۛ������q�L{���w7����2M�����io㤧6�N9��5U@Y���m���C�M��_~�ៀ�Q^Ցe��f��葪��T�Ç5ӎ���Q�FQp���I�!$"�驚E``�D�L��=
�.�Rj���@r#��L]��q�Ǩ��bx�<^���韘�!���	d��("������([ᯭ�r�Z�]��|/��m��Z�&з��,(��n��(���X�P��#��7%(��y���v0܂�]���(��R31�k$Q#�hs�b-�X��L&�O��geO�w� ]�8�㖺��!f���Æ��hM`���T��2��P�4%�P��Tvm-�o%���K��v�@�菋��֨�+c�z�����%�'0��h��Ю(���e�`ap@!4�H6�!L<J@t���+>u�>rU����f��=^8��F颐R�"E�z�|�?��R'�a�H�'���x�Q*.��PD��ha����q��B �vmmZI�:�����U�F����)Z�<�LV(�]��N6!��^� 3�{h��6�g�z��8�h�"�e嬓>ܕ^�I���e��O	���"j���֩ET(!�	���q�|�q�8���� z�C�9	���Q�w+�	�#<};ܽ�]=ۜ�[��.��ӳ='��,�w�f�	!| MM�b��{��!���HH��Z��O}f��j�\%ֈ�䄺�^�R��k�D�D?���Xӗ'}bb9�5 Q�!�(K��ȶ�p��=�(��[	�|�^�a���.>i����7���Y=��Z��aՊ��*����[=�s�`+�Xˎ��+��s"]q�M �7FDz��F�(<����#�u5��hYNz�MG�K� �r;>V�����Q-��EG�Al��(K��M+Y=ʚ#��X�������2'����"��.^{�0WVf�d�u�GEXi�?�*u�AV�)&E�A���S�֌cOھ;ekK����3�c)籤�H�q8j?���L�F�''\��c~g����ۋ��]y�x���[Tj^<����7O������������/?����O�����?|���ң�3�\��ޠ�d�y$�>��H�������2�-`�K����P�YK�!��\w�G��!�B��o�+��W��`=�g3`��Z���K���A���/�FD�n㦐�'`[���eL�����Y���,���O"��{%�������?�	da���9�������#�שG�]��+h�=۰EAa�'��A�v�Z��EXDH3��
ʟ��Tj�Ά����f�)`�U��T��c����ZO?Q�X����.V� ��s�Z�K~��y�
#��)��t���4aȎ�c��Ѻ�r�`���pэ"��G�Uz�F�2���Qj�8KWMRj�ǋ�\�i�Q.�4�f�����,�-�إuP�Y�ڨB��[����"v`-�g��(p���p�3K�����t��c�O�~?�V���nqÒ�RÛ��`�����(+;ԩ5E���0a( ��`>�1E�@U9�ֆ�rOAA[����޲~Q9�Y'�����3+��	��G�b�� ;��Y-�KX�eqE�$֪ٜp�Z���j,3+�UQ�QH!�h��H��z�9��MKmm���N�pt�XTƸ�N�j	�t�c�ğy���#�ࠇc���`�@;���ەe��F��L��R��ޖIqX!�ݳJ�H��o_>�I����B�C�� B-B�����ڷj�!�P�ѣ���2k�_�4�(�4�A,����k?1o�"��%B��F,+bE d*5�i�RC�!���(���J�V�����:l�D��&��|Z�*����Z$�
� �>崣]�5�Eb��&��Rx#�/XztN�`_AX���(HB�'ax�Uj����n��Yn���bM|��b�V�Ѣ�9�ٮ*5@�5B��ʎv	������*��u�W�tH��V��h}XI��*^׀��2�Q~��Kٛ']mS�'�m �ؗq�8�g\�2���c������ęt�3:��6���/��>�w������z�&�~z����'ߪ�����S�L�˟����Zb�������?���������o?}�����K����})���x�{"��VQj�\S�m�Ь�H�pM�U�rV��� �ȬW��leI�㭥	��M�d8)#"r�����¨-�]��<�l9���Rz���x�bR��e�@�+��g&b��+��@�����V���Ǉ
Å�R��';�-ۿS *�8�GL�P-,�\�� �����&z��a�Ǩ~��mC9��~�G[��M �	�jW|��r��_�n<8�$9�	�	�EB��dY�;dD��jJ����Z;C�&a�,L;���'�M�|� �x���昽)d��0TO�U �F�� k�?_���m���A���NJ�* �z��5Z��R�c��^��+�3ƍ��0�nM;Z�?�nL�Z�\�f<������1SS��55�uaCM�X6TF�Q1��o�!��չ��N�K�.@YtR	b�(�Y�W�b��W��T�=��r!����g�@x��o��U�骕7� ����]=;�G:�%���<�ׂ�>}��C.F`8�bpF�ϰ��S-|b�Ȱ��F@>\ê��- M�����؍�w�� !	4+d�=�)���� '�l��@r�հ��� ;i-^���ge��R0e+A��,�4惄!�M!}��cH�jؠ��&��!�\�Lm~\��c6���P��%##�D�>�2H�Q�dG?5�q��Sn9�+e�¸��:;��B����ݻ�ٳC�7�����*�Z��2��<6�M]J#a=��|�sK�`��J6Td�4:���Y���>�p z���Kf�d�ίIW���:�����u��0� �7�h���]�ţB�sB�C��	Z��x8YEA	�J���¬��E�S8l�g�E|n���n|��
'9r��� ���|]ہ�G��`7����>%Dd�/A�-k��7n���s쟁�>�GrHn�S�B�4b.|ؐ�n�&a��t �썘 e}��`�q$�8�rN�&=��ޣ	���T�y|��->1|�l��b�����o<Y��|�Լ~�[��?XB��y(Y����?H���ꋄ���������W�߽s!ye֛��[��=ǩ�d&���Ly�54�4��J��L�f���JMB�ͤd%�(�M�H�
Ȋx�3���s���z����\(q��i��Dm
i
$��4\>C(�(Ki�7����_ۦ@=b�,�(5BT�?�lD��:�Hn�M�V��r��/����RDd��eU.(�����ϊ^��jdP�h>�P��g����/D��;>p=s����#��=IWk��ZYSÂ��5���FN�we��q�	vW)���ݝi�����C��?��ӎ&�ckʽ��W��+���S��I���}oҪ,�LX�A��6��÷��xw�U��2����~O�N���G�5��Qt�Y��(��TNB@��h�E�����F�"�=6\�E@$PD�@�p��No	���8�7��6�`��@͑	d���2��G��g#����#?�ng��Dܹ�TSB��r�5b�/��Hg�l�q����W����_r������0�]DېPjh�8��.�>v�PL$�j=Y�֮ET(!: �mE�&�'���؇��Z��$�Vj��E��)+#�90��!93��dqHx(��!�H�_�N�i �m��R����i,��M���c�� �6G�h�ӛSj�A�F�N�G!V֬>"|P��7���#��9�������"zX��Bv�z�+=�8}D��R�E6�QPB|P��6�h�݀i���/IBj��^kB��?�Ԉ� >%8b��I��.㺍�����h�-��"����'Q��J�E�_�?Ϊ�V�(�Qj�ҊXӖ��O�g�R�Ci����P�}$�=��
9O�v'#W��Χ^>R������-�ۅ�ԀM������"���O��8�8劺���Gb�cSj(�d5�)o�F�qW�]��4Ig	H�����uq|c\�\��kjl$F�r���6>�+6� A#�`˽t����	�o�l��@nlh�~d(/1\�U-TL�VI�8b��%�h�H�S�u43(,A����RbFe���.|8 �����
��[�0�c������M�(8	\q���@r�ծ6�����Й>"��Yf��"Ҍ�=� �p����V֤�E��rA�h؆�*��]=�3��W'nMu\O��9�~��ṁ[�]�����i�%�h��b�(�S�Pj ��`�o;��`E���/��q���~�e�M{�
�g�v|Ϥ�-eo�r�U�KH���x���΍���v�r�������#"��b��oo�Q?1Rb��f>��sg�K6�Ь��Z� 4�b.�lP�Q��n�ڑ��+5�j0p4��#E�Д��V
�t�i�]B��9����b�$��_��b�GK g����F�#�����1e��NSʊz6��0c,�4$��霈)��itC�s�=�:���93_�g�$�KOڌ�n�Ly9��~5앨0c) ��µX�_��ŧlE�ғ�f�a'���	)!}���z��~��G|��:�H��`�R:e.�SWA�_��Zî� ����K���0y����h��o9���(=��BŌ�?��0�*�zw�`�N��1�Icώ��woޮm�ӹ�ݱ�8;��������7}����`!�� Zui-��R+2��5�EH3Z~Ś��0��Ś-��_S������n�<��'��>���>}����y=|EK��
�Eb�z�cA�%����F�}U��AZ2�'��0��8R7hT�Q/�M!�8^t��m�F=b�QV�7I��>��W!5'!�,1^%��7���h���9�����e$7���I"�⨩�̥٧�U��k,5Ikm�Z��5��Mi[s�ޒ��el�Ӷ�i���kʵ?�9��I�N�]�-�{R������/^}~����[��� �'P�i�k6����:����?���?{pu.t>m;;<�CQ�Ѥ�X�{`2ph��Ԩ;4�P��j5M����LQj�Œ4�E�i�f���5��zd�c�0B@�F�2�PXXJ�p� �9�,j`[��=Έxmo��C�j�RC7V�V�>�n
+�V�Q>��ӕ������J�*ֈc�"�_��q �v��	�r"�	$7�Z����'	�������L5g=������#
rT��J��r�����g3_M&]-){c�Z%q��l�L�UXM�qw�ww���݂����]w$���;�n����Q_}V�]}��SU����&����C���c�B���,d������3�n�`=�
'�q:���NErrh�;^+BՙJR�z���K)d�l	�U��-�3��̍�tAT��� !��죩���?3uc�G�'�ƫ����`l�wʖ=������Rk�H\4�8���l;LȚ����w�}jL�2Y�0� �f��'dk#�w���!~�`�!�2��h6��f�Gf�̻�dEթ_1SC��ǖ�dh�J8��p�T�t��~��u�h�O�0�X�.����sfu��c �X �tc�njj[��Gh�!l;%���[�{�O�uD~�,i��,V�z(����	��N#��3���o�7�9��H�X�B%F�ج��,1���k�h�O��~��(�&0L��"$�%�ki����x��_��м�G}O�Њ������x���k3^��L�5^f5��4�T�zV�q7h���ԫ�m��&0�XY���FP�8.�ɿ��1`#�x�>��$���E��Z1� �b���Vg��Q�U��F���6�؛e��M�[�$��,�l���ʃax�`gL��oV�SP
~P�UX!�K';���	�ק���:;�F!���>����i[���� 5�=�z�t�}�b����6a[�2�ҹ��st:�x���&;4����T�ė����]ˎ��.빉���j|�����OG��[�;9��%�ڕu_`���3Ћ|��7��~_�Z ��?����= ����!�d����A2s�/]
.3Jg�V,�����3�k���Ӈ�����A5� ��+�E��#gn3�?�1�.��E��hV�.��M�+��k+���T���,�x��?[��S@̇����nL��j�-�{�R!�t��^�G�z��LZ��W�}�1���0_���OA�
�}'�K�:bCD�S�Gk��nB�V��?-͵_��P~PQ�>9�����^z7� &5�:�p�HD��z��s�%2�Y�������M��ЖP7����;��ڍ�� ��Tb~,Q�Յ�2�VZ�䠺���+�~����,6j~���|¯��X�a�_Fm˅B�K.��	c��ۏ흖`���'C���t궄�u���x��?���\_���ā�a�ޫ̧)<�/�&��y7k��cw���T�N�lZ5嵵װ��3���l�r�ns��ŤW����[�׻��:���5"(��:ˢ�?n�@X|I�:�/�S���m��p�J�D�:Z��G�B�����,�t��cu�g����!��=��|j�����G${#(�K%@n�-���@2'�4�W�`��������|B!�y���^�[�Z"�J)�#osNa�U"pe��D#k=�$�ɗ]>��e!0�+�C�[����F����_���sr�'b4}J�a��mL�x��|1�N��/P<� ���LK,/��q-�Z�t#����ku�<O`����H' r�=��"��|�Gv�@�$Pj�(�[j�y�	��D[��.?Щ�e��IF��^��U�}d���*�2��?�{���;H���Wr7�#Ua��%�g)��!���c�-x��b�%��H����##�
�v�h��&d�8�~��ڸ*��p��$q+Q$c�P����p�l��☼)`\e��Oquu�nE�`��NŨs�<Lc�LLˁu�����9� �WRq���H��~?�涭W�#[���Xlo��`X<�[{�"zQ��_�;q��<�!�!&�Վ�Ռ�������_�X�% x�t$_$���!������ž�����p��^[�4Dep'uY��r$��(VLm���Mc5��u�SF��4g.�(O�@;�PJ��l�b�$�^��|�\��_7��y�Y�}(�(%]+W��ڧf����]HLo�[��ⵄkϣ j�J'�mW"��,��QlGB��sX*ï����4�F�}��?�L��b�.���:)�ᢚ4Z���}���!�J�q`�;Y��92(�1X����M���|f�v(�)84���G����V����52�i!<6
N~񯸰{#����߷K*������KeEU���`8R@�����#��%�W"YF��X��ꦿFǅ�a���;;����/bs���n��Z�Β�4�Z�q��^���]� �+'�3�j ��aB������e*rD%^<��'
C�+�x3��G��Y�K^��zQ�G3k��Z۴�Q��C'����u�K�X|	�6p��u��{�G�iIW�B��W%�FJt�"���EC�,��+��Ei�ّO},����kG� �5���&k!����>���[
��Ji�hRh�sC�1.K�&�*��|���Zuh�X@��Io�J�4��`1ח�"�\,��k<b���o���XC��@eHܐ�'������m%��%ϴ����*&\���>r�Z�g �̬�MtEuA"���a@��T�R�pU$�b�VQ.�㝮U
2v��k+���&d��x9ۼ�r*��V��H?9�-nM��P�o� XR>���d[)�[� ���>i&D�r�>`�V�xymǙR-�VUv=�q:D��](5I�S�Q.�fe�*:L�B�L�I~T�u�U��|g>��Y0�L���+�W�� 5�B@�(�r��@�Yw��m�ѭy�����+r�t>0�fo>)��2���S�_ @L��K~(���T�t���ͪ��44��Q4�*�Ԁ|qʥ� 	�r�ŝ7��ׅ�i8|܅��in����dnL�����+��L��������}#2���x=T�{h��� �R�,�/u�H��sr�3�ϸl-T";�a^�O�Ռ������%���C5��6~��:a��R��F��`�a�D3f[��QC�ne-�r�U�V�1�j��������va�M�Tiv�o�t0�*��R�,�xO������[�f���1 �\#�R�P�93,"b���,��p��j���D�݋D�\s�@���)��Xqa�_�4�Õt�TS�2���p��C�TD�yA�C'��3u�bEԍ/�0��K~څ!���|dx�\>2h1��g�DW�������$�`tR����y��-]�˚�,�����r��M�%�\�9��n���爽�b�ďW��ݘ��o^.C����,�V2Ne���4��V>���"ݖb��C�)�͂�/�T����N-	�Z8Bg�ԟ�QDm(Lj��i��Ě�El;����
��٤Iz RM(�4֪)�-�Wg�;����3�����>��,����32�}y��ɶk�w�ղ�0���u��Z���I��s�l�Q�mz��3u��v�9�%��%���ya��\��}L���2U�	�o:�#��|�?�	���;�Zo�	ǐ����+�C�~�Z���j3�ֶF���� ��o�XS/%���W2�20���X���
���
�����N��k��%���'�/�9
���@�~��U�׮��|��C?���G��/y���N.����,���_f�w4�&m&���� �˪X�+�3��I4��-�s�b�O֚�G������������N~P��:��Y9���肪�u8D\(=7
$yx�ZrqұJ�q�li=�E,;��W$|�h;�: �P�q��l�\!�X�Њ�.m^�xl"^&��}lv�|���R^;Z�70�|p}����`���e�NݢJMh�;�� �֝���XL1;l�6�j��lȍ���������b���$0�O��}��m� ':����f.�϶����l{{>�D�}?�G.�L��#6�^�ϐ�j���:&�ԗ�^����:�_ʥ)�[M��1m������x�PzP����D�b��jS��]qe��`��C��ӓ�������jH�ev�8���좜n�b�X��*�]�ҥ ���U�=yp�t�ԆA�N�����~�����}/�f>�tV5gŸ���,���$JB�o��x����	h��ӫ�|�Ht���D��Z���%��'ig�pj=>�KFKU�1��ʂp0,�\�!�߼�rU��peΟ~�@�%�?�|��v�w��@!�"Y�U��"�V�Da�v�p���x4��ZY��,y����,�hy�D�<.�j?��/Gӗ�n�-ܰ#�eX*��L�=.��<��{ځ��&<=<Y�����[��ZZ�OMB;=�m����Z{�% 	]k�ɖ�h��׿��b��%��K�X����{�8}�cB�W�L����4ټ)��"yv�x�[������8\���;��j�Μ�n�-0��ufI�5?X������I�'���p���b!��-QF��ѥ�heN/���{|��� '�Pon��"'������r�B�\d����gOn�J�J壼�ü�� a~^�?/9-����8'ttly�O� �T��1�>�a��S}An/�~�M�f�Eׁu�FŐ�,�I�.��8�cg��b�2�ݲI
*Â��SyT#��if����3�����r<!-�"�gl񺹃禍v�}���>K���j��Ik%S<;���<�G�L�6�i����t���ݎ|v��]Zj��O�pQ_�U3�_��HZ��zR���N�	ۧ�E���y9��hZkCŶ��'>Vu��/R�����T�~�I*&R�U�]B����G���I(֍��뚦��u�d�Em����?�w���nl��$��:���ͺ���@P����m�_83t����[��Sg�eP��S�]���Y3�S��,�K�ź��V����0�� Y���H�	�H�!��B0��Q���^Rs�H
a����D9^�f.#�N�W��_�z* HF�Z���t�*�Y6c�ݚ@�;R�H}I��M���Z�P~��'��)��˺��oڅ��ju�T#m��f��O�}sPZ[Uoo/���o�~����et7��}�-s�׾��H����n�����g#5�'e��Q�_����UD�z�G����N�.͇�<�Ne($��<�V[�մg �q��3�d}���j�cl�Qh,���^R{�8B$�����������B9���H�8/�m_�ݥ{��d�R��V�~*��͏��� 
�����'Y'�8�&i�"7�*���ӇCQ���-خ>��E�WϾ���&۹u�����M��@2.U��cm@.��2���3�'�g:�
]:�TC�4�e����Y�����Y�>dU��e2�<❞�cL��d�}��LL�`�5%�>t��mDɾ<����m��v�
3K��⿡p���1,g|
��#&A�pB�]#OMˬ����G���-�b���GG�����ݤ&����;�U\�H�Je�(��,� �:�w�#���V؈�������:�Lp����e�瞹��������P�_���Ƕ���uxrq�!<[]�p�+s�5+NO0�ʡ�8���G~����)�+~�	銂�����bc�Y�2��_#|��B��ؿ�~�x�B�%������~*�wp�Y˦�����>���9������� 6x:�n���yyL���G�F��`ë�/6��1�B��W!�Y�2o��=]�+4���X:o�*�����(w����~J��{�F����5����$E��{�5�ՂE-�00�詭E�yw�,� �޵���C�ѯ��k��:w�k���3X#;�`��[G�O�tC3�%�Y���N��\��x���/�"�M�>��	�Gf�
L��)��$����WFU���M�?�L�d����M����=y��(�iĦ/ۗ�qC�^���#���D�������٩�$YDk�IJ��d������\=ɆT����~ӗ톀/���v~�TO��NH&v�������N���9tR�F�C�<Z�@SF��:�/��^�3oNMo��v�b�oWq���<��~�<��G�	�*�8�Q�}�|�a�o�p����{�����ݤ��S=M∍N�s+j�%�~�Fw4��׍r���'�?�u�"���ݝ�ș��毶���쮵n����F���]k[Ŷ	��xq3=z^_����p~�f�vq4�����<��Na�I�@t���`��d^ў�M�'�ڝ�+sv�N���1�;�'/z��_xx$�����,:��}�:����&TP��2�m�=)w��-܎
��#g	&�����ƻC�͜�/Y(�!�g��TëG�ܺ|>�`p�e&T�
��^gʀ"%���q�����v� �
h��>�*CX�>�L�l�z�%E0'�Y�"�2��%�)�f����� m�G��i��4�����ε�������b։��0'1�6@�7r���۹��%V�No�������]�C&Vm�%���ҏ�R�f}�������k�[�O#�����~9yb��y��l<�O�F���S�&���z����q�G{WX�,?���0.U^��W�%p�����T1��+�k*Cd^Nd_��iP�����_s]ޭ��w��*!߷�J�j�Y�{��Nc�f�D.�L�����3|{!������c�¹p˂���Wp������H��R��V�#����z�|�Û�Լ��Y'&��䧕�hq�������)3���<�æ�C�i��%êB2@S!��e��*7-�Γ�ˋ���M�RҌ��M�kgy�!��EF����y/�еC��Q��Y$G�l��R��g��8�yR=yZ~�1BgE��;2D �{����-���x�+���Ut����]l��@����;š,Z*2���D�l���� ��5�A����r]k�\�Y���P/C8�z�bJ���Y�U.X�^�^���k��jFȸI���^��u�
yI�}��j��^>ܪ�? �-}�p��9*�7���(��kC�c��o�q�=\��1W������x���4D�fnF���`�r8�����h>_�5���o�y��?Y��S`�{[��%}Z��~����������@���?)�^�YF֭�p��
��.�(@�-\�Y�O��Yڀ�Ľ��/��M�Wk�< }gC��k�	�9��)zh�zj��̫X�P]�*j1[�U� �r����i#����S�-(8�!hd�+�c���~!�
�%#/CB�`.�/�蠍l��B���E��]3C Z�98�pI.�$QI��i��WG�v����su����*8T�Z@� ����% �Z�+�BB��yC�J�Z6Y�z�"��H��G~�[Ǟu@(s3�_5OT��-(�r.�ӑ���$�f5�oC��5�=����n΄��&.CavU�M�Ǐ �P\-����~�t�m <�Q?�᯵_�ݯ�}M��MDQ��_������Y�v��h�{7q6�_�}:�(��;Rq�)`��AjC9���bEΥ�x��q�@�y%�q��?+#Teƈ^$�7l��8�y#�(�:�7ӥZ֭���(4{�#�K�%J �k���($������*P"���س��b.�:r';���4�S&e!X�������eഔN��Y=��·q}�4���+"����}�*tT�_5�_Lj�o��E��*{};�,0���gY���|�:�Q���&e�ዜ�B��HU }�L��-q���3B���~� ~��t
|��l��s*�1Q$�蹯�q7�����^�u�j�K'�OYA�����y�h��b�%�D�?֠�I~�o� �����j��hj]`K�ԩ�K��y5玌�47�Q>�b>H�Щ7���{���Z#�&����3q�Q�YW��|�7ӀG��T'�~�E`�w�v߸�`�֓՝Y�&����+"Kg�K�òT_��2O�r�^?^�	�KH"��a�b�ۇ��d�˿�����Ek�c�^n?�Q�dgdUJ������b;�6˚�{v�Iˁ����o��,�i��VtpD�Kkɉ��3�P��7�2i�Mn��8��Q�5�P�n����+ϕ�>���O������;�����O�;�)��3�1�!YNw���b쪛�����s�������ܨ�I�⋸84^S��2���% �Z ��LL�l���|�[�{ytq����Y'�~����ֿ�F���R����`/g� Y���L'��AyLҥ� Ws�SK��K$�Q��(����:���;������Eȿ�	lidf砫9�-�S5�I2�֨��Ŏ� )�@=:Gw�կ��1�4�^�*�T�Z�>����~+;�f��<���{F5���P_3�iG���`e��k�u�o��3J���3E��D%G�L%�%�zx���ֳ���Ha�>�$z\�՗�S���@�uŐ%ƐZ�*�B��>t���u}���'�yz	I?�	�ӗ5+��̂CYj��Ŕ�1C�"���ؘjݮ�� ]y��=�a�BǬ�~H<�4p������!E?(�kc��iQ��݆^�s5*뭕��H�1�yy63� �(}����)� �ox��5:@�ٞ�ٱL��VwG�XN�%0��w}�:��d���ê^�+]��6)�}u���-��S�5�F�8j�J�N�	��W�gb��B����8�H����ԋ�t;�jQ pz)��3���_��z�'�bi��^E���I�@��Meo��
���Z0ح�f�P��&�>a�g��?�P���Uρ�J*�9�(,4���S����2l�.Ǹ����}o%��.�h#�$G1|$���>P�+���DJ_}cK�y4��Z�wm�V�2�Ԗf�n4G�3]��}���;����,��l�\!�[� Z6��quH�~5q��<���V���e��<�fO�Ⳕ��;�5�4��_�@r�͟�5�%�k�nHU�["-�&5���*���y��^4M���W��I��|{�ҊM�h�`��ζ(�r�/�LV��ѩw�j��췘Vg�O�_g���ZcM���k���̟��|���&�"��y�S��]�����*��y����n�G�~��(�=�4arJn��Pݼ�Q5�L�n�`ܴ��z�bݘ�
>$;xs���v���-')	 �"m��^��b yѴO�4�t	�t�k�Ab�����V漬�����=����_���S�/��Sx<qK4*�踫�R���_u���Ӛ�k��N�����\��D6���|[޼��|�����P�0R���Mj\,eP8�N�.�����v�Կ0����rm�Ж	O|���<�����,���`��[)o�)�w%�zӻ??_�֚_��W���ݟ�zMk�wp@B��V����+of�x����\����9��%�L�����m+�0�S~�j��q��g��w�F[b��[b�ή�����2uq��`��ǹ\�.�$m���SB���dK �H5�����0�`�}���������h���&f �<�<�*��T�_7�=I^o-�va�I/�˫����r�]8y�sSn-o�u����)ӧ�Cr���91e�!�+Bۃ\��I*Z�a��6�&��x�9��R�4�����~��oJ�( ť�Pe�ٚ���N�hq���BYۃ'�'��j������g�9|/V���k[z�xtu{�=����X�cj�;�Q�2��4�%������cƳ�dFE�	E~J���*�g�=�`5V �Q�֤e.�6��b�V;V���]������:$��/Mv5m�֨���Y������_��s� ؑq>�	+�r�b��_�i�Ŗ�2�܄�o@n��*:VD�C�!=���Ǉ4۠Q�X����c�U}X����b��l�����C�~}�!IC,q��-�Cʠ_�b;no�d�Ӫ�aT��\��q��	����b�����o
3#���h���D����-����4PQX{-�v�u �z�x��ӯ��n��p�����_�,e6�:�i2�O��^�r�z�U�s���d��]ग़����(���8�߂�1X0��h��';�|9��:����yBDY�Q����(oNZGڏ���D���_�t ��8��b`n�Ҭ�f�Ky�?���b����:�ؿ�b�F���ڀL�b��UݖE�hv�VO%��)=�R��}�(��.4�|8���gD]�^���^N���xՇ���3�~Q�o����'�O��V���G�\�y�۴�����P�\���	�X����k2�V��6T��~�^��aH��4�S�`�(#sx-��J��� ���dK�e>�, ��H�vi�W���w�j#���V~r�FX���u�aC��?��e���zghTlPkX�wlv5Ʊ	��V��5� �i؏��T�C�����c��������n����5�����_��)£��/��ý6������u��g��Cy��þi�W�k&���Х���ԇi�u�"�|�g[�?%�b}�ŷ�������?�[��\���s��y��W���>v����|��@� 3��|+?�Ɯ�R8&�|y>ډ�S}�&z���0`c
��	���s�E3��Np/[g)󭰘j�������w�&k���o�(rCJ�i�F��!bRt���%� wf�������i %����>�}�y�M<;��|�����J� (Qذa�?�\Y_M��Ǽ�ĦȲ8�����2�'R�b��"7��x�>|6��T���(l}/
/*���P*^j�4=[��vU�s�ޒB�ͫ����A������m|`�Ȗ�������tr�d���9ߵRBU����]�)e�h��a����P�(�y_�=�f�a���W&֡��<�Q�B�,
���d ��T������XQf�0�����J�{OV����P�l]w"М������mpz��~��9����V2puI=��u�� �~*l��(`��z��b��f��l�}Ml��0Ru�z�?`�ty�I�=�u&c�A��fcYӁ�����.1�o׼\Z���5x\%E5�eF`&Ǝ*�x�2�l�fB��ސJF�(��տ˦��Һ��Sz�g�j��Z8Lܥ8#�W��3�-XNE����ڠ&�qv)U��B�QL
"o�v��S�1��Bg�*��$��||>�(D��*�i
�X��8Б$T�΢ا�}"P�u!�AD_\˥
��Mt�	˚����oЂq�wXD��*��`��ym|�zY�n��3!/̒�<��#�T�>S�5�<�x�E�I���7�xŕ(��Y.�=�v�5_�Ų�t��z�G-��rMN�b��x?�O��{�L�j ��Q|&��'�\�{�%�u!~�!�T�/ݚ)O����/���;0�U��@��S#�ћ	"4a'��,��*R[gy�w6$�E�2j��KC�)`�+��o�G�o���ݟ�]�،�"���qKNd��)D�4LS�rQM}?��	|��q���y�]B�;�Xdj��U����U����;mL�W�����;oV��w������c��C�b�
�� ��?m$��Y�m�8,�,#��X1�p-F��@ֆ���7±��Z����vq*J���P����:+*�plxy�n�]�jh'�x���ǪC�|ۨ�E3]O��3�8��hs���=Ё�h�X*+�*�h6_]%��}j��P`��%���6c��ޥ睰���(v�p�2P�}+��N���B��h{��a�����^��ݴ&�q��W�K�_�L���_��^-%�~[L�̶~�76���j󨩠��g���j���TV+7�՛f�I쒤���PI�:ä��"���֛kN���
�4�#ǳz�M Y��?���4���AgH�>��f�?w�B���y��DV\rX`�1C�-`�}�A������)NzmUE��Pha0�G�ǃn7@��aФ�P�̓϶��	]ao�L�$|&)�p������E��0'־�ͼ0
�B��ͦz�$���!0����t�����ӏ�J5j�����Ο��qQe�W�#S�P]q�*����R�Q|�b��󪃝N���jf�����y�suwU���i��e6�=.nMh��Lr^!�'9�:�"j�+D�<L6��Z0�~��{m��YF�QLh|��R:��I�'�g��B����#��D|!��w�4�M]�a�|�<ٞq̛f�N���Vc��XAd�i��U�X%��8�ձ�)��Y���R6����e?�5ijs�4GH�+��EV�}˨�d~�J�j+(��]�io�N.���P9���a�&�
Mp�X6���=�;t]��+���a�X$��.��	ԂU3*Dˌ�^$1}خ�۶�ڍL@jJF�E���P:�b������9%�	X��	X�|1�doo�:��iEvi���Yp�(������,�Ep��y��P�z�Ց#o9��"wG�w@Oh�#����g����9w���un�b#��E�?��y�v�����?��/~�fK~�-u��  X
�^�i���HN�Il�8�=����v�u��^	U��h�b�A�N���O�!��|�����&����	xeW,���'B���F'�5�u� s-	Fe�f�^�V��K���έ�!8;��c��U`���a(V��D�^�/f	��r�{YG���/O��W�k*�g���ޞKy��A� Wk���UC|�񇖿/ܸ�˱�9T�"Q�3+,�+{,���d^4D����@re؅Ƞ�3�IT���X�X��md20����
L����7"<�#�A�����
���9g�S��q�Al��Gdqk�g:��d"�#���K�X۱�ҝ�:.��VF��v2]q�`��Tx�:��� �s�W��0Ł�Hwh��@���� W�{��NW��癳Gr��WR��Vmܼ��H,S`���{5Q��u��!k��!��{��R�3����bd;�ױ/1&z7�+x�m�w٩�Jr�B�
's��xp��8uë{]'{���mk]���5�a5H!��V =a+�[1���~J��I�H��HB����ݚ���k� v�'1S���QO�^���'4�؉E71�
;�p�yB�^)O���5�WS����F`О�Ա�~�C��xrv}��#C!:�ʢ�˒�ޑG%�f7�H�h�4b������k^EήJ���d��!w�]D�_Mj0�9����q�w����	����ZP1H���E�"�B�k��
�V#齃<*��.�󔠱[���b"��>�I�Z�7�(�v�v�9�3�_��?��g����U��47����΋��肇�a�t��m�~B4O��%�A�	�\ݯ��1�@��� ��gL3I�t�cq0��r��U��*hs���]8S���coW�f^�a_�iC����x��"��<C��m��G5ȩ1'ę���(*��8$�-�Sϱ����|D�4"*aBQǁeTפ�ږI㖧˜���Sx�Q��78l�����:��5��*��W����X~�!Jk����Ah;��C�i����"�DF���lw�6@g�7d:�3��5�m<�`Ç�`�5����y��ƄBa����]�	�3���U4e<��Ǖ/?�8�(�������͐:+��}aUh����S�P�V�rm+�o7�P�icxl���cCx��Ӳ��M4�
�ە}>gL[�)Z��c�E��0�z����M�J�����ZV��Q���	�&|��s٥�1���O���:A��<��p:�M�!4	x<�Klx��h��S2����Wuԍ|a�>�"�ӈ��ah�p�9��E�^[�B߭��|'7F�B	m�l���҇gg%`G`x�x�^�=oE1]0 �����']`MȘ���c�H�$+)Z1Ui�/Q���TA���H�R��9�*\=?�W|=�_w��6���<�^X/����0�t	��Q8��ro^�њ*�$/[�"埡� ���'����h�_��%�V}	Q*�������3 )�_q�"���
��'��nC�N��N���--���0�l���W&��d�\��V�Ѹm}4 �m�LKd��[ܱ]^�Jy �ƽ6�u�TuZY��)o��Ƨ�<���1�@�vg�{WA��w��-"?|R)��֌	L���@��^���}E��e���Hg�G��1�����?�Vy��v�|�0�πv�h,���I|Gs�Z�	V��ʄ^���E�NZ�%��YFT�IuS�Ke�u�~�~��d�@��O��3�ޞ%�A�3��옮C�С�.�ѿ��G��ɡ乲��ȣd�zn���@}χj�҃Fk%e�rl���*�5dy��gM+="�1{�Itb���A�
��x�Pq?�YĠ�U���>��\xR����!Ŀw���=�%����C�B�.�������ͫ�a�>�R�l������	��3-��LB����]�.A��� �	�>E�����$�9�E���-�Y�������@2|lF@�������Xb�����y�+{�:e�EB$�7�D C�6�/��!�|i���wP*����@��U`���@1c\�x�1"��K����EU�,�q�~*��y��~�7_=4$_;��k�:v�||cZ]k1��ƪ�
�hU���n�2�j��I��A(S�D��c��b�����3\:�ON�7�ˆr�z�����A���G��}E���s�u��Am�X6\�8���2��c =\PCn��2�F4kb��@�s5�]$� ܴ�w���Y��$A�UC��&��!g��r�iD��P$�����k�|��c\E�_����/��X���k�� �k_0�"�a�����cjPjfQ�Kp. Po�sf���G�`㹓��I��J�̅j��餧s��[�s�}:��~'����մ`��hG�q��H�=W8ێJ�K"���Z.z�O���'֖�����>�*O_ʈ�OYܬ��AZ-Y3��9$����99Ʊ���\F]�����E��m�p>)i D�4jLD���\H�y#wS3�v#Χ�q�A�\���h@'B��7�\��5�%�e��\�1�F�fo˲��T����i5��q _��3p~�L��i��z�7Ii�s�o���v�+k �[���M��"��#�9x7B�]���*�&���{V4~G���ͥ�����t V�
�]�3yd�3��'0#��tΥ�.A�{Di�E�)�(�i��l�2��T�����g"2v������Π��79�e�����V.z����d`狤� ��v�d{iD~d��ag�?������Xn���Qv�>��V#��H�� ��
��4د���N��x�����1�LR�V�� �f��&t8{��c
�P��ߦ���=��2��ty*2/����8Uv��;^���]��Xl� 1��oXG$��k?$��N�)�����1�X��H���A�γ㳑�}n��C�m.�⢹`�S�����&C	|Z@	����a(+�oa� ]a��C��W�$.�|��C�<��{r��^X)M�`��"$h�j�Wդ����Y��:�0@��X4"�-b�
�2Ǥs�n4j�l:�N;hYTݼOװh��!�%K�(�C��3�=�*��;t�	��(}O�jo��>G��ͻg��r�K ��A;0�!�
A�4�IxLQ���w�9_2��{��?t׾��'q]tй�m���E03�)����jd���ʆ�#�WD�(��raw�,�G�OLdՕjqKkΆ�=0��t^@�@P�&#5�2�斌~��7$|Z%M����6{`��k��r{D�T7��Q�_+��C_{�Y<��X	����Ff^��g�A�^:.�,�b:�vO#��k��g?�P�AC\��N��6n�����?� ^ `0�[8Itv"�Ւ7$�#�"(a�jdlj�D1���Y�-�ZL'��5�Jd��od����W�4�I�M��? ����q�JI��N���ub�L����Q^ø:�c*�4(8/��p�;B���ƍ-U˘�w'B���k,��:�`������7��ՊŘ�����䣭�R��2 �}˝�_\�MT��D`*�>.*��uLͿ����K`Gt�!0Pz3Ѭ�N��c��Ģp�cg�<�)��P��59Mb�2��"�AZ�_�6B����%���W�V��i��*�7~A��B\��sY%����x�D��"�+��G�M3<j�:��n��@��v��C��C���ǩ	�Q�rl��6���z�XK7�}Ž��D�}- %V-\�� ��.θ+;9Nsn��ާ���<�>=�4�d(�(���rd��)�"?ɖ=��~��$�����A��b8����6���z�^|(s
��Uu�|g�Fc�Zk�|g�U/��-�f�8����Pu�<�dn�h�ӡ>X�?D�W[]mqw'Hq/Rܭ8���^���J����]���;����1��9g�J��@y�!qI��>��=�,@�]�.d8+i��t�b�pn"�b◌����o^�>�4�ˣ��<З���w���4#����{�[	��	�@~?����~Щ�z���uԪ��t��К�<�K�O��c�G�ե� �a�\{�����t�}���?<��w�W��qN�84C8w��X�g��P-���1�pC� �Ko��˳�=�}��}&��Y��Y)��K]���>�a� �{)��]������l{eE4�����W��Ϙe6C�����Xap��_)oY�w[���I���|��M��� �F�D�I󌃂��y�Sm��������n:>X���b
��Kx3HRj��Y�~RD�������U�v�6��-`����6<?RG�C2�;��y����g�o��J��*?�����P�U�v�kv��S܎�A�w�/�	K����W��>k����D�q9!�X�Hp�q&��  5�HnI :��@��Bܐ.�?���,do��
�V|!mμs�8��Lb�:�gE�]�<�=�8Է����^6�
9�ܚ���Y�	�	��{Q��"Oq,ÚO&�ݛI�Zu�����:/H�����3��Fհn�a��ل��2q�@����[�",ʢ��ȋT�]ݴ1��u�?�Zo�Uܭ�36Ӵ����L��K/�.���}�F��
�J� ��	�Kc�psGw�Y�y��,�! $b��
���{��N!J)�������c�.����Z�'�ײ��]�%()�VQ?򷻚��1;;�W��sl�+��3�U6����R#%�Dq��g��㷷��uxtV
�'�Ū:)�Z��m��%���^�~�#K��_��盧Su��uL���n�?ܴ��ZrY�$;j�P,R�ؗo@���dU�l�7��do�*�����[��\�p��h��5�O��\��e��J`��ׇ׋�����vw��R��5
���5HHw���p��q�GAҒ�E�P��U�)��
t���F��c71#$ē5V��p|���Ȫ�����߅%Bm���b�M1d���;�.jO^Nm�
�=��La����h%�<K<k��ag{H�����p���Ӫ��)���G��������Q�D��ۯ�AC��룼Ǭ�F���Q[(Y�[i���ڂTg��ޙ]���D}�w6|���l��v�G��<�nzjJ�>�[[�{�3ȷ����Ҳ�ƭ����BG��.?n���2"��sN��~�9ܣ0��<��6�$�.����5s~\@/�U�?�MII���#+�O,�$�
k-�F+>��d���b[����w3�����pq��R.���6��rcd���������a�s����QsP`�������3��[yS>N;Ig�2�nE.,i�� �~cF��m���x�D��>cF�<v?p?ғV����37Lj0ЬqlO��n��L�[�����Ԧ�I���߹�Vsg�_5o_|����R���W+�*���sL����W1�׹����b*��|����f�bxي�}+ʿ�4��Z�jK�۹��S���W��ln}���F1�c��`@��{�c�Jh(�t�9^sEw��d�����_�Ќ���OG�]/`h�~�?w�� �,�����p:)Y����!�+�I�Uorӹ�/4�K�jWn=H�މKGDi�h9+O��T�E�+��)�E�5�h.2m~�!�nˁ��
7�,�|YJ�q�����e2�AP��4ȉ+�2���s�&�S5���C/r-|T� �G��	Ӛ�N��A��
R���f@?�rԡ��E+�ȷp��N�e]@�u�ر�Л�_H��EQ���L�(�a[eHa\7��M≾��q`||*�c��P��3�e5H�b59��Y�9Y�,��ClV�>�~o��?'�@���Q����0s���3@��#��X�Q�X�M�l��"�UpT�t"�7��}"�ne*�IH�i����`f�����=�, +c`d���W���s�C}�RMѲ����`�g¤�U�����U��9R���Zr�4�DR��6���lK�%,nR�2i|]h;�`�����9>G?^���jJ��/k2�N)��S�4��mi2ǣ�̼�~�9�9����i_��Q��[���h����V���-5L<N�E���o �`��aD�~�:F��[ܝ8��F�$)rc����f"x]�{կ�i2�i2�9ܽ�KM�|�,A��:����4?�����4=x+�6\������(#� J�?R�a��f����D��XuAf���ж�E2��DB�}�y3��pvy5�iJ`'e�� �?�0e���j'�Oi&�E������� bE1�~c��P�C�w�j�#70������c��h���]��`DT���a�@J��
�t0ݙЗY��n�������S	7�|��ؠ����>��	�~{V������&�t�pW�6���cjq�������y=�M���ǛE�<�AB����%(T������,����_�����Ǝ�7�G	2c�O��=�'�S��4�,EXcƱ¼�nvsV}��šD5\��9��9�&_0�$-������8m��SC�7���/�F��+��n/�*מ*/^�=�]v�'L����4�q�8x9�!+���p����ؓ�ay�68�xj|���ꭅ��8;.��v�-�i���֑����T"o���$8����Օ�ò��Mm20�%�j��%�
OB4�J>�F�m��7��%�\ �b�����a��Qыsff|�S~�Z�$y����?QZ�?8V��h_;9��g�*��t��Mq�M&���������3�� \�%_�$Y(\^�$������O����/�g��!1�T\ 2Y�3�ΆʿX�p��zў�o��N�
�.d�1�����Z�i��0��f�%�Kڵ��#���cB�S�����e��U�wn��:����]�`��F�;�|��J��)�S3,�j�$)"�ܞ֟a>�����ľ�U#���qbG��K'�7s���K<�H�!Y�¹"�'|4x{Or��p�EZNk:�hc��	�@��bJ�o�-֊����4���U1%_s%��T�{*@�����!Ѱ+�ǟ�A���p�?-~@���꣺��>R�6E�Q�τ����ˊ��7ˈ�� �����c{�M�F�u!ݟ/4��������a�_�5����@�� ��(�,���#�jy�
�1=��0�}jH;d!��5�u�_	��&�xQ�؏�Q@G� �U ��G9��]^ϑ=2��㠱����`�`��5�����og۔k���U�ь�M%���k�/�xb�O�FE�Ӆ��q9l+��2�t��t6�ø���h��/8��+%vЌ�֨��5�r'(�Z{��#k-�9� �es�S���_t\x���+���j?�K>�������ޔ���L�s�Jy����#������0�Nj1D�vJ�+H
��'J��Q���j��B�^HŲҙ��Cj�>I��G��S������#ˆy���Y\�a|KhC���H�3R�Y�`Kj+✜��.>����^u܌��M�&��^d9�]�aӌ�m 8�aOL���;��3i��H=��I�H����g�U4At���d���T�	Z�����"��:����6�i�K*1
�B_�ø�1�%����B��u�����(+S��}VGȜJ�- ¼�\&s*ϥ�\�H��ꊍ��t�z�gpD�f�=�����Dj��!�d�p��vƎp��y�q���?��7##���$���-7��A�ݼSE��?���c�+h�4�V��e��c'�ERk��j{���(U[ŕ縫��z����n}�f�vB�iB���2�����ɸ�
�7\)��ۗQ��(�G�����7�W�izv9��j���b�����X56S5�1]��\~?��x�{���|3�-����^O':���:_�E��_d��G���Yl��VNn`C}
�N|��[��{��8�/��<00�)�b��8��X����Q�X�z��+(��@�D|p஽�P�A�܌r������T�I
8{��nn�*>qkI��T�-cL�؞±v7Mƍ]��h���ȅ�f�������l��O�%B��r:z�~^�}cY���$��p�C�,���_�����$�-�+;<���b@���I�0�W-s�ZW���L:�a����������-�/��k�VǓwrK3lg?7�+/rED^W0D�����#@�=!gwe�:F?��+�
�l��[�*�8i�2��Y~��1yh��Y3�cs�ˮ� � �G��c�����j`GW���JS5�c�kw��DPm��@�������P9ڞZ��	��E�O|shF'��	*=9��o9��\aY���1Ix�#A8.a�_��PĂ��/����+ `  � �Y�1(����B����-�> đG��c;���U��IJ����	6�^ k1�e �<.��݂Ƕpp�T�)��d�b�¥�Me�:U�������}�acL���[Xm[ ;�`�P��C;	b�:���Cwp^�g�/J���S^��h�V��\�`�#QB�R�΄�0�v��z�}|�k�E���au��� v��]�3�����Fр���ζ�A�����s߇�rL�N�߿�.�ꩲE:�뱕���%=���r�$�~,&��J�4������dgUO�o�^#�CS���ƙ�+��í��Gq�j���WJjx5-�R>U����¥�>kX>2ʹ� o9��֭r뭤df��%�� ԹH��iu��N�	={�Jב�-���z/�+&+����,�]Ԑ���c�R�B!�NT���ˑK�g�2l� ���S��n&�d���Kǌ1��P*�:;%�)Rg�Wk���& B��]s�"B=B�~�9"Z{�9yeD9&R}t�ُ�*�ٗ���8����c.q���6b{�����ÅU,u�u7
��NO� *R#��<�c"Dbg�w~k��D�/,�� �G����,uoF�Zٚ�֟�5��5�pa���of��t`��e���sy^S�{ao�>Oa���>7#1�F�ة ����p4;�W�w�gڝ�W�㥝��^.�ݎv�����o	���} ��핌6p������],�H�?su���Z�H�����q4{�60�����<���UXLX�C�Rl �`�w�� IV����ܐ֪$���r�")�՝S��8���!���kUD J�2�H��[��ۂ����w����Dg���D�ǿ�ڀ���� ����Bѧ�M;����T�M0�3���"tS�ֲ�p
ѭ�G��yoC���G�-���UM`��G�+V7�.��P".\X�.բ���,�"rytz)\�wĮ�j!��_�z#��A��I��z8	�a�n2	&
���>_s-%s��#-���k/V��r�nƧs1׽{_��=�a�h=Π߸��~c�O���m��t?���G1�&{�A����Lw�
~q8NY�\���e^��wL�jl�DZ0sS����0yq�s�*{>Լ������4z�
��go`"�Q��Q��ܯ@�vq,kދ�g�X�H���ɢD[i[wx߂[�$�]:uO;��N����0�a�Aَ�.%�fB�q�P���h9�ç��Np�°Mb��ozZW9Ph�������T~cD�K�G��I�裏��F`��@�5�S�`��L:�vE ��{R
-�U��:^�.&D��Zd��� �
��p��Y����&��u�?�aK~���0�R�͐}��F�� P�.	R��fpN�
���e� �c�c�[���P��0|-j^�j�(�3�5��)���\D��ulj� K��(-V�s/MKJ�`�dԀ���HN�ƒW4��.D�`Y� �R�Vw�
�NB�����}/-�*���4�4�?����V�r��ѳ�.g�0Y��M�t
y���w1���<����mʬv�1�9-W���c�t(��іZ)5p���&bK�%�k:l�p�f�����7��N�c7z3I���Wr����@A�\���oC�O9Ͻ<6����Wv7;�N^,�-|}���W���z���B��ox�S��EΘ1T-�_�k��K��efi�`:ry&�1Ǘ�F��#|0Z�*���l>�D�%Q'����`�RL�NU���܉q壈m&M�6�q�B9�������?p���{��a����{L ��/���5&!#�*~o	y4� #KY~�8�4���YH�[Y�H��� �#�֎YU�D n]�(��)V�qQH+��I=P^�z@Z�^�C%�G�
bѽ8q,N����<58s+KZ2�� ��F	��ۣ``�F�ܛ�SQ��g,[���CB�_�z -��rn�������}�j�q���T���e��_�?\T;��ᆗ�te��R�D�����s���#��yG�cTT+R$S��#.�S.�C{��\����D�Y�#�;F�El��Y��$��c���c�x��+L1��aӛ�-��l3�_3c�2�}�h��`��1�}tB�̶R�Zfnes���`.v��n�����<�EM��m{u^��ݴ:U��?�7\��D^u�W�O���2�5����X��$���X8���^)${�C��=nQ���XW�>{�]*�C�؜�jcy�`B`-�����t�������
�DrkU�;*.�M��*$m�G�V�	���T�i+ݟFdC>7b��lo[�ʿ(����eU]]ve�`)[�nb�v���}�L��C�ɳړ�P9�/�����P�a�٤y\�v�C�<#�-��)�(��6�0C��\`�%t�à�^-�'�m��]M��dOj�5f%�����@TƤ���q����`]���r���Z�Ou	+N�T����)/}W�) QŷU��[բ�,U�I��O���9XA�+m��\I��W�ٳl� ����A�f.m��� Ygӏ��uy�RD�'o�����&	���1�ݝm	�S������03���C���l���o��x��������� ʓ����J��&7D#�K;#�SQ�)��B���=�!�Ŏ�d,�vm��ު0�K.F1Q�S�p�OC��rP"|�� ��eh+77�("� #��+�}�ۑ3�l�J/�2R8�y�_�֢��z(�.rZ�����T��=�%Cz�Q1��מ��y�˗g\v@:EZO�tQǵ�-�/1DTd��"N�2�yt4hv�F����1oÜ���{��z���ʈ�jmC��8s��K̂����8&ى�E�f�a��M�����?�N����{��
� ����	!��fm�f��paN��V#��}?b�4z_6���Czu&6N����B�SB���a�!�m�0�Lg�Y�|p���$�\ɿ���m���bd�yu��ɢ8�䯱����[l9ӈ.�M1g*��.=
�d@u
�<�~��Eƨ�=;PǑ	ez�q���R�H�&T���Y�@?�P;yY����l8������H����f!X�'8�4��J�5 =����Ӂ1����т�a�*�Or�:У) 2��'E!q�J'��`D���Lʄ�M�o�7�x�#'��b�L������]�#���/���ZK~��"������5ԗg-��q�gh�6hۭօ��b@�~D��p���l�^n��n�����%+�6ĹNB��_	�~�/G��\�l,ߥ������أ�G��6+CR�1�5{��~��҈�f��P�1�����3J�[��r���ف��2�-�O-[��vws��h�?��xo5����a�wu� �Y�_5�>;��@[�E<�L�t�̈́���¬�f_v�o��`xߒx�����͖�dF���0�;'���ڪ�T ٖbXtC�m�J4a�l�uY���P�#����B;��v�ŵ�vg���B�n�!	-�� ��u��׳T�Li/0\�S@��[�':G�sM��\k/F�f��9H�7P����"MTH����ǬՒ*�h;���zO��q��\Ձ�ɝ�[�
��^>��>o	���YU�=�u.���.�����26�|���ݵ���;��6�Y�1�F��y<�m��eQ��/)�_A5���*���?�=�(ݩi���o�.�ςZ�.�dAq=f��� S�y����.��y������H�DY�����һ1������B-n�0�"85�Iu�(/U������*��jW��ݯ�Cѿ����lT���H_�7�$��ԫ�e_�a�����]�Uo<������"��5,�_��^ەn�証$<H���o���g�R%iC��,��c�������r�龇�`Nr9���o=�,dDXƭqNNK���ĴTKׯ��������I�Ϯi�Yx6�g,y]�3O��ZP>Ih�$&������k܅��q��רh����ǎ]m�i��y�2�>S���|>K�b���t�
���l]Z�C� 3�l+>��|5ˢ��=|F
�������L =bں&>ĀC,XH���ϰ��|���{٘VVY)�eN�� �7���<�8Ͷ�<*Hr�� BM����=ET����^
��H*J���f������򽪼�IO=d���bl�vl�! >n��� N-�/®d��E~b
�s�d`PƔ_�	5,��:�b9R��Xֱ�&	p�h���2=@�"������iϻ�������dj}�TH�w��#�iT�z$$8���l�z��c�w6�1]��*ò-� [�\h���I<n����ѧԈ�� K�fǮ�׍�?۽t�*�Z�	�g%�;}��l~&�`�������k���k��'h��R��K��-K'/:nw�W9���������G5�I�x�
��Б+@��e$Z ��[涡�Ԭ��^�i���Y?y����&�ϖ6��K�����v���4���na�n��w{G��OV��N�vB�SO���tTS6UkV�]g��5�4U����T�f��*�\cQ���Q�%���_]�~gW��11����o����Ӊ���p�˄�� �l�f𥊾��p��1�@�����G~v'�AZj8IG�C�<�Fo�����mH��o;�#�N5���nd��ꤕP�j^/�b��eW���O�%s�*��-0t�uʅ��W��TPn�Mt�zX��xަ�S��G(�wO�@3F��P� ߉J�X�b�5�]|��!�o�6h�B�1��V�2����� y(�
z�2�]�M&�&"�&��d�n|1�E7d�t\�u��|�1 �4TutL�8L��������!�߱��F�?1	)~ ���y-����m]� � ��(<�_�����$T�t�7gǖ�wֳ� �M0�X�%��{��2鴁�t7N�5^���5>�&�z?���j�>��j����iO�p#������� ��X��� 'B��~��YO ��������?��c>�tN0���鿳k�+�6.�>"{/���,-����!�e%�m�n��n��mϲ� ��� �5�}�]X����_��ӕ� v�?�X����`��G�M�H�ɍ�PBJwdpt�$b����w�$Cj����Me���yGa[���)
{��#���2�ۃ��o�-�����!�^��������[�Oz���dȞ��nN�7M,S����P�"�?ݷ��Q�һe����!�\Җ���3緑X�͚V��[��L�l���Dp��xXC�Q��	Oy(ߍ�ΗɄ;�6p$�a���j��d8]D��塣��t͡j@ߛ�{tM����Ɏ�b���+e�u�\����H�ѳ����_�dy%���e[���܉ގ��k(cX���=��#�E�&{��~�zUgF�l��od��$���G�x����3�B����'f�h@,�i�5j�I-��U�d�>�d��"�h2ƺ�b��ȴ�A��T�4S�����n�~5���9�`Y��z�O]��i�(Z�J��ѕ6���Z�L_/����h������6�������~��0�,�/8�F���'ڴ��y�yF&�&�'[̇e�K�s#tV�6 R>�(&0�����=F�h"4��j�����'0��]6����I���g���On��:ű�������W�3c@�l��RP��G�E<�I���2�����{I��8��tO\���i��`"L�R�e\L�-+��d}���/�j�-Lcl.� �9�
�c2�֮�@I�P��[J�$��,G�%F�#��<��E�#�5:e��,���0��a5����2]�A�M$�ͨ��>��rT�|��M,��ܶu�K	8a��`�މ�,����U��$v�~���)����5�]�"6K
�+�w�m<K�*��p����v/���&l�̲��~����x7Q���a�-����=�L-�A�Q�/K*m�]��r��}�)s�c�uj���2"q4�j���L�'.�W&E�ɳH�̌�8t�vn���"7�o�Q>g�]7�X`l�n9N&s��j�ӱ;#~�!�T3�u�>q?��2������G8���0��
��"_�����2�x�X����	��n;Ƹ�`��AX�b=*۰D�t���V�2��f���e`�ۧ�;�-��?��Ӏ�����<Fl�%r3�ם�&7���rݶ�t�I֬jsHߓzn��U�l��t~�5u�g����Jz���Ĝ�ǍI����9�"v�S%R�'�<�qnN�;S���3��|��{�� ٥��?e�TL,�i���s�׃����b��?跋� �GI?9��F|a+a^�Ǚ�"_�BmL��	�K�la���ӓd}ъzp��B�w�P����MU���xf�Uƃ��M�a�6�#gi��5���B�I���P�{���AQKsh8����w���r�-�D�1-�;7��,����/��&�*`{�^{�I�;\7d��ga�����f�91��	��A�
��^W��l92s��i.-�1����{m#_�31[G��B^G_��p�R���������y�Ic��Q��Y�E��I�F��~�kf]�J]�Z����r����Gz������@ߜ��N@����4@�Q�e��f����ao������Ƕ`�)�6O�l0A�ԫ۔"�T�� �#����
y
YJ�ԔR�U~�[IW�(P���M}�5n�Knh�/�����r�z�@��w
�u�c��j�
���z�f�%��8�a�bj�T�O#����.�+���J&�}�u]���d��^hN��)���ZsJu�Sμ+�OpJ�L�:_fD�+����.DH�O&�����)�#K������S���V�^����w��J��>��d"�B��@�4�̓b�\Hd�%f�Q�f�,�0b:��u�y�k=L��l����/��w�@YZ���	;�0oLW;�M���zg��
���m�C�z��i�Ѵ�I'8�G��Q���ޯ�s�V���n_�*�k�Ή�i�-o7Đ y� ZB�����$t����_����0'7��gI�𦊕�)��vLv3�7JW�[��qc��Xn�F������&�ѯ��,����u�gK\]��	�򇇺NhX��ǯrpR+A�ιn�g4��(��[�J��iTw��c:��Lb/��q}�<�^�� ��_�������h��P*��aB�'E%��F�g�j�zG��I{'�>�E��
*�[q4m�8ߦA�b�k��)��O�k[�bo�y��<�,Y¤�$��D�}�h}�� �e3ܺ�(".���5ܭ��-]�`�P���C�dY��.�9��  "���d��
�j� �&��Ҋ�&1}3 �)���!ԊO5�֨*���dj��R�HU%������+ $�Q!�c�_*���=�����R�qW���>D(�!���&F�D+`ea%h-.�q*t�c$�9McN�#ҡ�H��rW�"Y�%��M����O�����P�|9���n߇*aS�o���o�Q거��br��־���h���5xe����@��s�iMκ�r�����I��=��Ջۋ�Er~b�Cc����~:A���%�v�����ե��ڴA�-v��%���jm��B>���p�3�蛬��P"E�K�f&U`�L`ڹ^��Cw~��d��������|�	Ɉ{)Sr�f��}k��*�~�m��Z�f*�͏-�ɺ8�>�¡�rf�����*�\*� 3j��W��ļR�P�QƼU�c�z�g�q5��#�D�<R@u���L˺ �T{B����y�R�s��Z��rkǝ�˜n2�㉡!�������G����Η�ܗ��^�vD_����4����/7�Ӌ^AE��ĽLo(>NŽo�{#��w���n�O�>�%�c}��8) 
��,�]C �藫�}f�"�����i��&T�,�͉t��&,��[u�U�����?�����Q#�U��d%�#�;���S2�$=�����S�)�봿`.a �0ƄLHv���vX2m�G(����m-��IH%��O���o���W�s��(z�j:�?�0?]���;/�C��n��fV�dS!w�%��|&`��y�u��^��CT~�\�qJ�����x9���ۘpy7�7Ҝ�F~qQ��pR�k���a�@2��yvv�ୀ��S�x��F]\��!��!������<E%�%�"�<�CM��҄��h@QIQ�Qe�Qi�Yq�yIl���f�9jğ�z��z!�2;��\�p'�o ʯf͸I�;��pM̐McL�x�	�2Bc�vLT�iu|�
�������_��`l�����7�����`(�
'�����T0��|�Ht�&��%�/���mݻ�%/M颳�e.�]M���YH�aB��vN�P)1�`�[,=������kBw�p�9���Ԛ-����x�j�:�7Q~ [oO:�~���D����G��5��^�������(Ѯ�]C-¿<�rτZ\L΁�R/��+�L�
,U
0�U�������>�:����?o��ɩ���ԅx��oB4cry�tJѶ�0O�Gg�Sс�0a��jj4�Ŷ��WW����Yk�d|�r(]Z�_4OꟷD)��^��	�r60�m���&�a�/�GgX;R��s��~���Y-�L��v��_��O��(� ղ� c7ӻ�l�=�j�zC�P��Y$��bP�Z�-�	�i��@�^k�3�l���xxV�1b�bdJ�A��|�8��U�f�6����5v]�Ȥ��i�{�Q`����.�9�_T>��ݎ�&��)R�^�5�T�;���&�����>gˇ�8EXe8'u˧D�~ϔ]P�*f�3�=��	I�2�,�s
S�z<h*�rE�
�,�3C�x�B�����[�_�X��;G^�)��ápTIM���T|���]tO}��D9���ZoM	I�2�0�����Epds��qꈈ�,�.��h�!�/K�9����dT\� ��|�y��J�YcF���u��z����#K=�$z�YQ��4qEd����l��8������`��T��5ڈ0&��S}u��Y~�-�#�?����!0!O���
b�J��Ad�N�C�*��T=1@�P�5t�������g��i[N�3k͔��c�Y�:?�4-�4����EN��k�o-�J��d�_#ɾa�_�~-������ĄԁŽu���M���㹹+R��p� u�BxT�H�c8��ş>q��D�e�X�W!���4������o��3�vQ󔓿�8t�>!��+�g�}��#�+�6�d�KQ8�ׅ���Ooo}����s����N�)O��=�)rE����Ƣvs٭�wfs����_�6�<o�(�W
�_��6�d��r_��>����m�c$��ʉ<��#A�Uf���z��}R��$�NZxAXMx�/�z��e�����i2K`%�9��tOώ�Aj%xqEm�;� �p�L	�����|Ut@_�Ab�T6c�Bu��h���ǳf�v�m��D�F��W~u�YMϝ+�GO�E\BK��Q?����U���j�&��f��5����0n��P��
����	ͬ�k�߫�|��z��*s���\��y��b؂z}=ǋ����[�ɼo89���n5
�^�Wa#=;v�8�2Ș�`�n�}�h���7��j��ʍ� ���9��Fwy;VjA�E�k)1CH�C8潛w<,��m)5`��<ҳ��-��.Y�&؟���ݳ�8��i��7D"mAp�m5Vv 3����OG)�_ul�·��|+c�u|�������	}'F�/�OG�~.x�Oz�U~��B�#�K�N���o7V��|~U�E�����(�"W�?I�ˊ�Z��P��5���*��jC��9�#3����`���oF�~�~�2M8S�>�Մw����a�&�ܹpNlFo��`IY�����Oi��ᐪ����TQh!�[!��ݾ��e8�4AF3�í&�4My�@3=Iᚗ�u��~Ľ�H��*)�+�"5.KKH|�p�J���b�B�K�Z���B?`�A[
�փ�L�`y�[po��
po���3w9ns�t:H;��J�(yG:�x� ]+�yc�VH�ҾN%��{}���� ��0bt�B�E�2bV/Eٲ��d�����i�}AR��g�'v
�G��e�Z��(���(��6%��q� ?���h<t�0��}c�����V�Sp���s&3U��R���|l:�;Zl5E4P?�)R}�V�W��l*H�3X-�*B��YL��B���`bg{�eC{��/V��ؐ�\2��&oh��q0A_4��ކ���;#�^��������Zq��c�T���e��g�[ωt��b���5�7Y�öT9�m�(���A���כ �1�r��Ps~ƙ/r	^�6���`��T�� �6�;�_���
.hX�rAh�ϊ��+O�IR��G���W���	��㹍��m���@����x�U���\���zt���t�b[��B�,p��.�R���
����R �H<1$}���9�����r�|2o�N�_O��IO'צb�L�x2�y�EIS>�U���	��E��Wue���ĦW�pNr��{�~��y�^)��~�e�o!x%6|�`����9���I�����.���T<7Ȃ��n�1�\r}Ym��V��R��A`�8��2��큸o���t�NT��Q78a=�6Z��q��x'��i���J��f3�W��5D�.���7A��Tuq�7���o
��)�}��>���������ę6��6��?�@1S���xW����`F�`<���J���9t�0��(��<��OT�ߖ��ۖ��SRWh'�ֶ�?��	c��IOmmB��l��	5��c�7M\_(��[��������":
0��e�T�|�p��
��v1~� �?��H[$e�Ǿw�)z�h,~5P����{T�� ��� �Jڸ�V��ǌ�.g��-����5�7P,��}�VI;�y
��NK�[[&��+��ͭTbng Q�k�������W���x)�9(}��k�|[G_��94=u�ێ�������و�3��j��U���,�`�l^�}V���? �nju�� ؇����>TX^,]>5��~�� �����5���!5P-SK�PI)SE�x�s+�uj�8pa	Sݸ� �~
���>9�K"�q�C���c"vʲ"h�qB�g5�}�������\�-N�vA���^��=O\�u�ȕM9�7 �Z-�@-&�����M�Q����J�\F	y$Vs~x���Y$�F��2�&*(�Ʊ��M��Wci��Ƣ�]Ŋi�g�1���i����Q��H(��(y[����cI�s�8:Hپ2��(�6%�ȵ�xf��ܓU�͋�eUE�?��]7�D�v�(�J�ڪ�����4}7D`��&�o�˴by����a�*b���h,8[��v�}���3��Ȇ����.>�&v�	��zJm��*�������� ��3�N��_���h�4�Z����(y�B�wdߞ��ⷩ�&�=Ch��"�,*����<M����ĻT�����;,d�D��EdbH�᭫H�Y�Aѭ0��sS)�d\7���5|r�죦
I�2��Z�SDg�,���x�����Y�H�8;8(�#b��N_ajAe�6����2�?W�M�MJp�����^d`����jL%tr��V��o�Ы��Y�PO@L����[G��}�޸���n)�ŵ8ł{	�ݡ�K��R,H����P��}���߽w���d�ʚ�9���y�ٳ�4��o������&�Ͷ��^$J\���`����Y��2E���g�?��3��4Q����w�l�A{F�w�E��>tS5qͧs������?]Z���3�\�d��G��s�d��뷊,���6;�Z¥�d��&|�y�u�{휶��h6j��7���ګ�������>���ս6!���N��-B�8o���/�jT��
��?K�:�Z:�NT�染G
؜�J��)O,O��~����|�3�o]��CsQ��A9�z�cE�^
lv���,"2f5͝����ʺ��,��5ƛ�#�1�V�1Tߺ���џ�.��=�}ރ����+�m���ȭ���k���)t �q:��Oӯ��w�S�i�l��M���H�o5�H7/eo���F� }��ϓ
�4��7�{�C�-�lp�Q�u�̖v��V��e��'o.Ӕs���j�uб
��Mؗm�ۜ9�Ϝ�nq�c.ト�w_c_Ae����u��>3�^=^�{%�w۶?�5���:��g���KPG�a��$���uul�?��I��b���{���$rmu���.������	�B�{�3[�EaN�%������A]�r vTW/ٗ���?���!GXA�v^?�+������������N?�^tC��|��b�U�.�g�U��i��!�q8�|s�Z���}�m����%�����ϡ��Va�'jz�����B;"�F[��3"!{�]�|�L�\�U~�t���h:ur��V�,ۭTt�2���-i��Dܢ܍�=N�gG���Nz.��@[��&?��#<\��U�2_n_�l"���(sT�~h3J�F'�D�!�?����󑷎;4�s�N��* ��<wzW3r��*S�j��"��A�ʪ�:���=�h��H�����a����+Z���v6UM���<��`���"i�D_��7ǰ���ȱ�.����$K��58v�d  6�7K�K�4���?۹,)�YR���S�/�]u�۬���rV��KݼJDH�B�o�Z�A\��J�IoɔC9f9�P!�Q�E���c�% ���x�6��j�+FԿjV���	�EY�O�s�W�~<-�r�Z�͡#��H��D��Qo��A3o�X��e�H�i��)ř��� ����ƙ����es�O.$9e��u�^Tt͆�?�����Ų�:PN��C�M����c)��u��x����������_���6*�4��	1��pt�Ȍ/�$j5[��Mt_:�hEQ㈔�u9خ�M�X���z����:�f�����@�����t!;&���W�����c�T��ޅ�њ�����g�
n��(�I����[�X���,���H���&�å����@��n��%q��'�)
~�+xZ���xz�f���g}��<� �8�..���}z .�y2��}��;q�g|�x�O��if�D��Vj�n���neym�F\�Hɀ�w����\L�j����*��ޔHX�G�����Y��fdt1�Ѐ�H}5o��U�F+��*J��]j��y;L��F�� ��HԪ�(���:�*�}�#��
I~Υ������I2�ʹ�hWu����=�Fy��j��!�&h��jZ��檥G�ݮv�ȉ[ǡ�3J1��TΏW3�çv;�\��s9���	yՖUc��}8�p��_��S{أ,��s�`إq��]}����[�)��:R��):�G��)��s%)D�a��ߙ���,>�͓�����	p��Q�1��{�+
,j�rvG�xM[��v=J���ٲ�M^�y�!G�/e�X��"�Ӊ�c&B�{3���?A���e���������*��)w��y�!k�>�J8���:2��!�����l��$e������ڥ`l�w�Ɛ�,��ʖ�%ZVv���ѐ�*#�#�Y�����$ ���֛���jx���ZBw8�n�	�_?�^u�?V�U���1o���	 �)f��9)\���V������v8��́F3������#9�5y�-x\@������:�47%���t�����5a����a�1g{�3�2Ί��Wm���5y��"��u����u�%)Z�!Z#
Z�2�B{3����/y,̵��s�[�x�=���;CHE��@Rµ�{ޝn�D�\g��7>i�Zl�ŏ\	.�\{b�Ҟ�G��6�.k`Ι�l�yr^:o I�����\p�����S�7�o�
�`���q6�?Wn<�;b:���]� ��Z�1�H��)h
���x�ϐ��c���f#�읣�7� ^�v�qz��ݻI �(l��<9dv(�{s!�Lܛ���E���
ɾ��⎅�|V&�l�E>'�[Ud���X0%�e�+���jl�.{���a���� �F3��l��rq��yw��2�x'/58�W45,�w4�SM�a���9�)��Z����q�m��~�����	_P ��Rn���T�]����/0e���U���v�vζ/�K��������>���kうW���tx��͈�a5�i�֒���D$�x��7
|Jt���!�2o.&ʌ���)*7�`��|�bA���z�>�����U7	2M�&��.2�ψ;��u��d�I�zQ�O�WLz�� yV�����x� f�Α~�u-��N��X��#F��bU}N�d��Z�\Bg��Q,�c��&.� N��]����O#�#��P[O�
��d�t�1�[+5"��� �<�'�&��rdw���<�J��QS�tl�_K�X�t��@�������,�O��|m�M����-e��w��x�{�c_����#�#����bj�;���FIK2O�;E/�'/F����`t��Ӱ*D��xV�Hb?`p�0�l�V����%��/F����x#�`c-k�O��a�y����ɦ�����]�}���[RU�\�zF�|y�/��Z�q�1�z���}r���H��%FE
�YB-U�w��b3]� �������+�Gy�?s�9Y�u2|_�2/+���e��5�Γ���1>SF�Y ��0 {+���k%}K��x����T�������2��KX��ŜN!퟾�O�l:y"��j�:9��0/�	����:����̚`����B����N��L�(�?
~�6Pw��䰫��\aǉ��zG�gy����N�s�~�D�������X���^����f�X��])��x�����/�|����ɽ��a����6oq�Lfk�$��|Z��<�dr������Bl�ʠf9E���SѤ%&bN@��~~dz����"���!Q�LP��P�O�.��ɣ���mQ�@��exu�Z�$HI���Y��o� ��Rz��%dnm�E� '��pS+��@�z@���������`��nPP/,���@����������>z)�5�\�|Wv�8��/V��`\z3�����°Ћ,��CgدEC�%�i{�t�>Δ���hٙ0��x��>�_?����7"�T��9r�<����W���^�ͫn�����Z�I��Y�von�n1�9Hh_��n�R��ES�*����<>M��m�Zƻ3R�"j��j�j�=O]?�cteT#>�U����:�s����b��,��N�g���<��d?[5�{S����BC�瑱l�+Ba�_�>���ޜs����O�"&ư\]�ߓ�DM|���K'!�D"�H�2*gғ+��n��%����"ݚLp�
m���C���ȕb����q3��'[`���ؽ� ����}企���o7�������-��~|�C���^�K�M�WO_xżW���M�! ���$���䵻{H���|rof�>o?e �������g
7�k-��t�Ϗ�N�g}7�߭���\���w��`EV&����m��G�
��]R��]��Z��Q˚Ḕ�t���)>��MP	����<��t��� -8�8��5>�B m��w+-�;^|h�gOE�`�m�Me7��;?����lA��Dm�m�l#3'�&���H�=�u���P��ݵ�ᐫ�`����a�1�>b4+��^��W	O���zӚڵe�+�p("}��0&�8T�$��x�d2
���'�4�]���S�r,�1��FB�K��G���K��_H8@	�)���YQTu���q��c�Ѯi����F�b� $s�����7)�*�k�a�5*ֺ��(4�=4��3Z�pC�2N��<������X
��\��*�HJ2�Y�S,�t'�K�@5������V���tsWY�A\���S�%����I�DU�1݂�p���d<�H� �u����Л�ET{\�]����ѹO�rT���=])I�[؉�~���95�os�r������m��l}�Nf��oC�T��*;�LƱq9/���0m|dD� ԏͲ���U�g�����Ń������E���&�]_���Z�N���fh8�d��>��>��/�}<.��7�����#�~U?%���]�'�<�ЭlRv���H�l�&Dʾ��E��e�v8�Z��!u�6�L����z�B�Z������W{����=J{c�����u��n�<�x�^���pP�W%/�L���� ���Ѡ��a���A��x^x���4_w(�F��,�&tutD���ؤÞ�p�[8�
#z%ϱ��i�g��r��I��܇�T�^�
dP�����K�P���X����Q����!�F�lònI�S�Q�DƀS�1�}׵	ie7��̯�#l��s,L��0"�_�k�r���D>�������ܯ1��.�k%����Z��]D�-:~�t�t�z����ޜ6{�?-TU�����0^E���۵�n��|��2t{&b31���B�t
������ ۙ0{�y�*3t֡h�Y��7̓�'��z�\�����L"�;��&��h���]�8aK_�f���%F	s�x/z�;L�-s�:6X�Yy�n.�Ξ��[�	糢��B>P�a�V�^{�T�-���|Vn�Pz��­P�a�Dd�H����2k�̼j��M�1�����X>g�z�pI8Y�u�A�K�#�q.�����%�BLś�<�E�Jب�l�����r�As���#�JL�g��h��m;CQE+[x�-Du(��. ��͋�����\ZEL�!h���E�H�����9��?��_��ڢڙ�k�[]؆������=�_�_v��8�����s�BE3(�T��F#��j}����,�w�Z�Oo6H�*��q�/ �cx]D��b
�"
��� (�݅�ner	���~\���f���ʎW~�1�\������=~���۽���?a޵OO�㝁Ż�W�y�O���A�����Z��K.���M���}�iaE�u�O��%Z���Y֧�&uȏK}N��I"j��7%�3v�e6���.~�#��6��"e4��a�fXtk��3�
�.�(A��+���.�X6U8n��K�P��RU���l=����@�:��	Zk�1A�ׯ�M;�X��Лi߭ܯKh*좄g(�822Df�p�=kA%�_ۜ(V�=���#'�_�"Q?'Z������MpZ�3�0�f�yަ3���V��Q�q�DW�1ʽ��"�řb���w�1�T'���QL�d��G��1-�^ZA�ڒAYܬ�^*h���0��Z�"q+R��QT���eq��B�Qu�1,]����=U�o�?vŋԤYLR��W��y7\��.i��n���GI}����o|OtF�da�8�lE�I�А���K:��sbL���z����[��']yc3�Mִ-���\�M�>dkl��qo�������W}�᳽����Z��=��`�,j3Q�J�U�79�����r�	I&L�\���F��m����e4Ǭ�"�4�d�|��S;�⽘SF(��}��>��B��E��ڻ��4����\�v���L��{�n�]�f�� �{U_6_��b�ˀV���H�ڗ2f}6MT6����vbB[,KڹB>���v�]]����޲����q�[4������$MD����+0��Q�[6�MG�wE�k�M�I��}���ȗ����Cu 2�e��Y��	͚�uT�>�o�2Sd�26��B�C!n����#`T�+�g[�,�|iHM�^�%�$qBzy����(\�\L;��C����f텤�u�uŉ6��gc�/Azf���&)j�O
����Q�z�=�J+���$�3��#�1�/S������kB·��B�^�'�.V��U��Z�l�~�֩J2��x�j�R&�VB9���}K��U�1dw�z��cY,@��񴇐��Xu�..`��������_ǝ�Q�� ��������~4h9�]͔K�k�=^.h�5ݵ}�M�V�r�ZV�"�����$z��\V��|1�#�w��#+�X�����e�� �<�z��}�3Am%������]��r�w<)�Lɸ�_^�vH;/�o��Z����ñ/�w�nQo.�֊-	���8��]�+wN���������O��	�Y��g�� �J�@�0!ŬFX�$�̘t�v�sF�)��t'N�-�ڧ�Ǯ����1�z���G߱��	�-�r=%\ ��o����nlI��|<��YM?ҧ��ҹE�$�L�S���7�����s�� 5j޾�c`��R�mF���6K�w��D�=���`�߼�sE�{��Ӭ�t����ܘ�>I�f ��(YcE&�E�L�vCC|�2�[9I���.�����2��> *�|#���D�t���ǚ����l���
�ۦ��a�zW�+��3��A4[�Ɏ�qE�w�*pC�{�t*%����.����#-���=as��6RoM�n���᭕Xh�o(V%ru�b/�w����(�"kV��1�	��8��)іG��v���X/!k���J����e�ʘe�Ӑ+���⩾��t��h�ke����bd|�ӭ�� U	V��ԓ�r@C�[*�.n��԰Κ"��$ ��������wuy��\zx���j�*��y�o���Ȝ��c��Գ�{��Ds|�'P8�c؇�Z`��t@��6U�Eƌ��S�Ts�E̜�=�m�颺o�����@l�67�
�HI Ƀ�Z���$a�^ �WNj�%�V����:�+�mh&�H�P��(��dHC1�(��3&T�^,��O�Wxl�e�Kk��QD����V���g��Rg
�^���\ZAa�`e�뼼�������E�ʹ���px'	2���+8�zh��Jx��$�:@�4����g�L�N>��?���M����և��}�l���a҂l�gNv�-3�|��®�'�!����Xg��$N��w�̕q�w@-��h�N��jd����������E?	j��b"�El�ն�2��	P�Ǟ�bW}�#� ��� d��I�r&Ry+�y�c�Kj�<���as��O)H�EV����0�)��r$�y������ޭ��D��*�⫒��R�H�pm>D�'� �����d�C*1zi5���7~�T_�!�-�sS��\(���v�X�B~�C�\-Կp��k}�~^���X���/�8l(�3�� �6�EmeY�#`� V�x�=�X�M"�ȟO7�M��'�5��g���ke��W#�qI[�V�]���0 �[�7d�-�I��B?�i�<��!Z�ߩ�2 i��z��h�Y����yf|��|���R�B�N��ؿ�U��*0ݕB�m�>�^�,lʸ�
}�Җ�V���$�G%~g.�ۛg;Z�ځ4f���.�%sHa@�.�T|&���iBKaS���H�H�UJ���D�rxȔ�AJbcG71�_j�C1(�6HWE�$+����5ِ!�6�v����R��7��~q��qD�ъ�L�����$B�{ӾQT�Eؿ0�sV���fZ�P�=��\��K
�.r�w��i�f9?:�fI��1�O8f�P2 /����h��L9���=w���W(�3C�-t�+�'�_�vCFQ�o�;�\�Q�Ox>�"�sc~�� 4�}�ڸ4b�;^-�k����oX���4����v�a��+:(��W�����s/�v�gVW�v�c��w,���]?��T��� ���V pc�kts�dB�S�����!�GAj��VЍ��K���֤��V�)�f��@�8��x�/�Ҙ��M�܌�i@��@�C/��5�S��n�!��e/4�_�:>��B^#K��ÿ�g �@5ʄ#"�z�t���:+�@�y�s��-��:��A1�Pm�d�<�(�/�Ճ�YeH¼��� v_�#�*g���8�R+TM�_O8������&���Lʂ���YNf����_�����4�~�!F֘�̄:������W�x��%�G���!2ǁ��7#��鼏Zie�.}����N�Ym�
{r���]6�(?�/��VW��·*�]������x�2RO�p(�v1���9ΡF��9�F��w��-U�wr{�����f�;?�v�8��e�`�_�$�>1�P�C���x%0Cv�c����i"�~�Cb���{흘��H����'P���-o�k �顎Y���h�ƈ뉞ǭ��YF�(Fr���L�(���O3���<#�`c�ˢ�N�? ���'Jo��rŨȚ�0
�����b�r�m�m��\iF������ez�na~��]�ۼ��;�jX�pU�X�J-�$i1RF��Y8P,"�h}���0�~ ����]�}�EVX��ס�\J����W��~ �|��CQ�{Ax[7���7U֮.�-�=��輷�{�&,��hR�~c+��A�n��ր�!��POv���HmIA��ï�ʠ����I���`��2�Bk�Z���5g���1�4V��8���MY��T�N`Xk%�Mv�t�}t�+}Y��7�Q d!U.�d /���h��x-�lQW\�X$�]��_��pn�!�UB�?��n��g���+g��f�;�@��D�"���"��8
���o�6�E��RڰH�IT �A9�l�1������k ��>���J��Ơ��'c�7��.�*��b��x��6|4�����m���+0�Li�rM�Dg�I�|��|Aq�ͼW>]�5�� ֧>>e��c���^ˁ4E)��C���b�M�S�M����G��!Oq�
H�������(��<{��N"YWA��|���>�yY��Ж��I�]�tc�kj����G�)t�XAY����1�p�YF�y��
�G�����(��I�#~|T���e6p�{��S �w�j�I��r[�M��G����޺�Wh�ގ�0�O}����zF
�� ≚�#tBXDO��:�u8�R��&��Q-�W�O�wZ���o����M��Q9qJ'KW� �w�-��EGl������$�޵�K�C��˔��ݵ���u��	q��o�#��~��KΉX�%�$I��:M��>��K�w���K02̕��%;4]�)��h�l�s\�P���Ȓ�Vցܑ'�3gt+D�H�8�f�1�pP�f�%<0.��zU|������s��ۏ0ơl,3/k�4��+!|O�J0 ��ح%j�6�Mj,S�B]ZR]W'�"��n����4w�/O�i�r˕�p�=�7��s]yҟ2)+�񛘞zgƗ�ΧT�R�P����-_���+2aBR��l��2�9���7m��������Be���݋��o����=6���l��/�ٻ�9��/+�۾\��ͪUF�68;�e]h7DJ1��<�un�=��Em<&"a�
py��ȘR��9�Iʂ&�Ś�����W�cٯ]I��[>L|�j��U�k�)��A?�z�]q��L�YTA��`���ţJs0I�⩴�~��ԁ<�1���m�!��#Ş�9I$�ln��]06�X�$��e��6�I�6>г��|�x�p~7�?����:`T��[j���h�޻��܂@F��J��G=��w��ƅ�{	���m!��tn�>W+���!�W�V����n/j,���&�{!!�wC��yW�-�\�a!{;���su� 
�,�E���O���m��B��-=�!	Ƈ��<�����g�P��]Z7�f0|�I����Pf������{��Umw��}�Ì'���u���
�E��r__����}?�zN�u��K1}b{�MP��4�k��ߦ�<���HH9Nᖽt&y<�ө�$��� ����5^�5��v)��f�����z�Q����*��W<K*�.>-N���P�n�M"���o��*��2�n��i-ֻ�#<\ȧn=���B%����^�3�r���v����	�8�K)Z�a����#�(�VH��B�\��ZR=���:��R�w�?��s�ODa�ԃ��-��&���סrY�u���T.`��7���fbآb9�����#pn�DS?��|�C�\�`��|��8��XmU�c������T��Q�,�t��J������f�k�fS@%fBbS�����JM�͢'Ӧ '��ǎ��GC�!vx|��Hk�4�R+ZB��᫹jR�U5?�nk	{2F��YF,��������<���0Fv���b�½��r�?YmP�W����2�M��c^�L9
���`��~C"�>Jmx�2f,[]&���.iq��YJ�_[���n��C���T/5gB��C D�I�����+%������ T��E���I,���qLe���\�31� @�[q�#U>�{�,�ԏe�y����<gȬ�8�#�m������^z���S;G�&����r+ͽ��5�����65�O�)��ZPH��3���	������2����.{{ �A�s�n��R��r������Ն2�A��G�9�l��R�nL�!+'9�{q�MĥD�H���1���fqzQ	v{�W����(΂�X��N��_E����V����/��ܫ9�L�fp�#�?GW��y���UF�lN�>�ٻ������:p��]6�cz��s�S��Af`hN�i������l#6��|eS�Mt�F�����=��$�����'��bq��o/���Q�P����K�>�T����.1ן-׬�c��s�)a���c)�u�[?X��8$�V1!趐��'��e"��?��-�$���v{zZ���� j�|s�h���SA�r�����j,$|�������Z�9�����Y�����mF����0�b���!�)��P���8���ļ���͞��7(��uz���DgDΟ��� kߖ�jփ� ��F�3�����ξdɄ�١�����_{��)�`�/ߴ+��n}�5��.Y�>e9cX�S�d�-��c�T;	�1g _O��+�X�Ŭ�X�A�V���$@�=bu�ćt���c��)�$����as��NN��}�U`?g��a�x����&r�~"Uőe�m`6C1�$.�$�5V�Y�01�֪G'��5��Ew�KM�	g�(U�o��$��q��t��G�K7NÉw�� �"'g-E(���	��+����.�T�!�A�I���������V����IxX@Ns=f��$h�P5v�*�@����?�W�nI3�������jrh߁�	�.%_��A����Do�������0�!�ş �>��L^����� r��0*�c��إHA�wDd碋�]�ߤ"�%�C}���Fx�#2�7r �#��E�M�B�P�*��5*�1�<2B2��c	Aet�&"�v����kW�R��Κ2}$`1+���s��;��s�ڐ nBKJK��w�XR�ᶁ��U���*�>��GeI}3���?�랿��P�.ːȊ!��M�� _/�)$�lN4c����V�,
^���!=
^BQ�ȹ�5�CW��������K<�G���i�~�GOl�@ID:���Nə�-9�����A2��Ƒ����S��I�Q�E�M%��gN�F>������xO{@G���P��à��P2�ˤ�����@M�~�`2��1�Xi&�>>��ਕ'#���EG�a�6E��N�-4G��/5G������Φf�����*,G0db����˫�I{� 踔�y��n)P��ϫ�q��~���=I��1������]\J�\���OW�i�)�|�����w��<,|�K���d�Mz9�Dív����w��<y
u-h�TFP�Zfa?]L�3}�uD	��<�/���YQy��ͳ��X�)�[�"�g�(�bM}u^�����rn<��y[s6`ۄ@PO��1YIu�W���_ x?Kp�&a�$��~��:�vܑ5?���V���T��#s��.�j�%�.5����{��h2�?=b1p�:�'��\o.[op�ޟ[U"Ž.�	?��@�j����-߮�e���C�Vm�J��vp���a�����?��V�k9�V������v6_�Z���9�t�Yw��m�wn饜����E�k�
��1曼�1��8��=�z�>� &�\G/�	��Wڨ�aV7ӞL~Ua^tm�����[�8.��բ;U�{AT�RZ1Ǟ��J�����ܢ�꺺�_�*�ĳn���)^G�R3�I�"f��dH�v��nx�r�������L�P�!���+Ѷt�#"���V���+�L]�N�Q�H3��^.G�/����D��B�D���ì]
]��0$�F�f�Y��o��G���������'-��k���:s�[���c��S��-F-�?�v���Rܳz�5���Ƭj��]�H� K�q��")��l�]lo�0Ƕ[����d�S+�����k� ue��b�&x�(q�`�	��v���hk��lFۗ�B��u2ׂ4��ө��t�z���������g'��xj,|݁�M��^���X�K���"�02���bJ�T9A�lA������nM24���O/�M��^�j���ϯ��s��X)T��/�����Wߒ��[��yb�������i��>¼ѵs���T��N��ȉL(��o��X#��e��VV����E<T���t���z��AI��]:���ed���3�nW�%��{� ���Z�Z%����g� 
ºԯ%�CuSݠy���|՗��m	��K�9�}9ό:o�6�/X�:->���]�;>+3�(l����f(<�+�2 -����^|����V�z曚>-B��+!9"�0OUaR��DꞄ�e���#xH$�e���8a�N�p��(�9���xϽŘ�T�i�$��1i,R\��ܕo;�&�]��������Č�}��/��a$w׫;���!�o+�K��⼪T�,��ƉlX^#h;C	G��1��*�#�z���$����n�-����g�Gi,�F��R�fbɪ<�>��s��ӥ���5�ec[m��x򖥉��hɟ�'�o"}���C��qH:�ϻ\؝\��u�e�u�l˿�Ŭ	��bfى��_6(c9���ϟ���4^#��v��:����CV�/���i�_�Jfѷ�Z+��[�\��W=k����-9���La�@��i�R��lU"�t��0��o�եo�\�┩�<�p�� ˺����4�uޗ4ߞ}����W#j�z�;��#��0�W�eR�����|�6������	ɪ��:1YTO3����V�6oC�*ޝC|�h�&F����b-���In'_�n�J߷��#B����Q�</�ϸ�Bk��.��֥r��F.��%��&f�H�`t��b8��WE�G��I�JA��7����6,��Zj_��T����$�Uu幔@���g ��c�hCF�S��θ��:���Pv�>��X��dS�? �5�@`s��E�R�ǙsL	�EG��REb�y��p�qw#TiM�̎�,�!�+.)�2-cu�;����"�T0�v�Y�"2�J+���a����?�����6Y?;�J3��N=�����V�dg�K�}�P�_��4�:v.�o,�Dxѥy@�;���$�k�×���������QJ��%���ҁ?wc���(�k!��-#�z.�a��	&e��G�}ٽ���W�3��;o���.%�K���tJH�|!,��dS����{�JQ�P%�C%r�!3�v�4q��.!9�97��B
nF<���}o����k-�I���3$������R`�z��T����l�S HRh��饗��ܔ�2{��Yo��Eh�5�N|3�r^����Y���SB��G�<p)�w�����J�?#����:�t���P����FU�9cR��T{�xcN�)��
&wQ��%*�z���R=��W��ލ҉?�U�C�@*H+r���aż)��=P���T��C�!Lu�#�w�n�7�?��^P��ݮ�\pT��z��K������j�ǐ��
f�S	�:�g�w�ʨ躋�˴(Ȇ|>o���$�s`]��1���cK�+"�i�)�������P��P��ڨ�㥷1���Z�ǭN5�gŀ���h�M&{?9[���ď���A��3�:�y�}�W<��+��l�7�p��k�/lZ�b���O9֑����aRv�\���k��yR�su�p��kj�Un��d!&D4���#��
V�T�$������g�����ϓ+�s�<H���O8A�k��d���7��]Z?�\T��i{B��������v���>��E*��`�s	����Ն=��hL���8%zfI6���-Q=[w���v��&�A�*���
���� v�Mꄥ]�t��{�fF/���pm��ۤج�w����0AG|��d��y�)K���t/��*|�Z}<��
��v۟�/�r�e=�j��#��W�b��^͢lk�h��^~M������üd_�{��E�)�C!G��Ʀ����@�O!{}��|����!w2�F�OP����v�M�8�W<��鐳w�"�抈^���/Yn�[n��j,���vL�l&nz/Wk�1�Y��z����yǕN����/��}�绉�P���`�������4[��{��3SW�b�v�Ʒ�X�䩘d��7����_�@��~��i�?�ng3��fAaQ�9	I� ,���묬����C\7ݮT��1�h!u4�^�<Wۈ�\�7���Z�b(T�q>�"7k��up�B�	xbꝖX�&�(i�VȬ�NcX�1����+�k̶_��t~��;ڕ��l��K�ܱu6/�L��\*��eRU�.�\��~F��`���<.�S���	�t�@(&�d�7���X�<B.����U#7(���4u�+�?~��V�b��k�Ia�W�UwY����v:v��Ǡ���Z�	{���`R���LY�3j�:�|�8�' ����✮��CIZ� +Kw"��̒���jonr�kW������6c�Y1+{{�
�-��_]h���خ\./¾n��%T)ü��4Xx-n�h	g+�ƽr"��4DJ�R�o�(�혲7�xJ��ϔk�G���������{
nx��U��#a���(�V�q�H5qR 'ΓS�co�B�Ц����|q�3l7�7�=;]�xs$z�b�Pj��a�
�#�đ?X�X�z�pe��N͖��	m�$q�vQ�%B�����:]�2g���d���B�
T:�´�ֺ��N�ƾb�q������c��u��f����.0�f��nRQ�����Xa�(V>L��6i1T,=�e<���#�uU#m�z�+�K��o�Ce,�-~�O����i�Kymݙ�C��xV�"!�d��o�_�q��Ż��f�Z�2���hvڐ!j�l1b_&/��z���9Gۣ�r]�F�;)&���~\��\I��<��h���&´��"��VaguJ�������t�z(?D�~��݈RϽ��F��E�m�z�آ}Q1�u���D� 3J*hW���n�ŵK`�,7)S�J cD�B(����p��
2�w-������*���2����m�T&	דKr�$� ����R�����2��ۭō5g���-7k��I��HP0 ���7�ge��Zt#��߫��*ȩ�O���w���j�5d���[��!����"�6�R���N�{r��̲>�_)N`�Gu�ć�I�Ћ?c��ߋVϡ�zW��͞�&�W~���j��j+�c.FgN��?NΚXo�n��!�ጳ���F��o��Sz2���\^7f�xH:h��f������Q ��o���Z�������0+����$J�ᇱV�
[��w�֥���
��E�W9}�T�uB~�棃$]z[��j[�hv�S[=�x�����D�L_�',���J�v�y!\p�_`�?$��$H�OW�@	3쉼��|�kLg;�ڕBK�Lt�ԓ���[��rR�Wk����ޕ(Gu�gb F
^�r�Q6��nFJ����5s��-~��x�Ț��Hl\��1b]E�L2 W=V���ɶ|�;�?��3�Ͱa�v)1J��h��=c+JQbƬ�I�7��*EP;ČU[���{S�)}������|ɇ�J��8��9�3�W8�'�.�'�����Yۂ%�.�=r=���YG0����9�?��t��c������d�[kѲMb�T���VZ�N��{�-[;�iK�Ѕ���'�A"��yp��'	�����Y�jdƝ�p1�x���gƄU%;���{L�H�K:��x8f���ỷ">uP���\3��@Q�`��6��򢩰T�r�8���'����Z�	�O�"�]kþH�y����yW�u��>��<Yڤ��;����I��u8���a9J��rY�w�-�����X�P��Y8��ֱ.?a�<��F@|��sP�b�Ԉ��-A��=�L`���I��:��f^�&s�C|�'|���f���]����1��`����E܁<���.e8��=��uӯ����m$��_��\�oz�n�3���2���H��}jA�#�0�z�x�v4(���q�ͥ��ٖ��j���^��R��<H��M���j��ض�X%�Mux&o�ڸL���jgPW�c��ԩʕ��pBIfI� ��;"�ޓ�l�nǃ������F�^���?��}�z�S���:���Ǎ�! ML�]B-c�J�<�j3�;�.�?�xʕ
!�[R��=�����Hs*�%-�0���}������V�z��ԧ$������a1C��9��F���g����i�̀�I��\h���}�����|�q�ס����e�%� 3`�X��v���ؖ�z������(���5�8�R�>��?�9�x<�f�\e{o��j�R[٫��� ��O�~�_*�ud�a�)\	J&�.u�oך��h�9�*�Tt8�?���{מ�/�5%a��zђ��(Fc�|��k%~\���uY{�fqIr֟o�����s�_ߗ��d�=JY��x/��f��~��|�F-�l�U�~�D�U#��C���϶o9L4�a�o�ա�Zf�9Ԅ�2'�Gb��1Q�MY{Յ�;�dѴ������Bf/�cR�0z���Vדv�0yۯU��sY�z	�ߛ�0��r��ƨم�C")Y�G�D�rS)�>�������}C""s���ȼ�Dz����Co��p�� �#�c�K�ʏ��y�/�p.,�L$�nVh��)N�:�	Vj2���q0'p���s'��AÈ)������,�&�)��%'
��n։/hؘ)�	����4,n+F溡�T�3:ӬQe�Ĺ0G��E�-�x��>���F_	'�0۷a� 1�!�"AX<d���We\�r?�^[��h���-���ӏp
:N�@*¶�a�l��S+�pۯ̪�d��8��[-��Fۨ!�;�5��Ci�&Ã��^|"��Ds�P���kR��'�q;���������?��x��q���s��ӄ����1�	�?c>�ЍJ��w���G���j���D�E%?_�hG;���y�t`��E|�İ?6�L��u�[a�dmma-�CH��F��v������5q�����8��J��|�.���D����w�ؿ���䈃�u_�q��Ś���7������wJ�P��;���CT��2�VL"h��������M�W�2���7�%��xG?�N6��Ҝ���T2�#�~W�4�z����	x?�Wۀ/ġYP�T�g��كL敔��+>M4����¡=������P��(�7FZ�TZ������@���NX?�`>�چ�Qڵ��)�����6͢4�H/��]	��H��3�d�A����#/[�ܞ���w�6)�i�����e�m�mB��Yh)��'\�/����@鳤�AD��1x_��7�K�m��lH���bK�1�.v;iy3����md�mT��?��B���������c�L�{P)��@����{�������̧�t��\������~��Ϙe{�}�6�"ޖ��9/|�$�-��qIl��vWuQ�;o��D}T[@�MPn���:�!���}Z'�����O�Gއ5�X<��,ʟ���m�<���)ƤG��MX[�l`]�Pl���m�]���&�1��`��Yc��h�+�1�S���e�}�ψ�'O__�<Ņ2����KW�3	���H���|�l�vEYl�%����������w���sJ=����ը��a����8Հ���Z+�?�V�5?�0����uE0�U�W��ޒc��ڟ?��&	�q�B�k�N�-�31��d�N���e
#���AT4N��b�?4��X1�z�~�������a����_"a�"���[UQ�`��|�WH<y�����bI���`�m푪D�ac$�v^ݸ'd!n�:����j��=C�C�)���}E�����,������Y/��3u��ht���_�s��~ ���[�L�k�<s�Mc�LO��Ok��}!txX{�psfm��C'�w�=D[_�;�ҡ��sUr�?��͖��{&^Z#z����=Br�-��GN��9�����h��"e�����Τ�b�]��UQ�2���נ�i�$��4}H���ȷ����uv� ��ϒN�ٶ��'�#���˿*-k~Y��Kg����=����	�t��$`����p/�&'ժNc]�bfR ��M\�z]A0DVBځ��S0��[X��d'�x [���oЦ�;�@ }��|����)�o&�l!~Fk
i� ��]I��Џ�E��Y�Ԛ���q�iN��e� E�[�����,��1�:*F����`<zJ�d��OY�/_���UE:�����d�-��Jz����{����$��H#��-b`P��/V���'��i�wOT�����a�k�<n}���#z!W0c�O���T�R��mʇ'H�(m��ͣ_s4�r?�ȾhsV{݇�B
���"h˗w��竩Q	�#��ǆ��L�|��>�=�!x��hǽ���P{}���#Cȼoa�=��Ӆqe��j�3�0�C/��ˏ���ڊ�QY�|>j�O�<��Hf׹��Sv�O`N����l[��HS��F|�(j�*�GT���p�=}z!�t55���k��K�
|��0� ��Z�;��1�co�eӶ��t���I�y��}M;ǽ��S��	8�jq��S��}n��YÆ��a���o�?�PL�ZnvK��4�$�ڀ7*������^��t�O���r�F�����|_��2U 9�
��A����m?������}դ4g���a�7N�AIe1�_^���Q�+��-��_a*�U0Ъ�eRkܯo������
i�m��OS�#�H�͡�k�v�X<m+��������',�a4��qqg:)�/�g�p���Y���%�ﻧ!�2#;��x�#�]����ŝ3ny����~x���4�7�c+I�ҥ�Я"F��
�n��}u0���zH�GT&d�\�[o������i�d��]ټ���G5�#��Ә�*��,�2�ozz�%���?������H�735S2�0���~v�?w��2|'�T�����ʀ���N�����"��?0|���������VI���L��۰����X0�޶�����o����N��ba
ϵ����������@t;�rsO������q��	i�|L��[�{�>$�ѽsjV&���V@�
��ޥR̈́|�����![X㳭�ͫ��vC��ۜiB�K%�,��|�/�\����+�>uWR8U̳�y�`�O���w��S��V�z��#�B�{�_�FR��N�p���O�����rԀ������QO�c���;�7᫭A�e��ՐS�ù5���8�r��ɲP���i莀̖��q܆T%�^�>�p!	v����|X�Cbxl��ܼ@�N5v��*Wf���_�c[� hvD�M~~	ݦU-�^�1Ř�c�+A�����Զ��ٚTr,{|)�7ɲlp{�u�r�w�x�{�H��Zs Uz(x�RE�*��Xj}	��H�x�Wy��Hwp���Jט�{����69��6��`�}�}1��x9�r��w���E�LM�ۀ�T�=RмYpR&��!`��!c����i�D�fl龜�Ch���7{ ������L�*�C�\��D�0X!�4��qW���a��@��w��;f/u!�*%/�=2�Nc��Bh-0�f��?�<y����w2����5��߅}��`����'���8&��N�z!��{�B�^c5b�x�J�A�P91J�q���)�K�G�Y{\�̖����!1�z���f?�ͪV4}F��_��<��"�R�"���u��Y��Ea:��JB=3����w<��.ÁY��4f���n���i��O�q=sZd�	���ՃȌA_�.�'���7���-��^�TE!�Yۢ1tH�3h=�.��� ���<��|������(��
�?�~�ȕ�3��(�>:M3���;Q�b7�a�G�=��/�-nֈyl"Z7M�	�3�W@W�q��pA�c����+�~���
Z��s�|�[���E�D��L���[���+Q�������?�V�XjF�b/���m��>0�`%�g�o��U$Ke�}tN6n\�k&�Da��,�T)�VJ0��3�k��q�0����l���vI��o�].�<s��m>5�a��K6��sxfcK�Q0���/�B��-�M�F��R���F�UR��}�����}%<c����1⃎$~�BY4T[�s����Z�;�/��u���0`;I&Y��	e��/H��wo�WUo��?�#�'O���]B���_-C�Z��~?#�k���G�^�1N�.r����Wڜ��}����Y�u
�O��c�z�|���;<��;������m�#�.��D��dP~��|�o��W*Ϧw�i
��ꯌ�<��lt���3��&%��2���[��%�5���S/�Qɘ_�9*����s�.)Wb-�s.|��R�OL�$��K���P9C�he�j��������u��k��jv0L0�k�rv�ò*m��o�͂u�R���.��w�O��v:۬V����$��UqY�ߐ�>�<ڤ��8��(��7�$��J�
��/��1&)d����㳞h�7S�;��ے%k`����bR�V�J�^ɂ¥�L�÷k�7�&Nb>J�w"��MX5�������Ag��i>x��D�@f2�|$7���`]��z��n���~+�8�۷��I#[ p'�X��x�#2ۇ�]Off�׃���2y)�	�g֒��b�j�D�)�e\��7�g�W�v��:�q��)8@�U��A���o����]C��?��q7k9k{�o�����fE��%.��E"����vV]�ҳ�?�&U�z ii��4��-N�.�g9�#��ŷ��zWB9�f���)���ЕF��O���|��ȫ%П1r���N!��� JS&�y�hoݚ� (�]�z�L�]��@y\�p�yAtC"Z]pA%( I�7P�`D!
臱ש;ܭ{��p4�t4��������qdd�����K��6_���{Wk�?�(��Zd�tV����R���M�����;[����y��Sܙ�]�?/�,����Mc�o��mk.������&]��XD[�p �7�T:4n˫|WX	]"'L?�]�.C2 �{J�С�hS�R=4-8�7x?�>��d ��LÝ�����K!ծN�q�{��pI�����˘n��;݅��sIS35^)ܺ箔�����>_�}��l�N�D1��X��-��4��HE����p���8��0
��փd�ecG�"���Ւ����R��#���*q�*���j��b0;%-=��w���j����
���^�ǘ�;"�4�(�iC+mY5�葤�hesp{\l��p&���ă�Ni�">x��C�V{~m8vS*wo��H�w-ul�k�l�D�=r�p�����k�qXڥ]x�D[tm��[Z����[�<Њ3���&�!JH��#ڜ�D�sĦ��,+����J�`�&��B����`�4 �>�&�DM�^�jn����طg6����R�[�s�`@k[_x������9�|HyG�,&8�F�4������I��O� NL!���iÉ��m�� IQ�lcK2^�s�e�F�j��	�|�6klٮ�1HZ�D�M�D��xd��6�8�����{�PТ�<�)	?���+�;Q�
���i<?��o�RrK:�&]��������9�C��҄�7ӁQ�-EGH4$�(�+q��m��a�� ���*N���̭���tٍ����8�k���&�N�}�-��ԡ�XGXa곱��+�q��C��#pz����O�ٔ
ko�\.���ܕ�gQ]�A�$�a+�ycCsk���![sO
�ɧ��۽�\<K�<�t���q���x�����3�_}�À�D�qT��E�2p�g����e\�
*���Wv�:�n�_���%�#�	��f��*ը^���z�����>pr�Ĥ��fU��¯�|�HS���1���m4��0~�M�W(��Q������1�_�g�Z<�o$�x�y�I����?��-���.>�b�!gh3���#^��*��{b�ӫ8`0'@� ��l>k���(˄�`P!�����&"���S��EҾ����'��5`�Գ}x��vON9���o�L���}�z�U�1�N�r�b�Y�����;Q�ם�[��:�<����,����:����G�$��b"�PDĸ@5��ys" ���^�b�%q/y"��dQm�c��fAn�aR�hv#�7�Z叏���'����"������������Ɓ��{�7"#��0�dG1�%*햏�eF���)#�Yǳ_~>�@�l��#�Z;Ոߣ�P��<TG�A�Ջ=��Apx3ت��0`&o���@
�@xm�B��=��Q!���B�w-�6H�����B(�`$���Mˬ�G�J���I�Al���y�o��%wm~Yu��E^�;�ă�̝�ԃ���:�s�}M	�ˣ�v���@xC���2��:(�פi>3s���r��D��DRZ�q�Ed������e{������M'��*ѫv���R�ZE�%��������f1�E��)�ȡa�T�!l2!-X8������$��� a����_:�r(y�Y��pF� >E���x��Ω�#tm�+;ͤ���2�`ٽ�Q+]UG�-D�G�^�2 8�.m���ZL���\,T+�T�6F!M�Bq���n�M�RC��� �9�mկ�6U�H��.Tг��V2/�)@�_eQ�x����uӥ�U�_��$�M$o`�i�,�?կT���9+d��eoY�����F��F�̺�G$+>����@.�	��z�t��G���$$����?�X��~�Bǌ�W��k�)2�ZI�ʵ{oUzV>AϯF��L�9D#_�#R�&�H�����n���������D��2�7�(�����*3Z��!  '���+b)����m��8CSF$�3�M��� [�>t�4�~���%a�brZ�������,�r�Nbp������e ~9p3��Q�uV�"������6�7!"�J�����.�|�3�2��S�����#W�쭓��9��a�e�F�?Qoq�Y���u�K�� ��?8����:���y�iϯv#h�K'a��@��m�6�u+&���M�	��V>{(EG��U�]��jz������%����W(����!G�vZG'���-���업��
�'��B�Z��,�mQWaƙx�.I!{E_pq�f$Ro�������I͠N���s/$�]�6^.���P]�3�V j�yH���{��K/p���,D��+1�Y�{W��5�ߗ�Ē-c~�->�B�	s�掏���u��뚙�r���ž�H%��S�I�J��ob�i���/�ϕy��&%��,x��X�1���d����/|�
�8�	�RT�D� zy�T������L��.͟!����o��Ͽ^~���a.��/<<��Z�YM��B��y��X���Q�[����<4��x��K��p$~����uc��S|R�?q|�
4��m�[���ADTnG�"h0WT�.׾�T|�2Y�I�{��F6�x�J+��� �]<��G��77�5�����R���o/��抂�Q-:�$��8�n!cX�s��|�0���$���e'��@���#*�H�3r����]6 Y�(���;V�p7ʢ��Ӌ��C�$"���DD�!"��B��;����V��6v+�C'�{����B�C!��bB
	���Gzz21D�%D�%lWG�gB"�̡)� ٩:��:Z-��!���Q��Q�J���LY;����tr5�~uT _n��ϴ2v�%�qn�������m�:��7��/��[.�j|���B��[�R��1p�x�+�z^�a�24�12@��}�6͏1C��y�o�&�,��b��K�rּ���+~�.	���b�ީu��!0q��5�Zj����랁�ie�S~�씒��' }~�r���B�2띿j�c3D��� ��N}�1�:\u�\x����4.OO��JR7�������+�x��Wmt!���y�;�S�)�âXS}��b�6�_�ӄ�Q
�T�B�-�6e�]n(������yS�h����p���]��ڢ��h�K$}�nv]U�掌��Sa*�����C}J�HXFϖ�ɀ}�����[�(l=-׋��K���
!*mdVb$��N��COFq	4���Qh���/�b5�F���������c!��V�޷OT�5��xE��/��S1�0����p��*�
U}[:3y@<>�d	5h�Ƒ�c���s|%`�U~�h 1+;3Lt:�u��	�x��b��W�t��CӁ���梤�ݔ��T �cS�O�r�%\���d�3DfX����fo�9�T�E�JcfJ�l1�9^#����[O�%�l����4࢝�N�
���7��|����Y��8��H�'���u��^-Fe�?2LE�t`��fE�����&��UGj��t���ɕS���w�ζ~�q��'�y���)�uA�o�yA���k�����I�5�_z,��A���q�kH4�tT��~�L����U(vι��>�o��[����(i(��T��c̦CUI,UYL�=x*Co���&�Q��l#T]
�=a�bh��G?X�
PS�sN�n9�]u����ȟ^Е��|�EX��ϩ���yr����m��	�R�5��C8Q�@�J4tY�~�m�+�o�>���`q�ز��I�`PM�����G �r���v)u�X����ą���s�T��A���+�'NԌ�!�l.$e�{�a�P߅���h�a�����h�����R�v�v,8фl�oԞ'��x��|L�r�m��OĀ3
Z�n1�GҐ�װ��:Oc��Ӭ��J�/Ö�K⧉��=�A�����OP�r z���c��5!U�!hT�Fk��&UB����'�Y?�5�iv�����{���ѐ�k����V�ڍޜ�Y����x,��'3��������$��P2������2�db��p�ds<�p��^+� ��U,eG�+��k����¿�í
�V*!�}�d^�z_
��W���)C���[�v�ƒ�Os��~�������އe,�B��޷�̦Y��;Jh�F�D�o����l��#�l6����7ej�|c��s"�Ȩ�Q�̐v����prdC=�\_���n����)~����Ru��[iU�A�~��8ʰ�W#�B�͕hʄj����-�ʃ����/����^m\�^�%��o#w���)(�>�U-o�Q��mC&�/qY�k�nYmfyw
���ne����G��o��9�E�՜b�\���:�|A���I?[�h`
A�2�X��.�8b>eN����.���7aQd�+���F���{_~��'�q������g����z���������3Ş��ȏ������F~��mt o����|/���B#������ӽSǟO�oc��֯k�)͡-�g���C�����3����=B����l���yt�K�R�
�ᤈ3%|��$����w3s,ϖ����L��O���ǅ�����ł�F�9Iqa�S�n����i��E]?��^I9W���CWnD�f��h�Nt"{�SS�b��c���L+��-Й�3q����,|H�VG���䧇pZ�%KG���}>���[$��6KZ8�;�B�cl-��H�!D��@1���P�;���~8���[�̻���������3��B5	�M����py8��������V�y�t��Y.psb(*��c  �5l�*i�Cd��p��q��lL)Z@�N�(`�򥁓�U��Uv��������G��2�J��(�^��f�L��+������DZ�^ ��ի�1�O���*���h� z��?	8���<kk�CU.Shs��M�����S%��r(tVN���$;�-����b�ϑ�O��6.8�?\�����������Gd��`�H����ϸ[."ßH�)0�QvH��3!,��4b�M�;����
�{&T�4m�jj2���ϫ��rwO�v�Tp���][K���!0T�����:S8�|t>y�U
�!���D |�{�!�a9#w��]
�����
⑦S�`����A_�Й761�
�:`��TLQ���A�.~�'��8�	��緖����(!�l�d�|��1<=8�ϯ�9�3�����vh��<�K�B���YiљC���̴mGd/�n*Ƣ4~�$~�<�i�C��Lf5]vv�l�<���	�vf��8���A�����x��ͦ����H62;KyH���d��Uw��d������I6����Д�nٛ��gO�m�NO�� ����YZ���W��J�:
�L�E����g ���惺�а�7cI�����7�U)̣��F#,c]
eu9�^?�e�����w`���J�яgT���p�qe���b`�F+�l��Bb/KNmDZ&?Ժ��
�,N��fYI���r����Z	��-ʈ�uڨ�dkIGR����OL�A�)i6F���/��� ����:�����b����я��#>�-��i�`��v�����Y�;(�E5������GD���ۥ����%���[��L��6�Y}?ˆ���)����(1y(�D�*�U��g_�+çRR��h��e��h�Q����Az�G��f����LR�Z�8aY�XC��tR�V�� �1���{��,dj�|��J|G"_Y�E
���KL�2�g�T4�+�DY�T�=H�bO��/ؓ�/�9(��oR��X�V�@R���s�][��7A���hu	�Uy�A2����R�����c<�1{��u�;mG� ��^����|�vE����{��~����d��)��4���~��$�=�#u��o
a,3��bV�ڸ�蘏g]�p�@Y�Jq�������ԅ$p��s��0��������
 �$*j���x�U����%��]�r��"δr��;�iM�'�m�~�K~q
�竴��$'�]��xֹӤ��9i�Aй��ۗ��Zv�Uw�|�� c�K���Q>��7ȶ� �5C4$_�f;�UL��Oڔ��]�S&�;��05�v,7��1;�.G���p�G�;�g;����b<ծz�gg��՞f�a�^b�]��_d�����w;��My���SVLCIb$�wt��d���{���{��<���ar���~����)��4�uG��P=n���8������<���2s��z�q@������*�0�Or@)�v
9�3��$�������ʶ��0E����v(�ʧmN�~�������s�(��]�V]�\�n����ɢ������.��6L���5����M�Ŧ�g�=b��-=ӄ���᱁d�*�w��M�V9�VE�V?�DXB��4!�c�L2��
�1���A��JD��w
�L�v�3�L<UrV"3X.)��0I�Y:�+�p�_��X�	��;x���a�<lp�Gw�̃�M'r�ʹ�5�6��y�+w��%��U�/�nl�^�,9��s}���78�)���gėf�F�di`qr�ЙU�;W�y+V�1�=��`��@!���D�@������^�XZ�2ܼy��X���Mw������f�C�|�P�J�Z �w�w�Od�N�WSY�O�����(�k�/�R8`O-b�`D0( ���:���0r"e@=}�S܉����=�(���O;jT <%�em���_G�GI�s�=�u�~����#a���sA�s�䪝��S�;/B�>a7�T�DV]��<�s�>#s�������P�To� �E���/��+S��������}s���k�_�c�UH]�a��;��1�~ +y0�lr?J�-���7���i��d�ϡ�6K~� `)h��/�Əvv�1��<{�c�2�X�0�m#;31�*J�ڥ�]���Qg�����|�$*&���f�"��U����)V�w�8�M˦��X�B\��P��ymr�d��4�_�"���6B�䃕��`-E�`l���E)}�6�b���S/�Sw�p�BiRt=����%��lCd�	Y2���#���OSKTBEٶ��ʋ��^\�����L���"w��:^�h� �b*��.��U���΍�����X�h���\;��Z�iDg`p\��bo~_����!�1����<;b:�8}�(D�����������@�mN��Z���l{[���m�[�Y�)(T��Db �(����e���z.��s~�it7�X.qy�n:�#,o>���-����ײ��J�]���)^�Z۸���;���5P�UD8`ŧ2���V������A�� <5��2��]��)�3F+7�ۦ].��w�	5�eu�(���L��L!�Z<�1�n����`�S�8z�Z��a���N��񥗶֦��-u��5
S�q�şJ�.��z���,�k���~�Ƚȹ���K�1L���ZZ���h�F�)B6Q�,�|�~."���D���8(f�@s��5�C�g��J]�)�K�F�Jm�M"��, ���!ͻX�ȊsL�[�kXH� �
�d�������+��`�P%�t��{�[�4��M�����	i��ģ�s.���j��w@��f��;�
L7���:N�ϸkӥE���%L�����E�ٔO��j��]����x��}t���S˼Ϭ_9u��W��2ҳ�;��_N�o̶*1�ףQ/O-�!�Q܆D���㝛����)��O˩N1'�S��Tʅ��E�e�6-�INL�2�Ems;m�L2�P*�j�����x��x����1(oz�Ӟ�T�����V�lw�;�s����^�*�D:�m���PM��8@��I�:8b�*V�|1�љJ�#h��dT�w�^k#�뻤������Ђ��b�3�ߢB9[V~9��� ��Ygl�14GO���_�)$z0a��>?�A��zi�L�T��I!/���DG<q�h�hi�xb2�O���|�
��m"��
���߳[�������L�<����1��K���ӌ�Y�}��*Չ��K�d��E�Y�����i��$�ޡ�#a�5�'Й'�Rߣ�J^��r#��� ŽaA�g�W��~������~I�ã��C���I�4�&e���{<X��Qe^fF�������&�6@��ʊg��-���L~�{������jV����p��I��?��dt���y�����Y�HW����!���Es�	I��N�%� ���X���hg�.�U���+\ѵK7��^��z��ۆ����44��ލ�Yw�7ptt�a�K���%�EǬ�A�ש�c�a�r`�R�"��KBB¡�������K7LL̀� �=a�	���>�1Bn�C¸��B|LH�Oc�$�ɉ�P�\=%��b/0�)�mT�T�7؇��޹�('�wo�	�0xAО����19�_��K�`��V�k|���Wό�D^RԆw�K`W��%%�t��ٻ��O�z����� Kc�HL�^��Ԙ�Am�T�s�+-����j����VvQ��~?��L�����e ���6��O)�YL��?�:vr6ܳ���v��5��||��v�s�o&�흣�Fӕ����
��wvT��E�e�NX}8P���波HrK�н�I�@�h��-���N�e�ZjD
04��z�[�b"�݃�K���m@�-�;�䓿��{4����X��W��eƛ�:���v���d��;Gܒ��z����$��X��@�:+󅌼O��Y��<��΅�o)I���Yʾ4{yX���	������Zn	z��;`����2�N�B��"#���F7I�Q��-��Gی���l����MPl>�%@v-"J%��L�6媙q>�ܝc�Q�*�����^R�fʥ�B����$�i�>�R�|��FƮa����RDH��XA����jاgL���n�
zŔb:���(�{�THc/��#������!��t�>ճ^560fjC8�da�Z�h��)�����F��kҭ�&�S?e��KӐWSʔ��?�(��|d�T����l��ӻ9���g~����ww-�r73.t�y}=��rw���~��XB�o�]|���@�Ɂ�lhE���A>�M�,��37W��dT�)J���06�<Z�pz������M�i����9���AG9�� �.ukEf{|%Z�~5���.��<����%���!Ef�X�ŉ�S�#���(c(�}©�`��\6ɯ��������������3Ԣ���� U�ԏ�ϴ�ly\?�	δ�/�Y}��P����К��[��^��,��;�b��R
�n5@��-�<���s�魲&'o����fK��{C��x�Y�nA�c�Jf���o���ݍ�Ģ�n��c�	K��C�OWN��k*�w�Z9
�Km추׭�E=��I*��FH;W�}�u�;>��h��	�;�$5�c�yH`c���]��܍6�� ��$0y�G�|��W2��i`T���oX7���C��é�*��t~�� t_����?�L�GD�s+��M����8(٪�9�J̦���hD�WO�
i&�ʒ�v,��{�P&�����N͘�܎�$�hg[6���p�X��.a�?(�VE�1�Ǫq���!䤤+ǁ�N��������M7�z��s��V.R1��V?K��z�gK�����.ʵ.����]/�)>9�e�GxH�W[[�a4������4�.T�y��.�)_0��hn�=�b��G�Z{���U�c}�'� y֛U��d3V6=֭NsT��#�c#���y��b�'9R�
�����Kl�!L� ��f�Z���_�`O����򘒚Iq�Wb�<�=�I֞���G>N�uUw�ҙ����6���1�(�H)��T-�P�R5�:���>1��Պ?d"�	MV;JF�����΄5�����1j)ώ�v�V<�D`�G	M���!À�1�
�̻yԟ���NND��9����I�[��n]��F�E"�Ok��}uoA��*o�#�?�n��ަ���ן�7c�;"�h7������ؽ�}�䩝�f"�����҅.����䚋9�I�c��!�E���W���Kj2x����������h��'Jq3pn�O��Q
�Or��;�7Lo�V�͒�	�>i6����
����fվ
"g�"����)-�7��v�3q`ߡR����NO��#����SOj�B9�'[�sU^?)��T{�J�AeS࿵)F�_Hl�:�J��۟�k�\o#)zC���|P�V4v��bA]�X���-#�UYڣ�/C�r����U�]�G�X��=�l�!��%�֏�,��[.F�nף��o�a�T	�l�?xb��r��,Ϣ�۷De���>��폞��`�b��o�*�D�#R�}�B�ʌ�R�r�,J��'d�L�T�8�	D?b˽���L�w��ʇ�� ��k��D�؟&M�	���2�1pF��S*X���rLq֭���Ql�	[�+Z0���5m}s������O9밗�;��?��|����'{6\)}j��|;�� s���̣9"��GР�`�I+� P�̽ޏ6�Y�����3M��8����Ѧɤ���W�?c88�y�c9�T��C�K�3�]��ݚ�&j��6)��[=�M�<�ǟ�v��$ń��JM��?���]��x�Z�����?�5����0��x�%���k��jtf/O6&�\Z�Gn�ޙ��Z���T���J�*��a<sh���	&y����Ў��\s��H�^'�3�b�1c$���8�*�%!P�]��e���.T�Ã����~0
us�A�?T5���w_�a-2b��9����TxM��Ώ����n�4!6���!⭃��xm�b�@�6X�]R�)P�ݝ���P�xpww-V,�C���>�9��_&��L����[{���@���^�p�@�����'�B�,@��ԩ0k��xZ�a�?zF�u�����P����T&�<��GR�U;4;�b�X��T��J�k�z���?�h�����~���v�S,��f�Lo����#���{H�,��</$���� ���*_5NM���T/�Ș���l�N��2J�����2Z�˓��1+���U����� �)�7Z,9�Qy���]�)����˝B%M�Q�ͩU���'h�|2_5�b49�����I�#���U�_���=�����uE��T�0���s�C˄�E�;,m�\��\�l�?*_�k��	<t5�?�g{��@Q�m���F)n�|�v\�귟�=��;���V���n�^f�;o8�=^�Qѻ�%e3������`p��7s���?>J2c��Z^=RV�yc\擲�}2����"�z� hJhibW�&��g�( Cf������~�4�����c��q��g)�X�=�_����~8��\�ǃ�Hh&��r��QK;�X�A�F�?2��ۿ"�HI�
;y��zf�hdfԚO�$�`�~/5@��0>���X*�ك����yj��+KPƃ�-��f˙D�	�f�U`��kp�����=1�u��Yc�f]�7wĳhs����ܮ�ܾ3Y�fŧg[��|��n�-�G�Vszp�W�v:E���/W��~/�!��.k�Sޞu�0�3���gtUm_m=1i9I	�y�e�m�O��v>�Tu:��:su�w-�bW���S)�Gy�!���,��˛�)�|S�m��
}�uQ�u��u���ȟ��r�-Ga�����0hf_C�|�,u��?k?��kd�\Ö�ш�M�:�R���ۘ�h��
�(H�"������cC,c�|44�7�DQ�	(��I˚�S ��d��W]�e�n��w�]Ҍ�2<�8�(��߯�H�:���Xl���M��,�)2 ��#�Ĵ0[��i�i�������O�F�ÿ{�n�Y�e&H�ۧ��_��d4{ρb�p^�PC��ޕ݅��w��&��3Um?(8����E([���hD�;�?@P:�a���T�c��1-%�ß���xI"�����)�1�1101Oo��6�B,@mmd���%g׫,ua	�꺯1Ӯ�D�N痗&� ����*!A�N�D ��y�=�EW��T����Xt�7��1�;n&�p�ǁ��\��]���Z���5�?=������E� �ͪ��Җ�����M��_~���X2����\�1F-�L�,�T�G�� �ON�6�����n=�����Tdz�N��L�o��H�U�U���" �����F�%X�/4���!O�W��MW�	��L2����ħ��:=k������\���.�4��%��c�Φ��Uvvm9������bIH��6⠾3�#-���T���{H���H.�"�W,�Ԝ���N+����U�g�<�5�����I+ݕ�)�؛�c��H�=�?+%L�̋ʌY1�,5�{ߥ��^�%�f�5WMy�v{���ҧ�-�����j�_�x'�{w�L�aq9]z���M2|���ē���LGb��И"��}�/R��ɛKXlsn�o|5�Y�״q�����3��&�2.$D�vV����Mj/�$\pp$hp�M�w���mv��j�ǭ�T�}fey���F��&X�V=(G��i�W�>$���uC AR�2G�]�2X�����y�@��C		� �+�j!���z75&	� ���t00�@��`V�uIO�k�p�lp�u�����添H��qt#x�%��.��Ѫ�1��~�v�}(˘�Y�ͭ�k������,֯�,b�W@I��q9�pR���(��fyNL~F��XV2Hs�E�\����V�I?C�#I;R侚�)�(CDX5h�J~�U�Q���f���H�X��,%D�PtJ3l�0��Z�QG�!3	.����RM�IA�S8�Fݠ�=Mi��A�Y�o�q?=E�2�+nrч���sd�$>#ޏl��?��U�0�8��4����CE�h��XS$4����'��eY�Ha�	��8���ʎY�oIgw5� I?��4HTE��Ԯ�{<�#�*�̥h� ���jl1� ���=8j��5~��yc�Cg�*�0l,�����w��-H�kD��ј!	�C�XZ�@�!��2�b�`����[~@��$�4	k���D��y��f]��l	�N0�1B���t9�Er�Bhp�AS�����{�>S\蝈2ߗy�O�?�K�n�G��u:���$��|�\��~d��qfee�(oml�kWip}���*��D����C3�*�ב����#\�?�r��ЃG`ַk4Я��	�.�°c,�� �#񫖓2�Ȥ���|l�	৲�S����h��&��Nc��v��,�.&��	�e���0����2̛�d�G��9���)9j�����
 ��o-[($��3�֑Y�}Z��N�u��9(��g�n���Y ����h_a�@�-S�#Bٙ��:.���ڴ�\:����� ��k�֫��}M��m�[�E�N��f�S�<��L��+{i*uV =������"��15���|i~�17}������<c}��Qg0�n��vs�J��̅W2��ܜ�]n�g�ďQ3E�k6fg�vڵo�^-�_N�s�=�
,�U(+�@ī�@�/�R��G�
E㻄,��#�jY��h�������x��=��ʢ��p��a|�I���y>��N�À�q�q��\"b����1�&���9����C*���#��~|ge���im���E;���jIn�k�o���N���L)S����@�\{�v}s�8 3�/�cі��;�0H���|�ճ/��5:�T�����S[��V0͖�Pѽs�v���jZ�.��
v���_{�����aw>�f����Y ��?Jpju����	v6���s�Uc��c�����A�ӛt^M�TV��X�En6Q�e)�ZC%��;Ȉ��F�u&���{�ג����G�a�µ�J��SX�\���-��_Ǧ�ԡ �F��a�S����{O�m��(�[�c&F,9!n�Ɛ��\'}�h*���Un��C�R=Q�"�J�����[7<v��tA�I�q.��ϫ��6d�0��Ěn�f����'|E�{ ��7i���Ɵ�jb�?&�"@�q��e"ҁu��V�̳�M�֠T�ѱ���P?��2P��/�!H���iAR�Yz[��jτnd�-5�3�H�����]YR|Gn���Uh�������tRW� Cq* 3�3+F��'�K�T�[� �`� �_j�c�⨋�Ր%lۃ�T���_��:o'��:-We���@?CB�������?1�6ߔ�Z�s.�$���O��a<=����郅�V����-�,>�4 �]�D_�)����"�b��XU����ݥn�+�6�Be����ub;˿�HX`�5�)�u~�cC��_���tp�T���'T�#�U�CH�p�$�(Y�-i���A�O�M)���+�@ J����5T��w�o/�N�#��z�}l�:�c|�H��*�f�0a�p�'�pa@$�AE3�X۷(
i&���a��bd���.�d�)A�V��E�VR��{��}�gÚ��������U;���ՙ�l~������ƛ�X����ړ���F�\��-@={�w+�zN�\�k���z�6�pc�Vvk�5�����dO������g+��F�nU?Ǌ�K��m��U�ۤ�X	�B���f��¾1�9DYĿ�!;ۄ�wnv��Y���)��˭�5܊Ά��)��c�nz�l�
ON���	%���'r�J��Z��^I�������c#(%}��'�ݢ�fm:�����:��OIW��V�=I�~]q���Ckb�m"����A������ŠA����$I��#��ߌ`��=1;xu�ؚ���{�?p7�ɥh,�naT��R�)�4��(��� ݷ��!'7�Xg������X����b���{l,�%�R1q?���wq9<Ă��@��n'�����[�9kO6 ��c�m�p�2����Fb��ts��k�q݇"��=++,��E��c͊+���@H�u�to?��*�
?��7���Hu�lF�1y�� _3�߷K�h׶U�Y@y,Ig4�2FW�z�w��p��i����7��ל6Ȩ��a��J�ݝgM��
^�%b��&`����W\J�@-J�"�8=l^:��"$Wn��,b��w�AtR��N���e��Y��2ƊZ�e�w
P�oL۱�=��:B��?�u�Q�n��
��S��9��B��.,ry4�R=������ ���v�W�nR�A:9sd~��@ (+bXW{xu�m�bK�R�z"۷O��VU�U��/�{�?�Ϭ�?�����zTų�H��@�BPf�@,����*�t�7U���/���_䛾2�j4�c�Ǽ>�GK���=%�o
M�౷x������5�u,��$�'ǰ��I��G�P�ŏTe&��K�<�BK�Pm0����c�U-�dH���[�c6�i��;�.<{�`����X�����|���f�DZ����o�$R����x����t(�&`��a]H��286��Jy��w�A��΋�0��/]a�����g�>�8Z���>��RA%p1�o�!u�J~�&T�����kwv]n�H{m�OP�_�K����:B^&�֫�Πя6��J�w����`��jm@֞����m���2��o����ȭF�� ���LLf5pX��#?ceF��-~�B\�tU)�~��-���G�.��@��7��&�����N��No� ��O����wAaz�����k��S���/�V��/xy_��I�-�9�l!{�b� ��.���K��;���oN�	R�y$�M��������c/�/vu�65�Ƴ����gCaLY�W�bu�EE�ǂ��T^�P�}�N��+��ۥX>O��ꊲ�����D��թvj����lK�i��4E"v�|�,�K�s�Q$���C@�%���ŭEc��z�M}9�"~D������x\2�^T�do/	��챽�۸��n�ܭ�3˻	��A%2nu�Ƀ�zD�DEŞ;�/��B���>�,�7�n�k���;��wD�0�{?�d�*����1BK���|�=�
��7��Ae�?�	��~3/e\a$5��	��8�["�n�Hry����)W�W:��J�����v��S_=m�q�h��x��"d����D 8����~%���\�+)F��9��{W��57���	]�vmO:[�u����h�:V�<n���U�"��V��Z����y%˪��e����z�RI���ڂ_.ӌ�1f�4k*�d�#Z*3<Q@�d�Mٕ(H�0Uŕ�&N��� U.u��d�o�f����$A�;��X��&�W�0��［}']�%��5	AK���a]�'��PH���wl�����\*� f%���Lʒ
%��.��rE���ѹ����B��PP��g
��Q�LU�嚍���>���\��#�r a,<*�d�D��SU�����j:��<`y&�q.gV���]?�[�/�N��'g���x�&��y_����}>C)�F��j{���7�qȥ]��)n[
��E\�/���P�_X��M<�K�Y�+��xJ�	#M��o_ ���� ���k[��lt	*
��D�6����J鶜[��g�����C�:&v�dL'<wG`f����i$T��ۼ�yE�B,�$d ,��*,;[��dK,�$���[�b4��&�b@���{D��CUp�¬��c:N_�"GP�)���W,��'��/M4z�C�7���-�C�	��,�$$�'p��0��'~�#Uh]g�E���S�Y�5����X�_AjBU��P�� 9s��֞�yIs��EC�'a�Z��F�L�V�c�t������3|)�|"h��7@��, b�0s���6O�W/BW?�
�{2	�-��k�.�`u{�A�ƒ���*�-}oќ�ӷ��_ʏ��,��y>P��=&5�	�^�4�����8���������E�̬�i�[����/�-渔f2z]���ҧ��j��v�dԳeԾz�R�W�Zn~�9C�n�A�v��(s�&{taa��wd辝�e�,�p �鹽���u�=��=Ʃ�q���L���<�����L���Q��A�ڪ��Z}����TU���6�̔��ð��s���Vt�F�W0��}Vt�׷�A�����/n���e���6F����
���#H� �ۢ'��C�T(�6�8nlV�yv��50��a�F���n]�fI�芫$�%V�EG�Ҋ=J|�K?��}�wk��]�4P�����Fo:�w���u뎶��qL��Ej�w�������'�E��MP���iީ'�T�=�e��y����$�2���_9�����KM-�&s:(�X+�����@��b����7֙�!�.�:�7e�U7ÒO�J�un�K(����Xs��+�0M�j���(�&���Q��a$-N��h�ݷp>	
��I�Xg�{���pHvW ��|�GQX�/F��G�=l}J�P�[HUKC�bT���R^=�aY��U|G�д�IUbj���ضCrM� ���gk�%)����̝����uj9mm���GB`qL�/�Z�&5��@�o��`�Z�F�Q��V�}�=���2M�S~m��}�I
 �i�Jw���_�g==�&�y�or
v�/���ڌ}�����0��U �iatF�M�����>�1k@;�5�T���,Wi[(%x�����]�t��T�%�~���,F&���H�J�G��O�ވ]��|��~��߃wh��L��#�7��vZ�`�f�%���Q�|a�wD��TM���L��!�s��b��[�����w35��#�G�\�+�K-�p�%��$!秸#�b�?d;3����аy��uw ��u���V����pc�����Of�j�-uU?�w�V,=�pdN��/��R����_�d�|��$�+Ҭ�KC/������C�2��rU�^��_�V�T̓~����l��K�Y�{w�9�3C�:��v��6���h�	T��o��U$~|�4�(g[(β����^�l�Cƚ�<|8	n��-�,$���ɲ��� Fr�20�
[�+&ط �����^��"�S�����9V�fՈ����?�z���~�">���]BB�N=:���{�O��i���Jhs]Q�4V�Q|���"��Ў��+�@�9ԛVU�ބlנ�v*�}�f[��}$��xn\��4C�f��s�'b�q<��޴�y���w�b�A�Z�/�Д���`4�K�BLOѮ/6�%&�C T-r$����C_�d�����M#Nm�) �Ñ�K��(X�٭�g��Z��w�%�Ī���R�)�ȥک� ,<�����pP&�����g^#�v�V��
A뢵�e(s���j�[	�'��Q��F�`�)��v��C�?��88�G�X�D3�l�u�?�s�e�R�W�6�8&�\Z�B&�N2�T>*�j�"����A}�����N��l#�������Ƭ�ɡ�fӶvt����㲝��3����1{����B� �͕t����׹��yHI��[z�H�8�8����"j91'���=.�����ڌ��X4�:P������Td���>BQ�����r���r��V=�Ի�����ϣ,@��OI����k��'�O]x���k��2cggy�#@s�aA�Y-����H��p]�h][Vx�r4��Ʉ�?�Vt��9ʋ?Ip���n����3]�tx4>�|��Ȕ�R�Rȸ�e8)�u0������n� ���8�s>�����b���Y��ڜ�}�� �#�!��
ƻ�s>�fgU�𭆵�#���뎇
�󑟢<#�w?��z�(Q�Gŀ�'�h7;ځ�o��`m�����1I]F��]&�=*�]0��5M����D�1��v^�9�Đ��W�t�*m6]�0l�L�J�"�O��)Yɩ(��(�psg�O�$5$X��t�h�懁qP0��F]�iJ�?j~�M/��<������/�O���+�����#�$gP�C�)�����YN"[Ff܆�%������%W`��I)�,����[�6����k�X�/$�P�VA��+�M�p\�d�#a�)<`�wI�.;�^٧��&�)��x��X[�<$�}��{�]��J�۠�~������N'��B���-ię33�Iwd��UL�s������8�mВ�V��n�P�3�ztՄ^�bּf<R��%#�^�oI�G2��OE�g	˱X�ם��4�w�Vэ���E�
��UrM;S�)<ͦջ����z�����A��B�� ͭ�:�Vx�aHF�/�6i�~X��vC*�iĐ����~�|'�W���_�}�J
�֎l*�HRGtOT��@��-;Ы4������b�tc�[6�����u��Z�Т� ��\�挤,��bDќ*��D�"�[��&:������JQ&��M^�ۊ!�۹��������J����A��,�WW�X@]7�߉1Pl�J��h�I9�4 �1���|7�L���
��/�Z������
������_�8�,�0��a�S���Q>�CMD��2bD�IF84��&.qȠ�ܰG�+�a���m|�g�:�F ��*Q���_�+&�%j���`6z��&�wlt�����TvBV�o�+fO� ���"���t(��W�0�x�A���QY���6�b�mU��I��;�O��ҭ��U�lk� ��9�pL�;OE�P�iO}'��DF짠�X�����D@��T�:<�Rܝrڋق��&���X�᯲�F�UA;�+����}��ڻe���l��+l���0ߗŭ���l�n���ؔr�ñv�6�/��%0�q��Et�xm��q����a"�5����J�r^|�F�����le��Z{���;W��3�`,�c�F ����+2��J����Rvm'j��of5���i��~SP18������D����z�q�r��k��V�x��HB�0v��C���:Ub���^̀h?,�l5��M�I�b�m:E�̡I���,�z�ฤi@ħ��\���
���X`�o@���*��|yso�='���)�7S���Ue�s���,=>y슰��"^J����o�5�s��N��|N��3&f��,�mW�Blg�j�� C�I�}s� ����_�c�z�]�(睤?>�t����'&�;������`À�AԃͿ؀j[�x�x�c���?2)_J��k$�]�T��
yl����{c�*��G�u�{�ièdPb*��z,i�(t��;Ո���X�8�n/�o���D(x<�~���3n��g��������?�|��R���j��%4_&S�ܚN��F�ķ�#�L�&���:���Z*�V�I��h�1S�Q�ME�#ٯ���C����̌�׻��׼��CN�P|������K�l:��_N7{����NSƯ�u�xͫ�-��~�!/F��.�R��smɦ��j�iMAߠlh&�ֈ�}F�%��<6Qz���X!�5�ИiDUu�-���Vk��{PB+ݏ���\���|!xg���(��m�<���4&{����5f�E_cN����a�B��?J�3��"\xC\ k�������Jo~;ro-�@*��(1��j,ـM�#�lQ�8�J�g?�z{2{���O�j>TN`�M"'9���G���pI�V��u �2�$�1���Oj�������p�o��V܂	�Kf��IW���W��;�v�T��S�c2PI) T	��fY���lS�������
ׂ���QQՖ�����b.�����M<�?x�[���^�� A�73<+��sY?� ^K�� �
��E�z1��LAs{��:z��2a"�i^Y��k\����`Ϗ�j}���Th`m��@���2�>���PЕ�쥞1�z8�+pO������>��4�ӡe=��	Ja��{+_�ԭ��&e_��FhKs������s ��3Ȉ��"O��;���H %Q �X���'tK��N.�T)���Ι��k՘���i��\xXM��2����	�?�n��\�n�	����	�����^�[u>\
r=LW2���ouz�t�w�^]�?�'����H���Bku,�����)kD_9�ї�4A��듍i����o�#���$�x���겖V�0���򗖃-���?$���>`w�����=�"q�  7����(Ȯ��Z�h	bbx��������+�\�=$AK��>ؚ��9����p05:X`)%y)��۟_��rjB���6.x���y+�d�nF&ӳ��(���RiY�shǦA{u+ϬR�d�T$Z�[<�[/��6�=��O]sa��q�1�}�%^��v���ݓ��?P���ľE=�#�sʮ�Iyl�G��H}��M_�O��HįK�/�b�
H5;6@���	5Խ@R��2�N��S�Қ-7UXJ�K\�P ��⨱�`a	�/m3M1h�p�z�ZN�6Z~�(c�Q��TmG>�[d��o���M������l�#����	�T���WE���x2xq�R��W�Ǻ�ġ�`���]F��7���T{l��^d�g��N�a���������~�].s���w�n�(��n�_�u�^�b&m�{�#���m�4�2r�n��
�hUK�aU��[������������쵗���Yvl��h�b��]�՜��F҉��Y��� ��i�K	��>=���~i�8a�7Re� �B˞��x	,�Tj���F"�Y%Q����2�L��^�x�4<���̒���J3�$f�4�[5�=�Z���L������-]-b I��+pu����q\FBL�2<q�e��4��E���Ꮀ-��v&ںfH� %��YCqK��8�7�_6}i��
��1�U��Ԭ�QQe���!|w�`���(�V�\5'a��u��+�@Pf�d6w#�
�ƺE/6��U	P>B�a�*��$���:8!�Q����w���x`��i
�6���@p:�M֍��՞N7I���]��]Q�2;�V�ŠS���r�nr�d����,�-gNY%c͕��NMj(>��e*k�k���P��Lk$�2��	̋�T_U�(�Bȿ9���'!�K"���������s��Υ�u^��'@��Y���20
����G]�%�F�� d ����&��d���
�V��u��г �<�{~���\�lk��<�����{V��ϥ ��=R����y�g
�h�?[� �X:� �ċ��J%�beʊ�dE���t�w+�ZT�tN���N�ϝ֩�,���i<�%<_~��=U�,�t��>�>��~���n0U�mZ��Ŕ'u������u:�J���X��4�Λ)ɡu����,����U�ե��iF�����$��� N?�W��}|��?u�l����}Rz	:�-�����=��/�r󚂒���vl�aK9C uH��6`�������F�5�tFҶ�͏W��=wngؗ��~����=_P߼SF�~�>"켁=�]L�'��eeU
� u�=;nGE��q�o����zHV��p� ��/�Z�ԧ"�ާV:g�bQ�⦊0πQ�9pк�)������ ���hN�����x��Bt� �1��:݃Օ�*�tu�e1�ZF����|���o䟱ߜ��c <ޒ�gub��ӯsm��{��s���.�m�9�\½%n��t����y�e���Px`L>����L2:�J\�YI����I]����u ^��{�qn�R�2�@�"c��G4�ޢ���W�jQ�I|�W>U�av�� %��K�V���՜z n=�*�突_���r,|�k���
Q�ѳ�S|��<^�
\�����Ȫ�W���L�yW$F����
{���E�\�9�8FEp?�,����,�a����7���M���[OR�u�?9)����ps���ެ���t�0�m�\��x;�P���q�QK/��S�O�������4LG%�=�vT�\���>���{���Zc�:o�0:=�G^�s�lͭ=��n�m�I�m0���?�ًޛ��w!;��y�;�;:^�ɠ�M6	r9��%���a��%Ԕ-Q��Z�U�K�O5-���8O�G3N��B�PT�o�N�"�2���8�C҉��N�a���s�G�-��>�P�*�-~�va�X� W��3��ʳ?Ry�Pߎ,���������Q�g�؀�=�H�!�.����P�nf���v)PCKp�*�D�X�|���Đ�a��o�µ�|����G)��A:�<m�f�x�|��~�_��T11j������g��*��6������κ/�}��\Ȩ�� GB�<�ײB;�UiU�Ɇg	���{�y6�a��{�ny���$!�ckl`a68�-mԦ�)��@,����g�F9��LA�ƴ��Q!o����=�&v��D5#�|�)��#)��N8�Y},ח�jө�#d`��dp�@&�vW 2hj�ru���G���Lsk�b�'9!t�YU&l�2�ͮ,�nr}�����GBvdm�-�&�gE��Bl��>V*ɫ���+�޼>7������Nź���Z��������XH�Cw7�`�v�k�EXh�C>�k�6h��Jiϥ��㋊�x�խ[�仞�s�%f���݉����K�/'�/7��.s�/n)kϝj�ͅ4AQ	0��r����bnM�y�x�_��������ʠz2`��tt���E;�r�g���$��^^硗���l���wm��JУ�0~k�* �JY>�'b�mwV��ߟ��ZaC)�w�
|�;�Ʈ&�~�"_��M4]OM�=^��OT�`�I�ѥ�ry���d��+�x��R�7��Wsv|7���w���D��n���L�����1(�	�h5k5mso�,��qU�M�!�&vY�I��C;\V�:�tBΒ���/?O�[1Q[Kq$�@xtX
��*�ԠKc���m�Q�|P���2�Q�6��u�-���[��/��(�*N��b��`� �ؒ�\�KBw<1��������޹i齍����YĜ��n1s�A7�\�̱�g��'�O"?R�3pg���:�Ȁ��%NO�JXȡɖ�&�#��N?��	Wi�|��6�U+��	�DX���/TER��čAa�w�h+X�k�Q�4�L7���k��5ךV?ܔ@�ke#_b��q2%����0��\#ș�I�Ƭ��M8���Y�@�m�~�	�|]�S�[�^*L��]�`���������c�3��>8��чB>�\�*��kn\}w������u.��
����;���/��'/���z��=�z���H4R�Yл ~����LW���^H/��T�yWĵy��}c��v��Y����r����
���Q��������ӟR"�=V�9�4�I�&��Xz�&Y%pϭc����8����_�&����?>�ZWW�G�B��;x�q�Iכ׶���:�����0�S`�Y<�7���Į��e��_��'/��1q�U%��	�J�7p��TNcQυ�H6��L8�Z7�j����-�eӷ��
7A�al[P����)H���3���/y����dG�	�ۇ����6���R��I��B�P���=+н����l�=�*�j�w|�Ҫ�fL'��0�d1�%���}��U��(��c��Y���83�E}����o���+sfgҕ�q��؏��.�4F-�j�}�2���a�������H�G�$�5���C	��K��O�nSR���|����~�����݈p��y31)*`gN��5֓�kE������J����S (59����BF.+lS��S>N礼.�7�(����ծҝ��Xx$^�AL�:���8#��C̯��h%3��P
5�슘����L�͒tEW2��d��m�(Շ���� �c0��Pv�,%޳���֊˩\и��<����+���\oxZ]�TEx3!���n����aY��q���z����e7�ŉ��O����K��ay�W9m?m;��'�j�t������dk�e��-��X�D��!_��?g�����6е�[�q�ۇ���0��T2���?���z�g�W��rKR�ͦ�ٯ<�~@��X���*���c�W���7�S���g����$��L�r�|��'Ы�즛ˁ�9e�Z��V}�V沞vR��j�_�	�@Bu���혢!PFY�
���L����L���s�����w�^:��Dh�y�x�F�^��p�|���l_��ZT� aK͕b���"�W�>,MvV���C`�_9\K��v����3�"|�[�dOp7�\u_,�*i�$�FU����3v|Xke*�1������&��f�����x ��J������EG1��:�x5��1=:16ѫ�2` '�,`��z�F�R���o�Z��J�޸�@̖ܸ�35F�6�P�8gY�!��ci}͖��\,�q}0������4�<���W�:�/V\�H��)+)H���|^}V"��6&+���v���v���Ym@m��Dͩ|:�@'�e�ju�*��l;����ȼ@� �^Ġ�'��� ��� CἪ.�*8��N���Ñ���;4DoD�_�����^l��໖�B_hh\FA�0�K�L��T`�8~�6��M
�56�8�<�ea/a'����d�����	��[�1�������\_�����f�0��Ŝ�!6�#��׬��є����
I�qb�CA��o��ɡ����i�2�-j{�?71�-�[�.�����Z|��E)\��1�)��V0�#�g�b��'���DRoįr���5���|WN.��.���C銷�5p�"���m��i><�
���`q��ˤ�:�^9h$f��]�u\H�5��VG��AĲcjvĊ�,�6@Y�欿��1���=e��j�ˌe��`���kq�ѩDt���]��_��z����fZ�(�g�R��H����P�Bەq!:Zq��9�{��aK�&J�v���%��ً�A��������,��g�}��v�Z�|Z�TB�j
��u����|"��T翃#<GH����n�.�c�m�	�����Byk������+�|+�[�/!?Ax2D�r�P砛����)0�з@���BF�E`L,w��B�j;h�����#�A>w�	ees��H6��[��ـ��<p�D�*mj��Oׯ�����^W��Z���*�(X��ܬ���r7@Uf@Ȍ�&82�rm�DѰ���?�Q��l�Ne]��:f]�����K�2)a�On�w�Ibߺˮ���rC���)������.)W�����!����������K�N��ߙ���d�h��m��8G*e6-�F�a9��^�=@�"%�}�L�1��`��n�9[�?���We�.v�������m�k�u��*A�}���$O��WmHb���P6���V�?��ߴ��T�}n�O�̩��l�6[P�c�g;��&S�aVf�+���:��а��S��<�l��&b~y�k�Xd���{4N1?Y��í��Q��ꥳ�CY2ci����!+r| �LabfuJ �����௭x1n��{���ON��ezKj ]}\�R4��F��B�6f�������J)�Ǖ���2Ө ���>�����*^M��˚��@WX�ה�R��;	ӡ� :���x}X�o./0/�Q�<�IǗ���:�Fh}�H�c	MAm�\Yz���Y�7Y���~qn7�'k/܂d�v��>;����X�=�=�{sW)�7�7���5T��K#\=��'`M����Dd�f��>�\I�4�ل�j���tI��b�T+�. %A}��G"	�P�N[�L��<3��Я���5ɈTJpU�z�5k�u��w�	�O%�|�_4s6o0��j兑��-��(j�M�����'Ix�|��F����z�<�Kn�c�=���;������A�/��9j�O�Ϟn�Eߍ��m<�{ Xd �F~{~F8�-�"��|�L�R����`��&��4��� w���c�ؔ��i\�ek܅���,v�;Ŏ�?l9�\���?4R�>�]����-+M���f�dђV�ff����ȑ9p��bF�GƟ�X�?qta�C~`��^8�z�t//m�E^�rv���%ԧ�ON+��a��"k��V�wx{o��֓�t�F}��Y�`7���"�����>����F��M�#�n�rPF�QF��s���6ت�ŇsM)2���v��Jκk���>/d'���K˖�F4,c���a0���D�E����հ�0�`9���6F���ꭃ���~o<����6�C������5	�www�E���;/��ϭ����LMM͙9��O�ӧ�(9��ꕌ�������[��w6~~��� �����^ř�n���_�!�?f�X\ݶ�|�#�$��g1���N<_j̋>M���/2����g���Ց>�l�7�W�Ȫ�__z�]�7�Gt���HYc2���Hy�%���;����Γ�Zd�1j�Z7� �c��G*J�님�~,�Nr|��g�W��	����5Vs����-�+����g�Y��ʋ���Uo8*MN*�����<�p��gz��F��
!��?+?�n���3!�o|x:Ϧ�K�7o4|P~�'r��!%j3��+�T�q����ꡏ��z�@��.Z�	PJ����I*z����=kL4��Z����y� �N�N�k�t��2�7��T�W~�;p��>ڗ�j�ճ$e�~$Cնov�����xI�Q�.f��t�м?��/���w-�TJ�����lv�t���&Ը�~�봶1�vRuF��(|*�������β)�A$��m���P��2�� �Z�����:�n)�7���u��m3�6~c�Q�j5�*�sõ��~��{����04,#���r�[�q���?�T��	���w��w)o���eah+�~Oď��9]מ{�2����+�ț����Q=�a=���>�����O����B��� k�V[����!�l���϶��+�U��ah�㳀C;B�_�C�����H�Ͱ����Ly��q�Ψx�C�b�A��\�^�[��a{���k����끵�LV����8�q\!ֲ_Uy[!��!�� Ͽ�A�/��k���_�0^@�$�g��O��~�T��8�W�e+	��ʟ
������۱{Ep��>$�:����)[��Z��T�\`�5�L��ٲh�%��&���s�s�-���8��0�!�L;o4���� ���dS$��հδ-��E�k�n�E�)�����%�W:���O��-�G�6�g��u	��f����9}b~%�mj�2�O�d�ٹ	ƹ	8�	&�ni����uX\��@��L����@^fg�dM<�>�NŽ20L��NN�TsS�	��u�V��x
��^.n�cI�eW/M.��Fs�6��=d&!���ʟ��c�x�'�Bh>7}��e�\��G�`4�V�?/����K���[C@2)�OO�Im�	ki;���N��@����|U��ߔ����{K�G��G��v�]�Y��@�I4eߔ�����'��7��,�%���_
o��oJ��*9*)}3R�Rr|��IQQTȉ+��!7lfϞ�h.wg�������0ej����T�}55�ނ�O�.�����i����r��)!B�u&��e����2p�m�w���,�Y�l��c������H�juY���c�"\���߿'���G���^�Qcؤ�I������n��-�:&����\�DaNXȒ��2�Z�u0O.��Id��N�T2R��fEF�����3��NٙO�o��\`��1fHRC�@�P�&l�/	K,ĄyCp#�Ʌ�����
 v�-+%`��M�X��t���U��eW�V�^�t�U��]t	�M~��7��+;[�%����oĘCaڧ��D�ZCɼB>�1CC
IB��{ #�s���t�2x�+o'K�u��Nz���{�>�_�H"�-���a
�-rBd�.��l��_CA�����ט�֫�S}Y �j��K���pm$y$ƹ�J�_7r�T�:-�b���\2��A�,�L� �d߻�b��Nȭ]1�~v��'q���5��Ze�7@K�m8���i���_����֜	�u����񐵸������}Y��yK+0xzp���n[��O#�RD�T�5��/�v���8��g��/i�,@��k���~���w�z4��!$8�<�۬��-`>?3�l]B�Q4�%�D4��L��.4Q�)�6������Q�&2J�ۄ�_Tpp�c��=�X�['c[��~II<�(�Dq{�s�U�F�<�6~�"����R)8jR"��"��h�n�v%�y���_pm{S�z1���+Y� �_-Q��̎Ε��]2
fe�O��w����$��Ѽ��^���/���w�Ti� @d^R#��FU��N���uro�@I"B�(���c��U����0h��ֆ���g���R��O�o.��a�y!k"G���ʭ%deF,Q���c�1���"��.�f:\xx������L)@��?p�C,���`u��L�7�%b��kf��q�C}r�l�O?����D���L������p:x̎�`�)J}��W�����o��"='r�.��O��"�Ⱦ��wo4�{6]a�m�����"�pD�?�	}Y�j&G}m~b�C��+���O���shZh|Vjۋ�XM��/G�z�'����H�m�����:F檡���G�^�ぞ�M����t��.^���y1�&+��::f-����Ϟ˲6��u7�җ:��:?�����q�C���G���H�ȳ�G�ɇ�?���%3$a1Hcw���Գ��ws5�\�_n�x��Aۋb�&R(e��a��j|qY���_�hߋ��"��U�����Ikm���7+��E|��>혠���_�����R����h��jx��t���\
�)�7d3:�m��LWAb<^���M�[Hɸ��F�b�t�	��l�W��5���3uk�!��+ڮ�%�����T�a��vL���ϨNڿտ+�n�*2m�-T�e�s&�����x:�E,�uD�>��?f	2x�xO�N//B/ϭ���흡�Azd绗|�
�!@���+j�H�u袏W��vb��%��Ɗyq9Յ�T���2k8�9%D]�QJd��YL�^2-�	b�/*n�,�#�hd��[��-WK�0ۻ'vK����/~��Wu&�Ym�?���h�
xvQd�����'��e�,�k�����C��J�>#x�!^\���C����j�.�.�&C��2r&���zk����I-�Á��CV�&uTfՇR�բ�&���٘'���0�1���`A��������I�b�f-@���c�VG��0t"^4	���:��t�:1EEQu�i��ܠ�Mss��\*�����R��K�Y�y ��}(����M�����A!����˶���#L6=;�c)@��R�&J~5R�s<�F{1A�K%_��o�T�(�(�[�ؚgR�&e'��I��o�U	������|}g��D�m����>c:���X����������b=��nx^I�υ�L�	��1���yИR�Km7�Τma?��d4m1~�P�P4f[fR��J�B���6X���B���W�l�_Dg��D*��3�_$�A��c����_�1h'�E�"��)��4��5����Zπ��DJ�s����m0�KXh�p:_]R �1�|��6������v=?�W�A��˨�cp���#�Ќ��,	א�\�Zf	���v����)��Ͳ��2�����EZ�����N����Z���b����}���F���T��n�O�3�5���d���SIm�T�*�1�6�j1��,${n�Z���T� Z�-.��$O���	A%����I �[NMN¯>I��������0��/NH��P��m-�V?���0��)iM��~�M���ĵ���^I�H��f:�OO1K��ҹ�T�k���N�7?lr_���<�W���C�H��v�!c�mҷ�QY+������QTF�F�A҈�2F�P�ɛy������?��˟N������#�� ���.��Ky����C����"C���E�@aR�ݡ�G;����i�����jY�6<�V�pψN��*�撔���X�}+�d
���ߏ��U����e6�tvR�FV����+h���[��B�Y�Ã������J�e�,�ͺU�;��Ԭ�p�_=L�#x
:�����뾾�=��&ly�6O�k����܋��8��	�+'�vֱR��-r�}�!0p ����kYG�V��.�j���Ȕ���10�0@m^T5[�5<"�o�t�&����Gs�`���X��VW�m[]<��^@�"�K$��@��3��x���QD�{⁍Nt�W�U(yYDs�KI�7�%s;*#Zu��}�7�ߙ�}�>Н�	t���:��ߎ���s��^�@gNB��-Q�O���ԺU;U	3��s��K��u�-�.)�����qYD�H��KQu3����y�̻+A�ޫK'�^�ֵ�6 ����T
���IA]����r���||Eɘ��e�ڟ�_������ޜ�Sp�W�8� D4)*Cr�{�a@��^
�y� �T|��E���ѥ���/��w��Tjmcy'�@�ߖ0j^225��Ջ����Y��~�:�5K
�9N�&!�A ��n��]���?�w��U�n��5b�������,���7�˖���dn}�ҿ��?���ϔl�E?��a2�"��������ǌaG�\�{�W�vM�Y�PM�1���-~��������t*�Ɂ�=�É�D%��^f^NnzAffn���}^�?�~؆�x_$���-���'���ٰ�E�C��pOÊ�#�e� ���B�������|߻㤊�����êߛA��������Ѧ蓆MFsÓ����������-�V}�׬O}8���p`�p���Br]��K�R5r�| �-��T7��K@��㏫Vތ�HҦ=�;�%�Y�Y&�ߑC�_v���5͹�s���L����dC���!��2��$�;���\
}w���ɩ+i�	�ϖ��ۭ+����y��n�#p�Ko��'� ���p�4�0>���z�j�s ������#E�����p�8a����ä	j�Vғ/�w�I��^�Q�2����p �%�̒����v5-�y�%2B�Rv�k�!���R���vn��#]e�Z��HT�\5T�?��������x���u��F���2������r���A�֒�����$��b�C`���<;��I^W5P�{��G�(�� K�S�O����T�"��s�}�ۂ��p�g�Z���T=�,寏�#�QG� |_��̭�-Ѩ��T@����ia���Y���=�vrBD{�������`[��b�t1zx�Ҋv���]"=��6M���H����"�R�kU1�u<{�&s�%[i�T�E~��([���\g���*r_��ցw�j��B��|ra����P�����if��N�W%�c\~��F������r%
yy��>C�by(O�Gw�����Jc��f��ݤq�FO��ݹ�[���d��ljaM�Y�#�����m��޼Ź��1��oh��7�A��Nxu�'fY� J*��£�E�x����eMZ�%b6��(�{�G�n��$ʰ��j��AF�o��:��Be����b�c�Mq ��%/���^����3�D�lkZ�-�Ə���{�ݕy���5���y�w�X����6\��z��k���̝�R$���ި"%?�l�_��!�B1�E����뿺_[S�0S���3:Nu�s��_l]�'Yt�,,���k˺�F���7gڦ^5{��.�e��������M�44�m����WQ���� ��i�D�nQЫFT��nM���ٌ��mmk����l>�����w�lfW����-��G��W�'+����c�Qv�W B����j`�ڿXd�^��̹E(���w"J�4�%�Ӓ�����#E�*�X%_7���^5�߼��7�K2jh8<�S8��Z H�0��`@B����8����}$���D��ͥW�Ӑ��1�*�9G=��0�/��}'5�r������#j�}?w?��(U��ed+�%�<�l��_��No�v�&ʫ�qH|�Ec���#���@���E��v~~^Y�><�!T	m��]|���\����:���湨䭔B�
���.�����MT%c��^��K�xf����l��|\6��I�yt_;�n�鲬���w�؈xz�V�
�A�ƕ,�Hv�7a��4+�x8��?<�:�oNvNRP0s�������z�9�0�� ��I��ۗ��N��'`�<1Q�x�۩�+5����U�f��\5�ީ>�Q?�JH���H���O�Ǡ'�"�Q�w����i�-���
*��Xz��:���8���1NC�eFU��[j3���ar K#�@���߰�%�>��yl�	@B��b&�jY��1�]����.�c��v� ����7f�t4.�g�;R����3䑾�?B��zQ�n� $�rk�|��j�W��d6n%�;�[�_�q������җæ�5�V�鷗L�w֎2�'�i��x?X�h�i����i�R>�+ֈ�+��]s�-a�ntr[�W�ʰ��wu���s����/��}�4�Dbn���d 8��܆�g=�y!�1��e-66��mCb�]}Y�sVq�{nZ�8�ɟh���S��~�|D��Y�����*����?� �����e�V����&\L+��RxB?� ����(ΧSt�,?�i!?�R��g�Ƿҥ̢�Kd�K���_�cNr��wt�Ι����G<�z�L`�h����`l"�W��؄.�u�lq�ס	������B��\mMT��t��p�ҝp^z"�&��Ҟ���n/n�z�|��'�鬖T"ҭ�<�DS1̧2��0�\���aB�N��v�J�%��=�U~�oQۈ!p��O]��LNυ�2�s��q���O�x�����w����<5����0ݱי��y7�������k~{oO_���#d��j�l���u������*�����u���~�_�5���;�ǧσ�L��4C������D;ӝ�a	[���^Y�.�����T���G^�t��������BP�Rw�*�kB�j���������
?��
<p\�9ɰ�SųT��W~ڧ�3�y6T�2����D{n��s�ʒ��0)���9o�����R%G��m��N��̺Y(����N_O��q��0���#cd��#��*mo���MT"`l��tJ�`��fm
;�wv~0֦��Gi�o�u������J�uj��*���s��/9�ӥ��
	�-��2����2 ���������>���b'�hіFh-����A,�L��9�ni?��eXA���}?k��oeN��8A�d�QbD5?��CW���X\Z���*��n��vۆ_�~>��~����%�7�!�dU��F*�1��T�8�HùT48�ʛ�Nfnff41@��ΧMZS�,)8��n�Z����~�,�ͣ�{@]�_nS}��6��/��)ا	ħd���
�d;V5�zH&�p���|��a�DF�˪w�Z��~���U�<��"yU��^��o�(8n�Oh9�ϰ2��a�h�A��Ca6��k5�O�X<`>^�.�]<�b�:����7��喢\l��x��~�,1�x���x4�+8�p��ãU�^'�`}�!�F�$��FZT�g���ol3�gxFF��7�zm"O�¨��?5����q�GV�r8y<�P�i�?�`��U��a$���;��pa��Pgʪ:����5��U��ka(�_�H$F��|c�"�H5Y�[�~���ʀ�o�cT��yf�Ӣ���G���+õ��P������L��	6��YMK2��f^�V`r����*�e���X40S\�N���U�-4�x�ܻ���V�nQ�eIiWi;/�?Q�z�,q����?���%;����!�f4�@;%�Z���I��B���pP���ก��^ 5�D�VF	��Z"���Rm�-���g@� `mQ� �JW�=���@����_}�.������K�,���~���U.�LN��.�_YZ2�J�U���ͦ��� 
Q؈'f�4������߃��3&�$�v���7<���_��O__���Y�p��[�β�T��8M(A�x��yX�؀�l|Yl�Y<s�gKE�}��Xh}=mE�V+t�t�q��H?��O��=	Nx?.�n.�0 ��z�}��*m�H#�dZ��l�c��*~��Є�\�?���L�
�@;�׈�7�U�=�Ȍ 0�)���E�wuD��/}�����7��m���/�k/�;k����o�C��H��Cǡ��_r#uI%Sп�yp�I(�h�躭�鄨:CQ��`�n�i�똒�qŠkޚ�4��i��h,�N�R��0 �m�(' ��Mi���S9)�|��\EO����?�]Ƭ�����*�P�-4>XDO��g���ʷ���UF��X�Z9��r�0��Z�9*!\���y�x����v��ό0�B;~�	�-;�w�jA�#�>�
��������P�j�G�1:���qV�R#9�O̢��1'���rt)�H�8�D?�RFq4D�ʋ�W��}a�$�d��]�Y���e��tYO��6Ђ�ծ?�~aP�YZP-���y��
�*0��H���"�DV���#��'���ONu���`1\�1�b���@w��U˫#��}�5����7�����eD�8�x�i��� �n	X��Ip�5؈
BKa�$���\Nn������+/�8w���ga�qڱ�&�����{ğ!��
�"_��b��FT�	�4�v�m!G �Ծ�k�`�#Z�X�8����p*e�m���6I_���li�	�nE
�l�nf��r����V;KHjI6��W�8!�3^d������i�w�8�*-�k���~���w�H�)�*1�j�ʥ��������@��	��	���X�x�n��
ޑvqo���6�
���rK�<L�6��C7��H�
99������FsI�o�UD�;�:<�@�P`�'��*���������	<|��	�c/�_<SYn�Qnyv�~�a�D�&�[Rի׶?ߍ��TN�����!�,�׭U�Â��P��������SK��Ӛ�k��e���K�|���"y����u�������p����3�a���d�NѦs.�\���������Z(!�Liϝ�]�Ǥ\��ݑ)(��IJ�n@��(��?/�]W��C/����ք|�?�%��uV񩊬��Ƥb�W�ͨP��]M�\��v\��1҃t��3[�z���]�f�Q��3�P�a8�{9�� /En�@m��@K���Ϙ��B*$BJ�R<���lLy�&$��X�	�	�"P��"m�C�y(���H�DR�G|Q�0b��*�a�j�E�������*a#1F`]H$g�g����V
���O�L(2�&�=�T�X�F�9
�nUh�������G�|A��1����b�/Cp�ee���khoR8��G M.����N䖱l��Q叧&�S��N���z	�o����Un`��H��������G���KH�^�5!I(�V�Q�n�
a*��G�����}�D�>�e8����[3n�Ȋ��|x��5���Ô�m��ǎx�%HQĮl��>1� ?�Y�%�vq�\�zɜ�����`�����0���q�\#7�ו�����y�Z1�U�W#j���5@��fTI:o�U����|�dlP �"7�>V�����zp�Y����_[{���M9.�1a��P�K��.c��!+S-t��f�GD{��{N�1�ZG#Ʀ87�ʭ,]���,�&b�D6ˤR{)A%S�]d�QF\���O�7I����!TT��j����<9�w��v炙�P 96�svn<���<����v#�/>�#429��x��y�H�w=3�������#3��� �Ƶ���A�'�����Vg�����4�z��i�����S�����乜��^Sd͝�����U���}�	���M7�1��2��|�!��\��)�K`=�������w��*2�6N`��"^egn;%��iG+�`�G����f��֠ə�3d,�����<N�M�çQ���M�!ںw�X'���5�QQ�%�����H��h��b9�X�q=i�HY��-� �= ��_��֑��$D�]�>���w�P������E�p>�K����&�V,����� k�䒂�d�����U�� e���i�[tg�����;��fw���L�e��̇�U���E��E��|ex'5qa�0p�c���8N��
 H�c� ���#���5Xވ���e`tȉUt[*@�/>�XM�n
Sn�6�TY�ƙ��2�D�%W�#��q�`=1�Xj�����.j��q�;�����^�u#˸^>.t6"+�1��.��cQB��_�O�C�����s	L
-����1��e��oҟZ^o��������"�C�:��a���a�����r�r��i�x����{d���]C��v�Ωm�b�o�e�ZCX��-�\0Z&�C�&`
Uv��)�������}�-��R�&:��B�Q���1g�\�S���9�x��O��_���&z���������#V�J���3C�/��1��H��C叅=x����#�41W�4�����a�.�8)��Sk�L��"�-�V}��1�7�H���sʑ�w2@g���jj���zsQ�A;��d�WU��lai�D���xE=6)@n�bT��Ҍ���*ڍ̒��'}w�[�M�z¢6 �2� =ٹ���I��抂����P<6��C<��z|'�V6��L��̏���������HEZc�b�c�������L>;F�M�ܯ��t1̇.p���z�kn��$���m2��:�-��hgZ?�f�ٯb��xrV.�@Bp4�!��`g�ƶ�ҿ�l紳(z/�9!E;�9�� `�d
6����>��T<���<�dx���ƦE7.��=5�>���;jdwy�� �,�R�H�v���t���`����'���`�7�ߧj��C�������퇍��Jv�-
�9�������近��~�ܢ��F
BB�"�1&��Hap�w�,V���� �.���,IY�G	���
�C5�`�����#�2[�ʰq�Cx����Н(F$�v9��y�ƚ#ۻ.Ů��O�2P��yW�J���e�R��
�c/s.e��NGd���u�U�}�x9�h�Msj�j\��h�_�q��r��@�X����P�����]�rӆ�%�t��沖{����Xuo~E�iʹ\��y�����1�:� ��)P�Ij�Q-p�0�z;����9���[�<����d��9���v� �z���-pކ҈��ƫ�s����[=8(4��3�%{��j��p���5q��g6�TU�%�ڡ���6�������2z���J,άn��7��p�\��CW&ޅ����G�zz�D�H�]��D�����1����7��,|�뛛M��W[�yb�C��94N���!eZ���G�?�B0	������ꋜ�a���6����9D��?��A+c�!yi��V�a�$�^y�t�P����H�S0e�3%{N�M����H��<7�m�#?���Z�+UwɀD5\�3�AmO1χ�����E��t��c�^���\�|���b�����P�'U�����:��Ŏ��N��������+Ӈ���{�N�R��9aCH'��*��M+\cxcy�<�3b?��m�e�[��!�l�9���D��K>m�	#\��־.��v�3�F��+�͑P���!���3����v�z
4f�m�Ȑ~E
��{���6�}���{ϫ٘lَ_jUm���D�S�k|%�V蹻���M��ǈ��y���v;�#��;h�%1����:�����꣺�{��W�+�c��-�F�4$�2Θ~7ɝ����fW�FBZ�3Rkeި���{�h2�^��:(`C4A�m���6�%N��v������=�U/�(!���(.�q����ޤP�_&�lܧ��O��D���S��R��l�~��,�}y�4���y �ƴx¦ 4����R�yo�<,�Uen3��fAEuSEb٤�	���ZQ@��nWa⅌�>�$Kw�U�8!vݭ|���5'W����'��&AgUm��ԟ�1}kn��^[�{���egm���g/'�S?��/7��3�m ����>�M���M����^rwM�&�!�O� �d���R'k�Ҍ-Zj���Sڋ-����8��4���5_�f�m���lQ��Cg^�eWG�\��d�E#u@I�C�#�!�C�KL�� �,�$�U�'3{�AXlP�9�v�A�<w!���@�]s4�ظg�`U�����C�$r�
�%d!_I1W�SxeI	1�y��?�I~�Ddt\�X�
A)�)l�"�
�0"�U�5��v�m7p��V�o[�Ԇ�2&�&Hcj�k ai ��쮿G;k���'u�;#���٤�M�� 4�+b��Ti�HBke�
�rXn���K��xh|�`�UC�?��+��e���ܣ�]��/�se�>�) �c����O?+wY}oY-��1�H���A\�u5�u�F�y��w|��CG_)^Z�h�x��Òj����z�v���Y�ܰ?�i�!U�|�<��x�}4$��S��Z�ZY����T4�ܓ"�~������3���:���ڕ�F��+��'74�F8_�hp��燧�'w/2�����_���],|���+���o#�U@��_��xR�LRr�t���$�Y�U��P�֨�7��"'�c!�ɊJ�YiD�KOA��~��0�����jI/���6z�����*���M�K}F}y���i�A�\�g��_��G���jw�i���r�j��i�_�ׯ�g����y�`cQ�?�I-�U&�?|���B��2�g�O\���W���0��h����o?9��%��X ��5�d�+��=p�dU����˃�K@Y�x\�0���樥�[~�e'D�'q����݇��ZC�i, ��~��Ʒ��(�N������'�q�RF7N��V������[�]�r�ټ1�l]B�CV���U�3����UOÓ���[#d��Ƀ����D�N�F�2rw���'��?�����=&%�M���${�G3���_�(�"�w]_���*����h�܄+��!�
��������Ð�}xUD>�-�V�(h�XܪU&�^�9�#���u�控5eS��D�1.����R�P�1/-�I,4�훟��1��8��vELR��	�<�s��K�?2m�y�[�ϭyT�yyۉ�7�z{j�z{�o������m��!���~��%tM��?�1܂��7o��	��qӤ��́Iŋ�^�(+�_H���+����D������Ʒ'E��iߋ��>8K���s��<��|H��ߦg��x�V�ˎ���o� ���g�.�A�=;�����TX*�p��Z6�j��ˋ��ǌ����+�1j���u��O�f .[��R��3�q��������:�-��U��h�T�+ݟ����~��
� ���dg$��ۇ�$��pC���:�he��������`��`��o/(�����Iz���o�6��.�*�����ÒX�;�ƕ�I*�7?H:��]�[���4����1�!}�a�W����_�{]�\Z��HwqWЅyi[��E]�ӓ����i?�ܮ�4_�v�P���������}i���%�������*����J]���>�ݏ9���C��L.����l/����B�9?��0 Y���sq���Au��sF-ؼy�W?;�X	�No��S�0]Ĺ��Z�HXӎW�.����5�k��mI3��G_��z���8WA��OCW[I��TI-p��=UG/�6��0�6����gʬ�V�O��|���mJN�U��*�s)�eγ��<<J��BOsӁ';t�;�N"Ҏ�.�l�d�]K�֫򎗍'�n��ÿ��76ߗ׷������ר��嗞
�Z�V���>_m���kI1�96;��">ނ�=�����|kW�X�ѭ��a�Ty,I�tk�d4��̚� �|b�o	jy��j��_���n��H��sL�B��na��#Q�KU���g���B��xv�����.���fLj���� ���$O��)l�
Ly�����e8�B�����s^ؑ���$G��ܛ�պ,�ʤ���q�� ��J:à�I�%�{�#���0��CK �d��Q�e�-�Z6��F�))�・�R -t�s�1�K�z��wH_�tM��Q���Y� �#�ubi��5�h�'sp����ܧs�ω��5U�3�N@�Oc;㉨Һ	%e������0�`�~К�>�&V�zE���ۉ��H������,V�jFⷺn���D���연��N�0ߺߒuὛ+���>���w	�Il��2JA!'����%�?��|<:p�V9����,�Lt}�LH�5NW���zw���f�-C��1���u����b���b	��P�fvWe�$mʇ8֌�g��
����D��N�2�z~U�̲��Y�۠d@<�
짗�9�6B��JE2J��j�;ɧ)d�:�:{��޻���7DИ��E�_�pBZ}O��ē��=������]T5&U0u8E�n�rq�s�Xt��Z�g�0ZqC��7($A�U��)ϗU�OH��]�=@��k��G ���&�1\��Իǆ&��o�]����Lt<��w�n|���}{X{���m{5�}�y��Y{�{3�b󱼍:���xY%���*�}Z�>�,r��L��IЭ)����1���'������ZÇc�1ܐ$,�4�"�Y�7+f�Kl0R���Z�0L��{����c���OJ	��]͓�+���ץ|��dv�8��ܮa��	�?E�b�c�ܚ��ss��Ӷ���k[�HA��!HXt�a��5�`WnQ�o��G����������]���opH�u8����M��kV����>;�f��.���:�6��ugUU�Q��&R��:H�!�'��>I���{��>����^o*o��ʥ�P@�4ϴ�D�}f�R���o�ɻ��ҽI����z{@�9��n#�jRL�N�֏a�)�gZ����ck�c:�����0	UJ��;�˱��.�7W��y�{1���K]��8ύ~n�o�����	-�?��$&��!�[w��Z3��+���g^�C-"O�Zޮ|��W:��|/'N_f�Zow��#v�<����^�>���sq4��+2��\�Hm�xB��x] A��I���-�*�y�χ���Z�C:#��E�n�	���8�0�Z�����,E�<8.��cf��7�FS��pJ��n��JD�#80�l܂S��p�!��W�Jt��QO��ל!����P(��~4���w�E6��Rce|r���H����!��}w�qٕ[)���ft����pȏ��N+4��P��i=9j���C,�6=R#9/�0�7P��b�f�H�����>T?�D;q����=&��Y8s�S5��6��[+���Hɪ�W(,�%��5}1/��=��1�\��wM@dVb����v�ןE��&�F��� 
��QB���ԘU�Ւi��4d�;����B!���'�|�
O:��}g����b>���D|�F�3Ӗ�O͇0|��a�\f�Yi�R����WC��.N9Ô6�-+��ļ%����29��9)�� 8P��O,tr��a�&Ds�� I��h��0���A�.�~	�{Pǵ�3��j74�.BM rh{u�xUv��scRfR��Ő.�� �.zl���# B�V�չ^����Lq7��HX�9l/�~�ph���p��	�RN5P��/ ����7��A�%f�F�^,D�뎐\nLD"����{|��B��ٹᆤB� 5��T'���]�8^�p��}�MGú=��]���4��F�I5�id�����-����b�������;�lV���ۭ����������|0i*�|�!O��a�#J#~J;{=�px��y��iYj� k�H��șy.�X?,�͟���0��7�{[b�ݞ¯�m�X�e���~S̉U���E���ʭ�0x6,>��d_���9S'�Ol�lא=:O�YJ��b��Z�Ŋ�Ui��s�A����@�4�h��e�e�S�b������,���it����~a�6y��$SS�s*;�m;��*/���X�X_k����z�u�2�}��g��U �F>�l�r��O�:wo]���8~rP�묮��{g�9��y��A͔)g3H�aꀻ��ר�u��Rp���h.+�NVQ�
�ы�9�2�3�
Z��J�7f���*�##�uh1��YX*R,���G-���-����5A�L��q	�do�,�Ź��3Yy�4�O|$@'8�E����n�����J�(��J�� �Cw��]�%�C��]C���p������^k����~��U~l^|�zI�d}�,x���#���e3V:����8F;ݮV%#��F��Y�}T�Q*^E���Mdps�����䡔��C��āiiQ���t�s&q�^�8(��xq� |��z�z|3ܤu�<�����x>y�;�i�(�3|)h�:*=�lN�0�}��~XIN��y��1d�q�� ��s�W��
%��!-b�_��{~d��j�L��Eu �Y+1��$t�b�G_�})Β���/:�3���� ���)+%0��.�K�m���a]��M@�O�	)2&LNض(��ȡ��?Ձ�:�V��Xh����@(-7yH�C%��o�- �w)U^�r�Ek}+u֚A�ṣ?w��l�TY�,5��:��$aɃ�B�0c3��h!j�BzŮ����I/� A��wk��p#*J��L#r�_[ȟ*Y�q�]�>o�!�� �w����!�� pq�$����� �9��j%���^���Ķ�*����:�����~Ԧop0��wY�c�W��qY�Ĥ1|�.J�/�_`X���{�O�b:nB)�cs��œ�&I�Y> �=ײ젎ClȆ�pM�^����.�C�l�|m�Tw.:���/o}</O$h-���_^�\��r�6T��_ZLv��<ڵ	sn�	w�������QvZ��P�q\HZ�([-��Ef�H?��Ԉ҆��o�q�僟_4')��M��S�� A��&��]�| ,��,����׍���,�s���h��#37fc>�K?�+K���D}���y�Z�������J�/`�[��q�u�.�݌��9�]��7`'�C�i�A�"Qz��:�N<�����Ĳ�����1H���h7E�v��#;����r��g$26���_O���� ?����Cs��zZ���O�М������6��1�`)�9�Lq'�+ڽ�����g�#+�6��Ok��˽�~��8'8���/g8��1�O�c3�"�n^��q^\�t_?��G�*}u���0"����4��eA�~� J�ݽt#\�
�"Ud%�m��mS�rH� ~-�����_�<��4q�qkv�cL�5U�G+1j����S���O8�w*�t�؀2��q�y[ځ
�B�REP��D��[��d.��Maj�v�i��i��*CE�2^�]�.آMEp6���X�_��%`�f��Yip�	�" ��Wg $�����������,������o�|�|i�:\ɋ��)��
��hY�ġs1��܌��x���&
�۝�	�v��]L���Uv��Z�Ѷ�,bSH:�ޏp�6C�����(�T2s35�+dZg]�J�㖪��Jh��Jf�	uy_�*��iFu}��Zֲq���f��M�A�|����W��b�	ǰ��m	2o5��"5��ft�%-�����?/<>]�( Q����ܛ���׫�W�v-�����?]|�}y�=:y��z:�J䮗<�?��,�X��ig��ǌZ@-\!��F�6P(C�/�`�PU��-��P$�d �w�$	�Je�?Q� T�y�t�����&b�ȋ�?g5���?'�*{�!�A���>�X�d���{��Ҵj;�C�Ε(b �℡z:��$( ��ia����_�f��TS��\��[�Ch���Ap���F��i�m
X#�2����\)ҲU7�u��}�?7�3��:naǇ7_���5j� ���WL��I��|���n{ �p��`ILc0K���V�tz~8 F��κ�)x��r���3Yb$iu}����F�g��D�K��5Z%9��}�����ui�a4�[�r橥�v���U�R�#qX�9OR�\� �扒8�x�@o|�p1��[+�$�-~?�o�����X��? 6��U��������#-�o2�{�3\ܓ�):���}�zeې����7���+e�f��C�ĺ8����i�=�[��T8z2f�����E_ q	�>^�N��i*8,���@�c�K�X����^��9�������e��j�N�	�ܮ�����{�Z��\�m�� ��>�J��	�SbE�Mo�{��*���v��Ј�,�]9X����
x�X�Դ��������9k����QR_�ԕ�.;O$:h�k}?s|L&���/V���� bI��^ wߍ"0���+�l�k��e,d��jSl�q�a�x!� }���8:���a�{��q0����bCZ�m	��1��l!�����5{5M�L�Z}c�hf�y��^��h0�k�pǂٲ]�����_�bm��9h;vU�P��=�xmV?�	gQeF/��V�q-�jC����C+4KB\r6+5�8���j11�F,8%j^�k��&a���|���mH���	��0Q�!��S���Ї;�b��h��M��p*p���)7��T�2Y����`��p#ڴm��X���7"��c��4 �yD{F��'�<{w�'��Կ�FĹ��U=��Ļzu�0��YcY����<�_��!Z�o�	��N\�`k�c���xah�2S#$ъ4��wAk;ZC��-����J)$�Y�F���2�5��]���ODQ�R����%�2����+�F�Yn(��A���u����d���I]�*��L�^��q���%f��!�_/��MÇ���ygo��<�K껝|��+��>G"X�����M+@a�d���T��q&݆/�f�7���ǎh��O:�N|)oO�(�nP>�'��͔���cB^��7Y��������7�t�L]6�j��f���� ]L�nvm�;S����>֏�]��#C�7�n�H��śx���.[�N��S/=.N<�D����w�pYdXz⼕�]Qc��A�G;��"L5�Sj������*�-M�J1p�}��+j�'��P��v*���=�9����C��W���B����R��]FME.�m��R� ���H*�{�������(؁TVo�V}�����
ߐ��e��P@~\��D�$~��%s���{'�ܽu�WL�yE�?�w�b��O6!�X���DD'�~�KLͼ�׉X�Sa�x��*�` �U8A�B�+����4��Չ5�����>fV��u[�uL�N1�S��y�|��dd�_@���h	��;���z:㞆�$)k��8��ھ{4YmO��5�[`��ī��Ǽ���.̵�+�q��K�𰃠���:�i"��+,u����뺒Vރ�aO���j�<�֥"�V�3'��L�۵�ÚcZ���gj��Et��_����g{��dxl������&-RZO+�SR��)����ۧ���,֜����*�����n=yHo�<��
��.s�%��������L�b�RN������`A(2�$���R5Qл@\��2�����Ѳ�^CE����"=����?�*KV���B�$�T��zE�H��$�O��:s�X�tqq��@�UZ4F�|'�=������>�x�fnF`tZ7��V1��ތ��ˤ��+��(��d�Һ	7��]�"���
����N�A	*ǿ�R��Q�*4k��N?��?��#?ףpd��s�rIA��T��~���((Le�g�����aB�I/VR����K)Cz���v81�w�S�1�뤷��5ٗp� }�?�:=��������N��GsK�U�-�	n�z��0�Yome֒�o��+B����vU���?�'blH�����}*��L�b�{oڅP��7^$rG)��Z�ƫ����1��w撙�PQ��r�S�w7\���QܒO����vJ����5�M�4��j� ��ț���Ns��?�G��8LgI��O�'�;n�~4�d���Z��E]�6��o[���S�9��Z��I�%~���à�a7q�+�P�B����(3�)�������	�A9L�%kkѳ	VJ��!�����׌&�r�Y�G��@7̮w,�w��M�Ww�Y ��-���AQ*��Z*����z���ȣ����Zg���J��*\L�)�����!|�y�rm��2����������g�R�īf��#��DN���z�	K�|������;��s�LT7?D�(Q~���c�}َ�<��'�����v�K�{��3�F���m�l��8g
�A밫�{��B'�kזzH>m]��%Y��uX���=�Yq�R��bx���rXe�9��aE�>i�M}:��S�Lum,�M�K����Bg��ɰ�� oY��������%A�_%�+j������<@��T�6͖�����OT�0W/�}S�N�!�D��.<���]Kǂ�� +�'�3[-3r�$�;)�����Y�8ݯ�Y�������m�F��պb��y�OYU���*˩�C%���.�S��I���6W��>T}�p;�a���-�D��AY8$\u^-� �9/�- !�n�**i{�3��� �ՄS��xd�FL,���IM����8�&��gHÆkjk{߷��h��b���"���6:���nH#����"Kꠦ؎&_�</�Dv�WW5�?����v���j���Q�G��c64����h?}�̋�,��6�uˀHBq����2Ov�6ߵN�C�+��R��R�A�dpՎ�(��j����Wp�.!��m;'�i���U�bB9��,e���DT��;�C�S�x�' +�w�ޗ��~����JFd�Fdm����q���p�>�r�f;�R\�؇�&������<�U����a�f�?H��P�_�q,bw;��"l�g�D0�f�=J�>&�>L�c[���� Q^�wd96dA��� �����;��D�JCJu�bc�A�\��jE'������~���LX5�YATCI�O5��:��ϼ�*��j#�`�s���O>cG���OQ W�������^�����h#ס%���r�?��ˏԣ�1藲���_[�Р�~e¯ĔS"7������]|���ȷ�A�Hr�7U	fB���J�ZF��aZq%�͎�0�e���8H����
���=v��}]@�� �D�\�|�ġ7����@�	�{7���+]�z JƖ�.��p�s��Iok��t��ݨ���G匪��Zy*���VKv�R��^�ك<�\�bu:�ح*^��%�	�0���Q�{�r����*�����
��5XI͒U��)�_�)�t���+��8sIGw%�j�͋:k �eǿ�����E�e�0�����ޟ' 2(�����YI���CDa�.���s��%��ˁ���&KE��7]��d���7SWK�Mܴ��;+�o𮲏k�z�Gg���J{mv���O�ct#F8�7�ܔZy��w�?_k~�m��}|6�=�m��l}��<�=~����o�~	��*nu(q�ר�B/�}j�����؎�VOd"�*88͙�A�C�d�
�gÑ=f!�ڤ)ǧ�X���?�6��γM}�6#fyM��>��)bs&�j�w��x	@$�4��V�CH�nPp���oS�F�Y"�4ךl��A��cNޢU'7V:�ی09�Y;ߧ�*�&��#�򇂆������ʸ���C��r�8�yN�K�J�}������{z�!� ^�b^ui��`��>�b���OQ�66�}����LD��7�K����+`�����v�N�K�ubk���M�W|Z�6�����b}?���j˼��"A���fBk,���Wܹ�)�[m䕷S�ړq
���'s�㪐�5f��@�|�1���<v�D�h���/bP	��*glRI�q��$g��6a����ъ�ATI�u"j#[�IUkot��G��v����;�Uܚ������N��V����l�������6]z���u,��Hݢ��G��X�Mn�V�pk���P��^��u�P��ӄ�3�l��l��gj�.%i_�[
2��S�v�n�_���^W� c�9�A���ou�����4s`���~���=��X�l������3�.3��WDdӬ���n:e���g�}W��ɀ��*fb�����h^���ͤ�ϐ����[D��L�Z�̊/�O�?�^�y)�?�sHP������>4}��G{v7!�O�#ts�����r)��pU(�ɘ����-��˃���#�8�0�F�Y}/�%Q��R��5�SI����ַ�����X�+[2/����a�u�G� G���4�Ec����\�P9�)�&u�__�UJ[����/()�ʟ[�ݤ��,�pN��dܠ0�K@���{~u�h�����0|��KWy�pР]�����hisag?�mHb�j���S���f�Q�"�v����v�ҿ[�k��g��7@�g����(R�wqŧ|ۍ|�AH�N��}',fu�,�}iЈ}��s�Y�<�Xt
�Er�9+�[P��5_�Y�p�;�$U��L�� �s��e��m5��ߎ�E������#ȑ:�0�$����!o��Z��3K��13��`;9X҅��7�M�2�"�W�U���'�-
�.�@�5&]%��o���*�M��w6��	��B(�F���Ԣ].�}�J\�E�[�8��t�/��b��k�[��.˺Qd�z��ߕ=Ʋ��0�Z�ԉ7p�\��@�l��a�Q]H���Rd�r(��Xx��z�����{����C�NFC|*�-J?kO9��% ��I��������K�|c��rJ��egD}\G�@���:�����*��W�Y���
X��99b���t���N��'k-?�[3{��P�˾������P5�~��Rž�z1�)��hL���ku-�� �z{->�k�i��+���&��T�G��Y������� ��Þ���|��sq̿��V����a�O�'��Ӻ�%WM����)RX�L��*�fU� �#��o���,��	���C��ӓU@KFHO��Ezl�������Me�3u�e��c���m��ҋ �u\�M�j�|�B�2�n\�z�[?=C'��ѯ�����ds�Y��Z�B�$��g��������6�"v������~歷I�	Ͻ|Y�Mj���k��;�u喷��$��'(F2�ʩb��r2qj	kl����Q�+�3�A�T�u�8�q�g�!�ˇh�����lL�C��~��XO7�_�*n�h�-��4�R�P������[#�*1z��w7$��4�	��w#�/e�?H��1��^Xɻ��%�??�s���=\�� �-��˳"Z�s��Z�6]PGL^�?�*/ۅ8��u�,���d��j��MWб�K��W��iݕ�q����.�K��.�z���,rթU,�8����E5IS�0m��|�9��0(��.��n�NE1����,T��H��Ux��9����Z��*�	�ވB& �<�bs�,H���Y��<���8ɯX�R\!ҵ���ӻ ��v(�Ю�	/�C���0�J���iߟ>� ��Qlʢ> �X���_�W�؁�pb�`?!�Â:?��Z�D�S܈*�pW#�h/-�f��IVUQ�q�_�Gl8�÷�N�i�|�*1�64�$AAM%jˀ��C�]�6^/����pT���k5p�iI��Hb̀����̜�{�k*��J)/j��=�vw����!.�_���y-�_#�[<v�#8Z���/�"�T��;;�zx� h������e��/Z�Z�)Z��_K���q�� �%.���SEA����TƦ�='�s؊�[Ć_������^��/$sM>�f.\�#� Ȼ�e��c�<�D�X�p�Ќu4��Ջ��U<]�L�Q�Ӵ�Mpq��^c�Ӳ��+��R�$��=Bى���\2��N3팞ߖ~�ǹ�CkMCΌ��~�·hc�r��rw�Yoh�o��JÃgPaO*�ƴ�r-�ӕ}�d{�9`������J̼�G���G�:��\jS����Fnܽ�[5�Y�vv���`c<�Y��^����%yl��
+�_L���v�rE�	!J�{(xԃѕ3ٛB3�|��ƑZ�B�E�ћ��X{ci�Q*��2d,b��؟��:I�n�~��O�|i��nYx�bU�@����ۼN�*ވsy� p�H,��f���t�_4RShv��@A����pj�'N��g�ڢ���xv�H(f,�W����2y|ʴہ�ʡ�c)�uW�f�"�Z�!���(�3��ipYA�� ��M������Q���:�M��q�ƃ|�|����U��]�R�O!�z�T��q�a?��'O��{"����*�UZ�O�x����fDl`� ��L#~)#����.l�o��RUE���6ɉK��4�|o�>��:���p�=�n��_�sC�G=�i�~ O��Δo��9ru�&�FtZ�jRGܫ{-*��4������P��0�ykS�w�kM�*��q�$�Ϙ:ƜE(�1�z�~-�&�kVw��{ȶU{Q9ߴ��WÔ���*�����Gm:n��ܶ`8�Mť��}P����VN�U��j
߃�~ ��R6g��F��ذ�RZɌ^j��Ga�O�+�m��w<�89�~�����X�L�o^���Z�3i�3�ٽ;�Li���T�[����i�ͷ���c���f�����EMbI�k6@V��/Jߗ�-g��T��?jR��
ݯZ
�wz�<q��]����k�+�4.\����k���ʽ.��Ig&�F�nF���-�^���^AyXp��S�x�ݧ�S�����Jhj��`��HH�+�m��U+��A��X�
X�N���L�B"��_�ǅ�֍j	=�Q:�Պsl�OA�X>�T
���k���l[ ��Y��Zꏌ��H�j<�8=���;(O=������&!z��� 0��έ�;N����FJGX ����Po�Dy�t����S��l�OG�Eh�C$��?�"&�--�;"���qxvI�>�v7���U[��_b�5�/bGRJ��'E��!��؊�ƯD:��v�Y��ђ�B��'Q0���q��rQ�bw� ��V���$p�ċ�1q�Bv�Dr����M�S!�Kc�݀U��q/���� \ �-��d�̣!톡���9�I�kp�ՌW"i䎚s��^{�`2d�&E�9KB�2>�j�V=v�L�j��{�H�����.ƛ%��n�I��⟟r��d�*H���Z����Ն| S�Ė���o��(Vd*	��`���w��?���7hѼͼ���<�$�[S�]v#��<
N����Rp�'c���H�ܖq�Y"'��t)B3�"��B��+�$C&W�ICqL�t:������(~/u��;��zq��w��_�[.y1\Q���A�c"�Y	�fa,�Hy&�4��M��4v����	����Ҝ�j�@G��Ù�m��x�?i�]��70�������XM�:�w�z�`z7 5�#zOxVv���xˉ'P���̊%�
a���8�q�s6�ӆ�� ���5J19����z
�l?�0�cr�����@�ӧ�ǋ�7����5lw�e���m���eZG��t�I�UHSZ�l�����I���BM��`�L�кa��Oe�s^d[���
��s�$sm�v�f̛����Jp�5�J5��f�ɋ[��i�&.S���jm�:y��M�j9^+&[m�&@EFA^;Ky��_H��+bWKEA&CW㄀�)T���G�'6����$�����5�����~_K��6�zW�#5�ٮ���l�ruS�E�	>���' :Fy��Br�b�!۠�#����	��D�
����w��_�0}�'��B[��j��c�-2�\����M�D�6A�>!v�����͌g`&ᴏ����o]Èj��N����_$~� �Ώ],���
Ud�$U���G�n8�����Su�U㝠2��<T���D���,c*|��i��18�= ��9��p����k�+���r���r�8U��Х�wf1�|y��K
���� �٦;� �xZ�f!��w���l�(�Vɢ'V�f#@�-՗[5�E���wF��6c4Mz$9�a����T:�JB��;R ��yݱpv�{�ם�i�6�T[Y�{�[���G��GW�r����VU�����&�l�2;%�!�#bKS��b;��A��|���x��e"��j$�WVūt;pF��m2Kڡ4��6?SdF]dpcnN"����@U������u-�;�����O���d�^�a��.�ԉ~Fs����}�)��>����a����a7�Ӵ��U���A��-+e�M�˥���}����ܢ��މ�M�#)�CY}K%"�J	 ɡ��292�i��i��tp��PO���Go��`$t�7x�x9�v?��?�7�X�M���̗�W�甇�6]���=��zž�1�����LzF#��`�h8[/5y�EA��護�'r�J�]�j��#U��B0�®ͪ���8B|��C��1�0��]�>b_l(���1ԻJC�+��v�&l�� �n,;�)�KQ0�]B5D�4�A3�n�|Xa�֐8���'Bq����F��8��TF��6vo3RV��S�=�����D�K͙	P����)!�F�f��P����Id�;�ihZ��������;�W�a5i=�י(Q#�ϖ�ȉ��`��j-�����%u�[�/ۊ*��|�!�c�.���1�xq�[ޞ.���������q]i'fO��TAt�	��6F��.{H8.���=�n@v�=�n-(yp�s�H��;��� ��lZ�<,e��MD���ࣅW���t�sZK.҉_�T�]��`���khɟ���̉��Ѓ�Ɍv�۾���B�j#�^�Z?��Y�.�_gr,;6�Ո}3�!+��(ɸ��8�qf�Be�;����;�B'���$�big&�w�W��n��$s
��N�{.%W�76�o\��.��dh#�}���<�A��8��d���1J_I�5��nƻG���7��'Xc�w�#P������`�]R(
�x3�R�v�|��.��)�,����ڑ��0���t�����:�/dc;��e�6�o&|�X��4�˾����X>ܒ?�r��l�kǜJW���+K]�Y��9��cng5[��G:� ��+�]#fRߺ#ѝ���+��������>O�3��s0B=kx�%�"u+�����!��!ƀ�m�Tp��T����Q���]�L���wbA���|E;>C�>��\�0�6��8Z��0Db�mqJ�?.����W��,�R�w���l�-������p7��A����,��FS�����t1ۋ(�?}؞�:��)���y��X�]ۼ}CE���D���dDյ*D8���C�I��M��c���\���}��j
�\1�*�b~F ��q���uZ�0gY�(�p`��sj��r���,�#co�L%Y��3jn���N���,�n���ݜ�ۀ����T�k�v��\�óft:��U^%Rz���(��v�s�L����[א$�$G����օ��a�$@D����#e�6��d;�I `-/Q�������|��	��b�;����{�g�(���Nwє��f�p͞��ܗ/9�|3s5�;T���K7�OΆ�0$RSR��k��n`��� X��ɏ�/T��&W���*+^�]�U٪�0lc׬�Ҭ�2l��1ٗE�k�OVS��8지l��'��g��_�ϔ�Ƅ<X_��۞O�)��]\6'j�XK�~�5�F�ps��A�a�ޫ� �L��Cf��y�d������o�X�|��^�M:I�SJ^�)�Nc�t@א 3HCT������ʘ3�O��ڬP�LƮ�b�|R--�I��4JRP0/j�֎���(:E���s��`P��ʳ$e'Ľy?(a�<�^�!_�l�TV�;�By~��()��Q�ba��Ea.��PCX'?�D]iv����$�Hȶ�g��I��g��Y%�<5�9�xW��$��c�����Eԑ������sJ[ݻ��������z���������<�rH0H���۬�����WP�η�wථ�u�K��������p+<�����*�} W#u����+wƞK[ޢz�l
C t�Î�[��̦r~�Q��˨�]YNf�N�q����Lr����U��b,;���|KO{d�đ��d��S�}NB�D��%�9��d`M�k��m�-��a��
U/�pF�LڂuN��{��l(������
��_\H��T��є�2��}d:#���i�����F������o�7��;�0c��N����nK��'q�h6��s��������[����5 ��j��}m��i�XÒ�N`@Δ��"6��.�h�W�?/ �Ѕ���t�K��u{��L���A�Uf�'���d^@W����MP}�c}���h����(����-���w<>͖K������Ӂ8�g����I��X>˛�Ik��
����&rB��d}�5��z�ڴ}�5���:^���M��s�C��,��7�v��-\��^��b�$뮖!�S��F[�����9��6��� ;o��/�b�ѝ�?L��3�#,�)�N-	��X��� qÂ#���`�7o��VY���ў\}�P:P ��G�>%p_3_^�)��9C
G�S�ư4[�!f�����nE�0h�}0��� X�~�x|bU��+�M��%}��O���z���ऌ@)�@u�%L���N���h���A���N�]���K���22:�Wr�$MĚc6�"}�/,T�HD��(�|}�s'}�y=*��(�M6Wqj<�e�2�v���G NV�Э�)� ?���@4��w���Ȑa:(��|!XV���CN��=G'�\��<�˙BN��Ȗ&�U+�?�/{M4>7��=yx �d�xjs��)��o]�����z�3tN%2o��&*�4�/ gC�4u�,�o���u+b.�����]�`�@�C�R1���n���'Y�#T��)͸N���	���q�#n(�:V�
�ѷ�z8�>������$��A0��I(�(�}�ۄ�6g=�o�<�����<���7Wq{Y"%�.7<����|�5���ii0+E)�&��(��mz�
 fi���b��5Ezv9������\z�=�||��" >9�f�%�ʩ��v	:�g��t{����t`~�0}�ff8�\4��Yrro�~���Á͐M1�����9��� ��_��W^&�x�r ��O�`�8�*��"�u���J�:Hq�=Y�T�ő�4�  Ak���])8[������A2�m[$ɧO��~���]�V5J�w�BG��G:�6�ʮ�A�,c�
w�e�:�w�u�wʹ	Il��)�e��!�+a1�c��D�CqV	��ʫA�� �2�ЌȾ׭6��a=����a�����YyN��\*_����j�Q:Žf��h�3���yp�<h2���]XvF-)ܦ��p������A�#���8�HG����hְ�Y�Z�iuEBЩM�]wA���=ǖ>�4i����K�?�fH	�ڋ�?�mi��'9����Zh�;�ƬI�#ֿ�W9 "ph4�q3��Թ�!��p��M���j�d�C�L��p n�����L�OR�Q;�=ӴvG
f詗���� �h�+ns	��ޭ�67�/��J�ѤDO��.�7���uX	��0u�csD���+h�]+�� �^��OqΜ�h7\aJ[����Q蠂zw��B& �y:�#i���#u�J4�6
4F�)�>�3W�A#��&>9Z29Z�H)p	7�Eb_z&@���n^QkH����d]|�G<ҍ�ډ���q�r��E���f���q�@M��#GB�M�'͇�>˚M��v��G6��W��n��Z��Y����b�ߠ$
���{I �Wf����uѹ&���}7�+~�s�2~�߁|b��mf�yV�}4��Tt=-VE�m�S�0�X�i�i>��ԳIF�x+�U`�wKӭ�H���?��=3�-���^9[�d#<{���6�ڤhY+�f����z��� ��D�6��![����B�;�X�-)[L{�TI�f��#��<��&�V��cg���àL[	 w"����^�T?^�w��|��Z2d�#,��h+�p.?����|�A���љ�<l?��n���$�~�Z��.&��7�������5�	J�Y�Lї����4e'R���I��2���*���C8�c0�d͒#I�{7r�ë#F�(�c�42�6��;X�m<͹���e:�+��M�Gշ3L꒗�x��5F�]�0~�7��K7��o��W���-/�s����1���tBC�?�p]���",U�}���9%v�ռ��)���$SE�}�v�7�1���v�����	(q��yn�����F7�KL���L}��1�^��q�����n�9��N(`=�]�w��ү8q&O�e9)bG-CE��l����%��Jy������Ύ`{�Ŧ{3��C;�ěA����Y��W�mO��c�r�$�`����$1�U�Z)Ϩi�}�Zq�`<��ڼ��`�/�(�%�P�1�s$��~���c�
�KN���6&'F��"W�H!�)4د}BU�<��(���Tm�<����L��h��%闱/6�u6�؈�������w�,Q��=�}k(�[�6�rO���񃕢�.:�	Pb>�3Fm��t�#�,A��h�bl�Ik8a�?���@3>6����sW��󣷞�lG�RL���A&�Z�Y�9@���UZi��L��'|3U�l�в���$S�9��:�b<�����Ȩ@hΛ�س4���oy�@�R�	ׅV��
KqI@�Ի���Y,���:�(#����xѿ&9uj�K�u�"�mG`�w�!�c�-�.w��2GI���$��a�>�er�o�s4�lx��ix�Eh��i���N�b	:7��a&�PB��q��5�����aҡ�<�$0���<b�����Zs���l(o^INɪs�y{:�*����}�С�[�� ^x� �ǜ����*��F�����Wn���������8�-y}�1U�ׅ�\b����C������a��~(�c���)i<T�_�%��d�����. �Ы�ֈs�����"��s��|�\p �?�.�鳲���6�ĳbr���Q�іa�3��D;|�P!x	|���3�׫w�xE�F������W/�N/�I>ҫ�9k�q���n4 +���z* �ϱ�/ouF�39����
�����gj]���Ǩ��*K L=���=���3&w���Z�TC�͙
jw��R�}s�mP!z��8�#�˼��̻3�Kb�C,���#��"���|I���3�Ū�@��x��BSV�V�̜��$5�� ��A�\�g�b�@D}[FV�ʭ"#�&���m��L�J�)��	����v�� c�7n��]��3�p_��<]��Li|ܾ fq˝}���I��5Lg�_a�o�m�.�ęz�V���"sJ[9�Č2���۲'cx��ǖ'���zu��xJq�'l��թ��
�d"��*�)�܅��~:���I/ f���W���b��!�LC�"�0'&>壢v�PDFB$i��YR�!	.�CBB�Ҫ�<'�r��j+E#I'Y�&���Զ��O�n��ն��LjR�K�L�o��h^y�o���G�~�?����t}�|z���lJ~�Wz^�Z�s�P�h�Wt��5��W�ԫgn��>7y�c�[;C,��~�@h����[�v1��R%���3<��R�.���+Bf S��++�D|gp�RR�j����k�g�2k�4.�R�m��n?%�#�u�+u.�T�N;󺲢50S1�dM�.%�O�ғ	�q�+~>o
�!U�Y�
O�<�Ƀ��ڪ��G�:�B�����]u���]X�6n���h^�p)Y���ư�>&LV��V�J37�u�t��4��NI��7н��dП/�u�&�[U^��F���lĚ���L]��2x��(�x@�����u�'�e���MOG_���է>�u�y�i�ع�B T�{��d��*��
:����i0��i.�Z�Y{�B_{]j:��Wi�
�u��SW��>W�Ќ/d±�|^b��-��%����߁�
 �Bn���>_�b[�v p��o��	�g����{\Z�.��lh��(��/FE�|F+���w��G�.d|��n��c���1��´h����a_�"��B�HQ�D�,��a��W�
��?d=,����R��!b�����F�Vl֜e���$h�����}���,���b ��Pz���m���z{W�vH]ea�dL�e=�i3�E̮X�_b-@[���?L}eP�]-Eŵ��.���Kpw	��^�^ ���58(��-����ܹ3'?2���ɳ�Z[�6��z��t���>L�����w����J\��2�����nw�& �G^� 0䛻o����gQ�J�*+�J��+���ڜVZa�zv5�m�9wY����
嘴�Xś�~Fn5�srMs���(�_*��'%i��[����nI���w�ŎEc�E�M�o������p¦r��u�掞���2����(�]��qָ�A9�%|Q��i�ґ7�bH����ә���i��^r�6�g}�?���?���=��dZ�i�6>I������#eˋ>g��j'�Sm�\8Z]���;�KQ�
����B�7<�[R9��`�'<�?Zy(fE����� ��T:0�wi�C���|�#��
��b#E�.|�vŜ�u&sn��8�����c!���80��*���0�&΃e��wFD"����(���,wv��P�(3,��,��oðy���h+\/���K.�H����ܞ$w�
��/��rΆ�'i��V�ġl�' <İ@��z'�K޼*8b ����CI�&�^}|�ȸc[d#�5mc�OY��Jah9e[,I�޳h��|O�R������v��]S#njߙw��q��������%�̉�!,i�SA�7ҧ;�K�9�841���0�d����Maâf5Н�]4��r�ڄ�>���B{��-'����{js�����@�^�����^�y���Q��W��~%��r�<t��Ix��Kn���ӳ��Ii`�4�!�	�����[EC���?�C�wak���e�����xT��� ͡9f���Tc �N�r90\ƈIPb�������o)[��o����m��q�A8��
���	8�b!����Z����U�W�20?o�I�,[��.Z�K%\yo0/�o�q�LZ+�:gY�h�uB�O�h�ˮy
�SC�i�Z�K����Wɥ������r�o��ɀO˛�)��#��
(��l{�'��$����ok�'l����pOg���H��_s)�f{�	��0C���t�$#mp��4g�k�#&���1����� �f+����qH�e:Uu��1��$��t�+��4/�Y��$P9��M��CU���ƧZ�_y��߇��YH����2u�w���Vf�E�OF
�j���X�/=��;1�9�G�8>%C���@x1�f=�`ș!sZ��ۼ�&h�R���|�d,�B`�k��=nRLm<�P�������#n��B5����р��Xx=@�uA�����ϼџ���v8���-i��f��įm�B�+�k%�B�𽗫�!�f�� w��=-�D*�u�A%t�fAp��Z\�NJs�l���c�K)>�t}^��a�7���7����C����ԍ?���n-���f,l��[�"m��Iz�;
i���	ɔ�͟����x��!@XA9~E��	�JbG�8>_:=8��c
��3�O-R�w/�1�8����/�+�����G���g膧X����
��(�i>41?g@zZ�oU�|�����h��t��rT���(�0��r��������j�����tC�JSri��;ʇ�|�He'��h�y��z�����O������ۉ�F�8���JtY��V�#^3�9{�ʅ�,L�C�v;p$y�,O̅�`�ܟR����G·�����1��~����&�Y�c��Q��s��p�ڈ�/=��JȞ���f`Y���{ǀ�[&8�Q�P�mbw�>+h�z��J/�_abn�" !��&�a	'�N}>��@3�
	v��I�Ǽ{��{:E�̥ &o����9�t{Ѳ>3W�	M� E��
U��~�8;$ p��hL8D��`W�M�Dߧa��� ��ш�	0�E�)�ǚX���/^v�;f�. Z�7>#YC��	��9.X��a�%���)4b�]�O��$�hT
H�2����Ƥ&��� ���#�=b�{��y��Ŋ��-���[�����(�=8`R`��e�t`�{�o�i�y������G�oU����U��OT������|�b�����}��O��תX���|�}7��_���������O�^Z���˳��Eݮ��J���J6���#�.���[�EF���������]k�"�.}��jx-Mߛ��Q�rTO�@ӽ*?�7;ޞ1eE�؃,�W�(���������9�l��=��l�jE	�A�>~���V|%H���C�l�wL]�_���c0��؂��	w�5�nƻl�����;�q^.wh��2�CcY��]�@�����t�n~�@c���MG0'
E*�iȢnu���=�1��*	�>�5r�J�5zAyp]�X^d5��&-�WPn-�� ~��=Zn@!۴TZP�MS��;�1�,�"uԤp>�y������W��<�[���1D|S�'r"����9ȵ!Cw%s�����'�v�m�,���m��ʍ�x���%)����y���$}8��n��7��� D��^�k	����j�!IE~�����Q=zjJ�S�G��s���{��~87���+t.o��o�\�c}���\�a�K��&3��j�s2^���,��i����,MХM�8k�r��c�R�Y��彈��VoL*4��8�;	��k$ތ��M,�,PK����h�����{%�L�(�6
1[��~l�>[�3�%�Aږ�L���p���E�c瀙�s��[�������q�vT4e�h�N>����{���n��୘�z���q���C��6i6��`>��V@أn�f�3d����r���0������k����QYU��x�lF
o]�N��8r��c_�i�^"��ڊ��(����@�4 ܶC=����~N�l�8�*�t�6-<=��-mj�[ɶ�1����C Gi~�r�xN�qo���h-=f~�R��B����^�O���d�	"�v�-�7UrH."+�Y�/R�ws�3lz���3S��]�+*��,�-"�:�uz��O��gr�EU�(�4 ���+�xqCf���.����_�������W�.�(�f�/���7��
��ώ	ag��b�0?k>�	�Y�e�+=[��ͧ��7�1���{�ٻ8�m�l�!��"���	�!m�o9Wh�t���zW���<4Wd2sWl��.~����k���08|cD��(�Ҁ�Ԧ�,���Jwa�2�_c�9x�։��5�/f��[���\��vV�R����b�+���P�k�eɩ���6+���΍�:����@��}�me��X_/1!�q��᥀/�֞��K���k��hF�_⛞�?���ychx���ה�K#Q��!�W
f�ŕY,��ʧ��j%!!E>Q<�A�
���F�tZ��U	'"tv����ۤ�V��J�`�؇�d�ML������̨�e>a�i=���_Or<��c��Q�$�U�dy�9���+&楒n(�EG�˙�2gW,�|���;�E�)u����çDc���|h�U
:by*e:N)��؛~����}���q�M������֮�'3x�<�E������4���O��/t(p�؏.��"GLg�4��1u��\}�;�!�~o�!_��GT�>�8Ņ��S�I�8�
�( J!�+�²h*~���Uc@��FY4\�q󕫘�Z�t A�X]�PN�׌(�JN��3r:�o�i@2Z�)M�H�M;�3y�n�������{G'�Γ��������E[ݣ�화�Nɸe�]y���S�3]�'G'V&� qu��V��$��^V~�����Nm�jf�}3#M�חm/���N����]~��3p���!�?�;���������D�)�mBec{��S�1h��X����)YAzP(t���]!N3�a���)�������<�k��$pթw	��]�Og��׉�%��>���kl��i����19aݪ�5�I�����ږ�Jhec>�����Z�*���ǳ�0���e1�=��/E�0t����A0T:f��ܥH=�nv�ܡ'��^�*�� ȶծ;`��n����ʉ`tXU������6����	!+�����M���G�����i�q�/Es|�yVɻ����%��~Qk�JP\3s��3FD�?�ـgp��{�6I�O�>���`�r����o�T!3�oT��^�!(b}��˙[������c��!`��g��+ĭ���k�MXrI-�4��ݷd�'p�F"�}U�Q*�#:6!���o񳭵��K��4/��d7�~lm�����Tޏp��͜�Ƀ������U�ȥ�UM��{b�fUUG�͆��S�C�-�q
��1虨��4E�n^�߲�� �>��~�{D��{�������k�]Bw0�LQ2�Jx;�Ȗ;G괪(�]��u�(`۵����5�\�Vux\�S��q&N��l2f���\Pͮg 㹁=��eq�l  ���{� ��g-[�ZgM�}�W�i�<�xf�X�{!�G�1�7�hz�<�
 � �+F���i�N��&�Ah!�Q���a�*6�׈�F�@cpƁ���<TP�PD&��CU��T݈�6�l��5�q�G�à�b�~(W���^�bq�[.!(�d�h���]�!r�&��.�ȟ�"p�o�k���)i�{�'�6�����i�����_I��l�7����p(p�������6(��j�d�Duo�08��E��[�枲�6�첪�X#R���?G�}kx&���$��I��}��kz8n��-��up���":E�ZL��({��rK8�CO���>�%��]�}�X�ߊ;d��wl���W�
Xo�./�f+���,���8�|�=�D��I�=Պ֊@�j��K�5�����8�
>Zkު�ɕh����TN���KN����t�����U*h�J�ۨĿ��2�x�cbO�JLa��M��$����1Q��q�A3��$�U�S!BAH�%�wc)�]� @��ߪ,�#a�7h��tzR�w��<��*6㧦�y
A�x�D�&5UpR�������(lcu`����X�f�����ǃa�Yp����������x\5C7Lk�ᛀ�O�gGn�vBߥݸf��1l�*]ę�O	ߔ��-�WI��F�k��v�4�P���ЈLQ���$��-��l{'郀_N�k��@�;���{Ju�� �����߀��h�z^��yAz�!qj5
lZ��_h�1�뛌p��7k��b����]#&�>֒ad�S���+ڂ�-� �֢(N<)�*b���X��6��sζg�ёe18�SbKڝM5! L�:*�t���й�q��}�g��N��g����ߴ܀�3Ͽ۫��U/�̫��L�c7�W/@cd�`1�Wj$��sv�t����.�1���аr��Y�J+ꁖ^^��Q�IkXWŽx0���{ikW͂�:��J��хAH����-��ϵYu����ԅF���g#�j��*�S^�$m(I�`�\�����5��.�Ǆ�ޫ�DR1i�-�Y:XeS���
��#���a��M[`����CS��tF�U�n*�'o�e�<���OBK��t�E��0����R�(�0<�Ы)��-|�Ь�t�<O�Np�'{�t�4"�|kI��'zǵaQ��i���7TY�|��>��q�ԡ ����1�]<]>�u���zX�@�yUq���G3�1hV�S�T��[�x��f�EOz3�������yf�ST���sC�̛��X��x"�;�MXpۦ�2�'f�I�V?~��]j�}������ ���M��wtgY��1h)p��3���-L����Y����n
�ӥH��t��9��/:�o�5k��4��r/����W�	U*�V�jZ��y�_��*�;�C�Թz�b;E��S��V�ʿ�*H}�"D�d���J�QZQ����4��Q{FEG�Ǧ$`���Nݚ��͢h�ȁ/��g��'���"4��qja2H5.�
�sPT��;��7=�S�m�ZMʬK$��:=|���IXpOe�g�FkQ�a���y�k��~������΢�[7��׮���p.߳}˕^�wa��)��\��G�o�>'�fWa'W�ړ�
�P�f�I�G��(]\�ƨ0Z�KY�}���6#W��L��a2X���e��'k�/�.Íp	�~#����"�nr���D��ض�a��xU�xXT���΁�,�Kd�9c�xu���1kŸ���e��L,._兿����ɰ�R^"��+	M5�LՋ�b��yX!�YD}�75����B*���4�8�z�� �DX�
��K�u��|*W߻�v>j|�P���3�g��ǌؚ��3�/�H�ň�.Ng.>�Z�B��Z�'�#%���@�ԧ����f��ʰ8y�K���$��BQ��)����/6m'�Mm~�ت�!sɶx#ʅFs;�����\��غ����W����qE����V@m2�)�+U�<;ю�{��N����Xe:��"��EyP�j�ɛj*a*i B'{�w��D��Q�l'3X'iЅ}�ĂV�C4�[��T�a�C��.ײ=]��N� ��f�P�O�&4�_k��;e�}Zrr�k���K�n��0��$v��E v��"���qܧX�"˴�P]����H�F�� 3�N�\�=_����B����A�&+�K�%��R����Y@ȁ�ǷL�6<�r�
eɌ��o�GG���G��jS��}^i>��0�<�9d�f7����c��U���4�x�t�y=���w�m��u�qfu��r��U��������/1U��Ƕ���;ٻ�M���?�t2IM��rq���������l$��L�V4������o1��:S�f�ﯸ�Vͯ$�rIN��.S�4,��ȱ�J̗���������9�ͯH����������������}f��������L�J.��6Eu����4f�D��`����ȕX�¼NW6d�  �vU��8�.C���&�; J �\[�I^(������C�i�"�|���D��:8�ٰ�� �>��7l�/������k9�L(�{�:����=��0�%Q������2����L�^f~���"Q�������z5,b�c�G�X*M��83b��Ś�������E��AŦw�X"u�U��n2k�k���|�ct��g|#��_0"��d��=�KdA�d<ZM�[�������(�#�)̿ט�c<��������CY�h�!���ӂ��B�W�E:SG��&�8��D/�"�K$��"Mɯ�m�0\���C0B�/Bb�j�W��}���nY�>�ū�,0�,�[��(����t~zr(G��^~���HĴ2V_�F܆�w�{b��P:i��������2	ꑭf�m>����Sz��l���Y4�=�~�y��w�rUV�H�6b����k����I�`!T��H��Sq�*X��Y��;W��s蜅?ف�_������S��{�nN�9�b���L���f �z��J#$��

�����m"G��NZ������i|�BN�X}���N��y�#r.�G_I��M��@_���K૔ -i��abۂ=8�^F,TW8A<0�W����盘�7B�&�����Q���ӑ����չ帚�~��b�S��	�-S#&��T� r��K#�v ��
tØ�rShؐ��br�����a�~�Eh�p!K�VG��v�a���4w�>��JPmLd��?E���)A�"���h!�롩�T?�$�0e�zwy�<-�4�J�Ei������@��9U7[޾��rn�q���"������	`�s<�C"�m��Q!��RD��S2κ�e��'��8�D�Tb�|2t>�?j��	��\�/FAPҾ���w�S�4�#���c��06oN�ݛ"�t�r�/xD��(&��G���^7�/�$�O1�diW�l�w-�l��?So�����#����.Q��<�o���U����s���hm9��?
&�����l�� �"�|��C��{��%&TЂ���R��N8�}��Ve���e<p�Y_�i�f՞0a���W��8م���@�9�I�3��e�w%S�`���K�	ʈ��D\�[�W=G�.D��7?Df��-J��q�V��d�L��Q��`Z%��.��Mۗ�|,;6e���P�	�~)<\�W���[/28, At��[��]y�f�%?���Q/W^ww��)�Q6��F�bb�2o�k��H�%"�K/��侂�̹�q�}ן�������6ש^N���6u���w>�x��
��ɛ��F��ܗY�U+{��<&�`.��4X�5��Q�s�&�'K@熘zYY̨�f�&ݷ+�W&�D����w�� L��1��w�qgP{ą�XdD�W �O�D~���,~�be�Y6q�Ub�5��E:*����Z�b�ü"5>)��O�خ�0c����j�:k�IC%2@���[�(�bNi��d>=d�4ᖍ�?FdW8Fj\�y�j��rmS������  �mx�ap���/D��2籄^G�Xċ�YG'cw[�j�~$�ݕ�����_J'a_����,��H�����X �1�	#��Z�~��|��!�Dڸ�q�7*��Zq,��9=�3=����R�$X�(�A��렲�(x�jϛ9`�b��9f�Y ��j�$�Z /�Y����))���QJ�+��,C���Ay�üpy���w���a�o���68N����������.�4�̃�,�������t��4o�0�SǶ�HR�=`#�ș͗ڣ�jTy�'$��(��iz���+��F�z��㟸F�?��Ϻ�Fd��Y=b�Gi+��B�%��K݃D>��pɚ����Ș8I��.<�P�fp0�����|O�h%��}��Y�u��M�%���&JX`R?M>ֺA�
_���BR������+�G� eT���&n�.���L!�ݗ����o�n&:���0���(,�ug���R%�g��Y:0��4��k*��'^����8=I;��d�-ȣ���Ӗ��H�j��w+�.���' �'��O<�zd�߂��f�ٿ�G:�	�Z�U�,�Z�O�28��FWK^;�+��J-���*�Q�4H���ޗ���p,h�`b�\k����Fv��,H"��"�w���`�e����z��O����k����yl}..��xl�݂�(�^�l�N~eǆ��>j�V"%�["��O�¯8y_M
�@u��;�%j���εq���$��[7��H� 5M�}�X����{8�'��	��5�����������`3�m/�b�P�ǵHIY���`˖���U&��*�ST��D��H�l	y �N�2�w��R��{��$=���P5��D�w*�d�u�Y��c��#^:/h�9�*T���AoT�m�uHj�*ud�k�bmh�DY5���] p��v�##����g%/م����K%V�,�Üxf��%�N�0��r���!4���3�O�?h"�����:@t�����s�Ů'���ʱW#��;�?���E�ёb�5�EDq�m��"$H��R�1�����a�$���6���V��%�OY�o`�����
��/+�ƩV4�Q�0�|ZW�;���*�T�}z��ZRQ��
IS��X.���u%H���f�3R�*�X��0�Y���{����h���[�D1^��
�sX(�ګ4f
��TWt��ļ}�k�gv�*c#&o[9*P���Mn^� �v�Uθ�^��[ehd���^g��D�υ���Osۯ�/�pD�r}T���Ȝ�G�>�t�l{R>L�=S�:����(r�=&�� Q�;^ �lg���o��MعrUL���+�ϣA�U#�E�V��L�[G=ȼ�"���T- ��,��m� �"KI^�i5��ӛ|��ߡ���R	-A"�=z:"e�J���D:�C
�1F3����#�w_>Q*��5A)���@�Q-ݽ��۶��S�b�ц)�$A�c�W1Ek��y���?�*�&�FAzy�$�z^zy����bP�c����?��G)���Nh��h�֧�x�¿j�8Y����S�N�.|@�@ZƟ�V�����.��j��F�毎q�{���ld=gz�������N������0ROn/��/&�+�����=����[׏;$x �mI4�N�\�-�H�C�c�2
���ZA܄u,E"�� ���C�O7?e>Oܔ��2�e�l^�!�;O��].T�Ŭ��cQί/!���g���(&��T_e���.g�G�B�`fG!E.�u��3<�J������̤c�T�҆�O�bz�n��w��#f�����Q[f�[��A�׈#�ϥ?X�S/��;fQw����G3�����&��:��F�]�ۖI�O�i�>�1F�?Ėm� R�[14\G���/~������P#�b�-�!6�\�'��GO �5,*1�{�ڒ?�k�Dm|kǪ���v��q]. 80�Z��S按�w��O���ȭg%8NI;�8�ӝ玵�^>�\_FZ1!�Q6�A����l2�R���<��{�H�� |
����{ZnT�n�i�Z!��]�q��<�qv.}q�_ ʅ�]��Pr<iW&L�ku�xK��W�j���� ���#��������H�D�X����Y�S�i�Tޭބ	@Q�� �^�`:��5gνOd���ՀUC��x��MO��n�F큢�|X5��b!���9���}yç�/�=�b�sי�[��nfv������:���A�?��T+s����b^#��k�:32�/O��:*י��P\��j"�C�a�l���+�������D���[�Z^��3%	�+ܪ���Q��ǉ'G�3
�z���+���t�0s�S���Y@�`�����ّ,�C��6��.���������3�m��m�8J��/8Hf��J��ǾS)�Γ����.�� Nmk,�,5�N?�[�Z���nl��������S�=��`
C�3��Ѻ}� ��+�H�1O2t�i؍�K�`��+�]��+E�����Q�����PI|�(�PJa�YM�����\$�����p5j���Ξ.�~��S���>�s�oޖ�"϶rͶ�:�ط�(߃�ֈn�ȥX2-J��q.�w
���1���֎C�QB埰���Z�M�1�㯗���TT賲yH.�J+A.�x�9�L�lD�O��_�{�+��{�8n����Dp)��k��+|0�a�4�o������n�`7i���k�tDz��F/E��Zp�F�Ɇ)�������^����1�=M&$�2� �+��*.*<����Le�t�z
�XF���������vB��iB�'0�Fྌc�9���܀獗�ɠ&���Wq�]Vb=L��~�Z����?�"�9�	��H�n���疠��.��a���ܶ���4e
�p�ڰ��ȋ�3h"�Dm���2ХAլ�`�"p��[�0i��0�w^�C7��Z�=��������4��"1��zB�R��[o��Å9�]H�c9��&�%A�TʼV�����@qxpJ�GWj���J�l���.�3Z�����������l��z^�b4�ybr�TGlYOO���l��SŮD�����
�D$L%2�hG�,�vE[�8_0���:��^���x�%�^=��s���\u�~�_(�m�ŖC5�{���WX�A�n�U7��������k����z�,��u%�ޘu��.�h�^�������%V;ݏ�)��]��eV�PM�Ft>w���Sq꡺�x�z��7��VP�j%��3�<�e��e�Gn�@��i���t���j���S�xng�&�A+W0Qr�4c �Z|��i��eu�R�v�R�˯<~��ނ�@\��1��vń��m�������N��%U���џC���o����fT>��^%:w#�1����I��9����Q�aZ�;s=� k�>����l���"t�:�(�ڵ��KR�[Q=���x�x�n)F<�y%!��rh����W1��صv\��׹Wcd�Fq&�&NҪ�w]�*b�|l)s�z5ް��j�_�����������G���1�.���ʚ�{��*?����Յ�(���G7���X���;Ο��B&�����15����Wō>�BV��Ϯ��1̈��E�	�wh-Mj$�9��Dc ��T3f�p��J^ڵ�h-o�ֶZ��J#h&)��I�UK�"�*�5Y���9
�-]Q��sB�����e0R�`㜢��{������������N���[��E*����6��}G��FI�X�k
ޞ�Y��N�i�;�N 2�nD��+�4R�@D�(�ý�Z�j:|�����$ ��(Wؼ��Z�k!2xm��F/�ٮ%�Ix�,��^�,t���X+j�+X�6|�S��D�~������*�%ؓ��7�F��>��,���I!�+�T,����d:Bq�]~D���8!��QRךC� �|V69Sp2���ZK��fD�E��?DM���#�N�A���t|�{VhR�o��&�Rag�}Z�>��<H*�5�����#�Iq=���]��	(��,6�zH�se̗�0�n`+���ݞձG)�7mhW�Z�<�6g��W��9�M0�����t�;�g9��(H�X����ý��[?�:G�V׺�K�� ����0��2�����"�D�ż��f��-4I<�-ũ�"��U�M��2Y�*�%�Y�k�.T���$�XC�ZgmoA���Q�4l�f.���N���S\D����� ��(����\�ֵ��CT���,�KQ�=�}��[T���S��g�Q��U����U�s�g�u���˅�K��CG�B���2oĖ�p�ڧ��92�d��'n@�do�dؕ�S/�Fe��y�<
n}# ��Ĵ Q���������}3���ɀ&��&:O���ǝ=�_�	V����e��le?�R�h���l�����L{���3�2K�Dd[�n��em?�-d�ɱs��+9N��y���XG�{N�1B���Y���O�\j���U߿�E�WUϔ�븡dj��l�|4�0x2����E��c�d��ʉRS�}�]�B�0��>B:��h!	gT��.4��PR��!�c,bw�QR�����Ј�b��(n7Am��f��v����Sy�3��J��#Q�wH�����9�$��e��p-���Ek:����n��uT���w{�����	��{�}W>@u�豀b��h�l�Su+`g�<�a�q���A���蘷�(G|W��SR���w	ق����8�i
LrM��F�u�R��U:��Z��<2�R�v,���M��t�HG>���M��������-S��-a��3�Yd�F���µ˾��č��3�*�֟���2�
��AX7�A�P5�d�� .8�[�l��HA�r� ����q����f�/W�f���i�2�ր%�p6��`#,}�M2�hIˤ!�g���+���cw��RO��,�t�#�[�r�m�������
B�����ؒ��Vlٻ~sa��BrY����6?�¬?�㴸���M_���1Fg�]�9]��Fj���&d�
�Bh0�*Gl�l�/�o룃*���`'c�{��18j�&��|���%�+9���l�//L��b �������mm��
{/�'}��=��U��y��Q*�4��vO:G�v�J�<�l-�3p[�GY;��B:�����c'�P���w�zJ��Ր= V���A�1�ɿ���ʿ&�J�s3`��zf���<�N=�~O���y�E������zB[�fa����i�_�D*D򍉘��ʤ1�R���$��7o���ާD͙���KRW���:J6���Q*�#��iґ2%�[$~��Q�����/ё�?1öq.�[�"A�5�/�!���t^*DӁI����)�=�'K���Uf}cm�YG�ͣ�x�f�8<�d�o�a�4 �b�e7����l xlY�9����T�����é��à�[~�0���4}�B���Hբ����uٖQ�I�g��u�ۗJ�@�i<OR;��E�^�&�_�+�جA��2�;�B�t�������o]��"��!������&��Br��nD�nj/�u��S'Y���	[U0x\������C�>b�[�0IJyvf���[g�u��	}��7�U$�R�lD?�R���rg�iX7��LH�?�TD�ȱQb`���n�[3��d�28b�t4X��%��\�B'�TXYV,�MQ��!��:��ЀB�$��d�bt-���8£=�rh�'����4��r��[��I���;!�S2�K�%���a��.m�.)	�#	��������hXE��á�����X�O4s�T�ȴ��~��� :�<�u�~C��]�J�Q�H��Ti҃�Q��]z]��(х|�0a���9m� �/D.�p�䇈����޳pdbJG�Zde�=�}�3�O��Y�]<2�s�u��qs��lz��x��[� udu����c�	��&͈s���֛OJ���	F��Q��\��F������Q�����C�y�C����������??�^��/2q��_f�m�&��;T�~�O�����9�����Zb���.�c������Г90�Xe��	�I{���Oe%�O��G�dk���m@�؋��U�ɸ��J�ɑ3�2�7V�5�>����ݵ'x���
��8٩���3��I;?w�ċiYM������7Zd���;���Y<Y�L�d���.;ޔ���w��ء{��yma�j��n���;Y=�\%�le+ğBEӲ�o[B�6N�(������?n"�ՎY6׿�.��KQ���Ҵ�W��@p���]��� T�~����ŀ�.�����j��P��쥊&�.#U�f�"��� #�r��e9��5�a�<���q�}�&��.�0��Z8��5�� �x�'�ը�	i>�3���!R���f}��B95*�#��`���PL�-x�i�ȷ\Lj�5|��,P�_��+�8�*_�����8^�h[�צ����]�R)iv8�KC�
�w ��ph�h]���
ϓ�-���L��ʩ7	�>���>����թ�\~�߫&��J�I-�W۹	,��/
v��!�eo��n:���h���$v�X�b�M�e��IgN�y��������m;gLHWhbc
&�s��3&�61'���+U͒�TTh�X��L�%!��<�"͂�cu�R��r59N���#(N_�3b��M�y�7�7�I��I_��^�PC[��	�O�?���5�2:�i4������s��D}8T��)��6����oc�m�7�Z7���?c�pH���u;�e�Q�Δ��y�@�AKY����Y���!p���#9�%��ĩ�jJb^d�~[UB}:vK7_@�z�>���R����˒��3����ȪZ5��o������y��*g��;I�d����L���"�	���ȉ��~`�N^~W:ﰉ��"����#���p8�a�Fڻ�L����,t-�����$��J�d&Z-�m�}�!�uw�6�}Mp����e�ͷ��L�����aTw_kA��ϊ`v�.�Χ������E-PW��ժ�AW`�������!�*@���z赎��u0�~/y���.��
��	K��@t�u�?#��F8�CTG����	P/��DB�F'�,�V�2 0ZB���>�DX`$����w�H�#������V�w>"�n=y	��f
�������������� �]�������������w���Ĉ?6��3�q�}�"�+�'k+��h��E��o��B�$��JF����I���{�X�,r���wC��$�<uLM�v��O{�iR/��nL�!��s >2�%Vn��:^���F���e�y���_��&��4��է˭��Gʔ�=)��ҐF�[�J�I�dIj�C���/�>K�a��L=�(���{V
i�T4�i�-A��X�]�xZ	F��5|^K4����K��SL9�qQ����P�V���,�P��8�,��C	Q0,.ؽђ�!�g��ڹO��>�
V�î�u�9�s'�ہ�վS���QP�c��oE�)���EQokS$)s~����\,�gY=�ٿ� (ʪr���-~���� ������Q��Ŷw�yt��}�%b����_�\m��{��O�s0b���A�h��*M���~l8��&�`�< �$���9IK���?3 	|�&N��e��#�es���e�l�T0*y�dE�t/�&�j 7��M�KaR��VE @���H�E�`(K�qj���k�SӼ_�G�!�p��멈n��4�*4�b�����b%d�S	��_�6 �e�ǎ"4�H�F��5/�F�����FqP`��V#��«lIOnO�(��a^0D�	��Wح�ѭ�[fڵh�HT\�?4�UTMn������-8w�����5Xp������w��?�\�Zu����~vuWW��fס>��k�n�G��qKZ�$k�D�ť��J,��n�
�#\�>i�@��Dg�5=[D��&Y�"��~�Vz�hwAR�H�rb�]Ϩ�b�TY�D�Ca�#jȼ:8}$��+X|� �*��Q�=1�����S>�\�JPd�l�Țӱ�5����Z�[;R�B}�b B�D�:)x����c�]��א�Z7g�Ze��v:�X���q�Z��V�N�~bɆY�ƾNe�0�yU����׋�����g5y=�-~6��o�1y�DV~2h\�u����w
�y�3�y�}1yཌྷ��Я�F���&�_���	LL��<
a��82��~�g�je�����m�2d��1z7)ew�]��MC��@u��JSc���c�_�!.���5��T���7�a����u:|}f��s�]w�f,��I-GU�O�kГ�PϨObw"a��}2CFfT�C�A�+������-���8C��Ur�+^ _	:�f��`0gD�I|�E{����Aܨ_6��v�ZB�io/8�-Dd����d�z�����n��r]�%+�K:�)O�����QWu�]��A��U�	˦�S	�Y��וǀE��={�k'/}�6�^�\�E��:�;��YT|���-3^B:O���������os|)k�[�58Fg���Fڷ��K3շc5T��C���u/b�����9�a��\Ih�4˹��sm�k�Ц�t�,=�N�v�����)��J4Y%�t�[O����i���En��7��<�+�]~�P�I�%�hkAڤi�ps�e#�8n�x��{�z=�B'y��7AR+,����D��i�t�t�`�������Q�x���'jB�TK�׺ V�;N�R)_ع|x5��e�L����9=g��ǔ,U`J���R�4ʈ�j�?_��m��aݍ���e�b�-�b�}�������`L��"l�E�g���c�"Qn��-L��c𛸏 '�c�e�t�����FIU���5O,0���Gss3�Hۗ��p���5 m~�z��zh�ǆ@_n�]�#����g���*��@���;�A2�<gu�Z҉J��s�*�2u<�Go���p�o����0�U��~5O4��5ܢ�N�y@������!hA�@	�.�.!5�J++Խr�j�;�_�9���J��m�����f��[7�én����mU����C^�������fr�C����}����`N���I�����s���g��󭓷��v#���?������Y2�]�:�ʭn���H����������'d�7�ThS�K ���궁+��r�U��,�$����� �s��7��H�?��eȈ�kѷl��[B$L����g	��r�QW�ݣ��S�dza��߰0��t�����-��-9�<����I��eϧ���l�OX]�ټ��|?���\��_01�\�:�}�����7W/B�$K� ݟ����#���	o�XňXˑW�g�k�TJU#�%u�Aw���]�\�a�Z�|y��Z�����R���y'�fjqA����aUH��Cdg.r�abi2?��|�Ⱥ=��d:�Ԉ���ʳ�X�5��]{D|5O�Q�6���e�E?'�v�3�W ;����x)^'T�5��H�#c""��+�ʆ����O����ϙ��Z���d���[��ײͮk����x^{��
��֪8�`�AX�L�Z�ތk�o@��k>XS��ۍ G.���`�R@JEHᢰ�-3�S���:�;~Q�$gE�y�(��w��F�7�˸�=p�u�9{jS&+`P��&uf�|��{��le�˔v��e�2>�kq͏��ݗ�{B�9c�!�2�]�0�	���e˽l�ߤ������[F6k��~�l嗖���3���;�����a�,&g��
���'�'�V��v#�+T0�P�D5�x �KD�{��5��t���V/�8.?�\�V����<��U�-��͢�Wv#J�V�+Y��4�v���d����,���R"�򊴜�$�ó慌�3�k�M_lS�<%�I*�c%˧��"�7rk.Pu��l�.��<c�����Tm����y�W�����L�N��g*���5���R�b�梉�x�
%~���Qe���"�C-W��
�>������<��WP&��2����T�v�V�uJ��ѓ��W'�F����c��c�ճ�y<ڀ���@�ǭ�!��̳���q�g����B:��O���=�s ��ҹ��w`� ���������ֿ�P����g��?�>��f��s����?s|��v�*l@ �������3����P� ��Eb�n�Vcʽ��.umΛT�X�!ml���<gy���&Z��
)�dx�E���;�ف<?�kU�[���v�~௡k���������C�<i1��]*�а(<sMX��,]��i�e������>i?� ������v(�Ge�M�0���!�9!_E�12T����F;��}��z�A��Y���h�?����-�v.�_�E�§g?��s�2.7�N�r�γ����kS�ǩfu<m+�2>T1=ጎ��X	�[���s(��K�S��`s��*,��jw|�es���<�R���Tw�����M�����,(P�~+e$�g��l�ډ��3�k�=�m_y6�2�.�0h�7Z��g%1c��7���Ω}�vk3�Ucؽ.��b1o�dJf��O�����n�Q.�i������s�M�=�
T |fh�ٚ�ʵ���Lۺ��U؂&"/$᫠5Z> � m�8;��o�q픀f�P�Ƈ�.&pum�D?CVZV�� �:�T6�����O��^+DpFz�������;NoooA<<��B�t|1!^؊�PG�&XZ��8j^�^1�9 �	붭�a��s|JܧE���	�>8��q>%q8<a��-�����w�'\��(H�W0[~�K���o7'[5Y���,�[�m�j�F�N<���p���p��y'ﶨ��INt�ךˉ��=����Au[��y�o7���~_/U{|��lq�?,Ա���z�l����#�6��x���U��o��o'��'����c[�2��ԓS��h�*V]n�"�>Ξ���,}u|��щ[+u��0V��_����� �1"�Sp=������%�R����n�Ǡ�M�'�=�-�_g� x�k_��	0n#�n(��8A9�g�J�l9���C���y�5�+wޮ�<?�gs��O�b�J3]�������(X�H�k����x	�G�6|C����'��˙0�$��%,5�FOU�?����[����͗\��m����Ϳ��H[V's6��
ag)���B�3O�U����� �5%H���0b�����6,��S����Y�P��aA=�o�s�]u�.7�S��p�3J�.��o7dԀ��$ ����3�/��_֐v@���Pпp�  ��hY`e�B�t��o��̕�w-3Tώ���S~���1��Y����j $l`m���:4��u-���	�JZ��E񋎙�^�����c��ŽTMB�6�mB$'[�+fh�L%'��	|�nS�����f�se�e��H�egV�P,�Ff{�v�Ă�Z�03��q<|$�n1�����u�z�Z��%f��iY�&�wS.�&M�#;2&�]k��W����`���E�.G�Гj��"��E�G�����������]_w���kŲ 9���w�G+���l������v�*D�ғ�O���Td=���-����^��1�"�����o����4a^��ç�j��#=�o7��]�?+�y"�2)�Y�ܽV�v4��3 ��vu�VX��h��k�[�	����wɁ���W%1���|�S�,d��-����φ�o���J�:vu�ڹy��k�۹h��0�a�Q�Ȑ���@Bj�f�u	����ю�s��"�x�VxeM&�����IQX�n��رj��U$Ǭp4����<��fv�(]���Z�L��葻��C��!Y�%~��hU�8a����$ Zn}�|J?��!,߯;��l-�W����
|^�x}bﹽ���2�]��h}v~��I��'����|6I6R�~}��� ���vaD�2Ւ�q�+9�J�iT�b3n{��(
��c�O2�-��l��8����ف�R�o4ʚY$����x�z&�&��-;������\9"�S�o/̡DP3r`�V�Y�)�Z&�l�j�y�wr.�Tm����2�q�k�ԐBT�@g�1"�n�֏F3��)����ޫr*�+ӬBlDԱS������N�sJ�"�̝��W��o�d$�}�o�8�ɥ�,�7����ǘ�������<�*���c�V��9»4���)I��յe?N�X+��Ծ�̓����<BI��e���
2TӠ�S��8:�
H��c��ߍ������;��ڊBQۋ�\*0�4�F�t���m�W MW[?|T��SW�<�H�l���_�IG���q�u��Q"��l�iy�1�
�)��%��sH<�ꂳ1ϣTh#�������Lc�EC�M��f���P>)��Q�x�n#�H+��JȆH�����������{�]]_@��}�(����~����!��������i��`p�i�.�©P�Ơ.��_V�Q�J�D��>�PA>�ʍ�dF`J��[������<S�鋲�`� HG� �SXI?ۣ�Oɾ%8����Ζ �LAJo�DAM�Sz�M�g(�L�Z>�Q��|/�x�}!�����-�b�����[��M����^�'���o�����뺟ּj�\�'��_�h_7�>�f�Ԅ�?��k��ݠ��<\���t݅�����7ި������f�acI���8;����O�<�����ۦ��+�¯��;�G_����%�w��m:����jo�9�s��>[�2U@�0r�h?�z���W���T�U��/��vZ
Tۘ�X�iZ-4"&W	���٬�RL��� Z��0ɖ/+d��*UCP��ش	q��JB��H�^�rG�J�����GN��X�1ڼ�mn&s'���
%���G|<���j���fYѪТ��w�ng��L�dr���cs�0V�˦'�y� �V;p�ʴ��l�ef( �clY�Z� ��@��`u0�OTW=Z8ǝ�	,m,�[١��`�V������<���N?ѭt�ok�6L��0��x}��o�kA��VJ!aSΐ�Y-����ma},(�/�]�@)B		�GT�n͞ǭ�W�����b�_�X0�:�a�K��{d@'�Z$�''>�r��W�$�`�0}7��0x��4��,%Ʋʴ�U} �Ҥ&d�Rm<� �E	�\��:Fx h>��)d�� <��:�v�k<���:�����9��� u1���7;�?�����>y���q��Э,�W�"��R��R�h�v�Z��B�: 4��GmZ+��_�~�Sb �!.ǥ*����r]�I�]i�P˧� t��Bx��������r�"S��M���2N�*m]`^aC
\%)��U�f�j�)�L}�+���Qj?��+G�������K��s����NqT��q���M�v�4N���v%}-����E�`mHs>�'���r����ҷSl%��l���uw�������vKH�mj�'A�N���~�ѳx5o,T;�����F>K�CR�>W/��Z�x��ѿzY����<m±�R,�@b�O�3��\ȟ�I�HC�wŮ�* �T���
���>0��Z�\��R�i�Rj��HIBJ�~`�"<Qʝ��`��~h�ZHG����"Y��?���v*����X��Bܯ���������wX=̓G�_�̻��ɡ9�oF��sx��>��f�9�'(��ڎ�	4b��	�4k-��O|s���>�9R�(�����=�����I:2W���,m�)LNMǓ��;�������v�N(��*�Y�&jֆ0�������f�D��p�
�Bg�,��� s�'�B���ӘP[��*������y��ܠx\��]T4��ys[�vCћ'��pI��EyWu�5úeb�p�]��ʚ��J����J{�q����[�B����[o��.��qA	"]��*��:�,Cd&�F�F����ʴ!f_NT%�耛$&e�ry�XEz�U�TA��©._�̌�ʏ�eOȝ'H�<#|�������9:;���KBF���Ф_���	ܬ���G��U��	�,GC�1q��;!�+J>��,�|��p�
��&?|<�Y��
.�]$«UW02�ٔ�@4��#�:���b�S�#�p��K�`-X�f'�ր��FQ�����M�>ɉ��i�O��oW_�x�
�׮����|dq��boOͿ��ź���{F�E^��={<��ִA��D���_2:I��ɪ{�_�gX_�L���{ZR���31�~}�����9c>3L�j�@IR����N��e6�p�N�����Q���o�f����K"��/~z�ۉ��:K�lc��������t���<@��8���>��DB8�G D\�NqN	�d����*�Nn�75�z�#���{�f���P���F �q9�nkp��e\T?Q��b�:�*<�����U�m��s-O��,��'�s>P�0��g[�����;���!�VdC�e�@�v���� lI��q9B(�ֶ��(a������^u�kp�-��a�L&���j���{OMI��	ǽJBY�=gU��	��PF�x�EJ64�����+j@��=v�i�4ϊ�S�[�n�
�4Lo�4������L�/�Ƙxe�js:\eY���P	�~|�_�Ǩ4��k�[���u�n��IO� ����o5��R�F����� r};�.�:�q�HÏ.�����+:$�O�>��y^Ӡ���^^�����e�U�����Y[��,;��J-%͉a��9�K�pdx�R�/�-�Y��|Yf�rT�PjH�����4�[��Vp�0����}���[�]�Zƌ�+O�<�]/�Фݸb�uvo����I���}�����޾�u�|����CB��O��|���@#%;q�|�e�7cH�%?;�E6t�a���2#G΀S��4>Zh�d�Lf������\�m r�Ѥ��`��a@ES����Rb��B�4�n��~�9��Ȑkc9�`�v��v��&S�ԟ��)�&Pk���fQxן��K��8�A�`��T���lb|��^?���!7�,.�=~��Gĳu�ZղK2��������nq[_�� �H`\5j��ȡF*�'UI�0�y���s�ݿ���k���1�yk���}����wzn���m5��7D���ڙ�jZ��n�Z�gwfv�*�k�W��Li�}y���
<mH>���VS�q�xv�1�p���"�����\�$��?3�yOqd�j��`T�����(�?e]�t%w�Sa�~�4�#
��fo�g����%F�"`8ޫmA�\�:���Ao酎H6}�0�!����g~���e-D������Wܢ�4a��8�z.S +��7[�r���I�3�:��'���Eя)��)9�L_�L�W9KS��cY��u���t1�����/��Sdf`�ª��?�R�.c��j�"�}����#q�/�͈4i�����F2�].¾E��o\�Ut
����V�6�S/A�-be���*/þ{:�lƳ�^�ӫhiē���Pp�+�@䉆&
p���ɕ��n �h]'E�/�����rtdmꉏ�=%�2�td�x�ji-�yS���M�$��D���b�P���~��%��ɠ�n���Z�[�:�Df���rU˒oI�����7��5�DA��jp����I��*M�T�Z�,�R�D��^�&A��&�}{{�w����~�+��>���"D!]�Ps��s��B�Q����KV���BʗX;u�Y7k��_�{^���&��a��w-� zj%@��Tv�@��O_:8��(sc즩@���˅��c.��(�I!���d���I��Sw!���L��#����b��K~��x�X[ �Φ�)�G�����d�_�U�B���
q�h�Z$ܯ ��b���!f� �#�U�#����N��փ	'e$g%�>�`!�)
�?�k��=f.�Hu���p[_�Z;��!��ø�	���$-��a.s����\$}�q.���t(�N<��V�-�n��L����5Y�9�6�r9�u�S�@���:�:|������\>^{8t;c��k��.��-�$�g�g�Z6vՖ�	���b��ߒ�2���������x��R5׽�K���%h6����a��+fD�徱 s�3���$X�sH���SB��b�b�C(��o���f��|-E�����+�������3��^��)`����<[q�\�=/pW,!jcj�X]��Ԓ�8; ��e��#�G0O�͆�ǣ�B�{�,ȭ{��Y�]�}i\3��dM���u�8��"a:�f�]�}���ap$�C�".r���W�H(@w�E��oDGM�:��k��6^4<W���c� �O�>W��<N~�����^�_\����d���Lvmj(�_�Tr���$xc~����D	뺐�i�U`�@QܾQ�ɪ��I�����@���2���$F>pxS�7{ Kβ��i�ǩ�ߙ���ޜ���42n���|������왚�3L�˝�w#{��_Q{XM�����������	�Yl����((�`�[�y��"���֧���[��-�,s��^JKRI;{+j�~�L��W �ɠ�!�(��Q���3r��!�|����0�ύ+�$�Dv���ֺ�0�r%����Mjė5J� ��p�Q�M�hͺ%� b~RK��oT��mS,���.I6Es.��Jպ��ڍO�8��P�K�7ǆVW�P�
�����2�j�k��'��^�UԊɛ/�F�|�A	�_P+�W�y�}v�w��*_�-��z���ӞP�۪���!�{����z���c��`S'?u-�ߤ
HfO��'gW�����;O=$��bX�W��MI�u�j-���.����wm2�/$�f����	%nV��Ye I�BҰ%," O¬��#�E	�`υ*L�#I�nAZ��Jf9�N���9J� �ho��ջ���M�� ^*�MN	x��%�m�65��b]}&�;Ƴ6�S
i|�B��#���z�^k�X7�K�*�T�gЁ�DZ��$�lg#��1>B��@�7ƝrZ�nz��-8���Y��1�T�R0����?�+��
c�Iz��#�&j��^,i6��Z���<�K��i:/���N���Q����]�����PS=�sUp���t��o�D�M0JQP��`'n0��깰H6"�hS>Һ��S��>��!Q�:Rn#Ʃ0���CCB��]��fJW@�<q���du�vtt��=���9�;�*k�+jk�����21Y@*��>cо3��$1��
�y�ஓ�)���[+a���^����h��}pw��d�]�%Pwz��Y��5JE�`$�&}�w2a�X��-��t���SSS�����:��D�������@��sa$5̊ �4��P�Ն�R��1���i@K�����EhY�j��)���-�����T����y�X��L�4�t�NZL\*���L�O�Rޕ��-�_3?[Cnj;��8->���C��a�e-���ĭW�͆�O��˿D��2=���t|�io��ήVlK�gk�e�����I�+���LT�Y2�ë��ħ�����D��m���ߍB�D%�����E��t�kX���@�|�LRN��;�����(�D��?� V+���o7c2�5����3���W��!�(�7�2"�s�lL�ꂪ�{��Nz]�����a�|���*�I��,݄;��,�i�-�c�]aFh� /��\��#��)v���,q�|����,э���*C�W�ٝ
E�c�	f��e�$4�.s�V���h�Qy���i��]���Ó�){��1�ls!F�h�j��	
�C�Oì8�צP&�����ػ��d�߶	������ǘpAZ�aN��1<��w])����L���b�f�J54�P
�`#�?�X�ɣ�۶X3��,�R& /�w�� ��K�YcT�8A�هй9�֎3��<`t���p_����V���2�Z\*�*^]�^�� b�1&8�G��x)8���E7�Mȡ��4d	:�FQ�O�Fp"��ɘ`��Q��5v�]0r$�l�_4��f�e�Vw<N�;Fg_��1���қ@A�.��B<��q�ı\U���e������OS�Z��-*$q�кLVĤ�����c�ֱQ0CG S�+��3k5�F���|^�}`��;q�l���[|����!���.jh��	uw�% ��^���9��E;d����.�����`�Б}��,����X���h�A��z����Vf����U?~$�g��E��6�,jer��aԠ��^E���z�Y
[�]$Ĺ�H��kw;��u��"��E�g�rީyu� U�.�y���1��8��'����O$��{�Hf,�`:p`��E;g�z̃Z*M6�Ξ��_KW���T�N�5���uK��EI�e�Oy�~�R$�,���a��ͅ
w�*#&(�A�~�]/���z/;�wV����ٿ�u��t�t�?,��vu�F��o[�Пj�����o�����g|g�U���?iG*^fj3'�g>��n�(���\��Z|�c�2H�`e�MK���(�&�j��B��.��o�L��1�
Ng��F ��Y�XEgk���������a .�d.�Fl��.����SP
���W@�=��y:kdt��Ԑ��z�	�Ϟ6isZ��i��4YGN d{[�kd��e3?��+�\�q�J�2q�d3��M%������wm�g��R��*u�r#��X��t��ԝ��|�c��K�>�I[&݉ӊeo���� =f&=N����I�Pm�f�Y��u�(���V&t;��y'd�ȗ�)H'�G�j��TѦ���<��Ƒ��n-i��]���kĴ�O��*�����f{.1�1�D2ᴳjI�ٓ
���dL�Y>�ʈ8�6"����9;:���T��9:A�I���,��o�֣"�Q*ĒWn�$���ù������C��9��i{
-��e��d�(~�q� ʹ��pN���+�/A$'�I]{��@�~B4Q;��@��n:�&i؏o�o�=�b��q��`�?�l�3�V�Kն�`�l�7D��H����*�1藤0Y*��U�;��REH�Z<?	v�!���F�I?zpI��h����-yx�
���B���R���n�>����4��.z}����l��v�O��-B�[��L=�O�u��_�|_��{����n��ޮ��l�;:ǎ��%TTO�ߨ�Oʏ�mM��~�ղ�.���m���X~��9��7�{��?�|-L��\�)]\o���οL����1��;~O�'R��N���g��
�춋�Om�`;բ�f�Ю�q�r�I����?y����:D	�P�!�T���گ�;n�C/�P��e^pȄ_C�`H����S��G�UL{�^bX�Q�k�#��4����d������3�����ů���+�-��vҥ~.^`���k��dݭ�4+���k"����1���=:F�wj5��Ӗ�O���Sd�G+�%5^��2P�Ȏ�3=��N��i�uY���F��'I���yhg�h�oU��7��lHcb?�J�� r���ez�Ñ;�����)Vd��$H`����׆���, ,ߣ=�^�-Ch.m7��%5K	f(��9%ӫ�Z�V.ݵg�[�O�צC�y���Wڋ�����~��yI�*�Ỹ.π�i�S2�m�lQCl��Z�8?�q���?��,g���ȣ�I&y�<~L[H�p{�I��z�����E�y��J�p�D�9M�Ock?R
��i 7��G]��ʂ�D*r*Z���%����Z��UTezN��D����R2��d��-�¡l��T֮��M8��������7Y=�si<}�͘9��?��0�k�!�o�ޢ��ݴ����\�8L���[�?�U��)� �!�ߡ��o��1�s	)T��ܖ�Z�^=��� �_ߌ�a{��0��/3���v�峨�^$Dg�!W)��!l�_����o��-'՗��"Q�#���*Z�T�d�����,���>�V�B���H�(j�f����e&Q\�@��2>L�����+,]SU�|��<v�L��t.+����ŧ>^���r�O� tq�:�����p��vZǘ��¬*i�V��OQ�0d���U%���	0�U�p*���~�|������p�V�N`���y��nuK��2��_�o=���>�Έ��m,n;z-�;��l8y�`��i�~�o��D�a��_�-���Ijzw���n�F2,% ��b81�QyJ�_�}��(����S�0�IQ�`�&��k�X[�Z����P�{��^?�%��g�EWA�x/v�.��\�Ń0��*I��
��g�M��b�O��2��UE�
luN{X��?�\����)ĐQȑF���\��wI���~6C��
lf.WC���RA�WF}Ac������&�x��a�<W�R�Q���OE���Pq��9@�Wv�<
~y�)|J_p���!t��p�=���"f6m�=�l=tgj+��'��$	���s%˦����2��G����0G~t�w��zZ�fv�m�i'�R\]�s�"V����	nu��:�Q���i�$�I1�˦[S/S���e��j���蜏C�Է���	��-�5��.ר�t>�O�\���T��`b�2ܚ�Vh�A��TG���v�c�T���ύ�|G�b�;L��4�.�	�X�fR>���X����	<TP7kW�\���o:��\?w'�r�#����7�k�؈�2�S�W*���G\���*҃$�&�6�;X�/�z	}!���)����T�%��!�o�˚��^��XY�}ܚ)yJ
)
��t�(��RX�+�x舅X�ˇ��Rp:��	y�l#{@@ ��I��]�?��C��!��6|�+gW��'�b�V/��Qvin�LlOP�l�[O���=jP�\ڥ��%^ �8iB.p5n~ǅ2ʜ/��<O���IX�������֍���v��}F�.p�DV(hY�%��r�ζ���{���EJ�����{S�`�]rAa�j�T^V咽�����W�� �qO�M�֓8����л�V`���E�@��<r����1�KS˦1ѭ]�4w�)����!d��H:ϩI{_k�p/ˮ���M���۸�/>'L������x�_͟��]�P����9���_�Q����B�+�-&}p��-�O�wU�m�n]����[%���v���s��d�~��ܷ�Uk���a�M[P����0�n�`+�����e\�����7��-�&�N��/��a�A֤٭����$�A��7�|�'���%�x��+H�bv1�z�bqh+Ζr+_��2d���'��@��mY��w�*�o�>�k�磌�i���~�.|� ){�|�wK��J��'��v�P5�!J��*<�T��N֯�(��.�L��ԫ�\st����x��2���������jI���a59=$��6����� P{�,�wao�)$���|�b�E�Uz�����<�F�v|fR�B�,œ��P�Q����6Ys���՞ēeY)X&��� O���;<�N�Q\�5U�������ck�ao�3��s~�~�0+I�`�%ȸ��rt�Ss���o)>f��#����l���3��5�u�1t�H3���"O�����!4MA�ҝ�jil����hrM�0���,}j4"�C0d$w�!�i�����$��'i� dϾC�	y��fx�=F�p�Ԃڍ�����;M�gfM�Yn�߮��v���Ⱦ��+�C(cj���4��bX�֠�O_�S�$�I�����C�p��a�&��C����@�t�� {һ2>}�z!����A��Dr�TK�
.K�E
��gk�	��r[Yu�":n-ǦT�-;y����,I̥��o���]]�J�S����<��t���#L^��w����>�������r�ʹg�?��W�gM���%�:��ݣ:���t�=�T?������c���mT͈�����mV� ٥!�]N�oC2_��-AN�j��C�R=Bj��R(�J�F�Lr�T�q���X� ��$�X�pj�,�(�϶�-gs��$\1M�hɦ#'��-�Fep���t�%�����*��M����+!��b���ɨ�|�{�4,� @�@)���E���K!ilw���=�v��j�N_˃��8o�;���7sz�>_m��w�,��wy�'e�y�4�}�{x^�_X�y6)�H�^o刽�%��M���'t+c��|��	(�C�������<^q1�l�:�B,X���Z8+!��Y������]��?�b
�mKc�W�
)h,׏�m|�G)��4�޵o�S?��"�h:Դ��8��j��׏��.3���N��Y@K|��uc{z�-�Z����c�do�[0��ϡ.��)O���|+�-��=kI��hu`/!�ʀ���,�����۶VM �a���1Lk)�������4��1C���%e2R�ВT��`����$��	9d����ÞOp�bT8jHLą̱Z��E=9"��e��=��!b��J��#x�̱��j�:3t�i}�Ζ�7���K˰���F����G���J)�����	Vc�עJfHW�ϙ7�`dN�]z�E.Xy�;��0�ݥ���%}��fL��ce9�A�Ŋ9damK��fnEc�<z���Fd�N�(bA�Q����xG\ TF���M;�q-��~i_h�B]�.̛V���_�n]߶{����i�e�Cm�tz@��"�"|[&�)��p�,�-$鶛����ۚ��.�2A�\	�JdYqKS�����,�!j.������<��t��Bd�й��z��A��j*m��Afg����w�f�� �
����/fD��ꨜ�3� ��q��"ô�!�����݆�݋���B�_��ԻW��wQ_��n�\����Z������� �u�ݸ�g�o���ӭ#5;�������U�(%X�#0ܜ��{�r�2)%F��DCX��Wq�wZK���j�JĤS�|�9q�����;��V���;A��#'�L�sX"t* ��w�V(�>z�0Ur�z��0�n|�u٠`���YσOR�/G�����*���O�!�#I��-#�~I�p��Լ?�m�֜WO�ܳ�:��컭^������5	�<f����� �H�S�]5��3����_#�������M���)�<�*������l+Wk��y����m�S����fĖ�U!�j����%���D˵8�����9T}��9�(Jk��a/;��u�މ�H�h�ؽ�b���Y��a��ohy�'j�|E�=tP'I������D�� ^��0@V�4�kn�xd�M����$�xu�G�-����l�S��!%��v��pd���}Be�m��;M�����վ��/������צr� 9Q�y����A4q�%���YIY>x��?sMvy.��j�6��ݭ�H��ҭ�$c�8��]����m9(�8�!k!%�R��CMun�����Juc�ٺ&�%!R���	V땼Z�k:�xf:&�<�m�t��N� A�hrW�Z�E�k���%��c|���7�rj���?�E��n�N��׏�/�U��wn�&�����N�Fy��$1�q���b��<e.4}"�}�t�����t���YY}��t�!H2;���稖Xf	'��l�H���&���Ri)5AgJ�۫;:�<:���g���X���̔6�bE�B�ROX�B���T�Q�3��3���e�:� 4h����x��a[�P.\�}�����v�TIX�*N�5���ʜ�J�V���j؛�v6�.�n�����`�q�_ܱ�1��f�'���������{��8ʎL
̕&���}g����枟�O��?����2�/��t���j���I �?�ɹ�򨺫j1^3�S̡S�� ��V6�V6گ��o v�z��W��]D�\aRA%��)I+I'7������d"hɩG��\�$�</�՚޾�-O�K�)~��o�R��DnR@�c9b�Юmu�Ӑԥ��!�ڥ�뻸��ث��v��2�1�����I	jY�紨S� ��6�M*�P�&����&�3��n��f�����=-�l�p(��귨	ަc?��n�?��|���"�e�����A`W�q�W��h���C�Yv��u�6�஍�;����kpn��K��%@p'H�A�;�%��~�q>��{�k�Z�v��a��$�h����'xi�C+�-�9F��m0��ʻ-�(��$�%��=����a�=hS	�G%��,t:[;ț��>��yL��9L�4�6���d�bca�y�M��Ԣ�P�'�WF�bSW�b:����bި7�TJ�������辏���q�l�%�@*��<4�J��,�3&`A-�AW��<���|��Z�,edc����7�E�����c���\��$�:ٗr���LÎ���y=�y|~Qe�È2C� F��@0A��4�3#T���Ҽ|p�"S���\���	qU�=5�TF�89��=H��n[*n"-by�4!��.��f/�����Lu�1�P���PM�,A�;�3�s8BD�z�)��Gf����<É�=�cf��·	��g腎3f��5ȧ�������:���Z�?*N�7��c�+�x-���]�x��^�5�H6�!������LFچ���MF���ks<�憎"�b]����}̐��[%�����QŽ����'b�d�֘Ґ��R|�/�W�>}�%Ɏ���=�����>�Q)�x(��&����L��jkR��^P�vi��Yq6p�B/����.����2F)��㵠MPM�R	��]�F�CNC��������y����!q������a��e�RQ�ߗ��d��v�Y$�9ɋB��bU��g� >��h�WgW��}47��6�c�5�I��cD0T6K�T+�$�]nWvs�>e������yKm�x��-�SE�J1)�����rvk7*%����=�ƽѩmLu��/��^L��O��-��/�#u~q��J�������,W���́ѹ�L��� �$[.�Y�߬|Cd�Yu"ZPf=�P�*2ݘ�<̂�^�R�z�h�T�Q@T�>_���W��7T�z�d��|�1���6h}w�غ��y7���lU3Mz�
�-#y֝V�?R5��p8���j�&�Q,��*7Q*�e1>
Lq�l*�N�%�^�]�tAh��0���r�3Vi(]U9$�jNY�j���wɵݒ��"�*r��;ʩD�����@V���\������#�R���c�I�Xx���9|�9Zvo��L:.!�j��"vυ{�98ꂶ_�A�k���q�6;�h�0�e�dYf�7q�MD1o{��KHҳ�E�*z�J�S�Keu��k:� ͐��&檛�b�Z��qy�Uj��L5�LY�MF�!{4|"�k�<���#���V���GH����B�ü�qԥ:{-DqIH�U[�r�s�媺0`y�oN!z+��:��253}5Zr�����̈́��������m$�C�p귗)QPV��=��Խ�l<��-�<N��^F-�<w�\��5���j�Ԛ�������K�0���dJ{�kr��PĉQ�쭿Z�xr]���q��٢�1X���'ϲ��R	��Q�LUFVI Wc��� s�WH��MzǗ��p�\��=� ������TY"�o��w	N�y�l�F�
�t���$+Q�dg�7�#ܗ�q/d<W��^�âs��b��un��c�����์�s�]�R���f��"~т@�'�s\J�?=�X_k���4�{-t�D��(��B�f&<e�0)Be�����Ӛy�Q���ĝu��3q������Qk*�p�~�ۆ��2%�J:�c���[wʶ�� ����o�@<9IE	"V�����=O�X���J��8���%��k?涖\�Z;lr�S�_�JX��Iv�[35PN-�̂�հ�1�ulm���P0�Dg�05��Kgmy�$� ��.��dʱ��#��$��I����G�Z�j�ʪڪJ1]��p�[m)Wr1��~$iS�f��ܫ�^�M�c�	D6�D�G���=�2׵?�
{��4�#_gE�[�I�eׄ�]UbO�8>	9BbwwWKK�FS�T���ʸNǅ�8�y�k������خK�[�>�IAx�����r5RC�8M��k�O��Q(�/�x��E�x��>��ډ}��
b����������f/�V�D�LjLyޟ9f�^񟶋�v����_#o���\�@��?��r}�bx���Z��}���"��zb8;��Epf�ёl�����=�q�2˩�������T�RR����3{����p��)�9i�~��|�u>��:S�~�X�+��q�X�q���{F��$0�gk��]c�g�ʹ>E�(Erwc�T�]Q�:/�釲�R��%����&5�`'�$�(�I���~-����ٌvW�3x�4��{��Ծ}��.�/��R�H���S4צxe>n�Z��wnɼ��GV/NR��@��������+2��N�T�R���h��K��.�r%��xH��T��	_�W��B�=�������ӰDa(�=��������v��7IMR~����
�R�x�7��b.��r�HN@�&���� &�m!�n������nC�Ѫcj)c��ư��%�Z�����3QMU5�D�s�����1+�`�.�(ˬ����n��}�jn���B	j����ҳӺ/��}�-a���eK0ՄG��t%�"��kQA�nH
e{���&�>�z������FN�U|�Z$2^��-�C��I.(X�s�-��ڌX�/#{
���$�s��Q兊��#�dW�O-س����(���4��Ym��L�.\�[�]��P��I�\viAo5]sG�wC�=fl�m�!�|p��
����;�zΨ������cV�yw����&���Vof��r��T��_E�T&����6qc��	��4��Y�t\L*�٧�(��R�'���x���6��LUT���z^��Ia����h#��&{����hc#��{e�f�~��ٌl�'E�O2ӆ����$�6ٻ�`��������� �<��/��0B�"��҇K�/���ϗ�EP��X0OP�ZD��/Kz
�s�wl��5s�Bv)J}��?3� �XKm�m�n�^*ٿ<�o�>tmt]=�w��~��t&d���U�Y���F�A��){���!�{�C�O�Q��Y�ۿ���G���@ᵽc�{� izP�F�ꃄ5S�hx0O/�{*"_�C3$�&��v��X�<�z���=)a".t��{j2�� �OD����ȑ��"�ې�
(�%�l����HL�WJi�6�fO��\<�C����a�݌.�SrX3%�y3%ǚ����~*Kn�"�y���#T'���=�r��5�9�[̸����5#�y����`�~��֨$]��D
�Q�lpfы$�	0�r���������5O�³��$æ�A����d
�J"5�ZNs��\	@� �����?�&ڈ�M��[��s}m��f6f��yʼ^�=�I�*����߇R�<s�uw����y�t�HY%�"���H����^�������-��La��U��>�F�$�|`����..��� ����U,U,���J��7P���!�|6����:�x�^m��E��%��ن@�&~�/pAMHn�Rq��o�@B�
�bt�97�����oi4��,�Ď� ��r���*�������x|�<B�c�y�)��	�A��M~�'ׯ˖��7,�)����fJ{'c�{4��!^MC�=QP9ۿ��2q1�G��1�^)9�G��0X ^~6tZ�w���
�C�����5���7^��|Y�t��o�n݄�T�i�sO��d�ӕ�a�O�S�N��ɏ�2�Z���D�ȫ@w ��Y��ɞ�����A���UBN�:��0҄�.���q��_ab��,�`SK�����7U�_�-dx�B��X��ߪ���U ���Ɓ���Z��6���A⁄&A1�#�(�?p�b۳��4d��i\>ͅ�%j�t�b��6OP�2��qbN��C��/ԥ��B����W�t@�?��.�5/U[��il�Y�s!=3�- "���F�s�*�	�+�f��C�1��R��M�H���jg,��O����Q:֎w� ��_�7m�1����"��Ϊs畷��d���7Q纪�K�0^������+�]�}�����%��>�(����J=��mݢ�[�c���g�kb���������������՘��]S՗)u� �T>�:�.�t�ǀ��\N�>l�=��blZ�!قX_�wX����H��38������lD�7'��}s���T�{1����;9ꢨ��1���3Ţ^�+zN�5�1`D2�M�`⥣gˣ�6~�#0R'�omm�q�a�ǥ�b�?��J�=�Jp�h�Q��E�p0� ��$�M��kI���a����D��}���i�o��=���Ǩ�MK��F\zI&�|ȝ,i𠎿 �tE��N����"̆G7���.��/�.��}�[��0D{�����#~MH��$�Fd�ɭA{����OD=�xR&��i�n&��n�W�%T��F���%����G2�(T��1`�kA�����'S�#����`+D�>��)�Z|����~��!���NS���=��ܛU~e�E�s���C�����\�����_������U0�^��'��A�E�	`�I�r��2��uL�D�ĵt�uyRt��9?[Q���u���u���9�S�Ugp�y|p��䧞���.�N�M��e7�w�t_���/���ֹ�U����=D��� u��6�i^�9�d y\Þkf�59��ϡC��Ȋ���M�3f�%΁���\�i2BxѾ��S�w]�
�=3 )iq:f�
�H;���x�n'_F/82�8D�tH��ZƘ�Egb*1C�����z�vs�e~��IC�m�P��[t���DLv���=�k���늰���xC�=�m��Eۼ�3�W{-	���U�h��m�m�=��12�YR�{fa��Ʋ�_t#�-Q���S��!��K�%����V@�����K�̮'��=��4�;���V�:�+�1�Y%�~E[��h[!�g���cU�p������ITO�<>*.���Ч���x��u�䝕,zB���R/�>wjWu�2�'j��d9j>E�+����
�D0�z_�eB3�7O��;������R7�	�1���_���GMހ⛵n��A�1���録f�z���Ra����Lݾߪg�0Cr����D��VT�f�"�'�Gf&-Ю�ш��"�B�K ��O�3���r���e�ҥ��1���7���ּz���i�\���΍�l�q�J5�Q���ň�2�K��-�33����aә 0:�+��x�m��������rf�5o��CO̕3�'{1���-��1����,.);��7Oa�EJ���LU�z��m���������i:˧ �SB�ο�QU���3I�Uuz�eݜ~������'��*�٪��q��e�}�.���%\���(��OAV�㋑�k�����W:G	�4:�?e����,���_�~�G$ �y�D�e��L,�(���*v����=�g>����sh��<h�/�L��M^��^�z�.;J�N�=)�SN�.A[I]��\�a��`���'V��dA��h���;��h"�~�)sƇ�k�?�w��n;प[E(��6� Wόtiר3�s��F��"�q#z�͔�����ʐ�f�q?/��~��Ԯ��'�QUcm��0
��؎����dV�?]kk��_�����a�轙Z,l�(�2�ތvtWJ8}�m����_Z"Vh�����ہ���x�
�/��k�\?���ÿ���O�J�kԂ��̾Ź�潢��؝��Q2������ٛ*
��s�0�I�BܢwޟH��ΌH	]-]+^2233Ћ�}�F�o6�w�l������ʓ�ഒ�iBx�^"G�
xdQ���SI��n&$n	&��#_��*�ӊ�[M�ǪI-}N�N�z���s�>��L���g��S�`�al�SqJo&=�n�^���g ���a"��.<1�����@����ID$pq�z��f_�Ҷt�z�z�8���&��ی~���YF����U�BE�q�j�H���ƫcK�T5В�Ad��u�k�"�����_k&.�͆�.5�\^�sR:�3o���P����������~�^�1`)��"j����RZ�Z��WЍ��u�P�j�dO󸊨~O�>�����X'�ǹ,\�I��/g��nTֆ�E(�R"�XD����#鑋�Βc%T#ړ��j�	I�Ҵ`��ǁ��6�y��~<p��-��"j�����$�����k[�h��68������x�
��-Uf />�����w6���*?�)j���?
\�8�����=L���l֠z7�6�̵�E$��1��{���}[��3����~t�>��8wdk���xب���1��C����r�ǰ�I^S��:H�Q�0Ϻ^��%�P�����Cd���.��?%�@(y�`P�sZ�p�����$�v<��5��M�Dӌ����Q�L ��<%��ևsT\����d8�e�$AH�D�p*}}�@�B������QK:��z�����,;�;�c���Ѱ�BkvC��nU�&݌F�X4�8 X�qpɬ��^
�\���O�	1uFH�x�Ǡ��]��7;��k�<"9�T�4 o^_�����sNT;��0}Ǿ�YB~�fJc*h�	t�|۹f`��-�4�<J��5v��1�X�������|"r���'$�
�i�F�c�p�b�[���R�*`���}��ח�K��.�f��`,t��]=,2���čS�剋G1C�L̚O�*_ц�p.5(�P�|���D�aIm�v�r5A�줐����ȁ�BuV���
9Z�d���;�e��$�eeU��ёD!V�v<��Z ��b��hou�klz�zW��F����N
�W��B�B9=ɜj�'����A��z1���6c>���޻�	��{hH�����&�e���H<�;�S��,�O O���v��}�
f��zN8�x����9�w���Q8)��/`U��U��)��� �}��?ӕV�ӣ����w��cA@ͅ���nH��yj]�OG���EF�M�s�����AM��N��,RY�`�`�g6�2�0oS����kr�qY��V0|+��^ۈ������MH��3���>e:�ETDb��6xR����͘��M�o-/V�}�ǹ�2|dv�ŭfK/rJ��*5~
3`��0��Y�Y���k��ٿ�Ф%B�d�:U�d�$��Y��o��7v#8>M��*��/+3�H�&#n�!���Y�$3E�ԂSW�}���e�U9ϝ������5m� /��|�Dlo�&�<x�U��m����P�Դ �\�5�9��?i��H�2c�5�_ȼI�F�&c�,-���( <����\�]� �Pb�T!"�}��ƞ���4�J��D���@��4�dG�&�����%����ܦ���Pq�sDd�-94\q��$���d�3j(�!���=6� A�Bc$��4=�i��hb�[��N�?�W ~�Y&��͙�h�m���C�)҅ ��Z\�T�7�-0�D�~$���S��1��ۧ}1��N�T�h��Si�$-��$j��䲐����lb	���fJ!Xhs��"T���g#��=��E�?|tH���8��D䝭8�I�C{����|��a��)ȳ�̴�ϊ��O�	x�;(��1L{Ȭ��z�w�/��"Ve�E��,y0Cg�I����#l��|�ӽp%�΢iZ�俗q¶��5�*�(�rPop�ٺ������T�~2\��F��1��-)��*��FK�C~b{�ň<��®2dƥYz�[�0��=N�Z�f�gXd�[e�c���¥�;Ǜ�������rz�Ĥ�W{&/ d��.�������{^:�n~S�1l������ |���9��>�}��pB�2�z������^����D�	���YIٝ��yzw�Y�ɻ�����qO�_��-���𧡒RC�	�m�:g�� z��y�:t�j�:�ʌ�&�Bez�/�8p[��4�`+N��k��J�L�BE:s)闂}��"d��;�����}Z��	��ɰ�D�;sm��;2�7+R�͇gf����`)�">Z.�nubG�faל�|`��G;�c(Q��F�A^�M�1ͩ�Q�B5J��ώ�M�؛X� u��a��S7e&�=/	�a�� ��8aI�u���jX�B[�?~82���><�,��_a�F'�csHUb��a))�ke|`.�(�r���=�2��g6�y^�ػLMD�!�E{��_���^��f�
Td�.h<��"��
�!	g1���~�"��}�]לْ�|X���dQwV�U��ЄD���欻Nҧ��S�_�-S��7���y,�#m(T#Ty�>�����GWl*Uh���č�h��ى��V����dNߢ_�_>G�&;��-�3�&ӍU����?��*^��s��K�2�T'Oo��{�so����a]��j��`�d�����:�~��`��)]ޗ�Y_iO^�WTh�V�Yռ�$�h�Y|Ȝ*��ה�O��j�K��n؏�����
1ʂ�d�T9{ϣmU�}��t2��\���g�*�M{Z)��]�����Ejv/�˻�V?B�a�e�Ԡ�� {W�BrAS�r�.�8����E��nƕ Jݍ�G~@��
8����l+	_��6� �S�
���f�*
��2�q5ɿ>M���n<��2Yq~~��x}�������ˤ�k�QDOg?�Iz>�i��%�� '�h���S�h-wTf�<�0�ǣ�,�zߴ��w|�<����v��Q��(%�<}cFxpT��L�����}yL����)a3kڕm���gK�LpR6���!q�˝	�|��}�����bmZ���`xN�	�J~G�[�)p����/���k��"�~����-��;n�2b�9���.�C�0Y7�:&��k!K�Ǌ���n�X�|���Ǉ�8�b�|L2��[�I!F�;���_��9�gJ�*	��qrdЈ�No\}�7*�H�돧�T&g͚�ZVݏR�����$ăDwz7�"3̳�X�	m��	ġ*���������QU�(�|HN\�gC�'F�=n�{m��Z��'m��TD�U��O$��|��	�:���m��4������*z�r�e�pt�L���E� ����o��xu���V�f�L�Y�;M�	����v��%��hAΩJ�����
����j���I� {�{-���4#�����ސ�����م�k���ʳ
"�=��p'lq�i A��4(HVl��;Bj͌
	��P��=g6i!�(+��``��e�K3=��nz��e�v�t�B�?C� u�۳��t�w�������4I�sH�N�fd�l��ڌ?�V�����>�7��d�?��/�w9�W���I�<0��jxd�<���$����%�m�g���7����C�R鎂p<>�ޑ�m��MV��p���~�#c{���Ujc���zUJ,�<��~ȗ >l���`L��:6�$2ěf 1��S��;5[
�jo�zO�k��g���A�T�Hmĝ5n��B�kl2��)DF��[�l��^k�[�/�@q�w{�,$��w��ó���vy�7*y>�[xM����]CB=ϣuA�7�O�=mOYW�LHDWl���^M������n0�L���Z׮7���[ޗ[�z��Hv1i~�ɒ�F�aj�'�{���?��c�����az�5�M����?�>V�ӄ5my�:�!j���gD�C� K)t(&�,�AF����.(��ڙ��˖C`���W�}\O��kT�,�q����5Y�z��pV����V����e��ox�ާ1�.�"p %�[�u�%1F�Ӧѩ*�� *IA�7�VIG�O���GU��ف�G�R�d����c��xeF]�f��]�����u�������ߤ�������ң�ĺ�k.(�4��#.Ӌf�k���G�K�L�=2��q���o;J�7p��B5���}�i�Y���н�s�P�C�,��I���uvZ�*�0�M�=q�������W�����7YE��Oߗ!��*4�����!�����R�c�f�Z5�Ŋ�]۴��T��bd����}1+ԏ�I0���y����I�@��.z�xO��}�kDޫ@�5����k�Y�_Bd�������+��������^�p4����e�mgB��v35��-NBN�y|��Q���+;�����f��"���{�bEKu�8��$=jS<T":s>�	�{R*�G/z�X$��D� �����DҜ����Lߊ����߈�T_��M4��-��/v���!\�:��t�0����P���SOA��ڴ1�|�<y'~R�����M{��m"؄���jBd9��kg+� yj�!6���I��T4� Stuc<
y�HV<AΠ���[��[�GW��|��[o�,��^�N��T
l6,��+�O�9v/�-KC��T0��'�l��%~�ag"�J��.������crj�)�9GU@s)�v�KVb])���2�=j��VD	�v�!% �Cc�9g� ,e�ߍ��<y��b��'#�����}^�Q���Kj��D��<��Ƿ��S��>��.�>@�|��oh�J꽁ϭe����˅��"&��Z�E>=W՝λ�h�r������j	���������S8��&Ҫ+k{�r/[��+:�Y�|=��Q���@}�ʏI|�L�N��uZr(Xu$0ݝ��������t4_(�1����q<��,�+��xm��Q$�!:'���XY��$ތ\���+�ج.w`�q׫ٚڰ���"��q.�#O�E�{d:<�ͭ�D��f�ǩn�/?ۑ����se1� ����C�t�q3\�h��y��G�:[t�K��J>�)rq3�+H��!���٧��~*������1<�wy̜WJ�B�Wk�	H���}�]z6o�{�xY���v�8lr�Yn�\SPj��ب��O��"���X�+�����{��[NDM�����}m
���!A��?��>.ID�ҏz,����HEF����2W��֣�OZ�rc���q�;��a.s�2�#N�����vT�[�k���5
������Kj�PZq!zf�N�*t�P�A�x��`�7sgQdw��8�?z���)��Q?�QeYJ��L�t-��4� P5ʄ�hj��"�f�S?�U�+�f�8#u�o<�Ռ1�Y��XxȘ
��U��I͌C�o��g�c���[x�/����R�+"�+y���N�l�L��|�$&̴�Ṫ�VfS��Kll��D��L�-�|�m�ii} �z�~�48g[��|ҚHk^Z)�tFV��m���D�I��ga��ȧ�iʼލ"e���hk�pP�x������� �#�!l諻���40�0HF��j�?Vb,�9Qd��=v�.-��N��)b�Ɍ�t�*jf��a�W�+r��2�AOX�J�iF�/�um֤욈�\�k�sȵn�{FJ�g�p�$!t�?�ţ��Mkl?��e`9ӡ�&V��Wh)��@'���e��]�_���m'��G/�s�������r�o���}_oد����}K�����Y ��.�ICV��o��'e�5M->�;��8��*�|r��1#@����K4$��V`���"
)ct�`!��pF]�kW-7��a�'�A۞?��V�=�����	7�W!Jj�L�|@�F��"NИ6�.�S^|��N�n��U���QngWPi���6Q�Y� 'Ǹ3`XB���5#<��'�$~6%�/,�����5�ت��P�a]��1ϐ�_X��ҽb�=��ݑ�m�'���5�Y�*^��6گ}�m�����=����-�+�Ce�E�ڔ��_ﻈ^��V�Т�k����A^M����]]��G�ήo������Ŗsõ����V�0�s�e*��z	]�~2�x~~}Z�_^S	~rٸm5~9B�����xa�f���$e3��ƴ��Ac�K�$��x�~��2��s�f�4��m�݂��:���ޡ�'g��4c9�����& ���[����8��~�I3Ǣh~Nê��20�9��q���}�"�u�<�N�|}���rK�#E�tq���{d�?�% �T[�&)��3w����y�a8+@�MJ���.��� ���c��o�>��q�)��\*uL#�W:�ו����
L��2C*��<1b�k��s�.�P���m�����&ҀX�敇�1��c��gx�lH��ċ�kvm|�J>{��m�]�
�{��a��̱Ya�����$�o cѼ#8g��}�O�8�i:l�x�
}l|��wD�<�o�}�Y 
�����+E���H&Y|���J�&��z����a��p杩</��U7�c�y�~ޅ�A<��c��_�ָ��b��ӻs�}�4G����͉�Oj�3���7�b��f�}��?E�&3�C>�	k��)n&c����� �j8$IR�Fꀝ�J�~�,)e7�dMj�*<�ƙ�&�Ue)�:�<��~gD�!��L%@�v1��+!�;^�`��OG Fƚm��L�6U�O�&�1�SAa9Z�bIR�z�2�_g�.h������\ދ�����n��5�#aC�����-�����|����%��]�ʲ
��8<);�+.�k���g�Ԥ�W�
$w5�iv;����("���$�fy�j���r�����kn��~���Pl[�^�K��<�z��r��Hn��<��.�O���AӓnE�Ћy������`��K뫻o9�7��A����Ë�ߨBWJO��Ju��~f��/�Gr»��o�r�P4�5k�}��5@'	�&l��ㅮ�����5XJ\�3���UF�]w��ϫ�?W��״��e�Iۊ����̋�}���Hb0� �&�
�S�%i�h���ނ�4১�Ly+���M��f�6���l�aj�~�OtF6d�n�@��Hе�w9J>�qT�g~vg*c�p
pI�<�As���N҄-��Em�4�"�
���tR��]`�ɝ�V�Ul4n�.9��{�����a����U�E�h����fQW�k�'4��iI�6�ڨ�s�A25c��+���!�Ӻ�@��^��Ӣ ur�	�����jS%�R�y��������rl|Ϭ>r��!E��j�����Z�C9Ǖ��ةʓQ	_�@�B\����4{٧�^�˔J���s�������]�
��r�)��a��< �i��ڄ?��r0�*Z9�&F�3���Re��կ8���{��Iw��s!���W�AT>�8T�:H���F�q%�1�{Q��(���č͌���8 ݁2��x��á��K�*b$И� �ɶ`n�-Д�`�O�JVm?U�N�짙�+ 
V9t%}�ˍ�;,��U)>V�K�5���p4~rc���.R�<f�/���uÙ����<�b�p����,N�l����"r��ט�aa�`��LX����Y!�:d"B��X�ѣR�����}}��9��.�����H,��p�R�on��%U"�yu-��3遧o�\h���eW8�Q�P����;���e�$t�Wβ�W纝�yS؂ ��smS�K��DH���-3�0r��G1;r�rۮ��	v�hCD�c�vY fk&�D#IDa\�5�8��{�=x�(6c-=�"���ܦWSe�Wh��.�ApL�ެ)���V��p�6���e{�KƖ�
�RyV�"+I��P����5璥5E} �˟�w�j���Dgbe�`b���+��
��7��N=�.�����E�W?����!� �!�;`28��־`���u�RNJM��{�.��bi�`�S��SykZ��b�Xs3����6#_H���'�-��z1ܪڻ=�VnO!�O$����}��	>���>�IW�Z�1	�k�>c�(�o���p�p,)K�PRv� �(�(���B<
�y�����k<Sk�u	!E�rt�c��Q��Q��)�y�����Cf
{4�Ҁ.������h����%s�&�� ���c4i���IL��iܢ�@h8�� u���8�������b�[�~G�ޑ+�qq�
��껎`�N�1��	����� ��ijf�1"䪒v���ߐ?���S	��8'�D�c�C̾�LpE��<��k3愱]��v�V�E�| ����o�C�l���T~.U��4n9��X���D�ȈdY���*Q{�PP�B�O���n�͏ޅ|����Q�W���D�C8KQ��aKM#��'��:��~e�!p���L��T��YaK��a�ͯK�1�L�S���N����P�w����>���f��V<ڰb�U�mT��.����OR$l�� p���@�;����*��8�ʊg�12zp�Q������Da!�`�>!��7$=�ަ0�ck)�$.N��{i�
t-87R&�W$h��Q�zRN{���~�
��1d�4;X���#:}�sd5�KQ�^Y��sD$���ޯ�KlX�4*~�E�~�����_�8iOM�j�;c��%ޣx�}�a�>�T�WJ�W��z�"�Mw��M��2�	w�%32~�?��J�.�0�L@��&9�ojt��92xҰ��l��W�y31����8>}��&�}N�R�rK�>��o#��N�^@�E;�;A[�d�O�	~.qb���2�O4/���ͣ���n�����B�^O�<��.���5^"K�����)��;�G/<ܣ����AA�d\q|�6Bk��G���ktj�׌j�������oi��|��"aj%Z��j�M�+oq��IE�\��q��^�õ�?F��<^��"���Z�_�xI(������I�'����U]Am��l���lF�;��r ��� �qQZ�*�o@w�{c����"�4h"��ů��)�����c���2���'t��ۏw���jw������Xk�4��ViyP� �:�ͣ���qWl�p��PbT�7a^�bq��0C��~�0��8��O�d���J��c��X��&,�?O0w�o5�7Lh`���#w/E�W�}��Ұ��k(�ad�a�%�j=+�*/�������s/{
�섴�������ye�&�-r��z*���C��@cdH���0*���?�}���Oށ��I���)n�< ���à�Ɖ\�X�\�;����/SFԙ��!��I��W���S�
�R�/P-Օ��?��*���>�����	�5i��=�Z��O�~�ݺ�0��������q�m��P9��FS��n^h�K�F�^�/�n��1�=w��������/"�/��p�T,jH�l�=���4۴�I�Z���G�Ӄ,�*�aIH�����	���ɜ����^Pb��E	��ڏ-B��+��v�qZ9 ���Py���B���c�펄��³:nE��e�� N��*�ƚ�]��^����G��f~z�š����(I2>��S�lX��.dw���8s��~R�2��\��L�$�Mг"���b��~0 ޽P�K�.ǅ7N�����㒙�Gt�v=�y�� �h�v3J�`:��S;�)��YS��K79�#�
�7������؁t���l/`��"�动�ZT�+]>Go�!�O�Ǌ���o����g����0��B��B��<ܾ|��w��՚��Z��z�P�<�e���&��¯�����|ҵ1<k�����}y��X\836���3=~i�z�BXX��u�@�!�=S���w^����篡?�{�m���<ﻼ���P��foކ�'ؽ`� o� -����!V.I�?�W����jp'��E����?��k]�"�h�]�Jm\�*ǖ��N��DH�j �ɇ�Rm�"��hR3j���a#���O'.�hJ� M��f+a�J&E�#PՉ�bY"uoe��>p��fT���? Z��hLaT 7bɐ�(We�Ʒ�ˠ*6�)��c-�~���X�T��8����x	�C�\x�u�>������N �����>��;�<�<L�|���h�u��uR\H�m:���|w���f�ͅOe���Dy)��eޭ�g�!m$�Wo}hIw��=�̬~�`����l�T�	�9������if�D.�Xw-��;ʨ{�N�/;�4�-��Ҹi4虥�d��i�5E�$�.��FEq�JC�R����C��js 8�H�I��(�hxa�P���
E�	"t���R!o�
��&FF��$���3��d��'�+�����#q4"�ժ[�t/�Bȿ���n�1�P�d��9�?�=�D�"�9J��-�x�SB�$�΁M��A�;T�
v<",���P���(����t��~@>"�� +�\�U#_�%R��1@�=���;1��p����g�N�m����xknϯ*�͡�7?\��뻸d�,9��*���������8�=���H7�1t���ݡ�� �В!"�t�Э�t�����~���Y箳�����g�/���]��g��)N�G)���~��'Í��?U��ag�Ma=��]u7M�<f4!�n�ێ���P
Ġ�;۪2�
w]�R��ogﯳ�
�ҸN��C�.�ƃ��5��}��/q�|�bv�c������6��u?�n�S�!����<��'4գi���{�}?X�S��)�mE����(l�5�z��R2!�)i�|�n$s���G{M>��,wí��O���T1<4�\ok���P^��v�Ѷ��X8�k�6�]5�rl�u�ڶ���$����t���<%�п*��V���	�����Z�?�Ѩ{*֓�e��A�0�#��Ty~���g����x���d�B%����E�Z/ ĶD���#�(N�L�2xI��	��<k�݌�i�tڝ��^Qڔ��V�%�k*%F��TR���⭡�0��2�ɗ�1M�_��y�ۨ�W�p�ͤ@/���C)p@{S̉���FG�r�����"���/s�"�k�5��g���9=l{o��
f�K��E����fŜ{۴���Y������]S���,�ݟ�E?�����2}%`����M��4��`(�
�
��G|��򥈈����8� ��e_X��[�f=� �s7k�:�7Y�P<�݂GE#��U����Dd��7�-RP{��y�j�w踧���L����$�|��}����|V��=��hW"��`���#WR�4����x�-1ő��|Ң+G#�t¢`,5n<�
��
�������!�%�c���Ug����,x@@�ҫ�L��e�j�x,������|������ �Z�/���pD��$�2d���+;֯���1T�!#�]P&�k���z6���m��nk�bW8����h��r''�Hn�Cspx~Q8�,��AX� �	. ~�Ҧ��[�c��b�zqc��Ւ��1�����%��w渺��%�Xj������?l�i�u���0~Y1A��3�!�Qo��w����?CcX�e�{��N��e*��:�����&75��%��Ǒxϡ
y�?Y�I�Ju=�m��3~v��)���g��
_�� ���y��R���j���k�O_�D�WQ2W	��>����;���"o�=���A��zB�.(���KL��U/!�T����L�R8��h/R."'sG��g}B����Er{1�f~'9WA[!�,��~�u(KI����ԏ�n[:9�(*N������%&�e{��6 �]��}	�Jeu%̤Qh��w��[
IXsw+��5���$#��1=��Be�S�L���������MN��RZ9��2�M�o)e��A6��J'��v�˿�gj��3���,ǄAx�!i��.g ��؇̻M� :�h�jU�����q�n�A*�{��A�"��H�aY�y�IWm.G�rXT&y�_I��������$���lL�@15�i�n�a��˹��Fp�g~I�x�:�}V�	a7�Κ!��"
����������)�څ���s��^��N�):�lɳ��1�j�u�JWӈzJ����;6�Wi��Qp\�k3y9�ex�Jx��l��5���}�?��H��x�1n��}�0ّ��5��ŜG��?��m�c;C Q0R0�4zl/�=���?��/k��gk���d�4��Bx��dP�N��,����ӫ9�NzU��'p쐰��	��p�Csb։7n ���a�������ۯݼ�`"��cE�禥�����r��c���rINR2
*�Zf{2�c6����	�"���ā�aH����0o0ax��$'��6f��Ǟ��.rtp��Y�\��?����\�{��op<r}?X%�����p��J~�)-�A��,��D:t���EEx�z�=���,�s~��v��9����]�̼]W�(׉P�SB�j{��F-mZ���Kb؝ŎN�U�T��JLdOS�Z ���"��icc��%T��-��~Ou�\M�e��Z<�;,T(���ע���y���uz4.��Eؙ�\L.2�">��]=.�����Ȣl����>�J߭d3u���7�=dʉ�?.m2�"�3�����8<�H%��f�����ʛ�k;�U��7�*����!?�!ı��!G��4��Ml�#X¶$�������^\�d$H�MiX���.i�a��9ؠl��N�>a� �Y��7��CJ����5�@�\�C�GK�<��l �$�\_�����԰��d�'~%���_}m���"a��m�����nE�/���()���5jgJ�*--u�Qȷ�� � F	3N��U�Ő�j��j��Z��C�Zjqx|��[�=N�k!~g���%ȇnҼ�,-��nq"��2@��9&���CEᖡ7����Ueu�����v�e�%��oLu����:��U�v���q�����bY�9�-�ņ�
{,+�1����i�n��{,��ʳt&���*�lBF,�#%A4|.&���Z7�����ggl��rc�X ��Q5�j����g.��6�.ޭi����J���y�#�a:)qR���-�|�7� ����u��,lPR�?,��@h`�M��z�+߱Z͙&�Q*�V�l�Q>�V-�Eo�&l�z��*�`�s{�eKܷ��l-+�n��E���zz���m�{�Y�P;��X:Vq-���
���C�Egx��GY�q}E�~����D8=�7(��'Sɣ������Gj�X��4���t_�
�[�6>�j�� 	��������Qo����N�]_o������3����uz�q��	�Y1;���C{�ڈP��@�G�_�Z��]<A@��c�'/�D���ԱmO��U:4�$jGg>(��DQx'8~�d�3T���F��~���
��^�
7�_��-�@�R��WO�jB/�÷����yn�P������0q�vd̪�[l�v��Y*G�B<,����atz�ben>uQ�����=~U=N���\hw�oɒ��˱zv�T*��j��ve=��Y�`�$�:�������q�;R2�B�a/-	��t�����ۮ�+z=O�U��oFο�e�=��g��*�`3��w�9�='�:��`��M�B&sT�&\s�x�1^�)�L��}�t.:�S����3MT�(5u?P]r���ڰh��[)�V#����K�T4��m��.�66��d��mc%����OcT���J8��F��2őV�Y��X�ݖ���D�V�WT�DȭF����^�!*�rt�r4P�㤅#��}�9�<�\�d �{x�{��;%�ғ���������M��*����.Q�;W�b6[ӨHu���L�^�������n��K�\�j&��릕Ǵ"��`�j����O0�S�ށ��]�m�íy���"{v�r�СI#I�<����4m�,и ���ߑ�����:�BqC�~�?2��`����O�<�/��î��RN���O����GF
���yC/CC,̍֩5]�u�Z:�|m�4�+-�5�2u�u��i�x^.�͉�u��u��(+���5�1V�L�&������!�qptH>��%��M�\�n��|��|��A[ꌲ����餬"�{�S���3����}����.C�]��֙�t_�JZ��Yw�K�/9r��L����2N�0t�'��#�&a�/���7��)A���:���E?�f��fG�*��`�Rd�p(	� ;�*���?g>��f:R�=�c�=G����qt���:z8c	����Tޤ��bF�A��+-��¼6'+��.��
ʥ7o���.�H�/&j4�St�)+a�&�#;8l��Z�	4����p� ���z��۰MrQ��PϦ�W0�g�ҞB�P6��~�ο�u/j&�(A��[��V�.
BwV��<2o,�0��K���'j�*o�5�\i��M�@rv��J�V�t�;-�����D2`�����,u�O�#+�X'bm��E�Ãfx�M���FS!�?'���?��S���>�!��|j�	�_W����w�e�N����A���]��&I)��AA�*��H$�0`q��8����D����Ya��ʸ�Q���`-��)Ǜ��7���UfOwd7�!_�%��i*�o(�����8d��xsY߇)�Z�۹���r\����|o��ϻ=�ϩm?�/���f���#��A:(�gF紺�����kc�Dv����$��!V��0�P����Jk�*�jZ%�ր(4�����`��WVo����p'��DH_��Z�(�&�C0ۨ�cf�ݼ���:q�L��ɀ��Z+p��}&v%k��UY�-q�
F��l���-2̞�F�aU�2=���T�(Ls��xT�}��n��5_���}�o��G�$�c�3�F%�!w�y|R�@�t	:^��_E�D�j�B ���5��;vu���]���=u���<`4�c���dt���_bJ��?�'O�j�^�kJ=��ο����W0�\�������uL��Y/�<���CW7A�ID��uc�tan!*�x�Ϸ߳�4��M��,���_�Rn�G�}F�IaHͿ}��]M����cϐ�6uv���A®-��b��!����gESK�5`�&�7��w��RQZy-!Z��=���ٔ"M�E�'w�4�Ƃ?&q�p�Ù{`�J��R���8���U����5���㸮.��|�郆��Ғi�jR��q&�<�C��*i��]�[���*�����q�a� ���ٽ�� ����̠�?@e�u\���z�س��ɼ�|���K�g ƿ�F!�ɼ���S�`t��SA��#"ut�(���������jf�)a"Z�GB#�1^��`�,�=���w�e��NN+K%:T��Nv�ۊ��,;U
�L��1��f.mdXi5Gw�Q��c��HȱH�	��ȪJ�����'�m�N0쓪�
̜	Ū�D�ؠ���K�qjĔ;-�h�걦��ܱA�p<Tj��5~����4Z_V�R���e�Nb�=��U������ ��o9�ԩJQ�FS��s<v|?{��$M��[��-������H0��g�b�A� �7�0�d�!'H%{�������d5���C$�]�S֞��,����m�Ra~��.Z&2[d�0Ӻ�p@7��N�/�+�tv$��
�o�D�Td�>�P&� *6s�s,6���C�����%H���Ɯ��<��(��Z�3ffSl$�`�䩛���qnv=�b��b�����z��T��?NA0*U\'�)O��ākx���Ѧ*��r��پ��"�('�Y�,���פ�+�B�+����Y8��W����k����?si?��T��P^4����/��xY��y�3�3w��������%y�g�D;�4���g S��%|-ǒ*���<��сY�[�n|���C��]b�^�	�1Y-,m�$�!�h��dv��&�ǊP�3੯�dF+��P&���6E�\��-gTw�� t���,�I� ��{�G��J{��_���4��o�ֵ��Z?�ziz{+=னꧪ�f�ji0#m��L�>����ld͵��mK��� �Q%�Zeƣ~���̑9~� �����׏!S�6���g���E���MAM��0Tф1�S1�!Z��b&/`�S�Z��?�q��h����f�zy�3������Ԕ�i�$��4.A�}�����,U�#��8�
{���{��/���$�cFdk�yt$����*����tX,Mx���5>s�-Z[w���\��r�,	)	��ܫ�!��Mk��c���H������U����Ԫ�|�\~���U�T�y$��;q
� |\��f���-@�Z&��X6e�5����7�/��W��.�E��&}3FĆKh����e?Ac[yؑ�|e#�0UE�ɟuD�W��F[���EX	���K����b�Zڦ��uᘡ�lH�Y/ղ.�x��\J���!><������b��$�m�4Bs<�8qs�}m��\�� g�锛A��A3E8D����,/}(�d��0��Nt���1�X�03��5c]��zFp�<'�!����v �M�mT�N�O~O�*�M�� �o�=�I�g��Y;=rҀ�О_�6��-_4R층8�)uF��᷂����g
���ށl�d�a�go�M���^Z�W8�N�F2�[�%��ؘ�|0ٛ����9XU�=�����\�uDs��&���蘌���{�)f_� ޼��Z�Sk���u�Mz�	���/��!��R�gc����}^�O����7$�"�1���x�zs'O��'O��nO�!�����X�d��(�%��x�闞�MWGD���Z�z3�T^Cy����AeC���8T�sYov��?������~��6i�l`o94�+sZ�e�}�����[Tb��yLo�� �D���ٷ�IIҁ�N�����Zҝ&Z	H&�)�|"SzFJ y� �GL�^���g�����j�p�)��gM���.O:8M����d F��ѩ��uެ��U);R��T��������MH�������ih�?>��7>09�ǝϊ��zv�ųK0�U��J}�t�it Lٯ
�t&�;䙖��3��`x���#	��
�gu�v�����HʠZE�Up� ����p�lr.���Ehs�7�,Y�dz�˳H���N����\~�(��.�N���(S�|�e1ƔU�=J0[�<���0 hZ)���/O��
�H��;�6_�HiT��`�M&+<�ٳ>�����mO埱��M���I�3̙��g�D�l���K'�H 0��H�|u�.4q:�=I����ě9�Cghl`�$���D S��,,"��eL���3K�L9�{�s��hp��غ`&�ے4u�s�ϟ��)EM*����)��JƼg�{$��],�+'��棎4V��&�#6�4c	�^�T����w�v�w�3�AoR�'�{W|�Y�K�'��n�v!�oMZwWb]O�;�o��h��ѻn���%�	�� V�r�KW�U��L�uq��s���}���P��9�����>9-�	9G�+�����ߡ�c���Z����q�#��W��{M
ط��������4���?Y>����Y?����`?:$#�S���� ��ĥ9��qd�װ��5���������2&ؚ�!����"^���ޢ¬��*V��p �ʿ��"x?�; �0Y8�����Ȏ
�J}#���ޯ�[���QV*�Ƿ �X]Yԝ�1���)��6��1�c���O5i)Y�J�k�I������a��[V�^��Z�ؾCzeǏ��F�_���'��\��J<M����JcZ�������D�XM���JI�z9MU�{n6��#z�F��_��z�m����y�ŝ���j4���C쫙��
0�E
L�����܄��#~�AZ���vbbb99o������j�&�ݡ=��ykV�� ��^=�9]''�ؔc�sۤ�(��(s��N�)
��Ό��Yy�oH	���LQ�+���_���6��#�����L]��E� ��k4��9o�VS�g�Vi�G�S�WaKپan����!��^���@0�*X��}�6_ �Z<�U����J7_��S�R�U_;}V�b�FĦ��Ÿ`G�A5Jz�������M�\�u����HbK��/x��]��_��L�?޼��R�oST�G��2�]�p���Qpm%��&>��|���`�6�2���Y��~ʒ�9AH0Vx̳ص��ǀ:�Uj�>&Z�����tQ꘴}�1�"mNϽ�ms�/��&p@��'�>a���e�+�*���w����F	�(mz��iX�H��%�_�A4�7߭������6��]����Bs�,gD��<���U��:��ͅkw����)���1����'� �:�����M2�]HǇ׬SJ�����Gz��A�_���Q[�������x�����xj��c����|�[��xN����ǳ#�?�&��r�P��*����9��o��~>�q3v����c���av�38���s8+��,�P\���*�Hri	O�E�~����JU��!;L��B�+l�E���R���N�ebp���Y�m<��Q|d=u�y^��aS���C�	��ZK�/f�q��DdrLw�Ij!Dq~	������X�1Jlo'S�mre���l
_i��tɏs�|�f�&�F�b��3�u��?f�|Q�(eg�/�����&n,s�Ȇ�y����HH(xG?�< �{�e���N�����^ev}E�k��U��<�u�q��ahbv���|��Y�8��5}x28�Q�{����js�Y��l��
ks�i��XZ #jA���[�f��+�����U��������7F'spG�)T�N8���p��a�O������] G刕Q�"����7�-!"�v�0�{������%��	����眺���O�6R	�x�C9���I��'--Ջ};�[�y��v�pSI��Z��U�a:T�g���Q��|��R%H����QA�S��(e�_�.�Ȃ[4C�}ZI#S��gC�i
�LPQb ����
S���>ɰ	U2�������G�y�J�?S?���qoR����P�ߡ�;{�)4B��R���Lr+��p��/'خv|�'$T�`��O��dxJ�n�-�d������HC0񿥙��n�!�2L��7Ɇ���q
��w�]K���i�2���#ӳb?/�"�jG�2����k�����Qm�H��SK�W�ʱ^�>�H�»�dL1&���?ĵ�CJ3U�/�9ԙ�;*�p����pB�P�);=�8�r�Ə̫���Z�j���rZh�8��a�>�z<����j��j��'��s�8.������W.:��n7o�oj�����%o�������L�(�%���[��q���=�\�U��u��봋�o�������E�r�x3��R:U�>ܕ���XG���̸�M�����*��Ww �E�Ȯ�C�m/y���,�i�s+�~��Mt��X;>�rXM�����8���4�%ˣ�;Ү�|l8���>N���k��vw�N�����Tx�����_����IM��@��]���f�(
���q�o`�Z�141?���=XRv��#��@���!�m�W��l�<�)K\�e��zo�n?��n�E�G�0KN�f�P�q�:�{�g���DY}�Y�ux�y�՟Dԁ]�'���69�+�]y���,�,C'��e�ABnu�5zeW1r3WS���ҳ!h�a!L�O\`�'NG��s15"�ƿ`G�;�#���Q��f�χ�s��*\Y�(5X5dgiT���2�q{��_g2�<��ӣ��\(J�6��S��rQ2A����2�r*
�qa�{��CY��ZޥH+�3$jhϛ��}����t�f��-Ֆ��J>��|�W��c��８��*��2vE�����Ҋu�����0�蛇*�+�J�y���;�,x(���٥P���>:2υ.���	�i���� )nO/��۽���e�:Һ��Ov��Ljٸ9{�T�	Z�e!��",l(3��06�E-d�����y�pv�f�-՛Q���B�,���WWtf:Zz'��ե�杩f.��V�1+�t�ϳ˔��Hh�=��3Gݟ��.��D3���pV�G���5۪���5؃^��w�(�]N��枾�;+�N����PW
Yp�侘��ά�P����H�M���MDH㜐���ǽ��U�s��%�?\���[|	h\h��k��I6��)�pzHes:�]�N@�Tb����c�}Q`A-��W6�ܩL�@�Et�����?Q�Kl{����&=����2�(����+����sSd@\	>[�II m�'�n��6!��Ҍ�R����L�`}9���蹒����hi`�~,�R������b��BSz���s�?�M�-�;n�e ��/��8��Tne�I3�+��-������_2�ҷ��V	v�#oO�GS���;���6�8Z�
�em�0=��~�����` y��'ī����A��hy�|�D��D�<j��k{'�*|2�Z._x"5\sm�[�_����UмЉ��7?���c�����̪��o��50J�	|~=��J��c�C��E���ӄ������%�"�o��כ�*�o3A�SVdT�O���'O�&������{���2?P�ΰ�Z�glb�2I&����jX���}����J�W���'�,�a���X��f��\�^Av:�~�4�xp1Q=��-ƒ:��*W��u���^�9��&�~ *K��đ�R� �+�Y�[�t�f0�QwN����L�F��wy����1p�G鏯sG�'5~�B��}�mC_�)� ES��7I� ���oO��~��/�j�n����ޚ���Rm����tٰ,
qa�%���F�#�+���/H$A������� F��Z���D�e��징ǌ��x	��f0"
g��ʵ�o�ǯ;8���*�����V��!+���5Ζ�C�k����jz�g*��W����a`<��-�ـF��4{Oo�f�^a�( ����(FTkѶ��q��O�{����}R�4�2>���J��&�6�g*"}m�=����p������v9]n9�%��96��WhN��"��FH?�2�DE��(�y���M
���~[������HRC3y�\�_P	`��"�P�U����u �wO��0��\�#��]�[�j�r���`�j��8�5�x~7�d�C����~邽|^��hN.��+0������x�o�OW9뭫7cb�끮[A���;a��?��s��
��'^�|�:|�����.L\��[�,�!��@)����!@�V{�����J��ź��?^	����2��)b�l;��n�x�ys),�J�Uk�x#�P�Ú̩��T.f8!�T��r�$nu�~��F:+.+�u|Z"�w�G�~��q�8ɉ��Bͦ�gp�fE�����kpL�B��pu�\F��59�ƥל��Z�6=G��9|��n�U�y }�@n�z��ȟ+ts/����w�0~&MU�П�G���I#����\tq�_�V:7�_O�΅�w��VLĻ!mw��TY_K-A�[�6jꮬ��7��W�aw�+B
��DZA��_�3>d%&��/�3��ĩ}0)S\-x��z^���&S�*V\$�w�#	q�,U�|YE��A�XΠ���d���|�	2�^ߵ2�h,�|Lq���(1�]F��^1ea��3Y�ɞ���h��k��[�<],4�TT��d�����aG�������c����=�f�X�^��>�;j��~����q�Y`?q�h�
{Wv`�iTDn��6��U�4�H��I>��`3y�����ViS���Շ"n2i������9:{u����Dg��8�T"(�ι�e����<�=���R��L)0kp~Kq.9��Y��9��mH2�P&���b����IM�%���t���[I-Cn�a����hRX�F��M�cr����щϰ�%ȯ
��o+��]H��B�g�CR�4�UD�
����,fG�t+G'W?A�Ijԏ�jp�Vm���mK	��?�e �'5�w���ਟhF�6��3�AhΕ��xŪ��.���<p�h������NX7<� 5>�5�?��҃_����o��YY�i�{^ �>�8��]
�}����9�2�T!�^��=M�
)4j])2è�ҵSY�'��fѐjPZ�n+�y�<}n��i�d���a]�F]����4�R�!��Qi��"���6��uh4.U��ԣ��H#�\,#�_�Ģ]{ǵ�~�4��r���H�E�v��Me��R$�N-Q��� M#b�&�=ѳ��Y���21�"��ߙ_J{�"��n�@�2�ݵy��B1��&�mev�D��γ�γ�θ�N��LC� �Ԕ��+��m���1�� R���N��zM2^�nc����q��_�k׺���N�������FxB��_�yn�kܔ&��ҩ�um�0���k8qhX
��1	��K��{X��U�s�v^](ќs̑H���,ls2�����L�W ��!�T�n��ɺ��(����)�F��ק/qXB�Ct��@J>��,O:�0�V4�����c�[�`@�t�bU�:�<w�e������وw�>ˑl��P���T�����Z������^��l��/��/<L*��8��(<B�H>&�^_r�x!+!�j
~z��t�+��"�l��qxƀ���x���~�����Xa�e��/Tş���yO>'�QAh鋔{��$��2 �QDһ��x)ӏ��#�NxP�� ��)�=�����rX��÷�X~�/���?�	u$+p6@Q�"E҄+�XI7�Y�؛����o*Z�%ro�4���s�M֩����(݋T�-&��n��yY��h��6��0�'x7_����mp�ư���Jwx�1e&����>6�2����y4eb&^r�����0T��9��6S���+���(���@�ms�8��O�A]o�����Q��$pC��0zB��Wi/ʌ{�b��1M��XQu[1bme���t>8{~��t�������}���2;��[V
=�W3�@���EI���A=�8��u	=N�\�<���uPV\�]=*M�/A1��aЫ&ⵔ���f�o�3UH�̯m*���_�%Ѹ��$���y^m ������EV�����Bi��]��|���|�*ݘ{L�������(�y�� ��M<L��l�~Y������8L�9Ц�b�F�Lk+3�ת�75yCt�2�D�?�h�9�%���W׻���Px�w'7�7������?�w�x �o	��]V���rC�8�3a2<1cܸ&��(U�Ը�4o!��/84�/��L��"�sT�L��.�T�|.!�z�k�D&�� �6��S��t��!�^�ًd�$⏓.N1R͌��P�O4MPK�+w��'�DX�He�����e>�pu���	Q0���ނ���h�>���s��Z��z�B�'�Z��ܘ~	� ��JIrB�+D�N�E*ߨM+���k�ә6���t� 	]!�yA�H�u@T~���
�&.}�����5M2P ���y���i?�3�|���o�<Z��56q�O}��*F��|��]/q��!(VD�/��A��!������n��V#�Q�,)����/���"&ֱ���*���]�U�g��9�ɘ�&�Nt� ��h�v����U<��E/�	�:G��Ҫ����t_
��m���d���B��g���Ҕ���ړ�G��t8J���ۿT�7�,Ϋ��6�����_y<_�j�K�������P-��T)��[��1ͳWI��n*��y�n���h$2[��:����M;4&�N����)x����V"����+1�XFe�,T�=A�/b�f4r�쪲��{S�qJ��M>��D"~�4�,?J��mO tb4�¾'z��H��ns�s��C ����a�	�kp�&g�G-��Q{rZ�Ҍ'<�Ç%�Zf�j���M���aB�?�m�m�S��3N�x
w�
u��\"p��8	3�l��Ԅ2Ƿ��D�$c��˵���|��W�X�2�'�l����*��&#�pSU�(����o#UL��'�S� ���8ƿ����Z �:�&�V �f͎�B�#��m�4@f�XI�F���y�!���lc |�1�ΔX��<�4Y�}8��v!A�S�Hyu��{���; �R�ͨs�������k:S�i0�%��5��?�y��:
5���f�[��1����A���y�כ�����೥��Ω߇W�܏a��?��n��+P�2�����c<��i��ͽ�u���4Z���-�-w ��-Jߦf��f1�&�{	��9�
#<|��]�=�H�p�zv�[P k!��XM��LK��_�8���	#����K�����|z�в1Nlm0�yCC�l7���������`��$>yL������x�1�
�ʢ����q��I�i,���h~L��v:�2��ve�e�ŧ��a�NI�!�+��Q�ia?|���w��.���W/!)IQiF:rF��P�!h�?6}�x֦T .@�4�;�L'ZF^�e �^jF�s�7㩠:��[��b���f��� e�%v�=x!/�m5�)�x>�,��n��mٷF�˲S���/p�.i�^�_�9�@/dZ��N���i��z���}9�Ő�A��0�21g_���D�a�B��uEYh����mS��N
�~���.��@���Y�;�X�0�!C}���g�w��(N�.�� �_�J�nxl�
qJ��DH����ҋ�^�i�2cP(����� ���ʻ�����~|�Ⱦ�0%(�Fڴ>�t.8��;�b�U&-��N�$�Io���/��j
��������XI�Y��$l�ʩu�ba�4�fPv)�O�P.Ы ��ϰ��)ͮS�s����F��h��p�jbӜ��;�܎���������8���+���Eﻷ]���G\U�9,�|���>�4�#\��elHV�g=� ս۬Vcp�_c����--�#G�w���!�0��+n̙�2�(���5�%�N��������s��=]�,���)��2}(hy=US�=0�qlMg�>�0��G �u�E=g��y��c���pâte
y`i��5`զq�P�:DGILKRK������.�f�F�+��"Y��"T�9mu.BRua �nĊ�.慕��\����T��ʦ��W쓾� ;̌����:�l���g�D�\�
{Ȫ���)���,��s��jk{�嶴F(z�%�	�\;��u�?�n9���A\?IVd��$V��B�I �/ ��ih-B���B�c�����?V4��p�3SLP��J#�9��AJs��e (��� .�߽K&�ӆu�g2��,�ku\��d�׃��$�Ci��G5�ň�l��L�������x1�/1Ul�1�gAd����f�� [���ep$��i0��&�"���9�}ӈR@��W4(h�6:s+D­e�����m�SOȩT�d���T����=�����]�x5Ž�b�;�����np�Cd(�Z�xp��������շʠ��~y83���^���T����J���^sX�Rb�1y'����/�z<㜆������W��/�R3�C��>�/����<o�@?��15-�H��\rG�#|���׷%@�����PL5�%��b��Q�y��x����j�e~ʉ����E�e���T�|��"3Cm����]HL��O�@�v�tF��6yg��
��mW�D[�\}�/3��� ����W������~J��ߘ��,2d&�k�L�9P�ɳr#�`��B���[W�P
�iϒ%�[��E��`�� Z/�=��l�E��S\t�8��
ZyJ^�S�vpb;^x.5���qQ��$22;e���H�����Z�)ώ>XC��nf��G`{��m٩f�s�<���m5GGN�g��N�-$��RW0����<���]4��٠���_:oZ�>(��9az)����瞛L�"�T�x�����1.�8��� M�q��@���_�A1S����BQ��?;,��p�%�I2�b��s�yE�e���h2-��pC{˔�R�� ]�R̟�zpU:I��m�S5����f�1�1��,���M�M%l��8��wj���c�8��L�����d!�Fa񻜗����ୡ
'��C���lb#e?��f]��K�����&�!70�?ә��������D����8��[�6(O�.�U)ͫ<�۲>�7�`��ژX��ai�;'��7��% *wZ0�d�a}ΒH&��w�>�;YC��F	�`FZ.�z9�c��+5"�ӣ��T��M���t^�nK@bh�
cI�*M&��!��ټws�P]=Ԏ��3�$���j�5Y�kgS2�
SAtғ\rQB4�
�Ƙsϖ��=���~Dr���:M����7N[Ex$[�i�f��t�mO�52b���a!�F��@���%1e֕+�.������f��������8�ov��p1i��D��Q)4)��1�����Zw�C=�l枏W'���s@b�y����l��x��x(�<S�����J��J*��G"�vH��A�_�D��vIy�HCnϡ���v�SW��0� �ә�رޘ^��;���s��_��;~�z �ܭam��K Jd9d	���S���x��y̖�t������S�	�9��*GyXD̿R�ڷ{����M�� ���vԗyԌS�K|�����/n�%��~�A�Xm,�K�^� ���"��(Q+eN���<v�5ZC&s��k=�x�d7�t�~{&���̔��F�:j�v\��QtN��竌�^�2<����!H+��U�?��2.�.��� 1 �(�"1C#������-H: �"�P����C��% )%zx�������k�}_�k���%cWOĠ�C���)_��Z�S(����$S�Y	H3����*���S��]���"�+x����r����n4'Z	D>���BIz��&��q�}Q��d���aI�P#�9	Ee�_}�н��}���`�΢�m��*z�`�9�F�K�:�4J�R�ʔ  v$oT8�ߌ,������D��� ��_v9A���I�`���zA�����8}Yn1M�w�&�₶зj,S�x�!�\���`u����Ʒ�����FF.�~	�]أ�n���+|x�AHٖ�&:.�F,1'�*�#\��$E@��@��i�K#(�	d+�Q�� �g������xrMn�)�SF�n=l}0�E�РF]���L�Y���xϴK�q(���Ns��Hw�Ӗϱ���ӯ0Y�a=��F�iAr�;ݜ���)%�5���g�w}�CD��.1�ͪ�X��Ut50n<���FI{l��W�V��nO�Ƅ�x��"��i�3���H�~���|�fj�mW�enlK�c��w��1��������|�2�>�
��x�������t��yPKa+�4�0	�g\V-FC�hVB�������	�$�zU?j�A�!��t��g*
A��yA�2�8(�ubT�9�U��	�$K�%:����*|�f�Q����n9* DU��jl�s|�#(G�)�y��#לK��� u"_�ǫoC^PEjҏ��
���\�t\[����_��52���t]V7^���^u!eП^0:�zq��8���;ELq`;�R�e�}ہr6}Q��E�l9����gu4?���w�q�e܄��^b��{�6�?���M�a^�My�u���/:/��-��H��̻���mέ�H���$�x��YfӀ��T�D+S�-��x�����?zG_�
9K ��`Q��%�~�#�,��L�_\��Hp9�q5�zC$�eX�Ƙv�Я.�/�mH�o�>h�zrB��7�,q�2�+��T��sV$�$�f�j���-5��U���#fpA8x�S&��(�Ý p�9P|�Rv42����z�ս�S���0��T�����tB�ئ����U���P1W�O�wtA�}~����BzUЍ�b�e������<���rj/����y���*�+a�,��ɘ^E�47�6�$Ζ���^���)	H��d�@]C�!���c�I�3F��T|��q>�C�QC�6K�Bb�]le�q��+��hƜu����1�O�R�e�%���;�@�9��L�JjK輪µ�/��_�b��$椂q�'чåߞ��Ρм�͂r�\:��K,_��Y1L�׈�}��x0*���J�Qu˔��ǎWc����(T�Jzyލ/M-�)����~��� ؟B��qj%y>kE*�������'c���k��A@E�$dr |s��?��J[���Y�������F����ٻ9�|f�ũ/-tp��^�����t
\�T�3�����'��j��Je���=';^��ݧ��z/b�ܫ�o�!�z�q��������cBluۘ�%a�-kA�{cW̼۾l_Ǭ�(`�FH��)�Ġ)�ԟΉ�2ˑ����5^G��}�����/����5W#�m-ҩ!��Y�L��_�� /{��N.�Q��~{��C������4>'Wº��z7�o��kU����Z�ƯC
��ctئ?�2jAΌ|���4҉���xS6.[h�|a⑾@�b�=Cm	+�r��3�)���մ,E	�A�T&_����i��ڍж�@�0�/ٿNoә�Y�.K�f��q�����_~�^���*ʃ�6��=�˯�o�X�8��㝱L�=H������	#���v�h�������q�h�#3��Bu H��7��ۍ�k��h���2���5k�ǈO�,/���!�,�0�?!O�:d��+0g:8q|��^���Ne����5�t4���{\���|�n���Y��!&�C�O�+�b/�H�����k�
P?����Q������_��کkt�����;j��O���ׯ�Hㇹ�t�~iyM��Z;Dw��:��@���l�/L!�g/�!��#{
+�gyLߤQ�����W'�O���90���C�YR�f-�᫓�/V�R <�^2q$�r ��r�&/&!�L�7`���������,���mi�́�!��`;��ފ�����$Ў_��)Z���d�#��Ó�=��!Ũ�rټ�0:M6�x��Е#'�Η4H�~*<R���I��O\��#�S֋�a�8bU k:�"��U`L�u���mU\G42��b��S{Hp�a[G�A�ј�ٕc�1�@�P��ڠQC�pl_^�2N#�դ�<�29<?nv�9�m�s]UY�,�_�����Z�Ӂ��7@i�J�SW��;���%$IE�<�j���+��4�44�O�^�U��}����ix��g5�C�@u\����}9��=��W�e�ԟߏ���oB�
����K���F��v.j]Kz�o����!:�����յZ���XS�|��9�7�x���ۭ���\�^�O���/�T�Fv�Cc�xvKZ���1����Q�ڑ|T���\�C7��jLēFos�%:K1f*��P�����K��(3WT3V���3y���,');�|tgg2�U�0�~�c/;;�w���^�*H���-Z/�7H�C�`orCs��<>R�/��혻y=e��hJҽ�Ο��=A�`-ߕ�����[�㣪iH��9tx�,Ciq?�����Ż��ڷ��:���:s���Y\}�WꝎ��3\y�T��0�N8��Y o��?����s"��|6F����ʂS~U����^{���)���R8 r�%SFQpY��Y�� ��vB:���N�]"��]��e���4��A�}N�ar�sj'�M:=ӗ�&f���<�?T_^2mX���b]����K�P�����T6f��8�2��2��nzOl���>�E��q��JT��Y�a0��8/ћ�]>�{�3����RL��-K7�\ڲ��T��.{���5�u:g�n!��$�4����#���l8R��lW/
���Vȏb���������è���Lw����ٱ8��^Qo*ٯi9ͿuQO`
�D���~ʀ�_�lw��z�L��fxd���4��x��w��T�i�xl;�_�k�{=�9{C���Z�9����!�x�l�r�ʧ�I��w�fϩ�ef�Ʃ�����P��bk"��8�#�"�Y�w>������l�y�����l�o��$� �o�yb��݋��a��������yZ�:H@�F�XJǤǛ��V�S�³�&ײ��@K|�!?ӃY�^T�G�\�1/W�\���]�t����"�6��f댫&�&�m��u�Z���l�4�=�eb�`#/O�7)����L�f�����=��Y���<˜v�JaJ3g�q,�\s���3O>��X��+[X��Y"�VSz_k����G�#�Ym9oA�Q_mI}�u�̌Xz(n)c���6��_1��]���{�v��?<h��+m�9x���~T^;;K��%N�FU�h��3ӅW���A/?l�\yY���D�{���nz�˱*�(�N}�+3.D�^�S36�(H^L�s_�C��	ٕp�� {JQ��1��JJ[,�6��]~{E�N��&��-zi���&�<�zR/�1�rF�%a�@7(^b���`��`Dzf:����G���BF&�5�8'�Ŋ*�T��.Y*��}�%�������(�{ݦ����ܼ��5�/. W�IZ�3%�	1VJ�;xvc��{G��c��q�7�E�A���MP�ݯ6��ta}�C���V@[�,B��r��B�H�zŧR�\����d�PK�Ca0�8-�'h�Q�O���V_�s�;��T|%��l����g��r�~�{��<�:E���XC	�A�B`oW]�+e�:3`������Ub�ac��r�M��l>%bW���.v<��sV�����:ƕU� )�,����,h��A�� ����ǔ�f��[83�@��I�Y=>nX;�t{��XR^wT�R���0Ċ{����fM�F�L�?'\65�u�dh�_��n�{�����@��4�(�(]��A_-�6X���j~S��c��[Y�m<�tn�'�1o~.�e��z7�B����",Ƚa���N,���������v��q������mĿ�~��n`0�r���t��d#Q**���~�'p�Y6�@�x>"N���U6�-a'oNܪ���7+�+z��c�!M�}.�b{�萑���3�D�/Y�3�AQJ��G�j���):�xX�S�G��GGD�a��r͝�2N�X��J�gې	�`p�A��8�"Y��\���Զ�[�~�Y.<9=���x�E^#GJކX��|��L����90��F�DvE�ݢ"K�ļ�>|��ь��"?�z�xY\ؓ�2�C�ݘN��$�g��̧F}{-���"��Kzw�����_�!���ߤ��9�25V� ז��}X&\�ק�[<)T��=3]�ɤ�By�f�s���k�0OϬ�D�U��/=�{/v\�7]@���
.��D}y��X8
,AOc�X+WO6_�W�Xpt�ymPl�.W�J��H�����b����~�mRV�i:<���3�~���s��>�~C�'�",����K�\�1�*@l	Z�3�:�gF���Y�J:�A���b>��}rb�2��0��~�(?�ne���ã�����pi`�������T��Ş�io.� ��<^�:}3�n�����=�V�2�bR\xִ�,hu�4L�m]��T��ĴO�������	2��B�i�¡��a���F�%��d��z�4��/T�pC��lM�@�؀.�d�	��@Y~�C�I���d���:�������;̎�2rwY��-�tq����V�c_�c_������w�`�l7j�j�/@.��ܦ/���=/W����N\�G��L��n��amJ�of:D�b��}.\����}���=Ւ�?�����k WDҟn�
ܧ���ͳVנX��b;F�3�,���~���Tm2�Ɲs婉��צo�/ ��!NK�V�q-"��f��,�:}�9�W5k�)���,�N��
�8�l���*�o��y:;3j�bVOH���Š KP�E�A���|���1N4�&�h#(���OB{�!����5g��2?B��Y�	���։#oK�d8�є��\N~�U�`��k%ђ/�b闔��?�=,6˶>�I��3�);aIkЏ�U,�����1��c*42{h���m�q�����t���;\=LX�_)�0�ĲBE�{\6�+	���	��Ёb��u1��x��m��*҂]R� ���&Lh�O��qM����fU�ژq��9$q?�	HO$	�SW��mQm����\8�;(���u�kCc�A�����?vF,�
�Q��+��������o�rLZuY���ɾI�D���x��ud�4�����L#SUU�U��������"��"Dm?W����}�m"d�����w�`�!׍�g�`�����uH$�0�(NvM����쩪���H%�܏\75*��m�x�eib�&�sT��+�qWG٠kLT�^q����=�Yt^i���E]��X��/��mf�usu�>	0ĵ��b�)~��pF@^�Z�s�3�����_Y�n�YABwF�
��e��|��^�S��j�+di�3������JR�q�b!�F����BcP�I��˻�=��ej��~��!���N����RQ�G��	ƭB��5t4���� �|\ש�(��1c�,�'��B�)2�X�A3����ڪ�_t�SH���nꤺ$��'����)g��>��{(��F1�ݑ���i�Y �k���;I���a�j�,L���TdɪVsNK:c�g�t)6F�};�Ё�e��D�D�I�/���7�y��oF�n: �1�h�&���tQ���7?�t]1[(_}��*t�c���g�^&�W��0xNmٺ�Txk����=�=�M��A��O��1[�9:
����5&w�ԧ���h��r��.n���������I���I���_�.�ݻwZt\\v]����DiM�5s�]���C
g7߃���=�cQ�A5��R�ov�)=�VpM�ے��k(�,BV��:q��:���9�F�FJ�HJj�íó�*b{T�Z�
�j����MЅ\��G�����
�r��>��Q�2��?+l���-�|5s6�#[`._Wn��%��^RPլMx���'4��߯�-��~*h�f$�^gR]`���Wy���d-�xd'�upò��G��PD���^�������v��j�IBtc�	l8���83�f^�.�{L�5�l[^�9������3���տ*txN��y{�0��mh~���.�y8Ξ�kҒ�7�uO����(j�&R��e:�Z7�P?0�iv	Y_ 8iA��kJ���'��>�:&�Ì�q�;lj�ޛ�����z'#I�6&.z)���H�?��&�T�3�5�������:�;g��	
2|ƻQ�� m�E�<<h �"�\�pej�����|�;ju��l�a5�Fkc����96�ZӚXC�.(��Q/3P���<�^����@�Cծ�Z��,B�I��Ia� ������pm;�)i���������,P��h��l�h������� @�?^\"����⫯!7m��O�6v�"Ԉ_�;���ߛ!�~�ZW-�qP='�g{nT���L��)*��j�]���|�1:x_t�*�\��L�
*bL��,a�h�ea���z��(����I��|F��VJ����#K{��C�6�F�g������nd�Ǘ��=)�ivO����=�T�ɷ8��8i����K���;��=��	�-�{���^RqIL�<��~<�%���Zѯ��	���=rx��,�OaM���N�^U��+j�9H��I�u���6VefMk�AޑA���[�ۭuc�[�z��9-�<�YJ�."0�[�j�"z[%6E����aX�]��"�A>ɯ���ˑU��˿V"��J��-��d��US���P�����KJo�1\	�m�y��\:�8��-� G����A0	��d���"J�Rݘ��a_���<m}�/:�z#L��Jέ̑GBo.pX�<R��f��Uㆹ����&���/$�ߕ��\���Π����鹆������X%���:���L��S�aQ(a"�{չ�5�_�1o��1u�2��b����]A#u�1a�(���4h�23��+h�fQʳ���oNl��^�zW�/�y�ت�2����Hv
������/�5�����ʿ#�g�;�p��H�|;|F�̋.i�Ϣ�͍׸�[#��,;V�U���;08���'�6��֘��X���ų�8r�)�Χ�z���9�\��e�
F�����6�3���<W���7y�.'�);o�������Ϻ�%�j���r��*�Z?�5eH�+b2���.��7�s�YO�ƒDS��2�V�)�^�����~����](�Ep5ԇi�U�ΐg����|;�&S���-�`^#b*&�������5���$E�a���X�G�X#�
f>l��*� 89� ����i�#���rTm���%B���)���ax�f��	 ���r´Xo8s�*ɴ
I`f���
':}qo�{Å�K�;����Pڦ��CQE��uev�b��PQ��j�B�q.)�w���B��0Y5.��ۙv�я�=�+S�
��yρ����e�sD��V8�ж܏�Ed��Xu�r[�L[p�+U��#�Bz)+g��3��3!���A��+�|i��IUz�LR�
Tror�Y����Ad��=j�T�$��'g�#����`v=n�r��&���Q�'��9 }& m�'�1C�~��½�v����*���ɮ�u�	�	d2ry�� W�\N��E��\F�M�]��r摟�#�wY�� M�u��͓���V��v�ҫש���?��l�皭����Q����d*�`!�X�!�^A���>��}�b�����I��L������x�����Sb*)�dS̞�bn ˚�7�cG��!=λ	���pi���˘L�\�S>�gh��35�+m3Dй���_����e��ˬ�4$ּb��y�������3�Ĝ�f~{鸶��8�38->��&ӳ�HD�C+�۳W�o3�.j�
�맪\�y�/��� ��A��<����]���
��S���4m�A�5m��<��?W�n'f��C��-B� ��}�]ws7��z�����_Kؽ?X���[����Ѹ��;k�(�/	��0��n?��Q�Ce�6�T	�{�JD�L��@5��9��v:DR���Y�?�&'U���m֕��g�Q��egZ�������%���#��| � i��.�����N��U�"eϿ̔�v�$D�y��AN��2�Kś�X��5�h����cR�=s����,T��z��\�WV9�}u
!���#�j,�z��7�����,{��g�������Z]gǃ��o�]������R=�Xxjۈ�ٔO��9O|�)Ǒ�*zl�=���nߡA��f����pSp�p>rOۀă���y����$/3Ƙ�GKE/��7)M��e�#eT�R&MJ�ڊ�x�x>09o`�����U���h|��xw��&W�m����c�x���}^E�Y��h�?#�ye��EL����,5��8��n(yW���B0b��GL��P�b�E1G�l`݄�<�ל��-S42�U� ��+ʏk�8�3C��?'H�W&*@|��>"��Le�Z��&�A{�e��Y�m�"+��6*��ѣ�����ʌܵ,�b/��X�G�m?��2�L:Ƞ2N﬐�"���Ai�5�CC��2~����h]:��QJ)בIl$Į�^�����W��k��ڹp��l��M�y�cT2�1w�r�k7��G �4uhśB�&�D+~�M��?u�/m�$v�
��C�Ъ?e��7�����?1))�V�󋾗�~�)rVM���˙o��|a;&����e��	���ֱ��~`M��v(���V�	vW����Mo|�7��:Q��b|#�&k��y�L��ߣ�یR�)q
됊���.~?��r�t��,�r��Q��F��[���z9�Ԇ�;Ȁ�i��vP���3�������8,�aƪM-��'� ��[�# ��X<E����EX,Y	g���5��ϟ�j��D����6,�� �y�W����`���B?b (��G[�v����+�dUB!t�4l�%5��\�F�ܒhd.l��.����qV�����Ub��g��լ����R%��Ʀ����,<a�F!�&����w�TA���
O�JacZWSL���Ȯ��E�r.�$9Eh{��.�]/����A���5��W}�r��w�#H>4�%�p$/���,�� VwAL���޺L�%���	/���8��d�[0��˟�	~�.�ʞ�bPjs�4�V��R���XL�]��_���S����%���	���){�'"�[9���=�`0�p�S�~�0K��|�g�>��j�9U��m+X������hT��L�itS���S'�����C�:�r�I��fA/�� '�6.�g��:7ϫW=^�hY�j��aIdK�E�K�[��%D� ɓ���=t�8B�$wh�K���;a�)Q�<E��h/��1����Wţ���&.�����Q��-3�����cn^t�9�]%��;�����N,5���4&�?�������͚٥�q8�׶֒C�b�,�&3������o(����	���o����kU�7oP��|�`�Kh]���N�u Ac�b�.���(��Pאd�G߼M���J5��}��{Ap��.�G5r�P�β����nJ,P���W�ߒ� kc���dJA����v#���4��(TS�[K�ovL��j��7�晘�f�����<��:7yblD�.n��v�O�'Y���g�Y�[eKҪ61�����[[�t���O<$�l|��t�)*��;Ӝl���. �ـ�j�Q��h�׽�JU�pOe��BM!R�Pi!�Y�Fj�j�%�B$Ր�lSR]���P�mg�O�MO�]�b�w畃z��,��U��T�p8�ČK�ձ&*� �2ᝇSs���삔iü�Zk��>�vs��]��o��_�����1����?�n�ݿ?,?��٘�뺭������l��f0~��9����P(��J���V^Y�?8 ��3c�� ��v��Xc�?]�s^��l��O�����[���r�gj7�U׍V#YHl�S���\Y0��@t��؀�+5m�~�g�:�7�tx�T����l�h��\���4�?@Lf�y�Z8���>��Z��Pۯ��L�M|>3��b,�Zr{\�l�y>�hr�)L�j�ݮO]�ݍ����������2���%}/uw:gz:��+����������y'��QL��<�+�K��N�bG��-�8��uy�� ���Ʊ!��ʾQ �D`���Ŏ6֕	�����z�^�{�=��� ��� ���ϐ� �?,��o �yi�L4<�S�ĺLwH|M�O�M/����E	��T�9~NEBR>�%*Sdn�s������X����e�Qn:Z��]X��kIX�`�]�h��&GJ�;��<�Y�[�6���0�����VQF���1���U �k��۸
/�oQ�A!m[���q���7�CPSHq�yJ�J�N�4]eFt�� ]�t+b�8k�Ni)���p�%Z$�����>��j��фw}�N�e���s�����}Gt��t43�mx�7�iP�5T�w3P�`Dg#k�
��3�G���ػ����iZv7>���Yuh˶QY��
D��r���<�l}m���$��T��r��-�F@��M�w�PG����,�;�� �47�)n:�_\��`���U��C���t36�3o�������j�(��	��i� ��*�{4��/�|��Q�p�ן���'�>��j����Ƚ0�;�����5�y�i5���s��Ĵ9Qfx�`pI�&�Ԓ��	X���A�մ�;���גטV �hT����}�b�{yNm��9QJL�k�"��*aB���鐌�9��dc�`�eyոv�a�@�y/ܰ-���{r�$����mvN{���ɅH<�}L��S=��<��;��M��e���wvh�k����'�G�T��4�`�W�oZvr�6��o��Q*[��ۣ>���
��?���u�W/��Lv�D�r8��c�5�5���XomՁ1��4k�o����oA�E�<VF�cy�}u��K�%ȅo���4+37����΃;�H%dq?���Z�Yu�Ω��;��d�a=yw��7E5��^��ȗC��?��Y/��Y��l����@ԸC�Y�oii�0����Ф>�U���N���3B�,�Te.��H�4 ڷ:t�U���3y��^}Ӆr��:@n_1Z�a��/��F��q���Ɓ���W�L#8�;Z�X�"�u@GB�mS�5��([Kv�����~!�S��MƩ�����Ja-�r{1�a��������&K��z~�z|U.��PR?��ʻT&gh�O�(T&7g[�}Z�w��	�9 �qQK1��Eh#��]�2���G�ڂ������x׬'���<?2>j�c�"��.DiuB���!��#���s⨆VlN�F��}D~̼|3���	�6g�#C^]dk��M�5�'�C-y+r��{8%fY~:O7���&Y���d�ݺc+������h��1������$�G���?o�A!eV��K����9:u�W[����=>0]B���W����>��)v2�C+ϕ�r1��C|_QR�IVQlQ�&�4��ѹ�C�+�V�I�tVY�hoX�*/Ya,�Ǘ5�*S`@��z��Y�5Q5g�^��_���S��8*w��EO"�xl���̌�jD�=�I�=8���w����{_�}w6���(�G�X�лm���ʼ�_��oa�m�ü����~��G���Q�4>�W�B�☻���,_5�՘S�o���'y�O�5�bM���Gw�b��8\ 	���XH��q�};YsAJ9G���`��4b��9+2�ԓ~?#��E}��)�b���3�j�~>����J�2W�����U�EB��
��b@�ZRD��Fv����/�8zd�Q�^CN�6k���~����J��^�Ou�?��VK�xw��9����`t?���`���+��AE�*O,�v'��QA�3���`�M5^�ѐ��$�O�W�ԸTp0:WU��Q��o�2hMe�IWr��$�-Ź�{�P��'��P,S��v0��&�Pk?*~V�D�}P$�6��ʹ'�d�X���a���G�����ݑ��ϝ9yH*XB���ܝగ�B�ԑ�A��/1F��,Ln��w[�M��g���\�t^�Ko6�-M
�d.lm��MTN��x!�ao���b>��[B�%�<s?��I���hb9��/H6������q^�rR{�Ӆ�D<����A���׀�G�=�0~�X'��ؔ-�Y��r��Dv4ۛll (d�ǽ ��<F7���֧1R�pAf���(���5�t�z`��Y���Ƥ�q���Mzs�˯��=4�҆?��'/jjHx�^���J0�A�Q����}��k��M�د���vK\^��P��k�+�iV�:'V��P�Z��Ƙ?ȏO,?�G�]D�߈O�^D~k}y����^�?G�͠�����qɫ>Y� �}�NX!�Ph�y��[�O3�q�i;�ov'�[�b���?����q�!Շz�a�׬��)[�͌}B��hiZ��ɷ�(^�;M�h�X�[��.Q߱�0u�ê��t�cO7F�G K�jf�G�*Y�� ǥ�Ot7%>jy9ǲ4)ZG�2��!���mw��<g���VQ�F$��;���&41�*x�����]��MB����SL��tY��x��8��Y:�&�4��E�~�`BkH�NY̰l�Q+�o)s�Z��a��E�nd��΋	a���"�W�e_�;�&�z��L�=ǯ:?��A��̀�����ā��5�I`���_�=<���}��<:�*����G�E������ԕ]�*3�#J\�-ͳK�{\'`��ى5�)�30���aK�'`�l)y ͼ���tO��~03z�CG����F~�
8�y��\�� �B�Wmcy�ʈ��te좈�A� S �F�nn�@���u�~�1;�_�w�@���1��6F������5���<pa@{� �[@=��#&�r��땉�i�`_V�w�_�l4��.�%�W+r�v^�Ero+��������b��D������w�E�eX	�wV��I�k6�B���1�����C7_F�h	�Td?s�A9��
��I��2ul�6�����|uHd�Á���	��xX�%�fRpz��ş��]�9w��τ ��ְY=���9��
�ZV�x�Mi_K���eb�h�v�<h,Rsr��]�H��{��7]��<�3��T����?%�*d��.Wn����͸�+��'��Uþ1y�z?T�E�3�2}�����f�e�� #>�k��|��	����>�0=;���!u�x�_C.��̏:S��g�VgRW�H�d;e^T�[����/�f��H�͠��գ���\�5[Mtt-�D��������R�l9k�w7��gC?�n��3��Л��!��?��~[�o9�-l��������q�QZ.	�����w<a�5" �0��2�����޼0T�Tөئ�V^{F�ڇP[��A{�������Q�>5msn�{����T�k���Sk�R!�E�j\�;��/�9.ń��{?m��n�Ld�R1W�����ڳtk��&s�-�{y԰��������F��ܠ��ú5j2���Tl%fM�:l:h��]��9��t1�����b��ZsW���of����y�W�yK�w���fD��zsD�	@��*膉����b�2��>|�M���` �(�m�&Z2�'���rFw9 �y�{l�-dL��G��@BS��>�HS;L:r�7�H2*�|0(AhI"=�z�/�gu]z�䴝wޑ�D����c$�|k:3�g��C�y{�� sIJ�[8s�哮�"՞7�0]�,��	�Wӯ ���q�w�������O�p����7m|<mBx�ɳ���G��Nj�w���4�H��E�d<�nƍY��[�˼�O~4d�A����7l�6���ը혠�>���J�Ӭ�N|�}��Z2��	u�M�GQ�q��mu�w�v2����m�-��?I��d��!z��p�ތ�6M��� ��|���̞�k�'{A�ˍ]�U<!����֍��ZK�4�M��~ib�y@�p-�J�Ou7����/2�Btń֞��
�[d,^� Ru�&sl�^�j�S������L.����MVc��#���(aK���90Xi�v �����G�b\|�� }Clo&�#�4\�z��x/5�/wS-$\<��cb5(J�%��}��l`��!�0�� y�I��T���X^���_��ՌYi�Z���BF� d ��I�Pe���4���SC+G{�!�1��UW�c���ۖ�^�V�����U9�.2٫-�.�~��̉��������۳�}�DᏥ��������?~��iY�첇��5����o�G��pޒ��j�$�c�N�-�]��k��
�ƹ��f�`�Hy�e��Qo�V�)f shi䖆s����>�bi�6Ԃ'H�
�ŨDbX���k���Cc�Fؕ#ٕ��'��!�34DM����+~������,�{@;Sg��D��_����#�����$���gU��lS�Y�R
t��pMH()%�����Z*�Fp�)`K����!�Z�ԁ�!�_���<6�-sV|Ơ��-ZNxgL����8�kW{^��~_8������#i�X�+�yy,�W�%���'lI���B�S[JU@p����z)#����U�������I��������Y4�:j�`�>z��� Ώ4�51lgo@H�â���P��0�4I`L�жQ��Rj��������YWE��s>&Ȃ�蚐0Mʿ�abj#$��i'e�߄�ro�(�{N�}A�2h�`ҘH��5������P0���C���]��Tt�p��d���c�K6S[���3s���8و��Yio�����+Ix-)j50bu�� �!KeGc*B�?��ڒQȣ��1呃/Ui�"��bE� QP/��3-��k����X`z����jgR.��J�@W��Te9�daU�SFsPRu�����b�w�S����#�p�+�qO��}叮�#q���{E񧱴�啡�¼7�4s�������c{�!�bE������M!��X	c��

�2���
����j�4g�x{�rR�iF��Ѿ2�Y+\Kѓ�+I0���>�׸3e��䔡��k�!�.�@4l�R�M�PM�29{���H%�)�N�ш���G��xĤz׎}B����^4F�N@���waP��k7进	L���3�Ph UV�j�3� �ܖ�? ���f��C�ޫYt��T������y���5"D�$���B`�Bi߀�6˿<�縩�z+_���+m[�t�>��6��/�tUQ���LdwF�{��5t:���f
mn�QDm���.g�&��4`��57h�x�7�����R�2���&����I:�+�ȸ�3�@��e6��u��������Ov�h-����U�&�2Ì��==̌qA<���s5���3�2�\B�1'��qӎ���6�ܱ�����3ƃqw��R��{�b\V�/w6�Eoљ�eU�mv�!ȹK��LJ?��9����$G*鞕x1<�H �X�0�b��^����!����M�3�'"��an�"  �=6�켭<�ㅶ`
�4]���/�%���	j'�� ��[��T��-��∎���/T���OnF�c��יn�M!����Ӎ��=a�9=qv��wR�M?I�Rk�.������o�ƿ�m�kYd�^��'��]�o_��f�e�Q�>6��V��:�%N-��c4h�:��P���ۛ�.u�Ӟ�sf������tL>ϳTv�i{�?�%�xzlhm?d�S�w}��Cl��ɍ����@��e_����֜�y���>�	O��߸UZ�E�Ԁ�=p^�j*�mW��'"��8����"�tJw�Kg����q����"ݣA:Gww)!H3�#$��kH�n	��%�����b���ٳs]�}��9ڤ4ɂrMzv��X�zy�D�*�w��ȟ���_��n֘�%��M$���~�9�[vI��5�rP1ZE�i]�9��g}��_E����!3F�g�L�3��.fއ�c�Ǆ�榭�[.�̴�Fżݏ���".j���w�c�VFlU��G��nsg���FRw�*�΍V�U���*��d�D���\����y���>��dVs~��)NL.]󼕚�S��|���W�[��ؒQ$I���VGC'�n*�C�@<nǙc�y�����B�F؛2<��\ ��'�~�1a:��)D�
Q�}}��@j�	��j�k(��;�}\�dޗ���*]U�]�����L8صv�.�о��A�/��x�͚ҧ1+4XL9��(��#��QQGbj.���zE�^%�׆�!Ƞ��	� �֠i�K��T�qR�$�,qD�e�wx��%�-���XxS�ֹ�^�E��R��nrR��5�;Ca8�њs�[�w��)���}8�i�5�}�^���'N}��|�/�3���v2�/�X�R_2�e������`29�����OhW����qR�U����b��}���n��V�d.�Y���X��`��5WF�Ǆ�>ƫ?�0�sՠf�\{�Te�`�{چ<���N�6w{��Y�w
����֔�*� g]N�����ЂRZ��W�7[bs!X�hTZ �*�	�v���ː%N_'�)$B��\�3���oi�MS����D���K�%Ew�46Rr'�9��=�V%�n�Y��n��t���9�)$i�C���P�M�Fs��?xC�v<صa���у<Y&?d0u�����y���y%
�$?�,�xj�rO�D;��h�p8P߿T`��m�}�����b�ޏ����]���^W�>�Z��+V[��o���N^�O/?���2��I�Ş�G�ãE�v�l~h�CJ�R?�~�p�MQ�H��]_s���{���a�_�:l�5�Y��/�wɮ%�mې��*J�2��U��.��ب}G�T����[4y�-�ߘ��]�n�h�ݞ�|h��o#b��)��6?��ʰz��[j������e�zZy��$Og;��v\h�-�DOq�8eҝ���0��rV�.�~¬�p/cts�Gu}����xA�.쾭�7��Gj	C��4�n�g��>�z�p,��ɂ��O�쳀i�p<w�<sP.�)T����|2񗬣k�Q�eNY�k!���nU�[�f���.E�q��(���v�U�[���煔ƴ6;�м� ���t��{�)?��P���$�A�7%^�A��__��9��Z���͚(�3�SMQ~����,�Lz��b*43&l	���4��������B/�Ɵ%�S��6�H�4"�'!d����Ƣp�4s��'ϯr��(��\�!�gL���T���U��Ljzze��66�����2_��Q8��C�,����u\r~�1��'�M���6�̞
����n��F�xA�޵' 8����"j���"Ěrd�&�+�?*�[��ͦ;DZJ���o��Xw7	,X8�����\5^��.�n��w^���e��pտ�]&���Ƭp�!#0uM�J�ya?\�;0�o���e�6�\y��׳t7m
S�64�������M����-?�5����J�|]ғ��>+���d�).�ר�����{a�{=��!=4���ڋs�q����w��C�ѥo�k��n,)���S�p-���
�v����t&���s]v�x��s�@{՟�Z������LL&�}?�%��j�-YRo(v�t֢�M)Vo�A���o�(��I�܅D����g��ڿʅ}.�c+����7�[�;ηȋ����5Gz����.f����o��SqEo*���;�������<>L�<<^6�>.�ܞ��-�&�8�/B����YM���]}:�7��
�||y�6ǃ�)��Z9;����$;�kh��i�2й�u^��~!��|GE��X��B�@�0�W���Q��2������I(��-��_d[0��B����6�ѪLk�(��.������u�\|D s�9vJ�<�Ʌ�^��>�u��T�	�
�J���JCA-k���|ҟ�sѓ�a�z!��Bq3���0?�%d203�$� m֨c���Ӭ%�)�S��Y3�EbW2����Z�K87܎GOV,V���� � Gӛ�zwng�5���c��Y7�i�*��Լ��:K��HHd�\2oz |4q4*�-���Y���:��E�3u�W��-��Y�I�Z��J^33�IF����#kzh��{]����+HP�����	
�I�̻��_@�cZd��n�֙��M�
d�g���ӊ��e~�>'��-���hm��>)ol��#�K�k�|�iIv�SbwJ~I�6�A�B+��E�q��D�%*hnA��T�<Ę��� +��8y7��ǲZA��ς�a�36��6�C|MZKH�J¤�)3힤͛I�Wn6(/�4� �'�'�2�2}�����j�z�0���eb�JIvV������1�H:A���n�1U�d��f�P5�g��"�/-@��ga&��ar��{KCyc�h��P.uvI�����>b� �l_}�6��p�������;|�.�����"������@{�a(Z,��L�g��X�Y������S���_�z�����/����ێ{p����-4��TT�����K��N-��[��0��E-�Ȉ��>m�W'xT\$9�k�]����ٳ�:tZ�0������4�8*h�[Á�i����n�9g�����x�pW�����7(����$��� ��]Ǫ���k��H��y��={��=7�/�qF�7�i����5򸇝���cx���Hm�7���y]F9M��`�NUֿ8��	���6��k������5cQٗ����=CA=��A�, �-���E��VV.M��ڴ�S���T ��A��@�Y8�N.W9�4]"{!h��sC��$P�>|";��9E�'�WW�@J��Q���kG��"��h�����sM���b����J�-��ˤ��qu��*�%o�7Z:�f��ˢ�q��*�[Ǒ��Ӗ��
%�O��L,�d�����{�B:�ݷ���%`�����u� �x��3D�&�)�&G�e��d��L�TU��R匲H��Ѝ���^�@kH���nm6�3G3Sm��X[%8E�>&l'mr�E����o����i��&���/�GΩ�����o|W�ϭVn���Fvk��,B�Z� �
pu�����q����k6���j��]*�����]��_�Eρ=�f�y�f%�Ǖ�"_�/�˵��5��%^"���;Ѩ���ke��R�N]�12�?�[�>������˓�����Fܓ�׮*�X�RPCE�$�	�&dډ�g�b|�;�E{�ח�'b	ݿ�rQ���|��K�.q�ܜp?$��$��$E��U���X����t�h�?@��dv�H	vd�uxj�G�Q��5*���@<(|.<UR��^`�����$���f�Ϋ���v̆e��z{G������E��_�s�S*�n���V?s�ܝ��t�H�r�Y�a�:�~N����P�]�>.�<�f�=�:�ݬv��<z?<��<�kS�74��h��DR?��k���vȌ��)��J�����E�-@�3�ݶe����Vc@�J�ؕ��E�39�`�fj�e�����AB�����ae*��@ם�������5�19�)�$V|LR���q�y�����^gK]��<B,}[��s��^�fW�w����-B���'3ͪm��H�"�v	d�z,I.�\�0�b|�i��+��+��v�+*�?��Xq":nw$y��ޥ|4�D�_����la����R�I�����]-�G�v!q�9s�la��kO����ɦ,3������V+��:�N���f	����3]���(�~DDH�6�����]�7�.R,������#}���sF���EI��=N��F����P?|�����<`��)P���P����Nk�V�j��7 t8�� @����<j�,���4k����0GX���P���)�MDhi5���5�gܡb柞As'����jF��U�3F':��ˋ��IM��Ο����?dMZJ�S�?�����f�Ѡ�1_OI(�Tv��Z]',��^v����}*� Wo;��	��V�c�KN���&3��+��w�ї�|7ڬ�\5sp�r���G��Zg]Җ�0}uL���4q�I4�߬�ޚ�d�5�?�j�v�N���K��_J��}J6�C��on��"��Ԑ���!�?m�&y�_�ߟ�Z�X~Jq�W���a�ǿ���d]��>?N�f^�M�:���%Z��b_v}cy��\	מ�@����T��}����~噄�����
VRԞ��b�i���j�re��G�<�xn\~�nq����'s��[Q�KfeG3�n\����A�I),�:���Qd^��EgI�"����jxPm2���[ީUi� ���F���l��v?�����+�|�m#��;�m�]]p���5$bT��c��P�'�ƚ!t0��J3\��?ڻ��^Z����L��o�5�\x�rN@�Х
�W,?깻�l!�;�sD�j��oRs���W}�o<;<��Rg����{�dd��wS�4{��bs�֨��Dx��d<�6t,ݡ֧AX3y�]�C���9�����OzD��3C��R����[�E@�����1�|f͡v}%A��A�d:m"�إ�f�>�Z)��XZ��$F>�g^�e"�S�]:�R�A�j6"O�f 1hM��S���Fb�d*��@3DE��bZ�E�
K�yh�^��e�km?��o@��W��}pL����6��C2~�991f�ϻ�)�Zx����|J�Y?�=fO[l�ҥG�A4�Z֞X����ݬ�5Q��x�/����ط����/_��xyٓ�
�NC7�҆�K"�bLYNb��ޓ������J
�T'���n�+w*Q?�>��>v�� ��}�*� ���2���P�9���esk��v|�ȓ?:� gq�d�^%�I['d�Y�Z��0����%ϟ���Ph�V��I�+	FەD�����ƮÜ��ZP^��l�����3��l��Z�GVX��7��T�Ub�s�ZZ�Α,Ah�(���^��꿭��Ψ�Ŋ��_�+���v�m���?��L�^@|�,]&�aqZS�S��i�\�n�{�7��ۻ�:\5�o�~�;�E7۲�����aA���W�>D�ݻ��Mz{�� ڙ�
��o�o=����&sX�27K������H�~�ݯ8(/��\�J�A��d�@����-N���!k������q�7��O�'��^�X5ܸ�)��k�~8�b�-��F ��������w��Nw����f�nw�4*��%�	XK�y�/(ow�E�%L��'�O1'���O�X6ivs}M�$�f�@A#U`,�L��(�ƌ������l��󅗛���?2�f�ԫ{Ch|�6s�Т�Vd.i�:��݊K�_�&�,��.1�K������e7t+��^���/s\V[5_/���>(C��.E���g%n���@�����}��)v�����	���	�ǻ�������������L��e������> �̻bj��~sqO9uQ����3�bQ��DMa5�W�(��婋oiR��r���)0��u�����+�SP	M�������6ٴV��ü�*4i�PM��Q&w�fi��.7%�m�d�b�bb3&����
2��aß��n�N*`�����U
]T�>3K?y��1��'9ĸ��0����^�ѫ�����ґeɦ� I���4&܁V"jQ�r�}��T�kŮ�>���fWĔ���k:�I��>b���d�r��ʑ�&ۃ����T���4x�$�x�]x^�|���׷��*�V�x����S_%�83*^aa���IʞM"#:r�\��4*�Z�F�f���Fӳ+��2Ss�_��q�D�T|�1V�~ir�:pҷ0�-`΍�f��Yc.����e�ώE��S���:���T�0.��Eh��}���~�C��\���m*�LN����0�f"�c���.{m.�Au�ה�=9���k��)��.���#��Kꑘ����scu�I1��jt�5	�����I�v���tQrqPWF���3��Ly3z� 
�,��T���&}N(�e!��C.z��v�3�_�mY��u��}����s X[�3�~��m㏓��y|���C�Z�� �/������ =�"��	���<H���=�y�/�P"K�~\��f��/��z�$�>�3f,�c��u+��t8��o��6�[�D
������!�� :�Q�N+MC�)�1��L�g��t�*�t����M�C4�_�s��,	���|<���<��6�[���:�4`���SSJ�S�ŐE����3�<^�?��}�g�X����6�L����냢�Efb��h�oa��+a�������+�mW��E���R��-8��ދ�/�?���j��N�}��w>������`�h~s;ys��ks��ԯ��2[�4������	�`���l%l��[���L��-����a�«���\�K��2����ӛr��`�t�w���,gIZ�����*���'��s��є۾[Wa/x:́�'j��H�B]�W6��n�mŢd��M���I����&չl�xr3����"�G�
�."���(�G�W�UwD;�S���$�i�(bv��,��}2�W綫�{�*w���M�9�39|�?IԶ"O/�o]HN>�+R�r��,h�;`bt#���w�G�=[
ٙ5g����Lfj�|��V.��E<�����)��<Tp:�"�
X�o�E9�H�D'ڞ�9�/呒�j��Li��36�Ȅmzrg�%�%j�ƺ��^4/;ԊrQD*ԥQ[�1�7��^�W�~�C��K���&��1T���i%�[�����%����NS��C=#������~�ru��ZU���)���TF�zFI�W��g$��NX�A݋����'y)��cL��|,��v�=� �9�5BR��s�1$|����qyM��W�CA�7����{�9q[Z�8��S���W��{�*}D���x��q����%G�!jK���(��@o���C³�8;�nm>���c��2�쿵{�5ַ���42x�`�����L'^�p*�g����	�;�0��)c|\�ߖ�R[�d@WP�h�z�~�Nv*�&��3�be`LE��}}Ѩ�|������������U�����d�^��~��������YA�2�?���dB���7[��7x�N�ـU���IH)�К�4�A.F�;L��*�))x �2�UR%h�|��� k�W��S�O�������H���/��k��]��Q����a���%VI0
!�j�4V���m��['���!I�	�p��⠔���Q��*�ti�i��"���6Z�Y>�r���^�������8�L���Ɋ�@�� �_/� 9���G^5�bdx/�َ�)�(�#��}�\��#��j���Kǲ�������fw��@���`��ֵ�a��]__{���8ͱv1m��;3�������՛ʎۇ��ћTO����s��^EX�u���}�㿑�֛�,�v�����j����e�
m¾��l&��1H�5��R�Kؽ[	Tb��	��A�7��IX�VS���u��!�,۵T�&�IJ2�SoP�s`���:��ާ�+DE�>��B{�k�`�۹���]�v|��;�5ʧ%���
����1���uOcBH7�ko������'	;�����?������%[��@R��/%a��T[�`	��1Z�O.^��I�����r"�iס���C�<� �j�AO%��~f�VC�r�=$] %zsYe2�m)��V��aM��/�t�vF�Ӏ�M�uJ�F���_��!tj�}5�3��j����Ȟ��QJ%X�"��1�%�3' �)����	Α<�ۗ�.jD]��p���W�rRu��[��B�y��<�&���I8�W6�	2�jmNyP���-.����Eg6��S�zPs�A�����4(w�2&5:Ĳ��p{����0Ң�$Wҧ�6��p�wگ�>�E�s��EMZ��vn���.��HnIg=��eY��[v�_-���	��f��G{��$���+�c�� 	�3<��D�E5��N���$�ƙ�6����I:P��C��>��z*nC��XQ
���7:�h���E~S�������P����}� ��-�%Fgg��2��V'�|����d���ݿ{O��eǕ��ʀ���x{��z��q�����o��*�Jh�qܐ�0[�����im֊�&CzP7yp*�<	�G�e�v�t�<B��Ö��]߿9[��Jf��0q?�Xی��8)N���̶�r\s^Uru7Pv����-"x��,Ȑ��F���nlíR�%n�G�;�Y�y�b8v\7�R����J4tw�����\"Jڊ>���j���V5��e������m8�ER�|1i�ߗ�#������|����q�X�z�X��X��~�;��8��Ud���u�xڿ{S��q��t��%�,W��[�a��^S���b��{_9Z*�$F��]qfv̓�xN3�^���>�X^�]'����~�R9�w����#[ ��o��ђH�Q��'��>��J0Ϗ��cA��b��JKg}'S�:�E�Eiߖh�Y���"ǹ�#�T�����Ǽ��1��#��+��&���rW'E�V�F�J�����Gx>�
(JW~�ҫ�}2���(�M��-�'���@����#�Ӑ�[�!�b��$�7J�!jh$aEH�h����Xo�0���GY?���Q��kI�]{���:�F�8t��-ο��_	yd]�ASGV�wu�z�ZSU�����ߤ���Ku���z���GF�
�pW~?�$/���~'ݴX�*������4t ����!ȹ1d3��Y�w�A7ʍJ�^��F�/�<�k���p@а�uG����aߡ�K9|��kK�*��7$xr*�|1�b���W��z����b��PQ|��b�{��:f>��u�(���h��GVMr�5�Q|~�tp�w4��U�b�ٻ�4�?�u���"���c��,�`���l�W�)$�+^�:���T�'�z'�A0.�%�l����O�b�xR@q5��Ғ�`ܯ�I�[E�t�%�z�拤�P����e����,�_��
��L��%I���to�`�a)ʴ�zJT�0��M0&��7��>�XXa�Aƾmw�6�Yܽ�~�,Ȣh@��a�\��R��h������UjNS����)���h����ɱ�q��q�����bg�o�0�?�~a��<#�����f'��~'��~��k�)>�Pߏ��Q��!���x�ж�p��Y%�nY�~_0��0�������_e�e��>�#��*0����eT	m-V&=�;W$�P�����Y�9�� ����4s#�qJv.%s�#7[E������$�Q:i6�>��^z4������3�4ol�֎Lq<�( C�&ͣjR&;��
<��\�ϸTb�Vqˏ��~�'�Q�KF���uO�%�0�u�C	�q����K��Q<"di�^�� 
�;Q��咸�b�-�w�2d�F�K2��+rI��%П��*�c�fFׂUY�L��+�#��������b��G��S��Ep�?�!��t��;��|\����i<��C��;�xr-��s�:�3_o���+b�|(�����ɘ�y;b�$BUFqt�+#zp�����r��������Fpą�99^2h��(r<T7����]-T$j��)~|x��KϸPK`>?��>$�ȿY~��7�p>zi�g�|K"��;2�?��7�o��uȒpy�"��=��D�p���!�5��o=[	te�����o�FY�&��6���$$�S�`]�1>ɠ�M�W�Q�Kݛ�ǈ�5�0�����zNI�~.M_������Js�-�
��6U6�U�v2�E$y��8xob��"~Q݃��lFӞGJ+�oE�Ʉ!ۓۈ����M�ɡ���x��.�xL�_��?�v�>܎=��#1��YǇM�U��>vC��?����v'��ûS����a˩i���m�7�ڌ�K$y�����i��~tɠ���E�
�}h��a}�ې�f�����1��"{+����Ј����~�ѣ�p�D�"�ist��s��/���� �6�Q�RSNC��M�H.�ԙ:輥���w 9�פ����O��	@&�>�������sb]`�E�bG�T�����G�6V�.�N��;��Ϊ���'�ϗ<��N2T���8��Z������5��%l �h�E�O�R��N&��-���)#kUE3T�Y(�\ly��Za5����WcW�E�8kڋI��\i�򓠸L�	v M>�G5ۆ-&ۃ��eT%SHO�`�y���4���T�C{���>��� �A?EK���E�K����2��HU��f�5\�W�Շ�-%�a�֟
�+8G�]�aӈ��4O��A�Ew�t�j�˖O<�-w5���2W�íx"b�4.��L�+SՀ��5
.��pH���i�%i�@v��ka@�5<�����F�|#��3����Q�_�.�s�/��0���8��s���1�"mu?��mZ���ϝ/*�C-wݢM�?�'���q�V�zP@�'�.Δx;s������x���&���m�B�����0x�?�>"�9��oj��	���h8��d�mԠ��5"P��\��׈�*3���L^�BXT�č������"�����߭סVF���G~'��J6ѺWW�S\�>����-'g���L9��Չ�E砕U{L��������}�^���7'�"�U_��w)T~s�r>\��vxٴi����9����e�̸�S�S]���>a㔿��'6�A��f%�P��ǆ�J ,A,�t��}8�C�Vz}n-I�gJx��ǰcQ���˪8���u�zO+�����L�ȅ�3���D��($���kzr�}��?�1�H�x��l��~��>�3�����Y�v�Т���TU���mz�y|�j��F�4����JF���Ǳ��b_�|�˕~�������e�ò�À��c�}q��H����|/�ḯ#p�i�~sȨ�n��'{&qe����`	q�O�!J��ў��T�3���S1Ю������ ��!�?ɧh"#�4�����;ȗ�nk�A�'T̕�N8�t߶�u���t�>���<���|3�.���4��i2l�[;q���6肑C-�NA�i�.\��+S]��O��a�d�YX~؟���u�� $B���Z^AAA^>�6�Q�p+��Zрh�C�K��)\���L`� %w��pS�T�2�XL�`�<�>��h@py�M�0׃��\��S�1�g*�v��57�p�P%�M��Pa:���p����mc��:���$��A�'�ݰ3�a�kT�B7w���kX�'��&�l�[������|�lxuE���&E��QI9:G\���S����P���/QGGbn4|-ܬ������_�̎��絖� �i�l�=ՉxR#�h�����n�tQ�%H�"C�d���\�N46Z�Hꔊ�`���=��L�1�w]�A�[�#9a�M��@Rҭ{�$v��kJVX� ��@x��jU���s��[��A�o�Ja�˽5�
y����	��>\���5?M�D�C�]x���B�`}^���r�S�	���pA�"�����)�A�b�}v����|솷?��-F']�����/�؄}L�ov�Ʈ��?A�A;S9c;�b⊰���������_��d�2���4�DƏG�=>��Bh��}�F���i�^��2���;9��̶����R�l��2�����;���&��`������#��]�'-�N��{u+�F|�{�C�"�
�*զ`�H��jբ_�#�2���v�Q.�%�2yG��uYNK��̚J�9b���]\?�ؑ�ل����l�-�![��b�AMQ�_(Pk4z���s<�>���ŭo�3�Hx?NJ|� ��(�&(����0	�D�/ �f� ����NC������+�T_�:sO:c�6�ug,��̧�j-�Ш�x�VM�	j.RY�aP� �*6�~�)�CS��Xd��)#%� ��=~��3�Lp��z��"�ֽyY@�2l8���
�8GK�~�����Bk���l� %;d��KGUp����-if�5��5T���ؿ�D)X���$�)���z8e 2��[V���1<�z*���3�U�IJ4�ԋ�O�u΄ɔ�$'��e�n&c�R>�F=RUha)��îU�[��KV������ұ&�oz���8�����I�X����iz<��9˔c�He�Y*u�*<YUؽ/�l�b4��L�f�oGd���A��.J*�&�i]wV��*;����h���v�1zr`��(��'�n�4�o��<����ZDhoiX���;4̈́d@i��l�c��p����v��7�$�����`�~���0��y���r��|�����'!z�����b���4�B&�twQޣ /2u�D i�#ZcD¥A�U+�§�JS���Kh�XYt+�x��h�fg������`����g����4=�tK�w�ܭ��J:v�o)՛��`좽�*]�p�6~Gt~�ٌY<o:��,?)ʍ�I�8�9mЍ��GB�5퍕~�y7LM���=�?6 & �Q��2����GU 1T^7��^L�l�B��]��,S�;|1�6 ��8�oX�^��v�!o`X��Sq�7���G�-���9�#����ʈE�N
:��&��O��e�9?	d�Fy�iAVHo�E�-!��SweJ�	N@#�˖#�:����&��#�Yk���W����Cd�v�I�x<uL�8gN~�b��t24��u�`�ɷ��#̢�Ϡ�M�>���I�K��!�E�e�T׫��4���0#��M���1�Lb ee���k��������ם�gzQ#'#����ϸI����L,�L��j��&0���������*7wM�u�6�������z�7����ai��;MyP�|�s�`�bII5#�����t2�F�h^C2�hP.N�XpL4�CB����Wj=?;O�Hѳg��ܝ�y|Q�����/94N8�݈8�na]Wt��/�_!]�� �(hpG���?�l\��yf�I0[&X�78W�e/bd�nٳ✀DJ�%���;��ܐ��cm�z���ʃd���m�Y�qn�6X�-t�$?7#������Lki#+��J��<i4����o�!終X�'�<mA��>n�`���!d%�f@���9IJ��K-Ohh�U���.�Ⱦ��~c6�|3yW����W�9��8�Z���}�(#o��.�?��Τ�1])��^і�,'�TťqO�����P��(�����X��N�f��e����/ �}6<����v=d����+2���	����[�ov��#޴_�<a>o�:�{�r���]�Fzp����׊���e�}Zd팭H�S_G���c��>e��w(Y���A55O�zaX%���g����{�
��J�eF�3lPb��D9Z��׀E��)/]`hg��Oh�I�4�&���8�죐�..:;7}��z�í��I5�1��y��|ō�I��#�t.�� ���9�?,�[D4ƙz��R!8f�6Re$�7�jz$�����:����Mvy�f6���̾��2��J��1Z_��PgJIl�|�:���y���>ӿ%X�r}��?�iᚉIo����<k�i��QJ�!�;/K/U�s8в1x�����Bu��F�݁��<{���*j��zlٵX��g�� 1t�)f�%���P�亼?LS1�;��$瘲AU��EZ�+�͕�Y���+n��`ֵ>U�Q 6[�O�����m&N��:\@f|� _�f��Luծ䢆�ڔݜ�ۚ��?[	c.���	1r>��җ�즾pꋻ�W+֞S{?�Q}���^٣,t�£?��+?�l�>��<�$���E�����BUV�G�tQ�{F�.ھ��hˮ֮�3�KZ?��6�������d�V�]���}ԵǼDJ-~|W���e�[J�4U����n��y����~�1P̆t=T���q�H��?�vK��h}0�I�),@A*L:b�D+PД�Iu�Q+��J�K�/Q�A�8��߿���߈և��Շ�ԕ+܎~WC�b�M#��zG|��)'�9���d�uo���m�Ȑݿ|>�����$���ۼ?��E|�p�%L�t��?�Ȑ���p8�Jsc�[1���C���@c����v��A����1����bI'Ups�5�vc֪9?�pT�	H�j2%(��Ծ�ֽ�ݭ�P/c��/�����%��Ja��S�t��T!Q��d�n%�G*)s�1
�uM�[���![������8�n�o۲�<�/��������mqyP�	������=��o�F{�OɎ�O;�����*m�(��eE���p��w��w�yx>�O}ߐp>!���x������m�rwX�q�5����W�����9����������w������0�sScqD�~�a_����n�T�*2�L~��I����Lh��-Eٚ���}y>:�� 4��_Z�m!}��H'wc���7]-�4�b_���lˌ����ZQv&�ŲB���kL���]�tp�wb��&|܀�w�b�<J?����*�wo/�������޺��Q�Y?=J;"�Mi��t�nl���~�$i��f�mt��
�zyq>o+��٢�z��q�w=���̯��'\N�)�19�[��O�U3l����+'�;��{Ͻ���>��6�#��q���| M�`�u$*h^�-J(��A���������&�: !�3d����t�F�~
�)I��d��g�s*��O&++�P��7�"�x�	P��놅���A���}ʖc�ˈo���G��S�"��,";����d=��n&x Q���w_w_e. �޸�&ȷ�o�c��Q������巻'�{#�\M.�[
��@����5��B](����#/'�Pd6D��+������e�4*���o�������]Ч\R��K�3�nAì�f^yK�/����m�N���.�"��F�i-xˡO��5���s���R��:�f^���Ha?0����o3�W�>�F��������r/�fO<��n���t\#�d�T��w}�+�O����5�8 "�"B���� _V�Z�u��y �n��pk`��*�zn4*M*ѣ�;�8��-������/�l�V����/��Ɍy�iG�&Pmt�.�l=y[�z2)�Z�c���IK`?b�@���"��=�<������ڦ��@_�;��O�?�&4ѾB!.:��a>}q�r��֚�-��6R�U�-:䏯s�d>�Ɍ��;�^��6W9��;�[)|u�������'�*pC�w��}���|j�����q��F.J4��4ۀ h�8	�V.CX�]��^SR��]�=#����7�غ�Δ�*H�3;,EeǦY|�\��kh��m#gP��'v�
M��yDU�i��:�!��Ĭ�c$��gX��pR�Qr8�i�FG����<f���c����*��)�ij]��k�f�
��%�N���Nqھqf�E�:ژ�M�e_�Yޔ1�Q��������_��$w�Δ�-Í%V��n���B�}�.����S��ȶo�=!ۇiE�4�������̣��B���[����MsQJI5�\���ܞ��|��6�zi6�c�����=������]&��R�'��p�"�M�5��t�'��f����ـ�P<��O�a�qo��އ)��}��4�/��l�jc�S�l�W®��ߡ]/@�,����t��Џ��l��aq����Ğ���G�7�9��І���}v��dr�8����uI77fAS���z2�svn��G���Vm�?�H%Pp��A<$��*�"̋�4��^uK��1�zC��D'�s��,� �Z��DeC�ͨ�PO���Hք�A��5B�ZJjj�'�~M؀�^7L�Ũ���m\�^�ۈ�o�C���AJ��ܗ�H��MBa��rru`;:��Z�����,���\Ւ�|�A�������1�?�s� �?�n��-JN���[���81���pP9���p���;?,�<�Έ#N`@����E���U��ն�����Y����#�۝����Վ;�Ǉ����ʻ�E#�-�Yb�셝l�ڈ���`�j!�Qez歭|�f�����. ���������_�}�lY.�92�K?���������5�K�R��Tpg+Z�������݋��,^`aq-��]www���{�L&�|ȗ$�<�9�7I�����7q7ˇ��,6Æ+��(�b�v:�)����?�j���H&Kw�~�T~�~���̟k7�b`�b5��7���� �h�$"җ�l[���[9�LZ	�2	L�3�JCCF�CC�3���W-W�-]��\(?%L*[����Ըma�
t=U&�ȏ\�4�"	!bV�ժ���n�1�T����Y�t��W~K˾�w��L��'w��̈́S�7�݅F���\���:�
?��a�x���d��)�;�L�^�_��x:��x.��B�W���M�f_��	�"'7�f�
�3�'� nt����*L�v�Y�<ٺL��~gB��Z~��m�a2�02���-uN���E��k�LP�·L�x,��k�]F����ϗ�j����{���!�Ux���x� �M�b����b��$k�$����m	3	_��2:֌��[Wk2G�T |�4C#	��tT:�9:���������3�?�[�(��MT?Kh�,OV�I��Q���]�Ⱥ9����� (W�T�(��Ϋ=�4�g�)��D���_Ʊ��L��ܭ��K�*����B��1�q���?�#��B���~� xwF5�X����s%��e�>��'ہN��q̔l�<x��8�����8����#�<0�썁�?w xR)%�Q'Z?�E�wv[�OQ0�iy���f�AK,e�f`Uնn������,>�������7�Ϥ��A�^/~���{X��i�L�ս�����]Z�=m�5l,�u����:��KU�$�Ӣ pO9�L�Y�L�r����:��T�-@����+H[�Ћ�-�J��Ѡ	G�	���F+�rb֟����%$J�W-V.�|�b�aq�Ox[4�tG��s�ݟ�o^���q:���� �e��L������Z��R9�l��.V���E��_МA˶⸩�j�G�?��#]i�����T��F9���A�T	�+�9��哌!	���v�.�}���U�"5��W GO�)�-��/tO&-���㿲
z]ƛ�g$;��* b�F���I�,2m���t�4٦{B6~|2+J6�� �%�Y��	��`(��8â4�!��D�zUnF����(�d�&��pSIDm�jԣA\?�ʍ�4��tn�0)�o��7d�sk!��������4<j�I&����X�������^�ўߏ�/��;�ӽ�4����*YIJj�ZT^�Iס���[�]6%�u���Y~�keYi��j�t��єue���~!�Մ)!����u�z��svFӢ]s����<M����^w��G�N�JOy����Z�p6��t6z	BP���j���dd#�`;j0����Ly��&��b>�:��P_�w��y)�.KN�,�Z����Z�HK (�6B
}����J��p��u�] 4$�%�\�:!:�����Qh�V�.�o>�|	F`0|��GY@n����M �yFt�:��!I��C2�2�$!����U������[a�
S�&�eE.*��56x�F�@��$TlҬO���}u�Zf��i=�"������~�V�i[�{7WB-�G�֡�zQ�|}H�n�=x&�����Q���-Ft������Kq-�
7}���M�����Zxh������������d�fatX��u|Y�b[�㇧yN�-	|���'���E�OO��t��E�xa?w-����|�=
����T�ث�SG��7��,�'f�~�H��{��$�I�~����`5���P�閭e�ԡ ��'_e/�YƅSܜ�6;#swFO�k�s�x$~#�qN���u�U�r#B��׳�1?M>6�}G�3�������a�nP�R��F��3����i/8]���Tg0��$Ź�cRPuZ�F��e*�|ȷS�4�3���p�����"C��h�i��~����q%��~i�z�����a�����:��fN�Q������NdI�`3�+T����� ����5�����7�f5N"g:��F��h~�$섚���m4j�i�l�N�����J�k��}!������=�.o��
F�Oo��C�R�S��Z�x�M�����'���c�t`������v�H邸�7"dYB��G��t��+젬Q�6�6jE?�Zt�_8����'!��Nop�����aN 3��ڡ���Azy���XZt�����o߾}EEE�
�h�]nù:s�d��|���U��Ј)>E�IB�G��*�9}	�@9�$������k����t�h�S��B����ѻ*t�&�YX���A���+��+�nV�C�.M/��>�תk�H}Y n>5����,`y1�z%��K�:�꾹�L�{�O#�04[�������eo�c}�A��m-7]/���	ҳ�4c������oK�pI�D���1�f�"f���3��W����k��D�Y�`t��{�e'Nb���	�~7A�k'V��(d�^����I��w�:�����J��C�i�ﹼ�K����i\�
ת�̦��JS(�Y�1�������5�u+��Mm�s�y����O��ڎ��O�p�ā��
��u����m�R�o��?3ﾑ�"͚i���t
��+����
�w�����hP��Sz����!��fH{!��B*�\z|�qsPsuFӅ��\��~M�lxz��~z����*�PL;,��t9�|������޲��Q��;w:=���L���%������j]lJ}h	��5��g��u�Z7�u ��O���9dꞚHQA��]��{%�d+�q;M�%�B6J����?V�
�12��͝�w�O��k�\t �q��J�&,�����te���2e,�56coQS�b	ߠ�ܺ�Q9�:n�V3�  �#�BS0��Ł�xN�d�y�ͅ�U��[b�<1f�3X/�3S:a��s��f�bѬd���l�������:�����|�ۍ���uZ���%	f�BcYD��c��BE��U�n�|�l�"�Bp$��O�Y�[����$���hn�ι�}g�p0��%�V��9�`�*�������W�f���>�K����}��8^_0�|^C덲�l
h8�w��ɥԶ(��Y?����F���=���/OgO9��S��c[����e���rYr�K�B1�7�F�e��D����ĺ�"Q�3�a�������H���\8�d#'�"����m,`�V�� Z��E7�����b�����q&�B�A� �89�8s��[63��f1/D\�'23/xIgp�`���8�iX!{���`r �#]������뇵�����<����5� }8��>�%�>4��(ǻhz���������/(CX�
�&��-�����()g̍���իp��w��:�Z�"��[���0�f,�z�kZ�����hxU5��5Q=wY9O~p6�Kп��YZ3��a�B��B�۸<��Sj�G׊5����!��٧��=���!�〧���ܹ��γ�����ˑ��X���g��}�*V��]B�tb�0f�r��Ԓ	�����r�������L�^�u��VN%�G=�w��2�(��u�����ۻx���ќsx�Z���~�h�}��GgX����#<�p���RY�*�fE1����^�N������|?Pd�Uy�qۙ�F�I����ċa�M����M>P�����cL�>����-�O��6ͧ)f���,�"�Z�ۤ�����s�s��4Rk� `���`w�$�b�Xѷ��� �C��nsR˚�d�y�EP��oU������5�\�OS#.�x(����L��Gj=�P�]�!�P��zc�qMUx�3��Hd��D4~c�1�����������'A��5M4�>�h���pf�O�3	�qm�E6��/�|n��o.�Nk�J�n�~=޼�}�z:?�y���?���xz�p�|���������x���nq�S/�/�z5�~�� �ܝ����|�1�TLYem�?�$��'.��U���H%��x��b˨I��JO,z�0�6z&�4p%k����9L&wr�}�3���fA,?���6�i�iY-/��K���2�(�a4#׍��pҁ~�M%	���Y����q����B��ͺ�ʠ�ȽC`�ho���+yQ�Ϯ��ق������*�+>�kd*�KvN_���Ʉ�t~�
	�
�ƒ���z�Rq�p/C%&�p�����`��Q�uE�}!��_��}=�Sv��󙅁���#?�G~ ?���3�3�6��&����(�(ށf0�bW��S������#c@�wz�J�g��}&]'�����E{�;�V�uI��W�r�q9(�V��&d��A'�r#��'{�M؛E����[.�:Z�W[Weh��6�l���RJa��N�%Ϣ��$�"��6'���q��U��W�Z�>��`�������NyG��UK��k���f�#ҙ`$��2Oo����Y�}�,��v�ϫ�7�c������+d���5�cM�z����$-~�:�ޤ��HvS#ɫ]f����}h�,��*{iH�f����1��������H�1�1/��_-� 1��O�P�޾.��Z��y�cs�iy�~x�a�t�(��4��@旵��%��4ŕ�19<;t}����s��$�+pc��V/��Qd���u�՜��gs�E#�D��2�J%-r��CjF�3O-g4{ǐ/[W�8w
g3/��IsP�.r���o
ؽ�c[}���p�`o�I	�p."x9G�8G��]�gݼ���N�7&���H&�,�
�D緬֬�K�5 s��i2>5���.����#�g��|�ە�}��}�^�٬K��P���lS����U,�WZ���r���, 
+t��S͔,*�|U�ѵ��m�E��Z�,��(; ɮ�$+��<xȚ�#��Ӯ�-��:�r��z�׋�\�x��p�_i[s�G'����Vؐm j��U��D��q4V�Y��\����v�e}��"�4K�'K��Y���X;��y�b6�N����#c�f��B��T�E_���DC�T=K���ݣE�	V]�����-wc)B^�f�g�)[��������=�G�1�}esw�������L��JYL�j�w(ǣ�MQڟ�FV��ԝ�C��7�dj���w�ztC��N�Y��>6P�g�^6��[܅����l�&��dDo�m��jK3���m�b h�6��m_�aY����T	��Đ�0�E�Ao��IBYp.���@9��vh�K���m�߻�/��ñL���D�04Jh��q�d�KR�ב�p?;�\s��UzylF�?������5�	��5Q����d�J�����s�=u$Cދ��	J��ќ�����q=�ӡ)g�n�~wQw�n9e�D�C�E�q��]�k�D���wuZ�fF2jZ/��Y���+��$|�w��D��0��n��.c�V!��l��ь��p_飪�W`�'d�H��_H��K��jU/g��.ٳ��3(��͇gș����n�H��j��Ï�Nvkl�W��?�����u��������*�K*��6�mFڎ�;kVr��K��"]y�;2ݼM� �4�$t��{�&��4�f��o9Z���0 ��F/KR���֪��}|��Թ��f�Wg�V����V��]���{�֖�,E=�1m�I��Goy�f�߹{�{qMm��|~":��m'�/tmq�~w�I%����m�k���Wۻ�g&�:�fVJXB5�}���]J1S���u�:NON�e�vl�r?G��A���:�q�Mݗ:�@C'gŨ6-��3�<����>F��'�ٛ �����olਬ��Nv�sV��4����$ݎ�]��k����{�������p�t�����͖�ê��n��A��cH���p��a�Q{��n�U����8c6�[XT��Ի�<j&��'�-ERRܗwP���Y9���z��J*�y;W�95��o�d���K�9���?�t��j��qE�'��G�4�F��ܢ�=c�Ne?@�����]0�K圦�%��ěI�u���8�J�����`�T�/����$���H��2��?���t�@J�U�yr�S�8��ri(��8��� ��E���H`����V�WW��n+il�n)��㻧��7WY��ҖJ���i������Ws*!�1D9��h&���#����)2㲹�2���������:��k�5M�ϓ?e��U�U�%�'�ro��`a��Q��i��U�3�A�2�E��0�T�v�MB�v|s�~F5*�ߧ��*��<��������ݓ��H�-�D�Ev�l��z�MvU�lv�S��-�s�(j���N�0W�;�\a�#�7*U�,G�N݅?#D���}G&��Ǘ5B~}��(c��lt@	F�\��(Dx�|����M��ηȲ@�i��c��є<�D�ʾDX�_G��z􋢬`�o����Z?<���ƃ��꿞�7��^}��יxO���V<�f�;W��w�+��^S��EP'�0��,��UvdAY��t5)k+8�ݜV�f�7"��0�����<%�S2<��������\�ܵ\��.ݔ>]��ܭ'>ߐ!�t�'du]���Z��`Ͱ���fn�ls*�9L�漆��.����*�k��'�u|*�u)���Gpt�&=�| /���ʵK6L����xАi����
�\����V�~�F�c��������� F�S���׉UP�d��O��K�i:�r���R�׽�dQ�\��P�lD� Z)4��P��nښi]�ʸ�\�8�_z/t��!x���}��X�8)��ّO�ژK������AL�>VU/)T�ë�<�n.����l|r��4YIK��]�X+-�~(<H��o���JOf~���E$xBo�	#W���s��e��,Ln��}Λ�<s ��"�$JXpB:'��h#�\����U�o�N�e,�(�f�QDH���c	C*L�¾�/�!_
���0�v�ĶG��~�(ӕ4�mYpt]ĐUh�L��o��ߏ�`�u4�ޡ�RǞ�pH��<�^D���"�Y���)�<ߣ��z�v?�ԵR�qڲi�Z��@���?4�a�������Sñ����0,0@E�'�n����	K#�4�lu%x]���K�ePÃwo������� \�J!�,��I��	��ʂa�Z]�́��Mƥ�G����ǻ���b��՛�E{�����1�3X�E:	H�ab�
	1|��^���?�z�M"��y��k���wL���c����`��&Zj)��p��IpL�jo��>��������EH��u@�{��+�ω��1�W��=�pײ�_,_�LT���CЅ;�f_�p�~ �'l���hګ���L�iL�0�&�8�{�TC�;��4s��<�:�D1�K����qsQ7�tⷒ��(W�Jʋ1�s�(�U^/���u�<q�D�a�&_Nf�|c�d�����-M��>sK��a}����#���a�L�4�����L��f`Q�(�(��8a&�V�*�����.f)b���J����=�S.��$�� ��G�W��u-����R�L/�Lq����d��݉���&V ������$�N�_��"�G����V���^1�a�/�E���������+�vu�7�Df��K��b"*H��ױq�E9t�ʡ�Y8S㎚�����0�=�����d����!@��p���xD��e2y�/���F���?D��N ���G@`����,"2�7�o)�^���ˣ@��Y+m�H��t[�UIy��8n�4N8��ZN��Z�ښ�.=��	��KZ���JX�H��;;�#F���rH�/d�p.��9��3~]d����w�Xh�������~��gS�۱�yJհ0V��6��A֯�����ȅ=�+�<��v��[vP��[��O�w^)5i4DvP�W�x9ׯ�R}~���2�b�����u_�ܞ�(Y P��U thv���h�}I����&4-+o��Uv�Ё�������
ы���v��Ӯ�f��L��T�?�^���2-���ށd���뢨t�m�?�z]=�3͝����)fC)��B7��jk����V��F�0����O�\���8z3������R�.��#�R�����%�4��6����ֱ����f\���=�_{�4�!Y��`�а��6ym�����X�@nq�����D�������#�����Q���Ւ��ڕωK��]��u�����Uz���8Iz��U��}�E_�ͦ�YZ妄�s��4�'���R���d��N�э��Bț�D5.ڧ�hvP����bD+�x��z�#�2���#����O1�l4����[�x�O�l�8�	���=�Ѱ�6Tf"�w��e���R��k���e@j�s���E��6�����(N������-�l�w���2�w�7�&Î|�N��m�ܾ�0o9��w�G�	��~��e[1 c� �Cvk?]4������9Y.���L��Z����S$ư�W*ҊM�Тd��y�U+�6;��+)�6�+_{>9��+�mx0V5+U�/��Oo M�@�MP��;�ht=����Iz���}��"H��0�o�Q����#	��T����$D��!.����M+�{�Yf��а�!�"����.�����04rr�S&�wp�	�~!��;gaU7�sCqs)�%\ $���y��r ��xk<�fI(��l}[��"
D�aN73u���Ԏ���\D�অB�c��T:�������i�K,��}ùBV�ۉ;V��������)ϫnV���a=׍ރn�;nw'3l�Im�J�(�.~�#�	v �!���O~ ~���{�.�2{���a�me/*Y�aO��ڧ�f�wJ��Ϙ�e�����Fi�G{������؅�'�������P� N����=}�1t�׳�Y��ʖ�Ĩ`�{z�6�,O�w�?�J���l��a�_B��L�s�q��d�ɶ�yA��u�{��#�����L�������y�ZC9�IDF�cJ��F��U��FG(����^p���>=���a4t�"V9��RUo��U���i'����K�vK���xo)���Wh&|�Fuh�
�#��ag�q��-���Rfs��{��[9�ro�#�IIr�P��G��\���i��1ZՔf��
�ʈ?�⭦u"	F`���t`���~$d�0;R7e5e��X�e_&WG�L��`H/�7՞?LUǃM����ݐ��Jt��)�Ώ�~62�n@��,}K�Q�I� Z�K+�.)��xrs
:
Z�G�����������a
]�/��zq��q_e=�F
5� /��,??�$�t[����@b<�{`����7yg��@aY��W)�d�?ʇ�4��.���M��A{��ί����!cI�݂%W6�.u��j	�	��/�7%���� �p��:�z~�l!�g��v��GJ]��S��XG�kX#gB�	�浇,���q���bm��)�a�knv'������T��8k�vT��O�����t�T�=<��ct"��d?�<Y8[ȉ}�G�9M�RE'(*;ب#b��d����g�=�:߮�|��eE�$mW��O�-�� �%��A�����Tdc�+E`�R��r�j8�݋o~�6�C��w'~K#�pN9.���Ey9Ok=Z�d;��a��)�)w�bժA*9U=ܵ]�+n���o4���ښ�u��N&F�����i��f	~2foY�u�+��w/�fh�ߟ^�o��j�Z��9?�i:���+֛��Aڛ��m�r2��6/	��
��.͇�	X  ��S�ѵ��2�Se����ϘP�����J�Ԏ(�7�.+̎�˯��Q&|�e�A��iޅ�T���6*\�s�M绐�Oo��h�����g��W3���SZ�YE��P�������x�dp��;���No�>����<��X�މ�jy:�����tp���߳(P����Q���@_'�)�┺R�H#��%��}��:I������[���Et�{���"��gn�����!��� �s�{��8�����~=�CRt�o�K������L)_�N�� s��\1���h\�D[r��CW�E8�PLM�ͦ�v����'���|�� �W6p�1�<�bl����(��O�Q\ct�vV�iI���x�,(��һ�F�?8]�q@2�h;����.���fr��2&�`�=��ӏ*#c@��4��Ѹ�9�؅��=�g6���5�|<�[/������<�]�����ރq�s3�8��Y9x�v}?\�%ˣR⾨`1�<����q�-!������RO�����:�����5S����Dq�(��fn�u����2���e=|L:K"_fe�c��$qy��F�do�I��~d������3xsܕg�6�o����Vj���}X=",�e������!è� ���h`�F�sk�n̥Դ��x�C�@����I�5�i֩ZX�W+p˚m�I�hf�orM�to!�B'�JF��D�N�K��(6_��s��X��q}]�t���������_��D��D��ն;TI*7����#D#�BQI��B�翣�}N}C��#p_�7O$ޚ�MU��l�X�d{�b��Dg���X W�-�
��j�R������J>�#���1O�7��i�n��r�l�f�������qDf�����e�?`�i�4�z�Zh�Ȥ���L���ާ�'2�,`Y��92�+(T�hW�?O�lOg�������'_jY�ۼs4&);&i�_r9G5uvFyԨ���&}�F�:�s� 3�A�\�Є�Ѹ)�t
4���I�{��7�)-]/����#uR��3��D�����
���������r:��s�R`�a}�z��@P�K���-�w�l���Tw�t�E{������+*"�w�?Ér+�ڑ�_j�}��se�n��,`d�=1'�
��Q����B��|��׿ERfl�y8����dd����uw��#�Nԓ+�����?&_���R.v�U����T����:?��\O����g3_N,�q�,�����r���7�]�Wǿ�~hW�s�wЕH��0U��X��v���a��g�#S_��"�/�c%�S�Z�v���u�PO=�D������(���8PcG�Ao8AD4Kl�T�v��x�f�h�C!��9����bX
�Z�-+�U�N�/��qIlyz'Շ$��gd���?�C�a|ߡ��m=ӥ�:ys��������)ԗ{�g+���8r����F�~�H�z���E��t�������D�Pe�&~��V�\�ƙ�F��>�J	�2�޼���8��?�T.�/�ͽ,���h3�P����&E-D
�J�5۴7�4��P�V?��ܸ�l)��4`/��=��a�!�-��V
�S�m�W�AT��5���nɇ��ufU�;��h��=��9��H�i���C�l[t0���u}�|����%�&y�=��*����Z��]�M��E����Ѣ�c]�=.?GC�IL��ӳ�i' �f�6ঙ4^e,N����T�f�v�.p�kuv��/3	���,����D��֝hkV���@ꀖ��C�7|IR+�p%&X$
�ӹ�we�K�Y2�B���_a����=@�P[bn�1j�1���f|ʗ!"���o���p��ע��\g�tã��pۏAH�haH��ćh���o�C��}��Ƌh�Ly�aߎd:�m�����(�0��l�-�&�!Q��Ϳ�D��7F���x�L1by�i��y��to�>F ���k���r�(���/!x�y�{�!?I�|F���)��Z�{�8�ah��-�����T�J�(o\��,ax7G6bya���V3�梱�`�`����%w��(��c���Z��Z����R��#����Y��չ�t8w}�ڂ'�H�о��lAӥO( qB��5̩��pG���4�����+�q��h+�e=��g|p(o�~���'���ƖN�u7��uD����������(��_�R������0�Z�PD[�$������G_�i�~��pFb,b{Ѫ�i<��!s&eR+��D��<���҆l�n��i�ЅY��H�&��g�����砢D�����������#?�����zX&��/��j���Z�F��yTn��/P$��l�-�0�|ޣt���,}�9S�~���7�3�4�)�������Q�:K��Xl�\p+N�|	��#m��iYI��;��S���qr�?�#PA8O�հ+�"����-�;Ɂ('/�R�W��MW>�y� �Oǃ�H!�
�+d(Q��"��8/1r5I_���4f�Eؖ�b^hpBףR0cU{u�������$ݜ�3�˓H4z�)扩��i9u
l2 A��w���r������ܴ7jz{�x� �[I�K�^����*�J��8
,�����x�����Gq!u�PA�9vd>�Di3(w	���'	S+�2��]^T��A@���q���C�OpEU©���n	�������Ur�D�Ҍ	�!G��EJ�����B^W������Sm��L҂uNp�(|��Ѝg%��+�a��J�a^��w�xa��]f9.�[?��_L�:�9ز)��-�o���7v����>�k̰_��*��y&��'��ds�$Y8Rbr^戶3&��y%;�5�-$��$TuYCB~���U��@~b���,R:Ͱφ�D0I<�E��iP�숤){�Щ����i	�DI�� n�ߠX���+:͂G�_��s���w�B:�	w/?拱���~���}�@2T"��vX�+	�>�J���ߎ�n�1�lj���ho���9�X����_������Z����|W�J��*��!�>k���oK,��5�������k���CDMw��U}��o�/��X��/�ਸ਼އ���Ԭȏ7��x�e���G�1��!k��"ָX�)+�5G����֏�� ٤ٴf���O��b�����$�/�DÒ"�����ѵ�ѧ��0�q@oo�/�(ް�XN����G�R7�wd&�Y���x�U��i[#z�U��br^aby�;�O����y6:z���ÂN�z���:��"�3��U���(;�@�P}��e��������9�:�¢�,�p��s��k6����
+�!1c�ėn�Y[F�o�;9/���O�	���W�@��}m�ۆcE�
Xs�#?)�,7��~�T�����9M0;6B
�����<��k�d�[��U@�(���@HO#��N���`B �V�z�@�n�ª����5��vۂTuL(��rR�S��%��2���J�&\}r����
�A�K���HgCh(�d��J���|G�Ă�*�yb�o��o4A��7�w?��Z�+���kYQgP�7�M���S��)�lu)�]���
Ki}ZҎ-����?�vs�_�5>�
=��<��<<n$�4�m�69>̊?e���VBgt�ᦕVSȢ�u��\��drO���D�؄���������d<�B�>��;�KƄHj���$�B�pտx�<o����a�}��%TT>�'ؼB�GN�,�k��_ܯ~~9�Z��z�R>t�e��nD��a�v�Z�ԩl�ԗ��T����l1lJ��r�M����&T͡zNyj�A{���IG��p\��Q0O';(e�5���6$�~�;F���v��uI���GeQ_�Nn����G�Մ�C^�T����.�����W�7��]��u
�S?g�N ��=�5$(Ğ^���e���ت�)Uh�-z�;��4Yp$D ��J㻾}ˈ5����%� �D�mjKO�VQ�����%�h�`��V��\Bw�,�}Gw���FD�V_�1�}����ej�����0���ˤnɚ�>W��,Fv�x~�Z��&]�qP=iFUmڢ��f��`z+������a��$%�kQ{t,sb�-�*1Re]%q3�ؘx�/�h�ΐ���;5:��/"!/,�d�{�>����I������a��-46��9Bڎ�i-�o	�0\����d���Jߢ@_�G��3���Ԫ���w����p>��,��c������4�S)24��s���ң�y�ۭ�ӵ���M�<�T�S_)���1	%�H�3cN�<v�#��MaH���1�7�^F�Y�;?�Y��[���1�{���b�c8�c�d|X[�z��:��@ts�Rs'�ݣ#���I�g���%U�GE1�������G�~�*�u!<�~�����@t<�=�/�ܵ$��� ��� o�K��gi�gGJF��7�'�q�])r��L��W��@� �ϸ6�	����_�����2{�w��Z[9�fE�q����]�T=��Z>;;����-�?���+�~->ufx?��\7�r��;z�ǶyZ��h:�g�k����W��Nb�қ�F�U_q��
�a?`�c�ԅ�d
_�2!x�M�*�m&}�\ʁ��@2y�ZƼ�kM&¯a�3��h�����d��vN��I��R�Bi�|��r1wf�~~��W@�q&�rV�9���An�Q�zYu��lk^lM�g$�QݮBmQ�z��w0��)�қ5A8s�oK����R5X���U�����+��-v'/"]�n�uZܭW��J�)
�/6�9���fS��D���4X
�����椪��92����s��C`�e��P���h;���0���	�}��U1,r�#��Q���;��~�ξKHN�(7��8S�ض��9趡��
;�:D���|@"���1E[���@�'��7z5������>oW`�Ӭ��>���f���p,b/��lc��o@ ����pP\��݃�eY�Hy�g�	�/�/Y�R�2>��Q\G��_&$P,b��ia䒭��Nr�e�@�*�2@|�5��.-�΀oZ�q�_,?�eD�� tYԿ��D���,��h٤+�F�!B�T��V�u�<�=�E@�J�@��Ӷ+3��B���A�ۚ��l��������ï��#]ύњ���_�{��>��6�J{D��l�fY�pOn&ڼ��+QJ@��F���#��=�����I�>������B��+�aϵ��0v\�� � 2m�)4��oʡX3�����s<f)�m7x��#[#��e��h���6����c���$�U���qD���4�=��s��}�	�G��Yg�W�pq/��2�lW��H+�\;�����|z�ៀ�3ZFl��n��N+>>����@LB�ij�������Įw���5;�����9
��n�W7�]doR+�(��o��8��2:���ȡ]�p�Q�y"Ql���zߋ�!��7!j2�6N��]Xu�ݫZi�h�ا����cE�e��b�%��)43���a��<�|]1�-Xe���OI��Y`�,)"����	O��rn�s�:Ep������� n��dr��Jլ��v�+�ɾ�y.��n����+h������_pc��rM��2��Z�#��1����[T�n�i��x��}���@WZ3Rg��AG��q�S�aw �ٝ����� �� ��I�������ǐ�8�߃?����_�1|�d�h�/�ɚ�W�1��Rd�@C�Nb�o��R������7�wL�"�֌�̭*��f�;/z�S*��K�����&���8M��2wk�٩�Ԩ��i�F'�Wq�?��M�!t�±����
�%ϱ b�_�剿in>��.m��crq��5���V���!��pɅr�*U�eJ�,*���12�C�P���C�Տ2SCk���({��ߵ�'_�v`< pB��i��:6��a�2�;����(�p�t'.��te�
\9wc';�R�HK�{���"1����w�w�l��3q����]���Cn���1��N��M�ih��z��_΍?	/�$N
�1-dx^y/ޮ��^�ڣmy�zx���s�b�r9���t���|5X(���R6[ϻ�j��r�~��p1H㳆�֠ô�;�;����o��L��[�a���@~rC���(�,�S�74&�l� ��5��-��A�אE��t�X�Ú;��x 7C]�>��F5&���`q�v*%}���>��_�ι���䢤q��(M�?�p?��ڦ��$TmH��2B�}C��/����Azk
����[ �^�KЩN�X��1D��i��a�t[K���T��N�N9�ð����v�/�G�� Q�a�'�^������Կ��֫ߘTM���P�Ӵ���I؀Z%K䷡�Gֲ�~&^�l�V�!}�������k����q��'Xiq��N)���{(���'��Kqw�Kpww����y/���d��w���{2�X噀�2��J��g|�
�ظ
\d
�����CO+w.!�e���,��u�Elz#�#��c~���$�Z�9�zMF�PT���q��� �����:�[A�\4U���5(H4a��u&��������|�4p�4���p+��w"�@��Rb^Z�[�2���mǎ��Ē7�W��4��B,��גr�d��Erн�rW�l����Ǯ�9"v)���\�\�t�4�j�u<j$8���@�uCB����~��p�d-;2���j�ǚ<�m���o]�ϡBNK#�ѵ��q��������*#��Y�����ߋ�[}�cڱ��('��M5'�͝��?�5���Co�uo��w���e�x"�F��_	E�>��1r%f�1<�A�U��S/�p�%�}<���Cv�)Q;7c���bs�d<uZ)QM;�2�k��)���	g�*�t�y�±��ɑh¦�\K��Խ��!�#���p���Q�sM�M�8%j7�@f�m����C�Y,��O6Ibn2�1�Y4�S���>�yB��<�v#�W�xۃA�?�����J��A���s����$��Y�d�m�?f�,ɉ	8$I�heM,�hѕU��I<���������+ _�'�1zK��s����*�]�0���a�+j�e�Aja%T9��ҟk� & p�V�,�;��"����n�ǟ����~D[�!	� ^���lJR�t ��ՙ���5�N�>�0ow�/!+?��/˰�gK�?q�w_yzU	���'jr�?,/�n<�і��<���ͭu�-��,pM��k�nR��X|��M�-��j���J2��b���ai���P�;�W��}��x��K^ǃV�c	"�����u!��Y� ���h�R ���g�Ӓ8|�{���@�tցۏ(m�36�o����Ʌ~�e�}��*�ɫ3���Ҫ���D����S��lk��|jV_�a<�d8�d�!��j0GY�P�-��n=��t��}`�R+�V=~�	�Ѝ3�r<�STU|A֓�eN�˜���Z�}�b��j�\��P�ҧ���NG�W��=�9�z�>���N�Xmhz*ӱ޵�y�B>a8�$]`�ɏdR����pz#w���Ƭ��TEڟ�9
��Y��c�Wgޟ�5%?m�zox ���!���s�|���} X�lЊK{��֢�i���w$�ʐFQ}�QI�=s'�I@�oNjB���"��|��3��d�ݏ;�_%�?��~ū�>�1��Ѱ��Ҥ�����E���g�J!��~+�n-���낽Պ�����`�C���u��I��AXO��?ܵ]3d	b�e6������1]b1S��������!�P��M���
��Nֿgi����"����-/���>^���ςp�P#r�^��5����_��}X5-��a�]r �T�O�U.��N[_a��$.�v7���Y=�iŢ���^��g���t���Ϩ(��aB��!�c�M�e8�$G�����#����{�ge7�
J�r�Y;� m� :-0)}$����I��~�7t�?�g�L�J锁��jV�ҙ�L���Xk�:;�A��Ƭ5����Ѳ�-�K�m��o��c3o)���y%�Y��Ӓ͛^��}���	&.�Է�( ���9U�l���D���_a�m�8<m��9�;p*�ّw�r�w�^��F�'oH6c���r�%)�`H���c%��ݓ����\1*c���x.Q�}g1N
b�D�cM,�4O�$e;ĒK���Z��)�&��fO��v����]�D}pTO�1��ȣ����X�]A[�YI��Po��^��)X�����,��g�9�7�d�:Dl��z�����O'���%_�<����̝o��V���ַl5yZ�f$b����h��X}������y�-�t��p�3js��2=�.7�U�:R��7��~1�#R/���!.�@4��*�-U���b!z��'sx�Ot"��QD��{;�x�Rx�m��'�5^^=�JJ��G>ż@�[�k���`o�1jn=@�*Und�����C8p�X|?�(��k��4�M���_n´���g��ro姄K��u-��. ���U�e�L�O�y�d��̋�l�ݝ|���a�!ͺ��b�q?�FeL������>Ny# W����Uſ�xh�~�7��%\�#�0J�u*�!������Ijy��}��
u�f�Gp�a��2���onSt��w3�,�o2�}�����~��;�Gq�tXc�Ti�ikh�P��}��uw���8S�0<mP, Ik<:�\z=����F	�5_�l-�5���z!#�Zιvז� �r��*#sN_��۾�O��%����XDi��>���mڌt8'[����[����7)����ӊUK�eTD���w�-���,U$�.�OJv�
�084�SL�7�s����-&��+��ܯ��B�\�.ecc|o[5_u����� \���g\ ��S&T:WV�
����$�6�;�f4�H����:�_�wձ@�Ѡ}+�]�o�0��/,�{[���U%^>��XB��\��C���M7ҏ����>��>v���a�yѯ��m}7:9�y�Rb��pMsb�{RȺ?��m�{�k�o�<s][i�w���UCJ�T���!(g6 ��}�(ڃ>Z��NΨL	�,���w (o�d�T$�E��cUs�@ ��I���Ԉjܶ��{��zΰ��|��(G.���>N$�  ڕ"Xa���b���*�W�X�)���P�F�g��qs-������̮9h��5���Ϛ�����j����*����d���|H��n8�Iwu��ys�Y�K��^jRڢ��'t
C�w4ݓ��<giY�$W�P3�����^~za�:�X��n��+R�$��I�E�͋�5�t7dl�.�{�K@�25z�{��lCiAyI��ѹ�+��'�F�5_V4�
B>� ��-yYN&(a%{4@<�/$o9�	4��P�P�q>�č�>��d -����߆�ޕ���W��_%=W���'��+��gmU��T
)�TU��ڇjB#�}O�U^����x��y���)^�|^�j�wc.�g�ᑭ綩RNC����?��#i*���E�Ȏ`ڠ����\�s1 J$E"�X�*�vQS�'�47(��� B8�� 9:�Q���=4�n�z3���\@�~X��p�l��?�XH��$!W~����3ҩ�XM惖�D������h�f��gO�He$�|z�d�FSfD��B���(�MT���<J�xt=L�#Dɭ�Է� ;{�A�f�Acy�����_?��sUy���<~(��#
P�l�M��� G~�T,�"`����m����&d��h�>�3�v[����z��Q_�~�o�r}H�|�;&�x4�=?��#�E�7��uȠkˬi�:g9�c=��0�|��*g�J����v��v8��Ț�������I���gʶdvH���ٚ�̻�s����(����]~����{�
��D^￲�4$�\�a�������dQuW<Z���Up�1A`u���X+!���F���SA��T���	��k~�[VM1e��J_pi|�T��LYd[1'���l�ջٱ�-���%=v-����Jmkh���ݶ�NBw?B*PM��&'?�լ�Z+��;&-��`R���p�rg.%�5��O���i��t�����Jp�r��w#���)���2��э����ڒcɲ���<p£�{?���&&0D:�tL�}��"pԹ�����[�����K$�|e��
�Zx�+f�(-�Lej�X�}�Q�]L����j�b��}<VȊUײDw�*���u%2o�1of6�y8I4��hkMfC'�9��u)�6���y���~B��3���)�/�	TUđC>��>��3l���ucSxl�|�/̕��;A+�G'�͘�qb����2 ������̤{��/`�c�d�9�z]�mt9[��:��̭&I_�M	��a�'�z�,߫�K�U�Tb�����4FӦ.L��amg5��D w���CLEb���T�����
;�D��h(n���	>w=V�{�=ez^�`n}>���;�����o�7�S�p{�<��H��$c���t����sT,��w�+ E\L����$�*RD���%��$��g	����I0u��xU	F4jJ	L�5so8��,ć	)N	2�ne��?�U�k�"��ʕ!κ�"�Z��� 𣲰�T�N"z�'�M܎>NcQP#LeD������y��/�"�[ǳ���%"��섛�a��i�<�<u������Dv߁�$JsY�� s�>����V��?¥�B�B�� 潟�gr�a�Q̺m�a���k�`�B�ₙ����ɚi͚Ꜭ�[�Yj8lm�����F'��=L����h�}����s�u%Jʉu��\������/\�S�3k��S�v$���v��
���p�LR��hl�h4i�7��UL�6��06��]�L�0e�z�?K@�e�����(Z5-���ST��X���àg��[d���T�:-�`��V�������ّ\f���C��Z�Y�=�'9��;.���&R8jE�:d��Dѿ4��*C��W�'T�f��<#K��R���+�~,n��;�r�,�V��O��!(�I�d��j! rջ����,���>=�,#Z��?VH���
N�U*PTf%MH��85�,���H�	(��j�e.�,Ӯt�]N�+���oD���H`Q	~m��5��#*'�:'.q}2h��|figg8hz�P�L��x����z��p6C�w_�w�tK����`��k3��cŇn��,s�U�=�i�R,`1_��o"���^���~�J��=��dSn\��^��De�	�67�D��;S����m?�y�@�=�p�UE;�3e'�&=p
x����_-�>�%=���Ă�`ҝ����SX<Xx�":`�'@ʆ�U����b���{�d�u��+%�g�fmR�\4�KYT���w����
Q�4�b��.F�v|�i��2�9��lT�����m�l���n�ZE�r3
�P~dbaB*桯�y3%'Rm�+�d�a�W�t�S�)2Q�+DOL2�>������JZȝ?(k�7�����q����\.vH���U(9��}�=��y����) ����8w0��zg,J�~���4c>�|�-l�lI�8�F	�.já��I���)���M�V��ָ�Һ�'�8��l�� ���`�4��V���|@_gRYoN����4�#+M%��D=<��xwdJ*�K�}�����W���S��g�^��G��}��-r���*��]���d5ҧJG8��0m[��*g�3��Yn���a�Cʂ�@A�R��w:��P��Ð��r��~!.�?[�� ��Qr��=��=kG30�u�.����LB'82V�)�� �&��ɧcЂ��2V��-��V*�P��}g�yU�c������U��mڱB�r7+���b¢#I͖��䈏�u:_eZ��h�1	m�M׺�|�7�BM)��P�N.�n�����}s������?�*Y�%�9ı$f��o�؁N��l��>�Q	���gq�Z���r�X�:v-@,�� �;n I �%�譢ɴ%ȕ�zL���})Ւ�ӊ_䰭	��d�4��(��ɻ]]#�hy��R�\Na�>�W���o���b|�K,���+�u�ӯ7X�2X��_��ִ"���q�+������~Li#�九0$�s�lķ(m�,ۢ���/זN�����K]����윩a\����N�/$�n�<gw�ݤ�?2��'�!=����Gc��i*;`g�&�����'G����Ǎ����)�GABH����ӏ�xc	�<܍q8�8��*qݍ����������qxĸ�]�q�k��c�s.6>�VO~�.=8��|�f�Y��Lw��]����K��yo��
�5^4�"y�F��N��J��D��M
��R���a��J`���b����&�Ee��P��~�!w��ŶfS��bYe���
�N�D�on���f�{�MQ�},]�ghg5�����8�I�y6��f�y�0�Ӏ����7!G�Ż��S��͊�ٷ�Yʕ�7m�-�*�#�v3zÌ����8��u,[�VB�@����r�,���Jf�ǲN�W1�4F�¾��;j���k��h�3H��XN�u����uƲ�����i�x��]O�ݟ]+���a$+de���׍�^̒�꺤�:[Tj6Fu\�Y�"ԉuoA �3a�tW�n��	��&�>��_}bV7���O�ۺ	��_�?���������W�ec�e��lV���+�X���f<��c�lm(�5%\����؁�����z��!Ժ��$�ѳ"=}�W�A*ړhF c�wVJO*�׃�	�����3gs�\�7�L�ݜ�?ڧ�U.s,Y��9�b��G}��e�g���׹��mD���6���lV�(�lj�U�zoD��C)�	O+�+�,��L��_i�۳o����g�{�M:?��S��X������|�^��ߵ�¶�<����% �".�Ct��C5�Hg�8�;:b��
p���~�4���\��숢D��J��*��cL�������2L�ٳ+h�c*MhU�aR�mIOxU��Uç��Ǡ�Cn��ࣦ���MN��5��[�`�p7��@],��NB�g#��7emq&0&�S2�
.�{"<_�������@�&m��ͫ�_�w�w����$�|Ms#Ӫ"�#qh$ǚzL��U��s�6ᛠ�$��v�u��Q���;Pn����E>�9�����^F�,ߣ>�z�Ѩ[nU��х����I"�X�ty���dj��B�0��"�[Q��Ֆf1�:cG
@ӕ�[aӠ
I�����]���D�`��2������N��+�e\_���hm�d���='��N}jG�X!(�wtĵ=V�ӝ�i!Z��֞ޠ���!��8�_��}8	�V� L�������6�J�I�D��Ϧ���]IG+�Y�iz#���Xy'Aq�y��y������Oh�b���ɴ@|ma�A(�O�H�g��e����bt>�U���`-ם���eY�w'c���v�{�E�W"Z}lo�FǷko"JndJ C�#�$�<KK A�,@EŌ������d�8 .!�r�i��˂�w�������j��>� a���a�i�E���(�T��!V����!�Z�AP��
���5�wI�J�<� ��M�5�whRm���8?ȇC���y�����:i��Mr���%2�𢩥���4X�-R3}��� ���+2#�1	~
!8�hP:j�RK�[�*�iAOpP�[a���x�ӈ7���Y�kC��|w��Ѽ��k��eC#��|
e|O�$J���938�a��ܔ�8�������L7 �Q�A��Y�С��b忾�Z��Ǫ��D����!�ݯ��աQ4^��J���z�[�b�	Oh��֚&�%�;�^��΅)��7Ū�h%�̕����
�G2��Z�0@:�u=<�Y��Z�Q�4v�qw&HHҲ�F��ԙ���I�<
�w fU	d�xU�1��g��p�e0�����C@�^��8g��X\����KAs(��}Wk�cq�3Ed��ʧ�ަ�ެ��AS ��3�����]����n���ޮ��z~6빳B���V��z�T��nMAb�o]qR��v��;�O꥚ӯ7��tL�r`ݳMC�f��msL�����s4�ջ����rb�Ѐ�Uo�;�UU�Q���x;��C�������SY�`���Kdz�`)ڈ�x<)��Q<[��{�o�W�C�������t�'������!��;UJBA�&6
#���S��G���"���D�����z~3Ýψ���B��q�O�"��Y։���@��
�MM���'=��2�W?Px�*�UkV�%	�l�P��5��)�sQۖ��w���>���wX2��!���׷�0�-=��𬚳�!�.>mT:R!�Mb�;��5�:�j25-`�{��}�傉)��|6��'�	'ڶ:j�e?m������f�g��dd�Tn>D@�=�?���F�׈�cj]z��0y �G�[��ٔ�	��1Q�n̒8-k��W����b��S�Մ��.!ה!s�-@g���n���Xrbj.��ժ�F�A�T��G��0Ş_P���ǲlTN�o(MQIIQI�E�V�@�!��e�c^�+Mh�md�����2�'��[�����l�%=ol�nRDgI?V�j��HU���pJ6c]���s���	l ӁP��	�9�R@-w����(�`>'��N���PA�q.ʚP��l�U�-�,޾��>�^�)h�3���ݿ��q����p���_A��,�r�HWM7:�R-�ar�榞�Zw�!����z�{o���ĬǻG�z�W*q�ǽ_�D�Ѻ��)��b����b�^�>`IhvqƧ �v�]���{�yx��T&ɘ�؟�rNx�~0u=Q�߲~��=���S�������N���f�?�*;�8s��c� ��z>�?k幽�^y&>+�^��
4xyx��{�i�v� c��t�7�_��<��Z��R`��1x%��	.��
mlR���RV� ���؁{{`�f��"�������T0>6�\��m
�e\C�
o�t�����n6Φ�Η��Ex3���v�A�������V�;WcgoY�ﲟ�����3�f��	�<������
*�&y�I��RS��s��r|�e`�cgd���U��FBO�a���D��GB"�x�GN�NE���p��' f��q�3Wj#0�6�*$�ko*�C:��,��GF����3�>�{�ڸ�s�<�o�`�.�/�8T܁�e�k�� �����L�Co��νB}06��T�P��j�<&�K��9�w�B�[,d8��>P�L@�7e5�4[����8A^ϗ=���GP_�	+�e3���^�s'Y��HWVg�Sf����4Չ�=! �<=��x�|����F�_�����$�e���?��ć9�[���7W�A�S�� C\0��3��V܀���Hm�ǅy;ٝ�x�{��P17x���V�< �w7R���Pm�����r�P���)��kq��ú�}]E���xx~]N����k?>��=_����	���r��ؐ�Λ(���~	�=F�Ҕv�$z����_Μ�Ҽ��Z��?4��zy�|�������U�b-�{�g����J�x�����x�J?�OKpb�-f�8^?�y��u��9����t���+������²_������jˣ�=EO�!\�_�~��T�I�L��H[��f�5���LN�I��C��>M�B��"��+ͼ+�l3�5\�KVv�<).���m��J҉8��wt̓D���(���^K�c��&�r]05NU�`P�f���*�P�8��bff�?#�0�3���lU۸jL����C���ⴼ��Z;���{�"p�
�����j	
p�YJ���c��뀍�aM�_��jwl���8��hY��>8�1B�͂`�+b��-��I�(C��WZfG���L�$��$C2��������������?�8��g������%������@d�ޮo����z�� �E)�l{. |�x�O2���[�g�6�E���ܶ,�	w���/����z�L��3e��K�����D�S9s�Mjv|sx�T��*�P���:O9������h����*�}:�nX��o�]�E���h֊���A
��&��u"_�ǪZ��]�
�UkY9�Zl9D����+"�'�����r�[I��R.�>s��&�*+��� c糹0hb�l���M�-#g���C���3N���P�8�x����T�Nف�K���g<{[��T�� �?��^�,���� �g����;��S���j����Z�aw��8��%xW��f|��	�yb%NLn~'oq.,0@�m<nم]�5��tX��8e]�RK�8��<[�#U��r�:�3�c����}g����	���@���Ȫ�ݐ��S����y*�N����qK���	���gu�[�s!�7u������,j����D`f%د��m��J�=\��G╷��r�$��A�%��x���L��x�[&s�kB0'Y2*�đ_̲��D�	�"}�팎����5�tv����]֙��,-/#�@F����0��0-�ݘq՜��>==����jE�V�ϻ���{��E�7
��I��(I���܅�5��o����������B�.�'B�H�����U|!�zd�:����dϗ�[JO[g�uQC%�Vc�`�f~��Ao�+�ueP5-�I<
�䯤��6�ت���~����m��|؁	��@�(�:��E�D�Њ�@Ą���^*}�_��C�s���8�vAN�d�08P_�d���{�K�J�<���D�q*^
�
��+[���lU��~��[QuZ,E������N�L7 7����s����>C���r6]�Q��kjNs��A�;��bC��:���{Nç�$�������e�L
����1��.�nOpY��Lb;�n���y	��Z#�}�F�/ق��Q�ǿ_�]S��}G���o��Y�?�ik\lu��:/�k�s{p�a+���������rq�4ⲛ�lc�e�M��;$�7�d��.��^)ω�cүv�D�o�@���s�������C���u��h�T7��׏S��x�9�}���;�XXZ���A�<��v�Χ�G���1;�*M���s�'
�Ͽ8?��<�G��>bV�,�#����i��⒵�\��rVA��j9�Rl�
GW�ʮf53����HD�q���l�$t��VV+9��H�Ɯ٩��F��ɯ�[�ヰ���%�m��i%t���¦�R�t�4{�v�8�m~�T�A���4faE֥%@ w�U5��c�h|^)#�!� Y��f|���)$�%2��h@6fFaf�σa���3�M`.��.�xϥܓ��$��1���K�@W:�.��@���^��Y<��,����Y��A{K!w���5[	h�쬘��=?�j5M����s�slop�^�lã�{g&p�c��b���ܤ��NкO���.4=�z��$�[�<��ᨗ��bO���J.�92��F7��ZT�C�wh�8򑘁����_���Q�����B
Σ��rO��4�&�"aX��Zv@�qi����^�
�����.m4YȈ�z\z�Ri\,A���F��!�U��h�o�o��£�Mv��JA����[]+��ߧ�	_2�B\�Ū�#�_�����7x>���0h����9�]�<e�I9�)�(d��fv���d��a���D���{$�e��3 ��6��������>���ir�(G����ԣ%s���嵹��}�#@Xh�q5�A`g�o�ކ�f�� h4��?T�c�#'���J��&j�q
��#�ݢ�Et�N�2��h{�0�u\k���r��v�����#}$x���M*���V�'�F\O��z�1��Ns*�O��^�ss��ը��$��p~�ٜ�6�DƐ��T@�k��~k�vNq\nd��9u��Y��٘5:�U��o@A	�)1���o�ˍ4۱��e���M��?��Ƭ>�S{>��ܴ������؊x�-���K.���]bD�΀��H(���91t�v�̀ZΚ�<Lh��(���Qm��F���f1��r:�rv�$�/I�|�K��*��[�Ăi�������'��ϧ�O	)>_��5�h��#�2�����`�bJI�Q8эm؀ָٰ+���3?�����`]Gfk�pb-`s�?d���.Eo@�m��ߙV��"�XH�P�~��SUU�Аpw�Ѓ��BzJJ�OC��!�5TF6R᛼iU�\)�fu\�
N��&}:�:�@P�4�yG�W���?��5x���!��1��C���F�)���>0��~�8�6�h�(^ǧ;��6V�������<)>������x����*��z'MZ����kbQA�.�6O��K�`p�J�[�ѽ|�oe�L���#�M�R-'���>P c���*MR;W��,�]���ر�Rhx��%���!�>�W��WiJϛ�],�N�����^�/z��`�<���5����&��P�$&Z�b-���^c<
9)�^�YW��t2?�R�����C*��"_l�VS3�ƒra˪�"Q��zǄ!!�~�"y�l��G�iJ-'s�s����&J�wc��1r;I:M��V�Y���P�Q7��Ce��`�5�f��0�M���OU�8u	�?�4ō��O=�[��ٸ:h����)�tX����B��d�>�cj���y4��i{;�d��'_�3����&�7�چcX�niAG1G+��.�"`¶��i�c�}��,������\x�I����q\��1���Q\ܱUb�#��Ԡ�ޜ�su��#��j�(~����a-W���Dk��\���Q��j4[�H�ExYbt=��e@����d@�3���r���^����k�K�?R�t�҉*���9�7��vK �vX�������?���1;Pr���}�{�e�����5���:��q$�Pd+�����ď�$�c\�;���s6�F�ޣhY,n�(��`[~����2����hs��12%B�����������,�y|D�X�튾�(�\[<"��(&�21�u�^��9W��M�г8��Cf�}�������/��Ip@�ʖs�$���M��l��_�wcsj2dԇ>�$�#ֈ}��� ��ӱ#C�f���֊��5���҆�w]��y��
���M��e�r�R �GU=����(��NU]e��Ƣ������di�>�K"���E�l@d2�i�7��}�~�#6'����9�q;�hmU= 1��̤��Ï�.��9��i*MfI&k��F���n�[��Q��]��'��ys�p�G�Fzu�8>¯�[�ڗ�p:b���f�x�u]D�x2Xj���R w _)��r�kՂ+��G�)�^L�����+��!�,�G�����W������'��4������[2�Oˁ��%h��`�( {ȡƲ�cf�Y�@�������f�����ɪ��[Ѽ�u&yWm��7��X�"�����F���q��~�d��⣻��+^F�JT� ��������W��\�K�����+ʛ�󋲐�=R�O��/?{���$�S�3�;��x`��ZǻTt\tlG��a�R1��[��"�G9�џ��
���a��5���JU�c5��5��s��L7��b3���K���h�����Ji�t�D�[Pm�������Z>��u���Q���h��:�ft�\ʈ��L����SlW������#�5|��ʴ�u���naPH5���6T�q�MTLK��0ύzH�T&o[�ͶDT���N��z��a�v) f�ء>xܲ�^�l����;ObAk���s�08kg'�g�+s�����H<�SF`�A�~{沉1���d����p!h4@jMsH�y�eV����͈������r�;�9iT��&�/Xm��cp��X_�*��z�>$T�?���W��6q�JO�7$dj�!@��Cޘ�Z9Z`�=�����њ���ܸ(�Ge�ϡpk�wt��i����M���f$�G�?�]i�x:��o��
�FGc�s,�n��� �W�X��R��BP����P�4�\��rZ��!_������(��!7"u�r�g��y=��y�;��yT��i/�������ɉ��\���'�p2����e�����9�fs�P5Laf	
-��1�;�D̯�d
wr�,5�Ϋ1���I�i��#��n�	G����h�����K��K�����1���o<�A�{�"|I���#d��4��D����аs��Ӱ0 ��ث*�x�������}��ˡF�5*���cXqe8<䓪?h��Y�sL�I�������(+�����t�#��P	�[���Y�'ڗ�NԿ��&�"w�&h����i����f���p|j�+�D4�5���J#��:����+�>}E�3��vZ��ą(&����v�ɗ�;.��@(�s/R�<��
��A@SŹ����\�0-	�~ӫ�[��+�a�X�I���Rv�N/P�ph��n!� �
G�TP������ž���Œ������0�zG�oh�-�c��4S�v[�����#��eJT��8�o��s �����g�4ȏƀK|��p�B ��`| ;A�-���3�I�=چ՜J���G�,�ʟqt����&7��(x~y�1=%t�.��!�>V�.V�V�0��3+MP19��z<.`�Y��W,z��J�z;�I&��5�|����|)h�b�Zģ��a���w��<�Ϙ���utD�M��G�撱ɉr����t�� [�ڡ����d�a��{#�z��0+�����Z�O#К�ſ�4�µ�7���X�Y���S����dɂ��w��I<Y'7��'.������H�%� _��nt�)l0�f���P6ZrtP�?K/1V�zb=�>�c#���3�U�	����toD݊����,a������z�ܷF.7ҶH����^p�'Q~�����}��<�*�5K���A�qA�k�3��n����<Av1�FrHOM������9٨n��֖g�/88GL[Y��[�B�`8*�d��w�l�F�i���C��N0�����F���,�.���V�2������f���� gtIU�lz��xtJ|�L4u��G�_�?���4z+k���f�� o���Jo����g~���}d:�w��r�v�.�iü�ό���>=��k^�r�w��Αi	���z貔Y[�ȁ�l (�� �G�HB4e�D0���O�g6ۃ��T�����#�K�н��{O��%�Q=�&�23r$��'GEòx��U��^���]�ZV�7���/��q�4*�BA��}�N	A�4V��c�{+�����	f��D
B�}����Cpm�צ���� 4^J�W��bR9���,`iE���%4�5���n��u�n�� x5�>Y�7��|�` ~���Yϝ�.�����IJ���}�޸���|±�Π���W`���] �Gn$�)X�M�*#�/�����˒P!��Y�-�8�o������F_ΐ���'�
�4�g�R�%��`�e]��g��F���uw��ƭ�E���0M!�k}c���#&��dg0q��q�Xګ3]OhჿyW)����,n��vua�7Pxd�A��/��Y�y4b�`���6��,Y��Uh��S?����>��R��\2�����ys��� ���֮�)�����wb!(�s�Ю"1�=J�{��m��wXzf�b����0��+���EC#��^�G0�| �[R� mZ�Ĭxy���^�z�ݞW��;�m���,��t�%�qHX!��-H+)�q��w�շm�55Z��`)�8?rg�Ḁ<�BK�T�G*9��S�I�N ����+B�\"�����J� ��N�{e�	�uBK)�?��m�H�V[��hK���疀�Ŝx��܊Msj+�z�_���Ԛ�����j��2>�H?n�H� 5�--i\ �Ykc�VM�TQ��܃�$9k�����`����}^C�~A4x�L>�[�����1Zh ��3F�����_���S�S�żB��� ���\�Mj�w���|<=��R���̡P���۟�}�G���J�06ρswR��$O��#,���L�Hf#��-�x�$�SQĜrK��+-b��`o���)��1�J$V�1:ngD�c�@��هn�:�V-WŴ���d�6�׻y�8�YjI?Sl L�Y6����������o,<g���5rr�!ć�#��4S�{`�7V6%�h���$�R?��vЦ��� �9U�ѣ��W��wx���0	3W��2Go���.E��9SZ�bk&�����aՂ��\&`�2ݔ9Oc����M��c����֥�e������
7��߬X�}Ke�Imm�2�իI<�Z-K�
��	b*��O��"Y������l�����V
�Kr	H���ݟ��5�|���Uq�i9����˘i���|j���sl~�O�GVX+�y��\����}j���H�b�r��$h����zG���HF���k����"'����F��S�.��V��pϫu�o�0%z��k���T@��S dgEv�w؁�T��a��x��b4���%�!z�УZ���AT�B�wb�X�)m_u��B����a�,���n����C�R�	+�Npw	���n�-��/��@�K��P��|��I����{e�e���R8e{�O��"iT1S������kgf�c���(2��Sc"iiL>�b^�ٻ��w��L�4��f�4���b{w��VS��cd5q��GsZ���d�w:'�	5;ʒ����*����O�?�]lסƶ����Ԑ@���@���	��v�jw����smg�:�F2��x(�y�=)����(�O��)/0E�:���@{nE�'�=�_�/�k�K� "�5q��a�ƛ�G	��/�Eܢn�7�1>���`PU�\cw�W�C�9�pB�RI�A.�C�c���K�aI5�P�Ex��%��'�k�6�0�)�(xG�΃1�ڄG�DD���c�E��I)6����x��KGdH.��s0/��Z������7;��h�g�$���iW�#0���]/���y�RH�?4*,�,>ˑ]���wF_�k�����cg��e�NN�t���"9:Z�ձVV�d��j�����U�Y�����m���^�c���$n��V+�i}l�ҀBk�q��:�R6Ԩ���`~�k�c��#���_t3;[�����w��b�8F��,�?9q]Uw?��_�X)�T9����{ʁ$51%xX��,��j���ew�3"�r�)�v$~���#p��߅6��+�a���)��Kh5��[��P{��Ƃd��}�V�+n,=�;���qm0\!��E`�Գ�>j�����
Lݏް�?�t�9��6�,���sq�u���59�P	!C�S]��9{>*�}9�ox��hx���2�g����Eݽ��2+m��6�q���?YB?d�(l�N~C`'���(�q��1}3Z�2�F�l�u����TS+�K"s�}G[j�ӛ�AZO���l��UJt��Dx�YG�y�2/���o��ds[d�S?����~�
�K�8$T�ȳ%����\c`i�̈́z�k��И�f-x��݀�sE
U�B�Н�ã���J�����Mh����x��L����&5����'�Z�[WI���U+�𙂨S�0<[���̀�6!��-�h}c�ki�^,��K��e����+�ͯ);	V2�J�Y�6\��-@�l ���o�#�-f�(ʿ�>ȕ1�DptAbg�_���&^'|!}%B�6����^�98B���F�s�P�[��p#&Q8�ҡ�Y��b�hGN��lxA��;H|8�ƞ��gRk#��"�;�CTt��qG1,K�%�r�L?R���?��7�>��W��緳9��Jd�i#0��������L�q1�̓V�?-���㾣ݍ��д����ì5�ۅ���ǋ�NW��}m���߯G|�g
������<=6�ۭr��Qq�yK�7�pL#zJjt�ĘI+f։��T)QK""����	��bǫ&j�A��L��Ok߈'������&�6-C>b!��ʖ�ݪ�X�W�'d��`��/�l�ȠU�{��D��sp����,�Ύ��@����X}�q0�0��n1N;h�Pl�iLr9�\BR�I@�oK�Ί,��0C�=��Β���@��kc��+>��~=�ϸZy�n����U�R[�z�e!�
�oU0�Fe[�,4����K��Qd��6�a����5��|++ڙI�L��q��Eو���j��\�p����v�6�$��yU��(-t�MTYP�a=^���1V��n�O����
ݓ�ݓB�?0��K�&sXTZ�\�5m�3��-�.5G<Ԗ[[i�3O�*52~����iP�Uvg-���w g^�nnV�
��.�E�`��c��%
F��0^YR�q|�T΢��whь��7�h��u���h��HϺ�<
�}�ѥ�2�!�I���UnT"�c� �9�y�+q�J$�X��@ �}r8�
j�'�߫-d���w����*%��͹�(�uuL��d�Og�D�������xch�
G��i�˳�.�yT\t�iY��2��S-'2!C���fVFu��k�L<��@�k"��&#��򳘻����U���$G�Xҍ'N/"�/Fn�"N���3�ɰD<{�
F��m�]5���gV�؝EnG֊�^��z��;�>�1�oFn�jQ���E��e�8p�5��R��_�4�����~�*b�L	  ��a)�C��s�����o^�����=rfD�6�QG��-�ѡ��6����	�4&^C��Iq�[�*d���z��/�6`��V���J��oJ��T��x�����l⸁?xܳ�1�u��;&�\�<;@��9�����m{{+�}�?8�=[9�}��M�q���O�}��Ί�ʊcG�C�i�����`�ZM$��I&�6F���?\�B�'��=֫��Ǘ\�J�ʣ������$=Q.G6�yg�+�/�3��N�GO��+��qkA��Ǔ˛}`0R��kJ�n@<]��oنa9A�2�3a;͆��n��o����ڂK��,h%p��c��o�?yZ|���oX���-�<���S8&x�.�zL�~d�3�1ÀGw��>W���G�<����q�Em-���EKJ��������!�h[�&EG�����[<#�Ś�ӌ97G��֐NL����>����}. �q��b>?��K�ݞ�����؄j���i����nV��R��C�qJ�U��u4u�Gs˹�;����6spew�Jl������۲6��-vֹ��I��5) �	�"\|.y����p��mC�&�eM����n�N��]��I�b��ٌ��D�1G����\.�VÜ��6nǵ@�	/ǟ~�?,z�g��lN�uj��*�W4��:�F��k�<�ܬ�≅.�).�@�O��j{J�H�l.��}�s��Α�j�fC]��)d�N7���h5�y�n�ŰA�9�`a�9U��C*��mP��!�ld6]>�܀=Yަ����P��	��L��Ȅ�|��[��-�$E �Nȫ��#���_}+���D^�L~��L]�{RHĕ@}=�s�H�t�D�?�<��{x�a�T=%�IÕÞ��T�:�d,kpږj��Ȥ���譥�dQ�TT��T�-2�ר� Jo��uT7�4���r�b*w�Ј�����x���A�̼K	����˘�h�f�Hh{(x�iH!X�è��^w��4SI֗) $.%	��sl]�t\������Ni�ۨ�S4��lW��v/�$̤�et���<�څsUJ�VK7���`4Ih@����?�󪶔�W6`��Zs�`�<�x|�J�Q[՛?���C*Aފ�Rj�4��3����5T�8�RSYUb�U���R�i��%t�'�h����s� ���P�q�
��`�67��>�ds����	T7����EJ���ɔ����Ӗ�Vl:�פ"a����2D�$iԨF�RKa/���j�V�.��ÞB'&#ȂC��fKf�B����x��'n۩���ʶw��lYr�'���d����M���(�i�Cu���l��cQ�_]���
N�8��[pL��7��N&�6��[�מ)��,�ʒ�p8��E��؀!2��Q%�M����K�H����j��ڻ����/w�m+�A�m����k��~NZ�6�)lS�a��8	|
cy��Q�o��k�._KP8>��&������$.p8��Ɩ��V>l{�����a��vq�P��Q��D�)<���P4S[Hݩ��k�k���^�S2�<�1[�>N[�w�>|Du��Æ��Qd���ipV1��k{ڧ���?_����iӼo:L�QqYs��r����4<��7J�;e�AW�>ڜ7�����W����{{Q��Y�� w��4`���#K!��~�
$Y�+�h��P^�T=kYï;��	����H-��n"tک/��b?eY/d�mԯ;���!�i�����:�{Lj���%0�@)A�������;˛4>����$�CeR��&�0ruSR'��K���8cb��?�]m��}�{����� ���${����w�x�Xb�?`BXY����T�@�����K�L
0$�lm�D)�ۆ*ܴ�_���"N|��=����G�w���q2盷dd5�Jp�+9 �}���
6	y�-�BԲ:]d?�Se�
���<p�
FG^б_��.��og�	1�*���Ɠ;Ǥ�m5Lc����D`���%>�� r ː"\�͑4nꏖ�_�� l
6�Ől�	,�v��z}�J W^��^]1�{G���"�{Wt�����&�n$^�2�k�:?�<P��G��G���Fv��:�?N�@���.~Ԃ!��	�ꮄɍ4u���-�?M�>�˾{�'�E�������{�E~�z�5��zg=���/Q�Y/_�/��8W~p/�y����+C���o,�Nky0�-�*K���j��$�徙��ϝ���b��:�ȤG\b���I��-·^�s�R��pp�a ��?�Jl[I�,[�)��z���
���r������-��'u\(b�[��{��� ��G��~�^#����d���J��a���v\@�C��&��un���C��$����J��O���6��Ϟ�w�'w��#�r��XiiyYi)�Yӻ�%u�R*'�ԫ�ED�Lt��¬A~�R3iq5
�ϏFu%��Ռ��Ж��"\�Rտ��n�t�q�:Z��x��S� ��q���ٛV������$<��:�%͔��<ú�T�}h��.��ۯK�� �RC
PQ��|�N3eS��21%��|W\2����ĩ\���ɜ�+?�i�t�'�{��5>��q���5|n��i.&qd+<�"qdyo_S��щWg��+=�q*����9����NU�/�vU-
6x_(�\ zM�b�bp,d��PU�{*2J��[B�-�_|[0R�g?V�<�J�Q�\w�l����	ۯ�T�1�������L�n��Q���hd�vR�S/Z��� �񥵴���ym�Ԯ�ٮ�}l$���+��7�Ct@�?s�j3HXPڙ�來�$Ul^ ��^(oN_&b��`%<�;�F߸�}Qc�aZ�y�ً����;��nǶ8?��g�t�8>ݿ��|���o���V�C�*4��t�{�2��B�j*�4���	w�w0m?�4�,�u^s_��L�>�����zu:�ճ?�+���L�a4��*ґW��c���	��z�B���֠���-c-�˗�F��?����C]��O���Q��<E%��ě����7__�D��7���96y>o;���[�xS��a�ߔ�
vr�CI!�������+��3���3��7�b�R"�뎑���S��{� �>+��dy��o���?J-:xO���I����
=��5�������pp'�W��#��k`4f�FQIZ�I�\�\^�̸�Ó��΃Ϊ�U���o::��a��Bᛶ7��'WL}_u���ҫ�OѼ�$~l&~h�hRy�r����oa�h�����n2*�'�?��@Źk/e6I�Ӹ��D^ũ�h��
?i�.��Y��EYj}�+ffK�W�����Q�@�����k�qXdJ��/L��{	{�p�Ù�����^َn�m[����Bc���n�;�w Px�M�^��J.��p�2U��vDh��?��nE�����0n��K���ǋ-����7<ђDz�t���-��z�:$�c����oW�O�V�c5�\:��0���GV�bb�"췺�J��Hk�_�E���xhn��ki�{!~EšQ���Ok��2�����gv��|�Vk}=��/~�Ǘ��s��F��~����l�jm��\�[�1x�1u���?��n�׼�%�3���F�����$aG�<�'�}�2�}꟥���p%������T=i��y��1�1�nH�d����1�3�N��j��K�O�scc4v�4 ;��ҍ�N�U�\Ү1Lw����5�O��tJo�K�Hp�]����e&�l����0�U�>���������>gp���_*�z�$��Y7At��&�TƐ4�HT��/GF��	�6bq״j*f�k$}b��y�r5V6�b�w��|�����0��gK?��`ז�L!�X�t"夏�������]6^���u|l@f��$D]c��tQ	�u[�͈A0���g~�	0P�?.����q��Ƴ,�ig-�C��C��!z�ǌīq<	��dV�������R(��>��!bQ�e��1������-������r�N�#�av�f��:єg4�l�h[��E0�y���#\��}�I>�p��s[�6�SCa��;���~ֳ���mu01�����ܥ<k���2��M��voKN:�2V�3rL�=�̥L&r����h�U���h�5�Ԋ;��K�``ݞyU�4 �������;�0-�(4JѠ���:Y��H�]�G�Č�Y5S�������)��a=w����6�w��U[�~+�^���^W���V��.gbgbı��*$6�C�744��N2��-���J�a���z���I�Z��x�n)�:\�\�9�OE��cXowW%_[C!���z�m���O�գ�Vi׿�cs�3MK]��E}W�?^z������.�D��:
��FFswi$�����>�R5(���K�%.��py-�f�B�*��޻�R�u���]��4�V.���:`%�5A� m�^3��r�o�?�Dm��E"r7 hK	� I�y�k����줊�&��:HPh�ź�~���I�T��
����3K<�)Q����!�9���[��[ѻ�賗�'~�ǵ������]o�n�ڒ������X����~�=�v0*��������j�T���r�CV�����^5Dt!|�E�y��薱U�k"խ�t"�F�#���d-r����8W+Z��X0�����ɲq� �?9������Hy��/�i�0n�s��C�T?�#j4����(44��\��쟄OF`�I��;;���[�鷛�^;ύo^>���<��P���~�boi�nk����o��?����g���R�����B���GI�����C.���[��BQ��9"P��g����c.D���P�QF���,��#x����:>;S�gb�U�@]*j��X��
1�pZ�Lk?� �9؅0������m�17P(|���q��t�L>�fA����"�P��뭢O������P ���C���VgC�n��f��rW6��Șxy�B�H�;����H|c�$
����s��/[��o��atg`�ԓo��da1�-�ue�'�⍓��o&�+�W�	��	��تGo�O(/�7-���䭌U��y�gs8i;r��T�kU�ذ2�;���Df6��u�Z�Y};s��4ZS�s��~"]i>���}�V "���`(�"��L�j��3�j*�lJX��B�+3JS������B�����9���-���D�gu����{�\�e�<�ڍG�{hޘ�눤{�C����߾�V��X��7N�M#��ig�0�/����W��:���?&��a���+�ެ��#8�-�K��p=qҁ4�D�:����|�udX�U��r����o���M��۴���t��M�x�0��ɫN�p�XXw��Ҷ�RB��w]%=���W���a�����q������gjAq��Wv�s[}���a��:�UG�n�����[Z��V��-���+{f�#R�;yw5�h�����s3�ȃ�r^��>!n��~��3<�����������뭴����R:m�� *ɶ�!\ޱ�r
�FŐx���[<�١֓Y?���.���rN��9D��N2a?*���g���$� ��������U�	�
�a����x�G�\CR~u�&	���7WE`�Vs��t�<����<Z�5Zl�i�h]e
[տ{j:3����,b�\#PK��28�0�vd�k�3Ю��ǵ�{�t诳,bg��,X��	4��꺭$��uL�j��U�YSyS/H�1�����B
x����O��۞#�Spa�J-�vf5�Co��J�a���݋͙h>�����������_w7s���=���<҇���%r!(b!������0Ok++�X֟�	���v�=��'��}�6^�C��~�hKz?yl8��p�{w� G�[�r���_���嗗��������x��w��Fp���w@�&I������ΟYqf:K�yB�Q@<{��K�鶋	�udk��T(�`���%���l�a���CK��r	;��Kpa�J�����*���%��%4(�.9C%�b��)�ؓJܐl���u��Z���釦|N{��>�+��!��~���io?��e2�x��%[4�y�,���,��m��ӎw�������m����'��nE�i#o3��~����/VTdMŇ�O=�����G�zvn�l-�� ���Ok��t��ycC?��I��A���17[��2��	���镨��2�D��4�H�s���� ���OšH#8�~�,�^j̗KܛD#�4��?��55�N���$���o�
��Ƕ�]i���}w�b�]��uɆ!�Q��SO�b��BD!G��́���~Db�U��C�/����N����B"U����!Q_/I�$���|2)cm��5P��:kIf�� �����ѼԼ�\χ��mUJ�0'�����f��߆�3i�g�e��p'�/�<G��a�^�#`���|=�O��e9�1����\���g4�j��h��*�F?N���H�����q8�8�$r��rVaݙ��X��<j+_�P���օ:kQ_�� >��򼏏dj�	���(wz���F�t�{�!6��|�U&�Sj ��M6>���>����I�I��DT��=H!m�9�(ݩb<aCk��$������0�ɥ�L:��Vd�2�ٲj�!���ĕ��F���{�Q!�3�G7�p��#��Y��ݾ� �UH��X��Z�T߭��Z��MH�����u��|��-�}u����t6cܜ��(�I9��Z@|:`��?zH��Z�Ϝ��ܞMw������dX����X@�<ׁ?l(�t�f���|]�h��>��2[��vȋ����.�-t��x��1��a��Ц�5���D��CȮRh\W�q>��w~����3���"�:5�>)ޤz�4������;^,��.�+K��%�����?GLi�F�<c@F�@��cZ�rk ��!j�KK�.<)J��`U�F�S"S��wq���"U��e(3�΅��:�!�d���g� ��F`��	׊Ԃ҉����pD���DJ����w�0� 3���2��d�,[a�GO2��ܜm{d����8�ό+������j!�[���1��y��l5���MSn����z�]�����u���B��/w���$��kd����C�>(������g֫,�.�Y����V�r�^I�R��h�f3�$O��(wp�˩����*�
u�Ŕ�[/�[�l���U�}�x~`�Wɓ��.\��C��؎�Q�����})��2�"�^�Io�㎕8.̳b�	�j��,"X"�m��q$�����`�ub�=����D����P	5�4e5�`$�L��R�*�M�+Ѹ�G��QnY-�ia�rr��R�ģ�|j�6��|G���d�l8�:����}`��tΆ�σ�_ξ4�;������]}�T0����r��v��
gj��
�f��]n2Kݿ��G���_j>nw1$�^�PN	y�����3���G.`��7�� �S�HimBZ~mi�;���^�@�;Y�x����U�;�R��B��`Fؕ��J�X/Tc��zt�H����[(B�lf0vMו�κ�+�tN.b�Gp9m����%�#!�~�f�ۓ��}��n�W�LޱV��U2���C�},���h;�L������Ǟ`�P-͠o�ݹYQ���ѬF�C?�9�P�̅뀳�X��aL'�wF��G�uX�լb/ZG�����t����:.�'��;�`r�JLg1��e��2���k����ӵЗ��ǫ��}����?�jXD��7�}ɋ~���o�%����5_g���`(}�Ŕ�:�XvP�=�N�3B �j� kef���3�h8�:��j;�l ��0]�iN�'��r�����	ۤ�t�
��+R�_���^c3��Sxl�:)d�<j|���(�|k��?��FfsH�D��-��+�m&�D���^������$���uqyXX��=�]�����q�������3����Pf�ʜ��\
%���F��8���K΢�;���ϻ����l6�/����g`��9�{�C��kWT$B�o�5D�o8��%֌!�����c�Z��� ;�����0�Jz$�X�2J]���3sb7��=���O����y�>+,U���9_Ys+g�'�JFr<��7�=k\�E�"�q6��c ��N��>���u�����D�l�5�/����s|�γ��ԗ�~&F�g)���Rt�)� ��Z��V��2�,h
�΋2c/��,+n�����<��u�	�[��B\�k�)SB��ud"N�q+aa���i�};�!P=l��f�p �",��Np�+�b��C����0LF۟�0�Dׁ�o�y��������*������6y�o�vҹ�%i
R��@Dن��ѱ�a%!�W�p�FX(��"��W�r�W�� 
e2WᆤU=�zt�+T=-����4�ͤ:��k$�u�$˕�����ÿc�A��[��>�F��{{��/��6��f��m���?�Nky8��f&#<���$�^���l��p�x�2�:��#}�'�5�m�Q��q�,5�(kr�jr����#$�&�G-��h��k�|V:�H(�n�!��II�ߠ���Dz���-@Ȼ�����x�T�[�8�1>�S��E3�λ��,�kw��pgX��Z3�����o�,�2 ����`�'jU> zB&F@����<X��� Ʊ�΁\�� ���Ȏ�]g���${s���>+�I��L�6�͙,���/)=������'ʈw��-3�p���2�DH�����'�'��I(�At�#򠲺�n��!���3
v�E4U��6Z��9�qw| qT���E��	4�����i�9d���B���L�����dB��DUe�cN����V�4'�?N��1�ܥ�ET@�]���B֩XU���X �����������g7T-A�@K!I�R��^5j{2��W� n

4����8/��Ա���I��5;r����׏<�hmٰ:�ܮ�!�o^̾df����q��|���څ�aFYt���VlQ�+�q��[k��
����kI^�SwFM��ּghf-3��rOjs1[zj����{4��=/v���������(o�pQe@e_�$x�f-�nL��Sh	����O"ZhBlW�p9��*����Ky�Yۈ����v:��*ʒ���2��≽6�?|5�V �OD�3(�礄�.	��%.�n%�eỮKʃ?�c&~-�,����(��^���D�c�Ek;��[�ywt���\��������h_�.�[�ͱ��֟B��3�I�2t�>��Ȯ��'�ːG�����A�{ ���8]L���WC���).Ɨ�g@Κ��VBP�DF��B+�(܁?
qGd~�DC y� wwgT7��ה@�����$��&�a�ὤ�̗��[S����7�n�όH��~�;����)��@��EuTff&����������@Ӄً3�ʨ9^Sp� B�-�_jՓ��ϱ3�Rp:��WAq���@=#}Y�> i<E�"�l-���0LT4��(J��Q �LL��Ʉ��ӓ��~��$�$�$*۟������v�Z�;�4��a�A�+�l?��<-��XwЮГp"��Ko��K*��� ��
� ���tf{�oy����<5j�eS�prρ�	XN6ݍ����FG�̘�F&P��z�b�z#�i��Z�9bm�?i`�b4J�t<����~��b��j�p`�o��\�щ;E�Q��%�ļ%9��!}�IjkΊ]�ؠ��]w�:>Ҙ:�k~"%���	�F.�L�qX��1r�a�g�<h����GŇ��/�X.��m�B��U����<<�bs��|�BV~�{���m��NƸ[L����5�խ�;�ޞ����}5D�j�@^�v�{�h����p��b��5bu��4�"[�T���xqk^���R���DߤG0Q��_sD{P�7�;#���j-B3E���A`Q�)�q����ş����`�c^�	&N�Ѿ��$�ӌ�XF5��x!���1'���īP����2��B�Bu21���ܫf�����fih�S�?�Ӡ���b\E�����#t\E�yL��\�%��D&菣7y;o;Z忺õJ�;k�sTYv29/�F��"�v��w���j���~MY}'s-0,�"��6Ԝ�+m:�@Ҏ��ۀwi+���d3��&���YV\���6�C�"��� $V�l{�֎_d��� J�d����Ƞܿ���b���HpEX��� H_d�4.�֤{�hEڰ�%��x/�N��KӇ@q�G�X:���լU�3�{��`�VM��J�^%�b#�[2�Qx1�	C�$�.�o�-+��p��_���o����٫���.����>��U��5mK��4;�e_��ҭ�[_��8fw� ����0�~Q@�<���+�=C�5��nמ%ٸW��l9*$��&@ŷ _� xOs�0]m\��q}^�;�7��Q� 5����ٛ���"w_�@f�b\I��i᥿.3�hM�M����s��я��]hB֯��`ǻ�
�F�ӯ�_:�kC�\�3v�S�Euv7I.�l�{<O?�j[��9����ډ`k���'Zz�l)n`V������/K��a�V�����4�x'���ٙ����/O�/�����r_���߾���n��i(2s�WN�0�٭λ7�ß��s`�ND�4֢�~�ܾ�>L��5��~/k�@�ʌ�#�.T�Z�
����Y���ͰI��]�=�booy���r�y=/>�v����������U\�`Z��B�;�������̀�o�_�����]���VL�=u����6p����@�W�)yE�l�'�����-��$�i�F������ pKO��j�bXi���5=�_^�ƮJ�V�m���(���#��S�~E@r^M@�r�҇��T�67X�T�NA�.�)6�'����4S���O��q��.�)�����[{�ˋ��X��J�R���/��m�&�;�S4?&�F�Wo��x�tdщ��OBp���jC��b��g�sS&�4M�)�Օ�=�]�]����A��}d��q�ʚ���1=�������p��A����?�Y	������B�0U������ߐ� $�����_��v֊�)3Wq�x`�"�G�!v�WC쩦�����+l!�e���vU�!n��FG�F<NWG�nI�d[
#G�Ζ���HI!�d�Gg&G��ײ��ZkѼ����7��?��m&�̖|]�]�<�~t����q|��A�*+8*�q�t�r��~�}#6���}z�؎�9?v�#����,V��U��������ҲBl���mK2s�dޮ����( ��w�����t�I� �KԌ4X���!�>gs��+_yud޵��{`�����ו�P�#�9Q�9kOZqeX��Ot���Ѽ�C�4�y��������kq����Tp�������aqw��~�.�i����o�Z6��!���:�)��5G�,�Rvk���)�dy�uO=ڍp�\Ou�"刔�f���&m�SSW�J��8[F��MpfOb���aǧ%X��JԤ�uS��7k���K�m<lS]���6k�ϐ�f�O�O���P�g��}��mq]��<��Xk����3��.[�ũ��t+2H�,
��KԄ��ι�.\�f��N
�bqWm�S�PT�cQ�Z%M��~����^� �ߊ@<G�D�ж�7�q��vz�9vX9�윻�y�}�jWI�����c����s�����Ǡs���������F{���D�C5I�G��":J߈��Q3״Fm�x�gLܒ��Np�Os�N@�z��i	���\(t�p�2_|�g���͹�4���j�4C���hꨓM�m���<:[��J���7�{|�Y�N�߿���:XI�G���<o���׭�g
��6�˼�n����Z��D�k���qf���\����E0d�]&oF���d��3:2�C,\�k�%^y�s'�O����~Ξ8gI��%�N.2�Q�I�-�_�e��p��r�\x3�����w�����f����P�}�!�95$ �Z����'��|�bU�9{�þe8ތ�z�naɏ�����dXZsh��E�����C\P%�ѫ�f4�+��������=C|������}M.�7c��m]����+��{�J36E��-����h��aѧ����A�w��s{;�]x��Nu���G��o���0�A���\$ =��7�o� �8�-���C�����_����l���ݫ��g������-uDp�Ĩ8�'�y�S^׵z��T�H����E��O�TPZX;���kZ���iC\��T�g�aC�
���:3vYs3����Y��g{n����q���Xg�Y�T�"Wy�RA�<h���YK�CzOJ������:!��2�yܐ�^�� �5��E�����H�3��SW.Q���S@��X�:��P��R@iUB-�vAԡ;P̝�9x��ǒ��m��t"R�S��x�V�hk�?��8w7�蜬��'S���H�L��а�匤��Rd��B_?�t���85�Od��b�h]g-!ݕ��eS�$+ۺIp�**ĺA�˚��)��UN��:O�h��n80����Fa���R�F��l_���R{yjޏ���Y�:�+��?u:�N}���u�g�u����"]/���7��^%��=<���L/��[2��e�}��x�j����?����%�m�2�p��fq<\���"��՜$I&�b�-Ly����Mȥ�]�P���dn�,��O9�^�h�9����|@5y�7$��#���^m��ru� ��,3!�1������bG��Nڇu'�؀x���*���Ñqߚ��Ÿ�f䡰C���� ����<��=��5TXe�M�w�1Z�"2�V�bր��i|��6�yD���zFV\7�Gf�l�i��\�;��I���DOڂ�f���F���sEnxX\�ת��+�C~3UOՏ���KA��W�������t22�q'����f��sS�U���ǖ���� �ܯS*���-�
g�j�qĥY�ʟ�g.��	�^�H�����j�����*KrS�y~N�%b�A�M4�S�9�G�㋻�AC���-:�9{�݁���Yn�pn�<�8^�)�i�2��-�c��84�}�nI�!�M��A�f3ɭJX��H(QP.��1؟-�&�_z~"/�>Ƅ�m�Eq������[N~/�:�m�H�t�%��(1nV���ܻ�ӑ�o]<�� |�����ں5��k�YA�4j�v��#���iui�__����SE�L� CG�r���j���ʜ���$�JY�8U{#��*o��#�<?*�噅���Q�!ӏΌz�fͤ�R�'�������P�o�;E������̀��o����D_f�E�}-
<���?��t	����<�Z�~���O�l�%/ ��%c5e���� ��Gel{�]-�	$��X�����S�Ρ~儉�hN��L�B	#��Bk���|���������=�,g@J�頰%p�i����ݟ��g�Ͼ<_�~y\����ls��������?��\�@��SQ�o���l��Or'��D)�����'�$.)��!a:�J�ߙ��+�Z������(���M(�� w�CIq�k���%nV���Ú�mo�i&WA恞���N�^���������&�i��ig���v�|�^����&�����
bF�:�Ą���{��Q9h�����N���.n�,�-F���t	�z?��T ��.qm��T�<s�Ѯ)�l���F�St#��T9�v6���s�b|3Ƶ�
��z�N����֯m��#� �G��ʌv%Rh ��}���0jȀ��[��kpT�����ʃg@�e����k!��8�E�^w�~m���s�T��9��ƴ�Y���%8Ӧ<�K(f)�a�qlz��ӆ/�5��e]�u��o�g��XD>��������nY����`���l_�m���\�t�uu�4u�s/��?�����M�t����x:�(�/��ҥ�,� !]�!�.�-,��!-�t�tww+�K�tw������'�y�<��̙3����.�b��}���LU���ӡ�ά�������4�6]�l@,�͍����ڹuCK�r���g�b�O�"츙)-�뾘i�9�����������`���(;_\ǋ�ZX�dHp�;i����+;��V���[�(̝�V�Vߕ<�e�\O&��ҷ9����4���F�B^Y�ݦ:f��������RQ�fc;d�_fo�9�1��V�*�E�ܔ�~ҧz#����x�H�4w���F��{�l�Z�D��7��f��^��_v��U�eh3g��}u�A�L@��H���=W������ki��iiӔ�b�e��&��}C,�,'"D-�'�eY/�`�+S���(���xp��Ź����%k.�� ˃Y�����Ňy6+�2��CV5���l����i�x.,��`bTM�.�ޖSޒ1z�3j|�j���:�[�Ke����'�����"�o�X��y;![�x�6Y�r��T���NX��u�ګ�w�:[�痢�?�X�c,4�b���RX�D���3�R��CQO��1��+�-N� {����U�b�/�32��Q�243��	�6ɫ r�*ަ�#�]}K�S�B����)%���X(��ۄ�mm��h�����Z%��Ũ�\ca�ݱ�l3 0�FoQ��UEh&QwQ�d��P>����J_֨h����U۔�KX.a�GO�ϰg�]�����YW,/��(�R�v�4 �[~���0|�ϽZ|Ca�2�H~��f��LP<;'%/p44���\��fd�U}��w�h;��|�"=3}�i�u���b����q���~��a������d��w� *w������!1�[��&,/��{fx`A8��ͷ�-�.����i��P�P���綾a�GӐ��C'GoD�Q�?!o�V�2E���������������Z�H�z<�n���	��u�[��g����{t
D�q���|���je����h��E)�z�>��"ڙ���;+�p��128A�������"�ux����V0J���E�{#7N�*S�T��Ba��dGh��*���9j�Z��K�r12��e�BEǾbb*��1Q��-��O��Q�� ם{ղ�����bU� v�_E:b�<��̃##c��#l��D����]�4v�^���zhe��Y�b�]��r4~"�ǫM��)eY ���઼�5��Bc{��F��#��C*@��D*U��Cb��}�
	��.atr�fdֱi�
�qK	�T�q��p`���@�W�V�8�W�`�^Y�F%�Q�E�Ю�u�Y��O$^���*���aH�°׽΁9�_�o���W��!"���O:�����0/�X/ٜK�\�]�G�3.c;'%�7��mN��֥�
���V����;����K�1r�9��j�(��[�ړ*�W~��v��Zv�|��͒�b�B�c��e�w]�<�l�r�j��i���vu�iaKb`�n[��Z�Օ}q�bǢ�:�R rk�30	N��gP��ᐹҗR�x#p�XH9��NW��/,��h�=�j��'���ե�h��Z��Μ��Í����"b��&��b�zQ�'�_��6�Kc�����g�#�j�. � ���$A�g�x|#���7�o˭ք3^�˳a���6��e��dT�n��M"N�_�]�g*�a��He�}l	��6�v[y(�֔f�2T�~��J ���w���먪Gb����z� u,�o
e1P|�?�8-:J��Y��2�H��&�0z���ac4�h.Y�v�t_r�ˌX�ߨնP6���7p��-�-�`��NiN���|g���㐠*D<�]O�T�9N�M�F<ɵ�H�[:XR �'������~�c�7�#yH��,����`%Cj�PYb~ޤ����֦�����Wֲ���$g������\��/0A�Q�{�L*��=r�����+��Ӥ���q�g�����G���å�Z+!�D��w���#��t��G4�?�����g�5�g��zc��k͸چ��w �H5�'SIL�f��j��ّ��jܤ���}GB��vh��hʌO�P��
�.pQg�&U�'`�����çc���d_\1�y��� ��u���f��,��/�*'�&�<�t�����{�ä�,O��z��-�m����0Bf	~��|^�9���s�|�C��N�s\���αLu`�wn�C
O�/ne��Iu%��m ��Ԏ֟(��d�Kp����M��ˤ�-��B;i�^�6)+��n��`��Ό-����"�ȴe\�s��Ƃ��ϧ�����X���ׯ�����G�3�6`�rc�·�/�^�uÑ���Nc;a����c�����ag;�w��w[��Dy�@�"N)�o3аP$��:ptg�dw� �����2�h��t�QS�D�8bF�����E���>�Z�0�|�q�ّ����0
q�T��u���c�9M�C{�[yB�^x���-g.�	+�O��>4=�3V�ʥ|I���JJ��YwHZ��E�5)� x�T�>�١�ZZD|:���P�X�u�o���cB�7�B�֨�z5�VK�E����+_��"j��	
%��\E�"k�4*�������
��:ӭ��oAn��a~g���T]��(E�/T����<#.v:���͂�7V��R���gZ����^��:pb��Ы��7\D��-N�D�I�D-���ȻO��3k����aD_�1ϱc��Յ���R9�͆oM,	1a���F"�m�YDӌ��`φ�R�C����B݂�mU��C��E���~�D?K;a~�5[0���h;f�<ۆu�����f���Rw��H�)�)v;�|l-�&�x)�?�ͺ>����{�_�7��]>��L�RR-ᵹ7��=�z���gS'Ըtv�Vpz��
��V�gǥ�FWz������y'7�z����Vv>Y��m533!��U+��k4�	i�D"Qܧ�.>)�r��3]�C�QX^��p�������o�!��[M
���i����9:�DQ~,@�^����/�Sz����z�"z�%���(�c��^��ϰ㳱��}e���� �N~����&0�Y��;�~�n޼�R(U�"I����
�|JR��3�P7}������Tq�k%����M����	�u��f��9``�����5����_g�zź/��_��e�M��ҵ�WJ��컆���*0��V�L  �J��)��Ns\
K{X��`A��<���(��|>R�&RԔ¯�72i�"C3t�jG��j2`^}�5	��"�_"��e:[���>���^M(���fu�4�'���/�{8V�aU��\-�Zj�p���j����h�R��������kY�j�pkY��I���	�di&����S�1�v����1�vW1���V��-x,����u��ޛ�K�1�`�����.��}���0%�T��`F�����QU�&�s�W��Y��V�)��Q�x�%uG�bS�������%V�BП���Z���	0�]9H��Q֨���T�}���D9�.�8ߕ��O��NX^x�k�6�b�4�8�5��¸]f�����g��SJ:��*�.��z]��+�vtX�&Lm��<ʽ��5vU�a�� ^j���y�ٮ�#�\ͥ�6dX"�Er R��ZdP�WY���G�I�����)�]�$+g׃�����˓�ˎ��h��������	i<}�ǻ��6��Y=SK`����G���A�EX(h��<a��k2gE Fa�ט��;�̀�ё���"�*�� IڿK����"��IY,F
�!8�7рv'�ą3��p�[:�#9�4jӭ�-RQ����<b��,|�
cceM�d�o@5B��߅u�5��ېZ�VZ+E��C��Yv�x=�t<���>m��>]�t<�E?��
��}�*����j��o�vv�~�����9�L��n_H]n![����i�Y,�t^�ᡱaK�ذ�ذ��7l��TCS���F��태C-��P^���;��L�1j�)��AT��DNP���l*�)B�ID0�8$��?��bì�e�P+��"^���QB�;�����ʛI^!VԽd�eGX0�[)���_��9�fuJ�䬩]���#Y�(ɀ�$�_I�]����qqq���^*Cf5�ߠb�E%	L&F��j��44��������]��"D�

굨��{�����G��23��R�ūCRuݮ�n��Q$��
��)����G<��?ʹr����g���1��؃p�Ѹ��h�{ j�5�Y�?�XdK��a�����SvȻ�=�I[$;�w����\��X�tPh](�z�C����)�.��7��Đal��2����h�?nJÊ��X�"��)	^dP&ډ�V �"����W��DB�S��b��X�s��!���.�R'��IW���Ȼ0z}�$��2l]�Jw�r�Jb���z�J�◨Q'�s����-);ۿ6Ҽ>ٻ7�5�������̽Pcb~\AuvJ<9I����.^�k�8�+�Ǹz��%�MM�t��Ϛ/��<��_�.���-U�4�S.Q�]d�5�x3��D�憠�<���JG��ax?�K<�.,{"��u�UxR�O�=���iG���/�/�x_z\L��֕��/�����&�e��dl��Jh�͚!�v�Pm�4�޵%����/��slN�����D�h:v��{fhXmR'�^J`7���WV��^���f�N����a��C[2��A�8ڙ���Ւ��(,3��ZB���c�,F �׿+�U�\P���Ƭ.�K~��Z"yb��������DY$>֍��U�DQ�B��N���]N��~������}�sl�٫.�w�&!��k>	��Кv1�}/ѹ>�jB�Ӈ�=���b���u�[4u֗S,��h�J C���YR:�05��U�pR��jf�Ӧ�n.�[�ZT�~�Q��3B��ק�N?�b<��E�蒂<���(Y �`�&�H�B5Kf���k�zz�tb��x���3F&�^y�|��aa���:]i����f/so�K	��*7�/Ͻ����(,m��ڳvYx����碬&������ߤ)�B�DJh�.�b���7��%V��������!P�O*�HsFt�v�Ԑ�x�2ӣv\��(.8�<a �b'��A��2-� �? �ʃc���a?���+���ߟg}]��X�"�#g/�B�'���O�K��%��5�щ��}�gy�C<<�w
��,7M>�]-��=�>��db�ZV�&�6�.�1�Wf�dc�ޣ�&o��ܕ\�e~1q!�R#�d��^Fށ���YL�����:o����:�lIp����z�\��6����}����p8�m*�&2�`�`ԍ�'W�e��a_�~�4�Q� ;J����׹b�������ΛMZfQᠬM��M~�0�v(�r�����)��(��K5[Q������ei4ͬ"d�/�+«pmɖ��T��˟�Q�j�@�hȱR�h1 �X�ny����=��@����e7����M�{���V�5RB^��Vqx��7i1��v �ʞ��]�g�\��R�$�������hiFW �N����G)j��/�,2�>�!��<�c��i�ֶ�EӋ����!���R���ګ��Ѷ�T��e��o|��ޱ���������΂m��QI��<�兝]A����ӈu�~�"�^z�˯^�P�kL�6��u�ۛ)�.9?<�Z����9�s�����^��	�US��0�
:�!�7H�Y�2B��������L*�|����Ǖܫ��8El�`|���ж���,�?hP����{���-Gk?�,���-�Rxbe`Eȓ��'%媏������8X;?���"�nSF\��y��!X��$3$��ݕ*8˯������۱{��������\���L�����H�㖾�ݵv�m���ʹ� |sKx��2���T����zK���0�QD:��XI��*A>}uu��O Dc 䒼j*|�jxnY޹/����K<S�A��%yVA14���Ab��%F5�N�|�teЏL����@Δ���z֦����~� ="dIY�B�J�!F,6ޯg��B���Z̈�ok�A��b�O+	Q5{��c��X��v�������5#�%�
<����B�k�,
X�OV��7�+Z`�C2^8��Z1��u�a��ַ� ��ҹ�a��~Ю�rq�y)ƖGC���@s�E���]#uY�N�\	9�P��wF��ބ!|�84�{ۈ^Xc�Q/��)��L$�M�)��V=��%��G��1J;�M��a$��j�{7Dt��Mv��ƽ%���D#���iυ/���e��r�����_3];�2�ڒeR�]J&ko����8���v,?/k��O��͝��^��z8��h�U" 0䢅�HG�x���?/��.{-=��Lxv�׿ �ժ�B�/[��A����rr�k��Fxy�eEt�b�.��u��ތSP���8:@+pg�k8ekx�5ko�[��X�)0h-�;/��U������e�32	�W���~�o	u<y@���ƚ�K w(b*¢�$/�ڜ}VI)K�"�a���d�w&D< �Ø�ʔ�=��(S��Ǎ�^0:�L��q(>�2P�J�,�ȩ-0�J��5
��ܦ�;���Ml6�`�1���*�
4Պ�����?��(H��~��ٱr����v��;�qN��Dz�eQtT�'͵�~ЅX���(㇬�h� 0�p�$kK=�~H����v��_�t/��ba��6R��D�5������H1w���*/+|��I-i0ߋ~`��)� �H_��^稉��/�O��N�v�O��,]��hLP�M4e��*�s��r[��q��0��
��P�
��QS0��տ	�;~f�ÙE=�U)�'�����ٿ?��"���Wz��S�t:b�L�$ ů� Gj��1��}��15<�E�6�V��Br��،��#��|��ե��������F՟������d��S*�����M��;6�=�'q?_�o+ �i�s*ne~N���r��t���[� y٠�f�7��_��@�G�16>Fm]�oz�9�._�K��Ro]4�j
���?��?�����T�;�2oq�J�����).(��f��-��x�hjr�-��Z�RF�C����e m��M�D;��K�4O]���z�h��6�t�nǟ��0��@���TPT�S1��2O���g<�Y'Z��7*��')H��k�%|֝�����0���������<�Ċ��g#��%��xcN.=�Υ�y�j��Հ����㧞a��Ow�����;��G,,x!���?�����dˋc�vC�Lp��~��HŦޙy��u؍+&Cn����8N�T��	��$MW�Z!�F_'ay����p��/���Nn~~h��,D-5cP�P��>�!�21X
P��j�)�)�rW�8�\B0�ɏ��ʍ��Z_[/ؚ?����[���.��_����tEu �����Hojz.-�.:�7e�)|���{>���4$�{V��p�K��v�3�{�K���7�u�l}�B���}�?�������EQh_��uHc�5���b�ѯP��TG���2�YB� �ɠ�H���:vb�Q��U�X�5��i�/�qX�bEՠv�R�ʂd�Y�~�ĤP%�(�+�Ǆ��Q�Jb������߽����WISCCCIIIM�ӡ�.1�ƍ�.���,����pnӬ�fp��^��Pu�I�\���q����"�'��K!]�sMnk��}�s<}L�E.����u��%ō���M��m�Չ��w|�ilz׀��-|Mo�H~��z���%�p�u��i��x��c���b�l���PW��Q��3��*;�,���
�r�U|'l�@�FDX@���z�D�02�H��2�	�L!��q#:<�F#7�-i�Ł,;W���YBz������꯮T��<kb��"�*zt	��=6�A|Od`���y@p�����	/G����������k�Vޓ#2o*���ձ(������+�ڶk���W�4F���;Vk���.����6'K��ǟ���e��/���u7�CvmT�r��Vxx�7[��S9-;r83�zFM{��eZ��ē0>�і��<b�x����
��k(0X��a �6~���Bv�.��`�r���p?��НQJ�_��h'.㍃�Ph�á����Y�6��/��ʦ�|�(���M-��젉}��	��3-5茋!S��d%zI�����?�wWC��V�lW��p�o�ܷ!�^L�`�J2d���3�1$���=�}0�fՒ1ߢ��ѓY�!RJ��s�2��4.f�������DhzD�9������h���#�U��II�Y�Ǌ$���eY�Gf�0"���,o�߫w�~I��_�+�s�#���ϊ��
���x�6%��Ei���
?l�#�?\"nQ� [��+��8��=sĬ���^�i���$-&1w�Hے���6�4�~���
A�7~!��A�T@�~ %�9:�o�̺yh��SxV�x'�o�Rả	O�Dm�J�}�Ns��q��V��R��V��m�\�录���;��&U�T<�}
H��V��u��S�<�jaϔ������y���}gx~��&�s�ZC��BV�GT"��J���֛Q�3E/���-�{,��g��%*�>���W������ڃ��E��9���s?`���-c_G����e���C���������·՞A�1I�[��hvF�1��'Ӡ��33�\x�M͉����$��g����� �}�Ų�P�ra|�^�Y y	ף�&gJ5xv�{��Q����?�O�x��A��7?T���|� ����e��0�SQU�Xj}Y�P֠8�]6��?�����
��X�؛�T�J��*5uRg\f�Ւ�0�	�1�13�?�"�\�hYn��tt�d�THh10N.2�����*k�B?��\9�逓��w��N�u�+��;�Ǐ'�OW�������>���+^���˱�ow��y?z{xJ��7��ş�5�o ��R4�9�z�k�0��H�sY�<��W�_� �V��s��t��9� a�������Nw���ūb��Y2��݀6ay���������_f���c����xR���k�V>�u�.=H��=�|�x����x|�y>��}�Xy��wj�^<,�gʶdB�pw�O]��BJ�Uι���B���N�W�V��=����v��1���:�}@�R�%yu^К9��ٵyZ�]�N�j������i�7S��n����V��^��_��`�}��ѿ�*�/�'9��j�*y�h�:(zh��Y=99�*rO%EE��np8<�!ȝ������"Y!��M�V��/�C���	/QrRUKN���ۘ���"�쾁�6z:�Y�{+M(��,ᬦ=B�X�{Y���$.��E�n0��8�ڬSQ������� 6���LB l���%���h���9�,�q)�!c�Xi�C��?κ30�`~���,�JGѬ�rުE���Vc��yNt߽lG&�,">a3�Ub�#�cZ��b2��<��h�m��49C�/tɮ-lL.tp>�{���+�mx�L������Ș���]��5�J�ofJ�O9W��QE��6Oӓ����#<���m�c'��mi�܁�W��+�o=�/�])�;~�~�q��b�y�i; ����f��Bz�����u��u��MKˌ�wz˚}x��Y������/��"�&�y#ӓZTgXZKO�|S4T���t�X[�A�ˆ/�5@����� t��W�l`��维+���h�����?�B��,�V���^�dĀ�* �?�����sk��dPK�1�(�Fds�"��(g�"v�R�UȠA�i�����c`�匬͜�8��p�JsN�$%��'��ǛD~�hI����V����ޥ(�&E�W��c��?0#K3���q�Z�U��~�#e����&�D�>�􉟢E��H�M�녛�֍�E�iq��X���Y��1��)�s�ib�&_���"Q��a�a� ��8�����,y�Z�\����+QS���y���_�|y!�[jNn	m��������8��9�f��M�ݭ�k�9��k��M�樤��
���� E��J-��a��u�H�L����S��-qG�����F\�$�@\k�mJ���B#3�%"�۞�$���NO��a�I-<�\�>YEb�s���� *�01���w�<��j��W���Bp۩�Ȫ���~9^�֒�{}^��1,�E��@:Ʉ�*��o�5ܿ��'g�������h��0s=��*lZ x�11WA�q�ez�����Rή�%�N/�ac�a�b��L����>de(��s9�Vz�+	�D�����HhD�z��W�Ş؎�jlSЫ��Z7q�ѽ�jǍ��]>���Yg��ia����g�TYX*'�M�}H�\����{��Rn�R,���a�&5�_Ua>�>�+Tޟ��*kiN��!dm,g|n!�[3�ǝJ6&��	7�A'@��pY�k��'!��Y�0��-.z�߀�K�
^�~j}5ch�J� ��n�o�7����K%�I���k{��[y�~�Y�x��9���-?�R�Żr���9_jqir�NL���� �\cHF��q�x��&o����Ӆ��[�+�L�8�ۯ5�O=0+\�z���Z^Ӆ��c�Q�#V���4ۖ�Ioc���ٱHh��cC=�P����b�e�,Y/�[�{X�t���v����9���p,����p��|)�xF����ɻ����o��(.��! >
��,�\y���3tof�b�̯���fa�/N�u�I���Ë�8�4�;���Mb#�w'B�V�#5�R!u
�N����J=8���F��(���gs���Z�52�0
�gà����<�|Ub����W�L}п9�$��2�%I���2|�O�o�x	��~F�LnRn!����'��ާ�^=��3��v��^�.��aA{���"Ri	�B�*��_>}k�p-��\]����9y�A@ы��lPp�$7a������cȚȐ`+�,DX����� �7��,V[�d���9�[�*�w#$�H�b�3"��.GZw�?��~�Vzv��M��& �7����3M�hY�����2����O7�+~$1�� ȋjT�������*S�Z*�=P��N�-xd��+��{�=l��D��z��R�_v�F�y���E�`4�����k?욪��@�t����X�w�����㠭A@ȫa�Ǖ_ث�q�q�G��B��g>Pr�*i����~沿����yZbd��������� �3PU(�϶��=rk6ݸ�k��0���L<L�ּ
c0�v���@���w}^� ���i^�	��he\vm���L�QAq�L�{y��w����w���c� ����!��|�J	�Mq�����pz6�h�mJ4�a���Z0�a��Ǖ�}iFR��-�|S�=�_� X5V�i$'a�
e���@�����Y���s˥	�
�xϭ��^���e����]�v�kz+iS
ù�kd��XL ��,q��!$3�׀t� :�Y�r��>;A
*�� ��n>�WS; ���L�q��D��tگ�΄�P�±��%���$�R6Q5k��,����%�'��j��P!��R�*4��9R�br����<�+>գ\��DP���\rtr&�z���+�5��qYP���`����������y�gD�١�O�Uh0Z{t1�?��-�z4�9ټU�y��m5\�M��ٮ��B�.w��$Jr�稯S?��P{Iq -(=��M�Zt�C}cI��D�QL�.��e����-�T_G4%K���Lt� z��>��3��8<�����" �r�ٷS�r2p�+}�b10~f�a�����?"o�Jߑ���'R0aT5��'R�W\f���i�	dU�?�;�����0���w� "T�WKt�tk`�v�p�W0�����=��L��\�❜l�_�uco�h<��'J���Zz��+���V�m�!�qf5(^8w'�Ϩ;�A+\���Vlԗ̬�e��Zp�v+|�{�c7y���*��mG�S��h�I��t�ۚ�|���=:����:.�Kl�tZ�[+9g����e����0�t�ʐ������]�P�8��~���)��?�%�!U�'O�J�q�E�C9��z2�?j|�� ���R
c���8`:���̦�d9�3j�66�K��6�����nU"�������C�X�,�/+��@	�˚��P�*��P�x������2�V|����}�+:no����)�ܜ,o�ds]�[lJ�u���y|�q�f�������|�^��@-LN%bw��}�j�CT��AJr���V����2p�R��E�n%oxU����[h��z/������;k,r��y;ޜ������)�?Ja�����4F���Ҽ�D�?�̈́�b(���o�!D�qZ��IW �rh�~7"�LP�	4�K	�PQ��#�9e�{_m@s٨�w��|6oF�ڝ6fy�2���gc�^�MqF����nw�zqh��E�R���+�G}r`~PQ�\�7vk~D���M"�@�E$F�ga����/̅����@���������,2�P���WI(�٪�~�/�fq��a�z���ȅ"A~8�ܝ>�H��#�
b	���43bq�+v�oblU^���a��#e�:�[���*��1��Li7Lh7LjS9ڰ�N{������o�U�\-7�5�֬��{E$�]t��R�.�w,����G"�cx}_!J��M7�Oq,t�u���"��q�~���!��auj��]o/���|��΍(��U̽[=�|���_�ܱ1OA�ҪH%���~��H=9WFig"��*���h^8�K��bR̝6?��U�Y*ca�yT�aE����>ت'S�t|&A����睚�+�AQB�,q�02%?3���LP�A�p��߰���A����I��D�=��򃌦����u�qB>ϮQ�_9��/�����)��viTf�kB2a����Ml%c��+P|����An�T�YXV�g�+�Hu΃�A\��d���AZ\�A\�����Y�#��w��f0 �g�r�̖ut���OEx����N�=�"�쳰���%��$�ehK{C��k�0f܆^O���2Q3[������##�̃D&*D�P��������q�EL��h� v���8�]+�G�E�bb;� �v_�8��,E�/6���aF���7/t��}�V_�k��O*	a�����֭��-�ypԊ��ק�#�\d�1��Z�!qWi"'Z�p��	8�3\�8�\P��)I
L&�Q8�k�6��X:k,,/%�����#n���>#uÁ0�V�sH9'��`h�RD�SvT/�R�T���B �r��Nc<�%������Ew�a�ȢAz�3�Cw.1<Zl�*Jb�:w�Z�A=��-�
�,)��������y7�T+�:S�6Xh�ٙ��[��8��N7��������~�k�u�I��z�]xo�3�>z�L-���C����|��V{S-=%+F�ں�e]F{���C:�3���o4_� ��KEߚȿ�R-� ��m���J�u��B���L=.Z����ҟ�Z��'G02u)��t���[�#�{ﭫ��̈́[,,.&�.bР:���B��߬��.�3U�dȞ2�Z�(D&3�
\�Ԃ!/�odS<��I�nh�I����~D�<���V��#�������ϱ�-\�Q��-m�A�-�xBlm��2��j쾻�r��n�i��ԓ�۰�-K(ǲ�f^�F���t��y�F�a/�����\n���a�a����q�������nQ��~��P�䲭`��A�Ya�r�q�� ��� ��7���U��}l�Ƃ�
8��h��;̔�YH��õ~I�'���{M��Xi=].�iV�;���*�'�g��Z�E+!�V�P��.� ooo���nzF�#//#�Ѕ&�ۯ��))��{�3�۬`+���Ml��~sη�BԆ$���NJ�ᶹ/�w7FS�&�m2������xX��	��B��/Ңߊ��F{.򔃀j�E�Qw�Df>��Ak̐����B~셑gb�cfMc�q��;�ѐ�@�m�b�8��?$q[��i�~<7�9�k^����s�#�2���ۑB�����W��w��I�D>@��h0�Q%�*& 9���@g_�-��ޗ���wOa䵔�����ŗ�9]�vm��ߕ<�K��V�o?�Zx�=��O��M�q��������Bn�O{f=+�;���-�����x��hHD��^pl�"��ن崛��o��6i����.mq�v�MW���������ә�ˍӧ�u���>vLW���gS��<�\S��ٖ���חw��e�� �彄~��謕����������=r8����FR �Yd�����W�}Vue��2��0]���-�#�?��~)�6yj�@�Q�A�5񘒡�!�:WP���K[zy���NX�@m'�bf�\� V�3o"]lZ�h�ݛ�տ�	_�B6�@m=�����R�~f���hip�%��N�,�G��_g?/15�dx�eo�^)����l��������E��!�(�o��� �C%+"D%�ankEA�uGE��MD�q��ڭ^�J;[����&�K��WrLd�9�� {�_���N4�Mؑр���ɭ���<3aEy�)w$%���n�@cVc.��}�a��K��%���Q�fA�|�]�>���v����<��vl�2F t�U�-�v @�r�Vp_N��n/qf�%�}|��S�)�[�q)�;�����Rh6J?���N.�����dSB��H��%졠8+r�(�ө���p�m$?�l?��m96���/��c�t�d��R�3�� zG����ø:�
��fKEA�^@c��7�W��B����~�0�I@i*X��Y��\�CA�����*�/!�9]t>���s�3/Bw�&�~I�� �����=�oY��s���ŖP��5�$Ǔ9���Pg��1bi�/� �~"�ʒ�G��s�6 Z�W��J��y��z+�V
��-��*"񁗴�/�:���|�RH	�Rl���P\I���}K���_6.������0�'�BP^W�TSc)x��DD���B��r�8��T����a����~���� q�x��L�\�����B��>���,7�<�Fqq�p!��0L nX=S���F >��~��5��*o��|K�C��C{Y��1��6�|@'8�-Ee� S�0����$�&:T�Lͳ�@����b��Z�T�����N���,V@ t�}|Ĳ4G��
h����ݳ-�i��:�q����@�N�M�P�ϣ����@�jD�鐷�q��m�0���jk'y����oe��}����Qx���"𗙉R���e.�w�(n�Bܞ;y{*z]��b�qW�w~H�l�;}i�������Q��H��k�0�ׯ��.���]�_DDT� �OLZZ""��a��� �Hf4�I}0����l?� i$\ْҺT�x=]��beX��}&�"��������1���t��$�x�7���Zº�>��A~�oJo���Ѵx`���8&l�5y�x�3 �_�9rpx�k�kKD|�v��SQ����թoP���3�~ �?0��/A�:"�o`�V`�"4��T�?��b��)!ȧ)%�ߔ !�`�J�)�OU�J�d�W�!��W|_��Ë���w���S"��ya��Uu����gR�1�$�l�f&��Ցn�^S�'�ˇ�ȱX�
�V����
ۥ�/��m�%Ǉ�=�6��{0i<��K�䧭���eɄx�v��C^�睇�e��<^���!�v�۱z!㇞��6����NA��>M�cL�T�7'
�.�ƶJ�����*��xk��ŭ�ˬ�2�J��h"��F��E���?�m����A�B��3��wGlaH��$��
���	⮻R�+8oV|?�;�-�I`wQ�?��8��?�)��~�D5���+����Go-�����*|bޅ�����\T�c�z�A�$�Β��F�&�+��Ϩ�2�K� ��K����5�󔄦����oz��O���^/�d��Nf+}M-�o�����D��D��	�A���Ms�M�����k���-HP��:%�0�g��0�0�(�-�|�O.篗z�t��U/Wt�k�4<y���Pu�AQ�o�'WI�XD@$�ki�V:�[�[��n�N��Z��.���3g����3���<����W�\c�!��a��-�'9+���c��g����%*;���D�Gk�?��aYB	�`T�,��qɿ5��l�eM�Q�VY�pC�{�B>�������V T�1���ۡ�o]�܊�/ܦ9��[�����_�q,��9F=���O�M͸������%��5���q���9��G�R��9�Ks̑�K�)����T�͒zm�m��|���4����BoKɭ���T0o�_yWO��ʩ�M�Y��c̎�֔���l&Y�]:�"����oϜ:(�?��fx��@MEU��fa���]$D��ll�j�g6�O�r�1���]Hy���}�I-e()ׯ [�-x�ek����G�.N�ٳK�iٲm��%/�Ԝ�ʼ
�[�"�,���V7�W��kRO�.l�2�����۹�ϥ!�N������-[�y01p�L�"�Вc@q�@�.�t6�z^)"x�ܼN����|l�G���@��o�����H�rY���Q��u�����b�ߥ�����U��#��$m�f�;q��s�]�Ԅ11V]1 	�k�H���G�h�� =�
���	�\Xr.ڑ�[�2��Jo��ǒ�q�H��6��))Q���Ǯ�zy��,�U�}���d)�ˤ���V]'!]$m1��O��tsn����s5�R�����:��P��q"}�\���jw�"��,z<c�ޫ^��9�[n���<Q@Z��b��K�GC]V3gEcsVk}����wT��5k���gu�0��-A���b���@�-ա�RV�������ks@$�ps� �u��Ǟ5�(�f�F\�MT��L���{.,Q��t�5������+���\?e�2i�ؔvEXY�T��ת���xn��вR(� @i�v`iR��)#������iiiKKK������8��KJ�z���C����t���������Mh�;:�~ f41�쯖���x�;H�J�u{@����!��s���D��4~'���ӥ���C:f�)�Al�NnQ��Nr��ӽ�{.�:�)=��q*8�͜VD�6ٚ�D�C4��C3�"� p�g�5òM�/���S���E��I?�,��-�yik�M3�c}�OMLy%lC_�� H���"1Z�vU�I�8��Wg�&����F�A @a0tD_�����b�W*��D��}�@�A�B��&���ĥ��% �v�KW
>���Dp��P�`Tj�M�҉�?��������pl=�����Ԝ'mӖ��l?m���]�z4�M��^�v>�!�~�w����v�Vo_�}?:J��|]O��pZ��~��im��}�nu�1�Oۿ߷�����S܏���͑���n/����}�4�X��by���������]c݌�	���ǯ>��mMs��U�6��z����{;�xq�o�.�?��)�ũ���>Mv�Yo��Cc���H�5E-Ys�J��l��ٿ��̱����|�������Bz��Zemr� >s{�[�ލ�uv�d7E���%�K)��&T��Q@󝌬�{��� �{��bV��$C�&�ƤNEБ���
u	7A� �K��4t�]y"�|qL�.V����ʿ���]�-�ͯⲏ�&��b{_�BD$ן/�CD/�"��kp�,������R��}k�(E;�m�/>oU�OH���L��_�cf�e���=@�A7�}3�2�N"� ����L�p�(� �����£��
������AW��$R�Lȧ��Tі���T�l�P1Rk�cY����	T����%̜E��ԩ5�
V(�2��!��I����O;��̪�U���-�VϜ����z���j��D׶R�t�U�J�N��Z���@���L>���bGFL�p,'����EC� �u@�ʋ��_�dR	CV�n�u�|����♤�;�xۧ��R@�4�+J�~y#�cͣ��1݅z�B���aԫ+�JW���\�!ƣX�ږ��� ����8,�k�P�*�6.�g�1�����6�+��-8:�yw�{�&nP���w{Ƭ)�P�ț^QjK��2ux����}�S���<޼���a�KQ�'%j8���n��ַ�ht��S�0�uS��-�f�G�@��d}��Yq�-��~���Z���p:cB#:�m���@��������P���&ʹM��r5+�K��b��:����9��R��r��Z��_,�F����<�ba��������}�EX��Yg�H�Ɋ�ټ�,�O�6�O�uϝZs�TH_-���G*ا�`���PK��G��lenGT��������f�r��s����U9���*4�*��	"g�Ӑz���#�Qf]��o��q�y��aK<V�F���Ws���u��D�O]��"���ʓ�Gm;.�,��n��p��QS��r�ײ�jH�֘^��.\�ֳ��>��Ƅ�(0��J�~�|������ʵ{�nvc�b���qL5~�f����� ��L� ��e%������<]3�n������;��x���&��&}�x��ULa��!�fex��_h��gD��꣓m����@	�9��v[k��~!���}����B�_ѩ$?j/�������Kr�@�q�������3���/���{}�?�����ڌ�n]��}s��b@�\Pk�REn4;�}�I$*=�x$���"�_p�:έ�(4o;�������2�]����?�O�r�c�#�.)fY��u5�9s+�\�VX��Y�Ā���M9n�۾|�pjt�'/Œ5f#y����h�'@�,H`&Ij� �'�ǡ.=���R���I5�d��8���X���2Vr���Ӥ��UE'{��5���|�c}Ĵ}��G��R�Q�!٥�#�d �@��
X��g���Xw��0=�z���#���쇿� �|)}�(��	a�ڋٝ3�T�ҳl��AD��Iݼ�B��k�	�?~�=	�X �E9#����z��+�&w e�Y�vBBŊ��FcܬZ�M���Cgg��x�C�-&��/VB��f�V�8���[��'�O?��4>.$�������\����τ�Z�?^\\�49ϝ�]i�{Jo��_�z}��ڊ�"6�wC��阘��Zq�a�����{�32��*�W���W�?�|^mX�^9��Iw����T�G��5��z�;Z��83.-|����)�3�]q��5�b�J�r��C�~�u�`"�X�pJ7/�e'U�檈����)8h%I�>�*{�-X[����lꈬJ�Z�N$w���?y��tA&��tdT���@������V>���־�q�"�cR�菲��%c�5�[p䃲�o���D"GGM�G�@/�[�OW�<m��w�`� P�rd>������A���D�|�A��-DV��Y�.41)��Y�yZy�f�R1%��t�M��<Ԅ���J6�l�P��9�����gč��f6G$��7�����Z�=:s~���vce�� ~�L/
��yD�ڇ�D5B�a��B��ɚ�vҡ�ì5����R��������:q%�&�@8$%�sE)���o��
z�"��!A�D�H='"�h�R|��x-�8�V"�	� uN�Cp��#a�5���Tr�����U��*rX#�9�Dd�5��4<,�����̀�����<+q}�e�?󄮴����<�u��R��}rۦ�C/�����,��:�{�9Z�\�A��mL��a�|L��,�nJ�lQWLw(tE&ϱ3V,w8��������R��c�IH�t����������!�g
���{K�xU��&�*c��^o�1����v�@'�N�-ԫ��]O�_n�H�D+�0�U�_H�7a�=(i�~9�	M%̰sN��e�S��e���e:,)!���
d�Ff�	�� �&���8�enq[�v�|�r4��OL�f��I�)1���/��i1{�io�6�G��I��fL ��W��<�?�,�p8ǻ wm0vv4&5\Fӝ��Ba)���}kw��|���M9�J����ͥlU��JCb�����c�����עn���NTU�t�ɴ��V�;�D�4���&�[&TpҨ´�: d]	K�O�a�C^��q �[C-�Aq�H��aP`u���d��:����ER���W��S���֯��dh�0�K���@�]����?��d�,��;9s"H�β����n��2���]���e�|<;���L�������t��J3�W[!�[��ge�����zl��v�7� v6��6z��z9��%AVj����a��J[@T���+�N�E��ެkM�} ǱnO6�6�qqY&��V+S�H39�Q���ޢj�lk��u�(p��}���W	��y}3�e���/c��S�����^Ae���K�V�賅��Qz~�@ H���i�!��������膑��+I����"�t�
�[�j���X���b1��<�B@ :oo(���#�rdW��ю�|޻D0�oO� �������Q?G ��z�Y�@�DڹoyHv4�K�H�L$�T��DC�gu��Tz���r��f��>�?ΈV,�����4�$>aTN��0�(XQ j�*0�4-�M?���z�>;����Qǵ��[��p<���Z���,>;Cg�Z{�{5S��v��ƽ���c��0��?���o܇������w�:���f->V�ypR�^iz��y	𘫯�9_��Z	V	��:o�ɯ����>n�L�K�:��w�]_븹Q�͚L��Ϭ�ݣ�ݱ��}�܍���b.�8���]����U����uC�VaPn���{ʲPCan�Lg�K�{f�Oˌ��FJ�+c��%�}�d現�ʻn��3նW�
�����Y:�F��~�VU��}ቯ>d`�-�JIuD�!�D(`�����ԲW)?kg�0�@gj�
�P?�������Ë��������7���M��v�d�6�0�؟�������,%�%��3��?��`�TV6�}(i�PX�U��/Ya�ɠ�D�V�t��L4����>r̼K���&ؘ�.�ae&IZS�9����p���mΗ��`��B#&U��!�8�2D-�p�����;BB#]���L��ZS��\:�ny�+���^�8a7U�������){8����3����wl������y�6x�����4���#*&?	��1|6-��}Ђe�30��?��)�/��j2�b�ޯ�+�aOۭ��վ�"Rt=�Q��h3��Y&���5��Tk;��c���F���Ӫ@ҫ�V��#؏c9?���?�^>{��m�և��n^�ǍM�PK����u�����y���@���BT[�t6�2g�3b$n�s&�z�Ȃx���"��8kW^|ɢo�$bt+��X.��c�h���e � ��X�LE�{��<��1xj�؅7ő��U�ĺ�;/�(�GPy_�O�xW@!W�����ˠ�(� )�ga���Xw�.���z�Z��0UBϡs����dQ]m�P��p<�]Aο�����i<Un��KJF��6�J-#JݨL]Ʈ�/���EL�/���bϛ�%m8�Rh�ڗM��S��$�a���m�otU
u�#R:>�ף�V����|\+�V�ϗ[Oem+�"��[��������9
�sƑa�jYm�=��_w;5��Q��;�B��M��R.�v��b$���q��4���VD�{FFk��x�iS��\�� tC�RPm�����s&�b�w�3��&��TxV>=�[�wɩ^p�2��n��h�(U �&<F����do��ҫ�x^���h�0�H`HK@�0j�������eJQ濇���{׾gG��.	����lKm�A�G/�Z��JF��3ke�3b�ޕү��� ��-8�f\��n�@���Phn��E�k�3Z�E�E�$���~��� �B��%D��ܰSG����U��+��/�+���?[(��j0lj��I�"�e�;���>>"�����N����[��T���Ut;����v���~���~��4a-�+T'YY��w��)=�8����v���YJ%ҜW��T¨��L�}=_��|�sX��*Ӡ�_��Ac4�D��.�!g�ɪ��}(<Yπ�M2���[CX�1q!��R�/���9h�ww����_G����Tb��.�BJ��b�BvN7̠E
�g���8��c�F|0��ؕ7S�\�v���t�[՚��X��q\�z����~�w�잨���l��վ�֭c���Cz��&��p�߱�����;�YZ�$��ߩ�|{��~B gxҙ�����)E��lr8����lVR0����H�ma��s��[���d��xţ�Ĝ�}�lO�7׾W�b��Kk�wd[�X�� �ȅ����SʛB����	sh�!� ����w@bqgɴ�r@4�T"����c����;X#~�d:�?� �� o֌�cr5�R��V�4�^ph�-~Z��`\������y~�	뤃�'��lV��H4�C�l���0Q\.��{�짭Ȥϙ��c-��1�O!n�'5|��A]��ӵH1L�BA����V,]\]�P҈�# �6�����uIw����:b��"���YD�4{&k�[�͔�������KP��@���f�� @g���<&j�i���l�aKfU�|S()�����
σe�[��6��b]�84>����F̈�^�8+N9)֠�E$�ʠ5w��8���F��n_͈�T��U{٘���R�U1�8ל�p���D*�FT��"��{ʳ��тj��p�Y�a��P��(K[~6��`'\I� TJ6�w�F6���T{�p�f�L��ٷ&����6�"�)��^i�ڗ�nM_N����������1����^c��j����U�A�]gB�o�����Ykk�&�ID@'�������Z�T��=�m�q��x �}́
aE��K;����ħ�E�;�8}��+�����+�-K�'l��&�����7�p���E�y�R�[A.kw4���$����ݰ|}�;H@g�z��[XvoZJ������.�r���Ck��d�e�ԹB�VT-*gH�\�3��A(�eG5�+���H��2zꝈ`��{C����b��U���b(�/�p��?�+��Dv~��_����NW�7|S����`7�u�]�c�s�uh�ڔ������|�lI�gb.�Pr�'�,��.�}ǍSMkc����!��~�/�lr�}�y�-�pgw�:�v@��-8��;���4��#P[��<Xֳ{wTl���ex�b�����}2�o����fmd1��fR7�=��O�&�]w�Ӎ�2�Ä�mR�Ae�4Hhg Z0D��ab
XHr��~�
��<�+�h�8Y����C/i�e_���d�[;vH�����泩/|>.��cm�gz�ݲ�=�e>D��Ϸ�B�}�ݛ����_�ۣ�@�����קA����K�ƙ_�͚ɪkL�j�8�F�3��Zз�$�6��R���2(��0�'��}K�����o0��UtW��`�����7'O�S#>�٠Z�u���0���������ߣ���!�q��Y��I�[����h�\��YH�o��#7�ӱ��T!����-W��D��%�֠����
��V/���N���g�sW���{���G l�ב�q�V���]�����*R'�Q��N.A<Ć��5 ,�q���W&aUA��<��U������W�zf�ߩ��x�S,�⁚�׃1f�I.�����h�xi�?����Pu31u��Ʒ{���CL��u���μk�fh�FuA������U�vH�G��)��U�h�zv5^���$���9�V`��̽e�b����=<��
����Z��		��<�uM|z��wy�����俫L�'E:'E���ȒH+1�34]�W�a�egf���&,D��lJ�=��`��,~�RN������t�nV�K7SDX�t��S���d{{)��.��ә׿+ՖԵV0��}����<Q��� [ʪVt|�c�u�4�ͧ�6�_�aM!��g~Amq(�!j�P�d;�z;��2����#�n�w�d8-������Cg+��� %����v�)�G�Q�* �1�VĞa�ʹ�?/p�P���"s��#�w�:0��; �q��U��d��l��n?s����h��� �B��^ �M�"R��)��	��B���j}4�����H��a��"�7�B5>�ǟhI2I!���%T��d`�"�xLb���M��w�dɔZ! q�ǭ̂�`9�l������Jv�e�LfNJ6��s��1UV*nXͺ�Z͉-��ϭBЩ��J�4]G��~e��,����]rӲ�(9��1����e�?)��u,�;3�T��x�;�ԃ�1������y���*�YP�H-�P�J����%ߥ�;7�G.����l��E'I+s�5�A�h����f)�sC��Y��#�6~�p���c�Yn�Q���|v+(X7R�ڟ:�WF�2[�Oy�Y�V6�1�y~�E'>jb�h觋��Zf��3$YE{Od�9��l�v�GdT���9�<�0�R�@�Aq�|�S*���߽{Z�)���ғL����u���N1�e)��Ą=-�\��	$	��z��~X<��}����bON�9����ȑ%A0O��e^ֲ���0T;D4>sP(Y؀�=H��,-٢�I����ӳ]���T�-�Z��|Q�)�l,K����H��6؊S�h�n���F���/3>��TN͚�۳�-�4uOU����?at��*֋�*���e��wG�koΖ_]�sj�G��X�""7@��^U�Z�Gu���
Ԧ���'�.����NF1�[��1��JV��x��y����K�#�$WtWm@^�+��@y?�J���X�m�5�c8��,~Fo���"��L������0�6��6���x�>;�� 
�6�D���!���ŋq��O��A��l��g�D!��Eu������/0��ñ@�y��e���(�+ۻ#���
��G��Ę�活:V�R�����|��ǭ��E�̧��̇�O���y(V��������������z��#]�#_s�[q�8�H�m��F#��F) ��z��{x9��b�-����u���"PyY.) 
+z?Ag�JClU꠷HHx��/�'���fD�Dj�
�cįQ������r�ú!u�L�juۭ�����ٹ�ona�  �XQ�i�C�����ڍ��9�L�#F���(�,�f��Z
i|���ԅ?2y]/6O�~�*���!l$ͩNjӢ/<\�P�;:۪�	�igN� �3(����q�I�K%C�J�}�L0�?�۫�����8�o��U��P9D�e��3]�$Ę�g�ba�1o|!/��ã~�Gg��Y��*J#Z�E�G%_G5;;k��Ϭq�����|r3D���A�Ȩ"!���X"P�����{{.w����0�cR�v[G(���.xOl p}Ya�0m�~7���o�1-��,�Ռ�.D�J$|��`H�2A���ɐ]5��(������%d�ŋ�Ec��,a˔���o"��1�/�#+cE^V��z'��>�O;NҪ���%��s�
H�*Ua�2�2��#��
]N>��kCv�D�4C�j[���9�AMS��J~^�{\|�:t�'��*LX�M�%۩G���H�a�y����$����)���?���R	��C��]/�KU��)�A�TL����њt6�%Ёq�{�!G�s?l��X���v
BYh�(�W�<�a|7\�a��&r�P�=|'Ȍ@D�k`yG�;C�%��|0���"P7�R��^-2~��ca�CQ�'��1n�Oemi�����`c��:&@˟�I��'�㨅����4L��D�R1D�Pa,�ʐ�#4��.���PE�u;i�w�)?�bZ��-,���!KS�R.,��aG)�1���s�_�I(��u��xX|�B�(��,���hm��;���:	f=y�y���KrF�c��ó'J�txQk֓;��G�����[�� (�n�Tù�X��*�,���:�r_��Nt�Z��w�
�Vwכ�֧Yn�c��r�l�����T'��wQŀ�3�$J:�.#�Os�:g�h�='����Q���Q�h  8��o�KIz������
����B� y�D����w|�Z������a!�{r}k���r!xR�������wW�G.���{�%�Ū�bZ�N��T�	N_(傺�[��-�n@��$<�Lʯ��]d��#F���=�rh���u��*��gl�g��;���ʵ_�譯���[��9�X�4׸o��WmF)p^-������)T����c��voԐyӚ�)Oؔb�I�S�nI�Ҋo[

$5H'5aV m9�Q�U���*Y��?䑒�;�n�-:�OQ�3ђ��׹`�����?M�[�ܧkZeT˙�33��2lv�9Cg�'��BC��U\o&S�}�y0�h�Ho)��彫K��G\���s)� ���(�i{P�ĹA�֕������4�T�����"\�!Di=���	B?����)��3�����C�&���yy��+ƀ����Μ.�R�����WV��U|^&�Ow���g��z��B.��r���Ϲ��ſ~����O������g��m��V����g�S�����`�tu���:�<��ś���	]sT�� ��>��ܪ����	2�'#����[�
����S�Y���V�dK-X�<mXН;��R�!A�l������@�̀�ĥyY���!K�'\����9�Qկ�/E��h��`��/�U�c���D�*���v�q���|�w^g=)��� W�o�O�)�
�:z
��g�I(ӒO�oz��P���t�OӐ$��` 8��Dim�����0���y&���Xlhw�p@�HGf�3ZI�@��_U*�4�t�5OyO>�:��r;�J�3�f;��o��6&��8PYۈ�(����GV�����X�g7����'����q��ÑgX��JE��:�4ʜ$_8�@�R^F#u�&V���ƷW�N�i�ԟ���T'bӆ��I���?�m�j�����6������β��$$4-��l�@�!"J�L�щ*�z%q��D5�9NC���������Q�g��gg5N���N�g�)	��n0��R������}������A������Cp����4��'�Q�O襉�LӄiZ�&��j��3j�4��6��zǸ7���q��eے|��"�+�r�&�$&@8N�KD2����i����s�xi8[(�ʁ���L��~Y�Lskf#=`X0dz�$�r�R�&�Ryh�X��|)}<fQ#�D%�fw���K��Y��K����/F)KZ��G0�J��n�*��O�/���i�d���f��U���l�I�=q�>��(��2V��]�zzp��S`5e�����F�xA%*{+I#�bȒ����+�;��Ŏ{&���W�����u���9e�V[x�u_h�ߺH���(3�G�0{`��Z�-qM;$_*D�������n,�J�T����r*�p���L���o�Z�T2�G����G�F��U\-��N�
�+��E^#��!6E"�	w��	KV�Si�>���DLb4�Ώ�6,(++��,�QS8��jp�t]������������L.Ec�$w�Qz}0�Q�J�qN܊�7����v��E��j�LQ�T�B�Y�K���~A�m�|���I㦛K'IN�`7�Z�[�Iz5���KQ�?||�8�G��X�5p~�x�)����I�-�o< +~Ѽ��U��WL�ƫ�������X���1&?�O>��@݀�~�n�LZ�('���๒�� ��r���K
?�����g�����ϣ�Ώ�������5����KmG�4,�-��].��4�XR�Yw7�~a�x8ی.7�h_�	�J�[�//�\�]��˞�?�zk׼|�K�;n6o!!?�v��� 1�]�b�����=ad.b%Q��#�V=.e�}Y�C<nn���S��3��h�\��=�wp��<�Xu���R���2vG\�'^�μ0N��-i�������$}5��?����I `�����Z�6X@B��L���J�>:�o���i�T?����e�o�jc��#�vA��m��\���#>��G�d ���d��NB?�K���X��<Fc���7�����X[�oX��0f����IYY�N�������N��l�����-k�c�����W�����@N�5�O!m�W��x���zl���h�Լ�Z�'��:�� �������PEvOၽ�4U�_J��wDYL�!�s���@>���6.x��D�ʢ��ja��(tVk�F��o~���-�)�C�}W����
���M�+�{����^B�u#�-?'P_ᄩ�V���vJ�|��.�F�&S�3�fff��7��@�x�ԞDBQAkkkaaaE뻨_\�Kn�҅�ju�MPH���M��jL�A�s�8�e"�Μ�9ǈ���,҄����S��x=6���9m�U}3�?��XmFH
�S�*ϓT�H�+���q�٥i�5P�.���XM�4�}*?���b@��!��g b���,��X?oܳ�f*}Fx��hH�k_�$�Q	o��T�z�X���6Û|�]�?pPv��Vi!HD:d#H!�9H��eg�|�[s��a��+��gP�Aw���#�kҽ5��n���J("vyn$�ˮI���Pf�� �����S�ɏƫ���Ɍ����I�Y}� � A����z&�4�UV�.��I�����M��zzefӺ�R���P��<�!D������O��߇e���c����#f'��S�~�������$으����9��IF4��[��������:v�\�j�}�zȯ#�[�X޴.�gf59�X�]� �Λ_�gF�bR;�J%pʫ�
���l��L��sf��gpfP�|MvgN ����X�������OoXG�Y�¨�~��M��i�G���{��ء��?.iK�=G�j#�$���J�ѝ�I�A\�I�a��-����| �m'�mo_�c�S���$�#���h�~�j 9�հ��x�kU������y0\��P�l)�ᩬX4tC�{����m���)N�T�	��~O�Ȩ5+O_�ʐ���#!_+���œ*Nk�0~�A�ą�I ���A^���H=�*�[��RL�F�U�(lLm�������
B0�:Z��w:2<EI;�_�[mM#T�g��P*U"j�4K�!��U��I�M��zD�G�p֌��y=|����PL2Mg�u�K�'Pm�O�O$���D�<J��\�J^w�Vs�I�L�
��@�����9���N�,w{�kuC_����s�$m^��'�_�q��0�ԯ�S�D�7�?���}	ۈ��f�^����h$�V��9����
�iKdW(�`F�%_��d�����r*�,�;�Aa�I+/�e��j"��k�ԿX��haI��Is�T��*�<��ğ0Dy�g���6�8l}gT�8��f�3�n�B���w|~����<�;���<�{e.���8�!�T���XRٯ3K��ٟ�M;q��~�_���4�Bj%�ޱ <Y�ll
N~
5M����W�R�C�Ȑ$��?�}N��j�w��Q X��!����
$�R�ô�5K�~��Ik��@y#P�`bJ�EJ�/��p�� Rs�ߏ�M�婇um��rC����lW�82�+Y��5�Ҭe_���x,T�MW�������Hm!�vS��أ�lY���Fˬ�֙�*;���Y�z錿/f)rl��D?�Gv��[C��9���7S��	���'ۈ�#o��I����=5V��ӆ�o%z� �e�/���Ղ4�ӑ�2�^��@Ʃ{�K�����O�Z]a
���m�/��n^	���!� �Kz����퍘wY6��$.���WBa4�zC�<�|��:=6O�����l�߷����@
� �2��JV}�N��>�m\�����z��+�=��>���R|�ݻ���o?��o�<�.5B��ee���.ƒ�u;4�բ��Jyc�㺌p�̬��lq��`�����@&�����.Fi�,�
8�/�0���n����/y�p@A�پM�bD�6�rʏd8�{��wD�?��A���^CY�� ҨH�"K�,VTO3���mG�n�
��p2SQ���T����n�?,^9�8��OlVŏ����oϠ�"��F��:$�2�)+K32��G�����*i�����XR]��h�mf`b�;�%���NhCKYo�Ϯ~:��N(n+W���n��N�\W��g"��U�O$���17KHr�}�˥�S�����4M��B����Mʟ��
-*�����uޞ���sI�r�RJ9y�*my}1��lF$P����=��I ������TT���(m�],|�/G��bD�������'F2�!������;�.u;®By��vT^�	*?�"�F!�XMӼ@ߘZ%��I��Y6���n�q " X�4۹�N��s��c��j���?��9��S��6�k��~�h.mb�tLPv4�Q
�I.�L�R����a2�b��-o�os��_������}��=��=v�;�M��i���>��V�!}Ň�,��j��숅y�=>��Q���9.���������:��c8�<C��m�>�ߧ�'����'�;���v����>F�
h��!�U��>	�<J�����+��-G��V�<��F�:�ۭWZ�����}A55�ϒs�1��8�w����}��L>������؍pz+S���,��F��$���J�x)\���$*�U� ��k	�.���;Ǻ�M�m-0Z�
9u�@�����Z���
I�)	mHw��z�ؕ ���*q����I�����V��H��w�-�I~��ąF&�7��1֜/��d�~U"�1FBQ��Tg|���h��GT)�rؒa%C��jo��`U�%f
����ғ��4�k�)��C
1lbB��g���_O)��$�@��<���JO���+1��&YG�����z|B"ꏩ ��`��lޟ�c�����n�U$.qy�_�D��ػ�17Ċ_pT��� �am��0�
�_�	�u�b���(�������˚
�rfq)Z�-��~CM�>6����<�Ϫ���"p)��T��l��x�
?O���1s��J���4�BsQa�!�BP��ě1��K+�y�Y���ѧ����׽�3q��2�P���@F?��b�K������OC��W�#ϵ��U[�SO��F-ʲ� 7�� *��%�����A�bO�Ag�0<o+���L�P�Q\�~��O���[i��N�� �e�]F����kP�����dϓ�*�PL��$�,Lw�R�N.�ow6�Y,Zѯ�b胐�9+Q/��kB�v#�W���1��,���(�U���r=��.V�f�WYn�,�
�d�-M̸�ꑏpc,�$2�$��Y,L-DM�8s�q�)& ���!<�݋����n6:ʺ&�.����y�5��?E��֩dEK�kDY�0d�DR���	��z\�p�
O�l�_	ZD��g �i@j2���MbG�B�a(�n�d]�u��QM�gLPx�঺�C1��H~*B:rIWl�@��s���)G��l�H�t��%ߊGF.�ě�eSMFF8�磥
5�m���v9#A�*�m��Ep2��2["���W;�w��W-�[��Jʦm���g8J@�2&
q���\Ӥ���4�Բ	;{'^���|>���y�֙�1�|��S?�=�>P�S�3�#N"%B77�Bv����\�N���C���,D��R<��1W�dI�)�p���"�Mn/U@(�@a��b��Yz�03�[� �p���T���s�)��*�u��G�b[�`۲ݷAvy5g��f����_X>��l�El6Y�VR�F+�z�ps?��N�i�� ����k��t�G$��G�X�Η}�j@	��T�v�׶U'�7 "�*�"�CA����f�8ܿy�_v[�h�c!�ͼ����o�d�}����$�Q��;�7x+�YSJU�T�'�)jZ���@69դ�Nwm_�����O6��xU���~a�$A�Q��� $�|�P
����	Z3Q�@�=����5�"&W��Ī��(��G�t
LQ�R.�VE�����Y��a���-��K�����
�n��n�n;�B��J�d+�R���ҿГ5i�^�6a�O3�x^%������
3}0Ͱ.@�75>��>O��'�^m��Ze1����˨%���V?`��eњ��6�fʌ�l+q��Y����tT
g���* !�6�����Ú��>>j��#��G7�FJ7���iaԨ��t���$^~�{��v]�s�yι?�Ϲ���B�W��|�s��p�T.C-h}t�����$����Q=��蜮�"��ŋ��S=u���T9e	ѵ5�Q�Η��ޅ�_��֨��c�'|�e���h%�>��(�ŔsU���sf��u�gIUU��Y��%#Y�蓞S�3$_������VM9x�窖�o��i�=��.�����*␚��*..�H~�}�لg�܊�B�#��������qtx@֮�*�nzw+S�4@,�(��q�������R��;Pl�Ih����oR��P�<��7��	)�[G���	e�\��	�Sa��+]R���wT�/��Z�t�z ��Ä�؜,��a�D�~�?��tݩq"]������9�{�
! ,R������d��ē��DhX�1/;���[� �
������zn]��Y$z�S��"u=-߯�o(�(�]�c��Ժ�:C��/*�H��z���I>c񾘩U<.?U����r�h[�@C��æ�"��9���e�K� �UU�jWF�w�PLZ�o?Z+�w�t�g���J­�t'으���0
{�U|����H#��6��y�S�[�4�dfJnϧ8}
�"b��B& �8���$�>���k�Ҽ�:�$ݻm�dN�4r��Gzx���]s����w�q+<���&�b��QFH&�3X�)��:w�����]�͔� ��k)Ԏ0zF[�hD��&�����D��e\Q!*"<UG
�%5��;L�G��|=�^0��L�l	�#���R���3��#��@6#� ��X�݈����=\#A�s��HY����x�25_̚�]�$�-���1m��N,�8Z�IQ d���~� �%Y�m��ue�w�E@Ny�0hϩ�LwZ�I>D�F绵Z�h�>A�YCzڏ��D��jt�j*kŌ�N�F�5����W��V��OZ릗y�0�X�gQ&s�PS�+��8��,���]RY|����2�"w��P���j H���;�H%9���Dw���±��� /R' D�i�����~�6r�D�E��K<1Y�Ycl�D�����ˀ��"��_H��P���u6gES���_[��jq��'2?sdG ��ьl��$��t������7%��7�@mS��O�'�3����x|�|LI�����ښ��{9�ZD�"*{�A-y���}�mʔ�Q�ϯ��8H�c�������co�y�3���E�w��	�2f��GQ�R��Q~c�wbb	9v�%���ð���z��-;���a4�� ����vI��3;����kǢa�i1���p�Tf�~�=��� �1~q_A�_�`�df4��L��Y�����a��ˮa�^̷��*�6E�[�:���<>K�775{\����IUN��fiN��>.�?��D.Oo�3E��.�E��\�l*�W~��Ỹ�!����S�)�HZ���;��T0@�M�VS;��\��t�1��:�c��;�ϦP;hZ�5'D�;*��������Ϯ�"��!Y�K8q�� r��O2�/�C_�Y�*��U�ųY���Tq�n�P����j*�
�6���荖pl�|��V���)lrL�	䃦�%"��dy7	�%on�IB��.a����7�UˬeǠ�1of_I��_�L?����c�ig�3��j2~���1�` ���E�{�/���R��_L(ٍ��Lh��i�ҸSK��9�!<��R;�H������)���e�J������JG"w��:N�u3�\1=������3����Be=��^�b��S��3�ڏ,ОC;$�=��h}�f�m��������
��s�c���(��u��l�:��_T������;��sM�G�4����
,�&f)���J���No�~�H�W,�X�Z�G��T�YP'���ׂ`#v�3Az�

�o߾����(USQ�.�}[5gW���t��'�oݧ-..�^�w���]���_��糚t`Ih=��	$!?�n��Tl���1�$�4H�R��)dk��|
�+D ��PF|�+���D ��!������=�1���,%b�
�0�%%�!�d��� @dX.DmE��f5T@)"ɗ����Xm�"��X�^70�
�b�Ǹ��[���p"f�q�fw�\��[�S�ݴj�]7
�<1�:.�2&�<�4H��=2��	�m`��/�*�v�z��!�����[NP�v(0x�a��U��X�X^>W��yA�H��B�ŵ�j��c������#��v<&KT6Jr�*�l������m#�p�<=��x��D�~�3!�9�ڜ�ܜ���%7�S��6��/6@��
B� =a;���~� �Pe�R��Y���qH[���݌/��0�%㿎��i"��#��o����;�'�?��=�{�k�,�
I��L�پ�@<u
�|�Y�08Hk&o��=
:GT��"���ȩ7��#�y����=�������Ty���P$`;fpvP���N� ��sV4�ST$
���ϰ�3O϶����B�B�Tm^��􆔿�b����,,DF��hc^��Ӣ����,�.w.Vv�����h>��W�p�B٠C��j/���7�3?$���:,�{�	\���}щ��-��I�W�9R�8���#@V��AA V���lP�gbgM�I��'2`��'QԘ(��mq&>�/� �R����� ��x�:��v�����ޠ���
-Вv��[6�H���S3�%�>L ��9⃑��y����.1�H���7���<���w��/�ʋ�aͶ��siN���r%��x~�'�TW@�����R	�Ép<g,�x���]�q�kK�1��X�
���e�����a���_$��@�EzUQ���Z9�쳳�Js��5��^N!�aتJxec�/��
t�����6L%Pİ�ZJ�;ϱM-��j�ۄ����q`ァ��
�������e&���-׃�LRiY�G��ФL���w�I7y���*�a���/G
E
榗Zd�PR��w��_�W��T�ij�����5{�T���U �����OD�3�m�b�j^��M_\�<%cAA�Et�v�� ڔ�H]��Yѫ*���P5��^�WM�����(�wC�u�	�O�*���V~kG�+/Y���
�\���U���+d�SB�Ȏ��Q���.�/�?m?�� g��� \��8�B��E�m`���GԆ��'�1sF�PY<��Lz̓�i%O�H���N�C�-�גDڅE;١�+�y�^���"�0aмR���[�H�O��89A�Aj�^��3���Ѧy���נۡ�ҏ'��'#����TmP�V�&N�%�5Q�cc������ڜ���2ʵS�q�Q���ig-�f�GSQTL�r��	�|�gk��hp�c|��r#7���#j_����-���ht�)P!���/!�&�{�C�^Ↄ�Kŝ��֯�U��l�^�0��Q��Eo[uf�$�J��Da7�����2H�FC��ErfffZ)99v#G��k�Ȗ�}Jg�ttЇ�f��ߐ�)�<�_!!�i�,Z���<� *�|�+���=��׌\�9+'��z��U�{���5���q��ś�:�ʪt�_M� ��c�1l�ݗC��� ��	2e�h�«O)��Y-��5狱�-h�+���s�ކ�O{��>&�l�VV�v���#�c��b����Y#Q�L��L�FA<�3�7�VQ{7wy�LkA���J/�羕�a�`���챊*�ٷj�:
x(~��4�0�'��y���f�'�p��3�WՆ�S��{�?fK���X�͇����3�͉5򐜅JWUI9VY);���I_�����E���Ǉy���󇭎���^iPW`���ɩ�ɾ�ղ����ގ6*���Ӱ�?x̹(��|ة�n�	�B^W!T�Ik���iJU�D��=��1�)7�/.	���|C��o	J��xTS��b;y��#�I�uE���O-Pf6��@�d�XZ3ɬ��h&�0wY�b.��Yz���W��mB@Tw�m� ��w"��04y�fm�^��n�;�Ŧ~C�5C� �)���'�D�����@��Y�?X�Y�O��=#����j8����fvH~����X'%�]��>H�	��g�p� �B���L6P�j� �k����1saz,x���>k֩�{ˠ����ҏ!��4&k���m��!+e2"�3�^��&����BL���y���;�;3?NA|��R��x��S�$�>X����J�J�Eu���Kb����4"�� C��>95�����m!�d��RO��ۤ!�������B1@�а/=�ԫ�`w,67�gʔt�-Ŕ׹0X��ĬR�ɉ�U���Wʋ[fs ���0��_e�r��0@k ���6�(�ؘ�s��Q�a`,d��â��o�ᗷ�������c���z�-�P[�A��ݗpH��*m�y%e���1&A�Y�*����#�U5)eG� �d�O�P�tR�Fux�X���3���G��&���T�K墑�����g�����Q�2���C�h=Tg4���h��;*R��R.��פ���Ro�	���B�B*�rS��X'uOu�sJT�m��;�إ����<C999��>�z~��;T-�P8��{�Xn�X��������Q?��*�;Q!��y;����o��_xھ�V--i�V�4ꒂ�h6L��b?��v'ɶ9G��g	��4����ÊK����E�����H q$4��Ov'6�$����;("es�\��f�
ֶ*J߶�����>�0W$Ǉa�Na,0�W���cA�J�:��L,�*���t����ȶC�̀��'%�Đvu+��T�+y�p�����)��8�[H����'���*w}ԗ��g��f?����W鏏oW%��v����ػ"l�Uz{U�x���et	���Vԙ�7�cYft �ȂW\��
�o��Oq?�#��Nd �	G�9է�A�������A$G�s�j�=���'��;\ha�p������#��R��=E�~J2{6^� �.�0��KGL��"�9�"F���`䁠$��Ĥ��8>�����\�\���C6�k.�}�}�MTi��ttR�؊���م����׎륥�;;;���{���!���6����������X7b-Z�x���x�`=������I2?x�O��L��2�X��Z���kK���(�`����,��.P�>�C)Sm.��Ya�����'�5�i�kԸ��W���I�މ0tb\֘[�����Y	|�Tӱ��|Y����3�0G|��8]�e���b��`
�u��z)16|�?���ߡ�ۑZ��q��0����h�����&�@�;�8�:��:ZqW�a0����bkrn�g�!�WiC�c��V���r�?��E}������{_mv��L��������_�t��w��n��R]�>�n=�ҝ�#��7g�n	+mm'T���3o�k�X�j���C������z[ץ�%���i�a�.0BT[��}�G/�7Dw�LH/	.k�����A��!����e���ޓS�=Alл4��0�F��"�ӝ��k�|��B1N���nH�H�ZT��59�j���@�Y�i��7	$o�����o��2]�:`��լ����O���C<1��≼|� 5}�)� �v��o��|���p���7�L�r�1���a��g&U0Y�^I�'k2z�8�6�E�����#�e��E����<�,k|���O�c�M�ٸ�4�K�����_'��[�tH��3��I<�� =���Z����!�316Jaχ����1��q��0��p*Z�����-�t�;�dg�@1+t�.����WH���:�~��|u<��<׽L.��1��VѬ�`��3M��Z���X�XG˵��I��'� ��G��O�h�u�&w�B����d�~�7)$[�'�/���}*_�w��� kx$�W�`|R�~r��B���W�H �%0��JR�00�"W��+)"0e�YEO_�\C�8vH-nL5ZGQ���Q�Y����C���&��j����0*bu��'�2��XI݄��<�\�c���/�9�����W�)`��Z�v7$�1�kD��Ɩ٠%00Ez�ߗ�OD抑�*�<7�a`Հ����ƨ�;����3*f�
1�ز�·j�6�����y鹃5L�4�w��<�q�Q���A5��L�>3�q���t�!,B�*��+%�e�#�-�̠E �5�q�ډ��SCvԲ`�rK �3k1��g$�C/�/�=Y�<���@Tz������|ʔ�i������_�:���S6.�5��̑�~hȸ����N�9�Z?v� �C�k�w�[��eO&�: �0����;�c�J�X�0� |��N>P��!iU��)�诃��y'�%N�pH_1��M�Ix������������6����\yȅ��ያw���l�wlfnG��G�-�y �z���a"� JRYy�_Jw�J��rF3��T��n(���9�/�퍖����8���M[c��l��*���y�MwJ�:�*�A��u勴�荑�O��^ƒ���O��ļ2�=LK9NO�,	���-�O���k�"�0��LS�D�v��9ӄV`n�9��&'�������C�:�6�X�u_uPԸ���:� J+�I����U� �y#K��DEO�����h���?���G�Ϝ'�WZZZ��������t#��Hb^OJ���������F�k_4,??���E#���0��	���ͳ �˩H�a�O�y�@��-AZz�*@���_�ۍ,�J�9�����&�7O6�a`$k��K�hi���5F	���U������9x���{�A��gK
-�Le��!N��3dRw'�r�h��W�������WzN#��GK8(�շ\�v������`��"x�g�
�$�p`�� f}���d�SM�*��f� �_��;Y��\�X�酎���t�Sa�C���0�|�����۰1�����t������:D.O�H��e�$>����"�����u]������ϗ��Z�x>�������u�>���zδ���n��-���
���i�����bӯ���t�U��'���2o?��M���|�e�4���蘃�@Obt�3#~�y��	̝���ï?G���׏'od�H:�4~�i����{	$����,N}�Bopm��Qg%o$
	�=!W&̜�z~�b���[�0@�.ɿ��;�X�Syz��y�V/B{:V^���@��Ԑ/l���#�lv�s��BPI#F\�K����SHX$�Q�HEfO���$\gO
�Ta�5�~Α�$���t�/��Q���W%F	�O�.���J�z�@�tx��X��8��'ȵ�`�sUC�3ٗ� W�`��.��O��L��F]˂��e������O�[����hH��
I@�=�p;A:��ʞ,� �'�Sd?2qn��u���bR����{�i�a$Bl٦��,'q�B���"�%3.'���M����f�
��n���Lv��!s��X08p� ����&���;�o�hC�0������FM_�N蝅�)�*�S
�=\��YBs{��P
�C���p�]q7��$���a���D������A�|�C*���r�n�*��Ϥ��E5A�:��>{.�F����?�O �3��s��u�{�`�8Dd�F��tA����y����{��0�R�F���uU�4}�tJޱDr��󺍽�So/tn�q/��$����������n�#�������e�	Z����ֱ�{kj�ߔf�������$�_�q{�+1]�����Q�} �{7n'9A	[#��Q����;��%A��,*An�lr�Q���Ӑ��y�!��:	���>:����Zt�iM@�'��e��q��~k����3
co�^��u�Wn�d�މ���e5&H� j���ڐ+�p�amK�C�.f��V��J��,����2�� � � ���ˡ쑆&�^"��(�&	�g����l�I��{Hh�0�� A%ֵ�,�3>Q�8��ym�=ҮQ�_��J�KeлbG��m\~�W�C���֯Жp���������7�?d�O��o���m����I��_�k8�KP��r�����$5J%9��B��5%9��l ]�`�D�6E,�V��v9�N���H�yQ�Z�4���u�{v���?Μ��K�tۓ��<$�AZJ;��PAm�����X.�Y�K��B�x�R)�;�^�ac[5ޙ�:IR#�
�^��x8�_�&�����ɾb`�/�*F"{�{������JJJ����"�][���8|�V��뇿]P�3��a�ev��h#xk�i�>�NȈ�⯽'��_k�RdҼpN��Ȅ�.���ְV��?{q��f�8}��1��Bl��  �����3�n�J-w�3�" �O�4��&��k�@������ǂ=s��^��#��^���-���F��s�}�<��o&���O`y�?P'�_o�&�����X��E�FU!�)���uU7��<1�R��5�
6�����5̡t��_̍(�\��ʻ�����s�]%����t��-���7]��Ś�X��,��Ʈ���ι�G��U����kc����ǃ�_�x����\j�������f�������h�}y�BdV��r�n��������׎9�c��YΎ&�O�n�+�T_M�|l�vfC��5���A�҇m�и3�9&���?�b���i
l�&�M3��I՘��%ܻ��*U�#(�&�fy*}�0~����0�Γ�Y�5@4�B��{��ؒ��s]��p��x䎹�:f:���ݥ��e��G�	��t�*[�+3�ݡ��*1���G���������ÂOP�(L�R`�!8��J�la�&���YRsk���:2��m��,1�q�R��`��8����d��护;�%�����5>�T�+5W�/��ZZL� ���k�r.I��D�^ �(��KQn1!
Y���a��4��q`�����i~jB0&�Nc`T���N����d57gZ���4 ��|B�t�L�s�r�i2��k��K۝D��A��A�8Gj�~b�80\*5O�Ɠz�-��
?��S��(�g���x�,��B4T��{�<�c/忏�=W�}�����B�q�{V��-q���쭝�1T>OW'h�׍��	C純� �+&l�6���#)�z�N�#�UX�)>��ꑓ���|��q��M<=^�������d��1�S���<��D��F�c����1�~á�T���Q�o�����Xt�î��G�9$O��2J�Ʀ:xt;\��F�r�J�Ba��	;�y�@��P`�@����VF���^Ĝ".��rg���R韇��4˝!j�<�6@5}W�8.-�7\W5%c�u]���$'�fo/��Ǣ�^��*��������j�������������o���������N�&`�����"�i��ժ�o6n�
�k{c^��h>:���6t��|vc1��n!,Y��f�����e�?E�dT��J�Ic�G���VbDp��˴�p��Z�$����4��P�n������~G��x��_l����o�5�,}�=۱�YiIQ�(���;!��Ut����>�Ds��Ia�q�E������b�A[R\]P꪿�p����ࠤ綤`�5��c H D0���YZ�é��hsBFV}l����n~{B&�mW)����SZ?X"kw7v���IZU��|� {�G"��'�⽒�r�je����/�nޒ)�C����~*6+Y4'��A�,��/�&;����h �r�r�!Dl��Qט��O�H�uї=�} ��B�_,$�q��*�Zo��n���ż�㔔!1�co���8j�*��P�;
|%g�J����KJJJ�׶33�ߞ-(�A�@K^^��I��6��|6���'7I�Ě��l�\'�����ח	���)|d�4��m`�ńuƖ���;�MX�^�
'7��} G�1>��d�y`*���f�`{~p�(�`��	A.)xD�_ �������m���5���X����m2#�\[�BD����&|�h
�b�W~c�_j84����S%}+�(_�/ÔIZ+}!��Y�תj�0�R�H.�c�>���_����M��Y���k`g� �����O��˃n'�]�����j�����������_�^��ǊХ��{�����2񺙞���ꋢ�	l~��j=����Gᓁ����j��1�?7`�/ݷ������\q���.,i	*�=����v[uh�(����p2���ڽk�{]�����,��/�F}�4R>�|�}����]���[�r�o�O؏��*�F%��N�+�kߺ�hG���eޑ�_(��r�����aĝ�OL��.�`6
ݴ���.5�9/H{˝O���������mM۝�g��8�)HRcA�H�(��C�����QL�6n
�2��֒²^�ǩ��L�ϊ��I	e�����"!���2��2`j��[�O�M�Ec�4���˦�P`��d��)��-L-��A�>���q�O�����		X"1�{C����q�C�J?��_�����!ÜwG;�'�Y��҄&I�;�&}���A���B��3E�-`o
�0��ʒ�lP��;��L�)�f�3I��0h�0�B� P0|�
&~�7�[�$ʈFF_��rV'��~�����,7/��,ɺy��}F�����Bb�h�Ѩ������!��Y & X�p�� �E����I��(�0%3�2Y/(#-g��s�|����u ���M�Tzy%@�3x��5�5z��/�ub���&�D�cT�`�v{���j��W�����T6�?	g���E�g���֩~���am���S��M�Q����ݏ��5��В?�q 0#�N��X�����IB0�Zuk��,GU���2��VT�G� ��7�j��"��d�z)�rzɻ��-�c%���cY���;�N�k�����=<72���~�=!�~���eq���9[X�Ndb|��9�0��/5���[��kv�l�aB�'��M�vSv3�rU��,k��U����M��ta���gM�ڨ��>�+�������_@�N�/�:w,V\��\�gC �[T�����ͤ޶E�3��D0x��8��l�U�����ܲ�%����)�j��������CN=e��T3/�׵�ܯ�Wع�[0W	񽴠2 l�E+2ʂ��b\��@=��/��53�2���� X����b����Sҩ^NئG�0<���&ﺾ�,s�f���H��t*�yK��1�=3jϪx2g͗y��c�>,�T�ȕӰ��eF��^M�C�0�=S�H«Y�o�uJTH���UK�T,R���(u�iM�_"F��U�H������-���>��:\��>�ȶ����ǟ�-���R��}�\k	lW�&�{#�4��Y?��;���2�Āb41�tg��6�����`�PHW���N]nʩ�_�O���#`$�G�3�d*9��ٰ�/��[<_`�#�~�w�Q:���e���Rk�g��k+��H�尭5���	

B���v݅�F�f�<J���m�#P�nB't�,�ajac��dB��	��1��e�&*�[ZlN��r&R��N1�Y�I��);B8��?�m~�hT��[%�4J^��l��]G�$>���M�c��/��9����d��� ؖ�jQ�`�^��d����9���P��S��nx�W&���=0Ax��/��{fW�lۗ*�[n�2�U+�B=hz T}e�5&ph�L�c�-��_Ke�k��1 ߮P��$�.��<��mQz������ϝ�ކ�����m��	��fU�EU��M#V�;?��̶E|]��ـ��4�t��8I0��t���x}���.��Q���u�.�����C�
�����7����LE�^�4y�+�e�̻5_}%55o�2�p���7�^�y�8␳z�� 7!q�䶖V�:��ld1�KA:|}mh�#��2����5�n�B�E:�̾����҄��|i@5�r�FG/ژ�$U�ץƘ���uczS���a�-�::�d9����!��]��:�a���Q���Mq�k�j�}��B���	%r���2 ���E�)b_b��9������nkB/DX��pl�j�h�YzO���N��3]���Q���_*J��PS-�O��>A3Z�	Q5��ı��ƱH��0~�
���;sW	�Jl�Op���L�j�0�E��5	��b�=و�7C�-H��Jza��y��7^��4l �]�6��՚4������^~05�Y!�k��h�,�V�����1��%����1��^E����1����a����.C��6_���,�Q����&򗚀���/8�t�gP�����}�W)ə��4-P�k��`����!�O��l�
>�1:X<'���_�b�@C$t�v��	�M�����[��o4v�AJZ�3��*xG��vT�(��@\޲Y@ ����g c�eِCH��r��ͦ�gmxߥ,.���9c`�U����`C	�}kg��"�k/���r��5�_uG*'k�n.�^����+cʞ��ӓ!Y�B�-v�� �Z�C��e��؍�_�I
��U�����
�[NziVE�L�l̥0FSt=evK�9��UÖ6�:� '�H��$�3�t��$Ǯ�~�������Ů���J�g�G��bh�������g��Y��՚�!�9H_G�ˑdU��}[?r5!6Q�Ĳ�tG2��^{���XKj}���Dм����u���+�r#T�����,dl��V�=��ǚ��W�t���@����������_��/൹�5�<�w8��g���ڦ����mMvRM�?���<Ns�ƜY��c��MM\� ��3�M���Bn_��sv}�&�d�,s/���5���xf��E=�2��f\^5�����qpv��a�;M�����!�ĴȚ�D�P��0z���OL�����eF����U��*d�߉>~s����lg�*�W���I�����O�����t�-�G�v����Y'����֜E��'�7L�>��yh�&�,�QaԚ6`��o�$��B���E�{��.+�,�EV0ޢ��<'oe�٣vY`��{<�Ћ���sd��(v6�Y�89��,2���(��0��K�����B����;��x����fѾ�������ï����_-^��a�>6N������KTd3�ܶ9'�_�K2��?�Ъ<W�A8l����M�+H����� �� ����*r��%�Mm�y���֌o6H	Į���u�/!|�[��48K׭��������;c!�9���"�Y�Eඬ���(��>HB'o�P������Z��J]�T��:Q�+�'i�À�������Y�-��/���vO//B�2�!99�[\�;U��b�	�gj���q�����pPe����g��W
x�c��	�؃-�`rZ�l"��!���t2����@ϯ�4��p}:kX�TC�;�#l ���<��.��]���߹qQ���$�N��#�0*�.ɂ<P��U�>���7�h�j(Q$k���l{��/Lޓ^$ >�َy �hc��� Q�m�1Zm�顑����U���Pz�ٹ5�R�ȿ�Õ���Y�1S�f�1}ڟ���j�㞡u��e��{�o�\���	�c.cc&˔�^�A+��MWD����d��[�p�s�+�����Y��ɚ�T��K�?�&��~��W��w�
�Q��tA��"��a'�"��e��τ�~�>���8@����j������,�U�s[[��2���K��5�����<"s�"�K��@S��ْb�ƾ�1U5������>�9�w�N��fk���W@���|2��"���C�Ok$��7�B��HG-��y����J�b����a�q�~2����q�
2�f�8�ưrh�1��L�I�(�a�BƮ xm/y-|� �ׇ�����z���#h��q*>I��m%#�f�9���j��=�lk׾��~���������p
д����1�Q�T訊˝G�R��y�@K`"Wd��T8"�-�r4�0�!C/���]�4܄����	���o-\A���0���*VN�k<�3����gTG�TT��ӿKx;������<a��eo��Q#iF�7��韛�)��-���m�a#�C����T+F������ yZT��丧jh��r��P'�-w��b\h.+GK�#:����1�2,�e"z�S��V�x����g�<*��[P��p��_����L&�Q^0��	���S�X���JuOR���w$�����F���A/rl����j;=�Q�=�#��E�j�3�{�>-��&Ìc]� :JO(��ȨV��B��7���b(:Y��5��D�&�	��$k	�V����"��۷�����@?�
��*Vs���O���r�V(��83�
̕P�W�e��'��G|hO�����eF&~���0�:���#��=yzJ6�+�]�	�������RZ��f���b�M��a�g|c6k@��&ԯE��_��F����s����4w��SM�8��v������x����mdi^ˀ�U���H�� �ҵ;��U��+���ƃ�4#�T��DF�m	Y��;)?#sԂ<|B���j�c*�|�Tև	uJ��Cꐳ�6	�='�u;�_�̠�FTC�3��_�}��>�ߊ�4~Rˇ'�a������t�qn���`�W��x��e��F`�KY��\Я�>��Xr�B��1�@j{X�	Q��pף�G�=���W��`��7G�\��$V�nz�R��2"េ��Qm�dʷJ���3X���@�H���D���Ȅ������YQ��˛���o�5�����Nt5�տZ{�}����:�β����e_��� �/2���,F�x�K�wT:&�T~����[�0]�������� M��'2�vJƕ�a� ��hp�%�p"�Z9(ǡalzB��B�q����U���e_Ch����������^kۺ�齂�演pX�&Iu�����	0��Ly<�TN�����$�	!��߿D��6Y111YYY��c���66{��ES���N����p��L�T#W���{	"���ͩB��'l�A�6�?M{��*UE��G
��x�Z�5=�~�;�#��Y���f��PO���� Oc�D2�rn��X|�?n_Tj����Y�!R��;��`@=�g����k[{�tC3��5��\�k����U�̿o3[����ڗ�.����ۖ�u��Z��q���c�)S�O�KhNi�/�G�ZX}�w��X���|�2��Wm�mڵ�Tu};�q�����5���a���߼j�j�W7=�t��Q�?�~1P��x����a���Q\Ͽ���-f�.�n�$J�~�w���vD4���l^o�a�3ݟ�B�y�?w���Z�-@�ͫ��������q�QN�!�C�l\���|,�b�!	��諂���i[ڀ���F�$����>�A� �����`��&��&Ɣ�x!��0�tf��a�����k݉M��iߨL(4	���j��Ei[�N��`�V��/��F�L��P�+ۭ���k�K�\�M��
J��&�SO�9�~Ϳ5w���C�{��8&�Ǭ�����nIubG�ǜi����,���.d�2�{��o8�Լi�x�:���=pC�� ݼ�"m	�� ��0@���ٯ�� ���7a>?�x��z�.6kAxDw0���>��>400T�wr�a���~m4��_ɯ��{��#ɒ�22'�~Xg�Q�<g4nk+��Aܟ��1���
	)P�e�G���ajV�i�fPA�gr���H�P��Ӭ�O>ŭ��!$й�G̆8���W�fV iR���
�N���/���W�dr���/|�^!�=�C0 �s������^�����}�z��\�<�Y|�5���*�2����I{q&1�md`�D�{j���
�q��DU2�B�_F)����m����pN~��V(�r7E1��,���a��d���J̇'[4r�q��!ét�9���k9�4�7z�t��a�Q��J��H�M9���啞�P��E�3���#�3�_LԳ3���w� qS���`�Pb�D5�2�}#یѷ��-(�9��t���p��Qm>_n��k�K�;Z�whq���T��,����R�k��w���s�ZO�)�&Of�}��{o7���}��t��	��K��p���������~��N���%���@N������-���Br��#t?��z�����+̖f��K�6�7�"�9@�o�0�I:4l�IYQ�臄M�!���5ygbV6���i��z܇߶�^��E��L�M(�0���(Xf�D�+ݍ�|H3�_��	�M�iK�R��I�9��k����9}��AM�h�H4B.�@�N�B�{)�h���Z�L3�<%v1����O��@�����̌)��D.#J-�4_�� @)�Mں][Y�y�������P���RiS��Sʙ��nC*x�iy��&d��cj�xtJ��GNws1"�}�r��@\c��:t�;������m#����Cd�n��ӥ�����ܧ������[�3�K���C�84hR�K@��K!:� �r�dۛ��)9�G��_��<~�ވ	Z�TĐ��q�+7����fPIA����PK�!n�,��Y!>���%�ҵ?�Ӆ�G+����m��e��+6��n1p�����6&��4����E���%���{DD�����B�&V�yŌ)OWgg��nkk+����{p�%=�����i���3�V��◶��Gߞ�)��u�}�����Z������a��"���q�۰-�B�r�^<eG �uI�yI���m8`�<+������yR �/~k���*�@&��0�=��F9x^�}��
� i&$@{R`�MmPo����u��j<��r�o�K����1��|��/��M���}kVo���TLf��+��c�tR@�����-�C�oฺ=D�9���k�����Q�g�[R[�U߼����������VIC�K�߀�q��0MϞp�����|��NԊ�lSM�_n�������2�۫ʼ�9�;p]�ת��������xKn��[�~40��b���PcsbCU�H�]�f1�^ ��Y[�M1�����N��\��(x�Ӈ��,���:���ɦ���X��@a?�e��8���2BxG�fͦ�EO7
.aL�⻻	�+X"p��]Ic<�K�D=�-����M��f)���Lb$��K��'0������Y�@�e�Z�,�[T�v�yZ9kS��G���qS���L-X��Z�ØA���2�����A*18fT����XbR��rb�a�%Y0�����9{��#/��і@J�
��AGZ\���F��CP�����k�N��JR
�=�Fi ���A7���4 f�(�c���+�̃t�[&��g�-�Ǟ��J�oH,_��~�fT�F��;�PQ�])��u�tB�
<[�-Ãl�L���	T�ZF�Bhu�������<�è�/��PZ�cfe�䰱թ)I�Xl���ֶ7�mߏ��.�#_��E�#��k�/^���m<���#6,�L�!�t:lڊ�&����#���Y6E�B=�>��W'���_��A���V(�P_�$����i��䌴��7)Ϻ(?y�fƒУ^?;V�F+�=��|>"٨Yӵ>��oj��5��Z�T6t'֌1}>%}��C��y��eio�Ѹ<����XZ:�2�׋wD�u2�,��d>?{��C(��^����n}����o��&��y�oP�O�Q����5z�ٻ����o�R�V����9����!�uK���Jߜ��'�_D_3��n�q�c�?*v�Gom�qp�Y�ߔ�.u��|v+*��n0
��B�~ip]�>�PԸ�x���wN��ah��ɖ�>�.p�l8��\Z����^�S��F��^e��Ɋ����j${�bH2LZ�Y���sb��J(mH���$��v
�����;�������3��M�0�Ͼ���|K{���3�P��� �����-�%��诜��e@���E�ct��g���x_vB1F����5�G��㊳���Pg�əE[��#ǁ~��~�m�����ٵ����~����vm��ac�AT�L�q�~g�Kdo�X��_�k�\g�l��9��;,�sd�u���߲���Ģ�آ����5��*�X�c4����F��g���� a���v��G"m�y��3��i�@�N^Wׯ��}m)�{Q��,RS*>�:RS��$����L��hp|�%������i�":a`
5^�����7k�o�a=�p��]�@ T�n;W��4"$,,,$�uFALL>�Ǒ���TVoP��fff8h˅�����=pyg�{c���nF�r�.��ǩ��*g�8_�-�qb���^�r�����K�����{�z.�M��M���X7bX�ۮp̙<���T'>%[�n$@��m��r��Uh}л@��a�_��� �ɛ�ؿ�ޙ��	��˘�';�t�T�'�7_j�Śy�ǟ��o�\jMjF�W������ %��Z�6o�Z�6xw7z$\`���j<�<q��#i���`���u�AYƪ
���K4\V�ڊ��j��D��l�X��Z��Ϗ9���l�o�Yi���^��s���O2��v�{�]՞�O�_��Tk����'�ɺ\y�4������'���3`g%�ٛ�����jRL�jך�e����kU'�.�_a\�bG�mu��M���-���X&Vx�� �]n	���L����ad&����mL���>��?yR,�[<��	7�J|@��Q��5�5��;	4�'X�x,t�ҽ���^�F�p)���P��*f�w����c*��|��к�*:�BR��c�f�&���f�
�2��$����U�ߌ�A3��&�j�FJ �\�b�=�.�mMx6Z+�6c���P�q�a,�?Hd��Y(cȥ'��
^7�+��e>X�)����A���S�� 4�j�!����0�k1�- �h[��8�`Ym3��*y���������&�@-{��I��ѓc�X@��9� (,�gZ (�@q��f,�y��NT�A�����8���{zRa=&���&����Ԃ�`�[J�'�/�E�;��W�6��v��G%@�߭%É��U�r��"�2�Ԓ�?��prGߨG0�������!"�S1���Ӥ�]�p'�毯d������E:豰�[ep:��q�8ND��"��O�נ�	gO������)i,�X�g��QE��z3����r&s�/&AS�&�<��H����~���T#����-�^*_��%����.
ˌc��y_$���1����]���,��������Q$�t�:^����\��>�y���_�q@���������-N n�>�����o�8���27��8���Oyz�.�U�pjXnO4q`uw郞 ��a��s�U�,��K�fs���&����.X�TW��*#�����:C�6��7����$��t/>��bu)>�?�z�z�䒸�PT4���$��]�ƿ�>��{x.�j�W�+Q&+��$�!O���M�$�� �Eՙ�2tތ�N()h�VQ���#6pl�EK�)c��z'�.��{)3g�u�;
Ѿ�S�KZ�\*u�h(�&�cG�~GM���� ��r�G��v�1������Mq߃�'Igd�����6�=�rx��4z8דy����������;S%g[�^ ��YE��w�4��X~��Ëg��u�������y�{�s�J�LE�rR`^J��� <��ν鹺�S#R��x4�@)�����H��!؍�yO����������J֥I�UgM���m��GW|{��&���Ka���(���������>�^HH7w\0}��]�a!#)i�Q@B��/q`�A�.����0�������L�\��ry�m�ӄ|��p2�8��蟧)�b�_��1x���J�F�]n�\�w>i[τ�΢��Ԃ�������t�
�bJ܇Ki���"��5PB8cj�m� ���fi�zW1���[ �爼��èֳE8�S���r}��ݹ�F�'��W�eEV��ʻ�����k8�b�\���m0�o/[(0��j����"�h¤�6�����b,�֡��a�ү����f2Kk0GQ�~	��4{�k�!���w�~2����=�a�m������m�*,�+m"�o�b�w������}������oZt�#�����f�a/3�Y�;������F�K��>�K��E65��������&����Da�S��SZu��5u@��9�?~X}-��B��$8���2����~{���,���b�8���<D<��i'!W0"�#=�_HA��/�'W�ݏ@��{8�ŋ2OwtI��ݽ)��f��T�)�u�#7�ƒ���'�>ݕOI]��o9:��xʗkt~iD���J���8�C�`b�θŤm�s�
�	|,�2f�6n���/3{��]����zX踔@'��vb[��L \��C��&O�>�ʃ�&Ӑ��fI�gO����y�MiG��D]\5�]=��h�qo���)()����;o6^e�'��W֙W���V��fV�]�(!$��$(�Kv�U�"LI�yB���r�6��6�$����=ڇC��QƬY�VX�>�C����qкF]���A�>������b�w�Ǫ3��h�ד����dr��o��1l�%��٥Ɯ2�**�=y��6`���vV�1�G/�(i�P�q_Lb��>��Z��ql��u�}��?Q
ߵ��?�B��<|s�^�$7�$<ݑ�ѷ���n�ӈ�pR惇�`�t�[z�fwG��� ��"k�)�9�v��e�סL�QQΝ���~㩑\�{[[�=�Ɔ�u�����EW�9S�9I�'���4��
�B�?���� �9��59[� �����I�z��9�����2?zw���
�j�$w8��`�]�E���`9�5i����ѨN�ˤem2t%uӀ�����`���\��4K~p�?\q���klR���?���L�,V�Mdr&�S�.�(<�dϩ�X|6ӥ�o��P�H�Ng��Н�N�ɕox**j5��P.jQ�0IJ�`� ��Z��D�k��'E�v9#lF��_)\Z���G�DIFa�S0��(b��X�Q � ��πx����l#�;R�vcc��2.��;�λ��?'>���jP�R|[�3[�'��-Z�-�(���NKo;JF^��GӮV<�>�[�٭0�[��]0�N=��8�cs)��*��גś�9�香��~6Y�=�3V�Դ�Ԣ��:��~A�v[�
ЀLM h�0�쯅3�2( �K���K5s%1��$�N-;�j�����g��q�,���q4�y��4c4&�|t�w'`��f��f^��'����E��q|�C�ػ^���ԉ��m%_Yv�Ǭ ��0n�~	�D2���233�&H��ֶ������BG�|J%��Q헑��4��c���W�q���ܴ�|Ե�� /q�g�o	��h������>��Y�[�/�+��j?�
l��V.}�P��8��;����/����}�4a	�/p��Q2�����1��Ty,Ƽ�r�~Z`3�"`)	��+���:�ӉI���P�f���~;���a����.��k������p�H����FL~����;\��,' ?���^: wy�A8��665�ml�-m�nnTu��s�M�!��P�re'�)����Ԭ�un�8Tp���?g3�0tt{wp{Q��t����ߢ��P|]c�`������������Z����SD�5�u��-��g�5%��%�~Y�"�s�Fz\C�)��{M�@E��rf�ޱ5s����2/;�(���Wlß�@k�E��x�ĄI�P�Ix3va��yZ��@-�X��>�9qC�`�'&Bn�d��۶�p1����Gn�����ck7��>��`(x�4`S<H~�[лQ3�[N������I����7���aT/�8�������Y�,7eh��Y��l\�$�>��^���yB�w�̘!ښ?�i_�s|�I��~%��0��JE��*�p0@��x��w��ӨWe@ؠM0���/���?����-|[�7ݍ���/?���3�%�SJVH�u�t�a{��V��X�$�'�l�VO�o�y�2��mA;>�\�H�IT�<������f��K|E���Г�~j�z6�r̄�������>?ó�ƅ6�(�pCӶ�8>Y+� + B`K�[kcj�$���ЭN6��M����&����Ra�x���@���E�ݮ�K���W8�ȯ��Y�L�'�#|��,��C�p����
�Ǔ�W�v]��\�׃��nfS[��,ޜ�6^�h�]�.����p6p6{���ߙ�����^��1���]o�B��h�nڭ�[����J!�����E�
ENLLs�2`2v2|n���Os��l�u{�##ջޘ2�Z��B�F������~�*�7�;�G�)X����s*��M�^8L�WLj4�Q[�G���X��bU���R[(�ğ.��c=�TWzy9��^�b�r�s�Ť��H��ӽ��sŷ쎱�������WW��-�������D,<�,<_���7��eҍ��i�+]�t�����['��sҐ��F�ILz(���m���h^b�� ���{��Y�`�E`�H�ܵOG���f�_�.�G�-�$��x~,�nq�0[�iihw*7�"F��6yG!�<+@�b�(�_jL�.V���`��IdL��*��^�����Pg� �D��D��׸�ВV��t���U'��Aly������A��eP��P�)C��~'��n7F�o�s[�V��|�S���������,���%�kv���R�q2S+���ڟY؟��ok6@Y�׋Or�Q�]����,�E�e��Ջ�����"?��M"�r
C�W�����M�V9�~u�ϭ�L�**��L�w3,��p9���;��'kxv�5��g{U!�"��pkI�m|Oy���B���Ȑm
%�Mn�����{``m�lJ�PܰqŌ��(��� ]Rq�����ec�/q��<)�Z>|����קN��bW�2Ti�P�ȶ


��;DǢ�Y��&;|;�&���k�/Ij8�06���5�m'j�������L6Fj��ȅ.����&EEeõ�:���n�B��"?�f�>�����b����`����v/����4���zX�̛��1�T������q�u��q�^�?0��v�_˦����V�S��X�©N��̱=�]���C4���F>�8�
�����5`M������ʶ��]�����#��;��������z���"�|aw���*��5�u������$�����I�Sڻ�軑{�����[�ۙAo��ۋ/C"���n�����_8A�������T<��f�֧8���Խ�J�ڕ�<�m�R����o��z��^4�z>a�a&F�������l�c�Ӷ_�����+e�#�-�x@N�H�n��t2X�'�^���� ���#؏�¿&���$�9a˳��7rDt?��4knF�`0!k��囐�|B��,XFa@b/��n~B��3�!{P���~�`|�:.���iT�<�A�D���b9PD�iBo=Q�r�*W�I��E�Ri���;f�O�(z��/H�6�`��8y�ˣ(ck6!kkx�d>j	¯��6����Ö��!`����k3�ΡB.�1/3C�N%5}���e��_�н�����5L,!�O����hP�_ ��UX��jP�A��	D�ld!a�X���[Jh�+J�6֭��¶d�����ֵ�����_|+k�J��f�"�^����Y}�(N�s��s`��J�V�#э�a���d!�a�2��u�W�Ɩ��o'�qֶ��Yl���}��V$e�0�����V`�d]J�ʍ����f�Z*�[0�~�e�B�e�uF�#��UL���ʳ��-,y�7�"��X#���d>���n�(Ú�����z��&���-^�a��;K��w{-�^�g��=���h���󇦄K|��*�2��n��o�#k�F|1-�*<��r��>�@��]�EE[�`=�n=[�lF�7VV�Ŵ��./?�o>G0~�������釰�/�_�!�QB)Rt�{���dѕ�Qd�s���X�|��{����x�Q�6â!+x����ȟU���uC��ή��BFN657J3UE�Rs�w��S��%񳞹�����5�lۏuE�,��m4��͖C�Ө*���79�6��r��y;^u�aٙ��TI�����t���,��]φӛ5����S!��2��"�n%��]&�5�l�N	8�l�z�����Slt;�J��iO-����Z�oħΌL�uX%�ZI�p>�hA�?��0�I�J��kzƌ@?�mH��`u�4����'
S�y���`'�[s.r��_L�SzM�K��i1��2�|�w�^��Ws����6��ڈ�������2oV��f�3��#������m�R?�D�=a��)�ѣߠ�UN���c7nR����@���M�E$W1�*���p���wM��a%,ݿ�qb���|Р�;W�.[�y2��wF)
\3�����	�ѹ1㹘~<
L*t�V��)!w�P߷fl�HPRce�?j��|��t凋��F����XzZ;ھq��"���].2(�H���Ad��/:����\T�=F����]���dM�^���s>�B�[Z����>����Ǥ�w*���L��ld�_�tz�֭/F�J	蜖%V���{� Лr�'@`P�ߝ�ϭ���3�R�{�����e�z�i��O&͡*���3�4R��H��>�e}Ie:v��"F��,<���R]2$>'4!��<��xr�}�JkD;��Ke�?��J������d��	kj�,��O��E�ҫ&9�O�_����Y�i��Y��O�}� �v������}���5�����c�2(O�1�n���M@��!{���$��)���nk$R
���G��Gnwv!*�Yㆧj�����$d(���yZ�෸gY�`vn֣im������@�P�F�?ŉ��y�a,W�0r�T7����@9��H�P�bR�Z��YVҒfU��˽ԉs��f���g�;�	�z�]Inz�-'�F�k:8��|��/�mZ.��r3I98*�����J��j�|�W�����ݛ�:���lj]>��Ϭ���'�q�������\��f�:	�Z3�T�F"T���6��t^�}+%���y�Y`��(ߚ��ʷU���m�0i�a��G)�B���xK"@xd��O&J�iK3��K��)��IFW[y���,�iyR�Ԓ������k3_���i��������XfdRֳb��W�)����ػ)�o���9�F;�[zI���|�V��Xd�[���W������$��s1R
�ьE'���>`\+%�C��?�t�E0S�^ӿ�0Z@˩c��CW��s�J�B�Wh�Q#����旎h�?���F���U�+\p�e�G�����H-y��z3b�h�����V6ac˩<�=�հ�2,n,���l�od��0B�Ĉ���FE�����%SD�+ⶊ�RDcH)��8���$�)D��*�d �cB��q
@�����o�
��?��	p��b��~ᒲ��~OHM�z���0T��(C
�W�v��g��F)�*��Xt���`�y�a��?qN��w��=��=��N�P�غ&��q�\/+�D�������:)i���S	;`Ewk��J��'���"A)��pD�ݖ^;��k�T�ަ������k��m�p�'1n�@��� l�	 �8�/J�E����
����*�(��ek ,{I��� �?�h���eh����v�����q�,/�Cx�O�f�m��/2K�F���$��Ж�?��A6l��ث6�>���`�f�
�����9���6��v�Ty?d������=m�(�e(D�C������]�[v�Ep1[䰽�3(6u�=�yfP�P����q7�t�ڿ����_y���L�o֦��d��ڙ�dr�i��������ݗj�N�?��T�q	����=��@�?��.��EN�\�ۅ����a_M��qXz4����ȼ+�Qũ!���o�s�(��SH���%��a�������l��~����3r�p��Q[1G�YRL��9u��Ef���s��[����3�+��p1+��O@vv��ޚX8bm��k�;L��X�;_n\���Bɵ�B����<%��)l-��V!R���&�H���Ʊl�'pL��y>�e�q*l�
h��i&�o·;C�C}�^�^��oߨ���֋�W�����}|�ț���IΉ$������U&��gF	�-5�P���Fl���{β�� �h'�)���0 ��r���A�xzl�H�Z�T��
H�+|�>;�7F����s� 6��q"�N����Z�i��UD⋈��n��Q���+t�f�b1�f�bM��w���R��iJ�)KT�
,��j��߄�����Ҹ��uw�ӷJ������8�5���G�'9��F��We&vǨ�^1��	K!��"�F!�z>a`5�Q�[@|�i�v��S���V��%��5��>E]�b9��!�;�Sͫ��'5�
��MDǚ�+���N؞�Oz��4mوZو"i	��%��������.����4�c��E۠y�mG�p�WO�p��Ȩ�e�_�,˒���%3�G�kp��:���v�����hK�e�;cx����&��Lc��|	|2d�e�ė��x2J���<��2[�Ҳ���/�;y�/2~�(PgIW��,0����Nf��`���! @�0��r����ھyI)���+���D��)i$��P�[��u��Q���X�Ae�Sb/竓�q��4�˓�$��ƀd����\YNFS9����	;���LQ�^J9�~T���"3\��qĲP�(�D�6��s��p��*DR��yS���_�h���y>�;	yʪ@�1#} ���[�#L6��0�ju�
�	�:����/J:�#�@��+�z_�Ў�T���D���}�_�Q?�tj�sW@s�fsq���Iqs��N�Z�`� Afh*�� .v:�k����j��k`���ԛs�M�d�ҟC6�kT��U��8^�N<5��9�:�7��;�b �Wt��=�H�h@~���ve��nK�.��~���ki�b�\���x�*��y��oR�`��sg(�V�9��mf���Qs�Ve�Ne�Fc�Vi�Fi�����&�$�T�����xC|۸�~Q����+Pvp����"�ri9���q��k��u��7�j@�t����b�<Dq<�ߐ����BOg��#����N���c8� ��g�e��h�/Ba�:�&"�@��j�)W!�����7_�dX����C�i8B�L�wd�D��i�[� �5wO�Q��8(�_?�i�xL�{,�=cE���3_K뗢Y\N[�8J���_����hʛ������v�/2���������`����b�H1�C"�p�2�+�|�kJמ�V������}��a2� =H�8`�L�%�wN��!��n�n{���%�[�'q��_�-�K[*KjY���C�̃᥃[n��7oؕ�]�dH-C9ҙ�E�4��^�3 �e'���-�tY P(����"u�t�J�V�hI���	�CՑ��H��IY񉹘�7��
��}�H�	DP�C�j���4��zV�g!�=g��M� :�1[CŁ:�N��$�
��gc�A걓4��o]}�C��9K��	��b��2(���cI�e'=M=)0Y�����,��?�P6�����Z�:fq��̞�0Į�Z�!�+�FD���� �����}zwܥnZ%i�y��.e���Dc�킦{�T�b/��Bǃ��Nc��i�[*9'X�~D�/DvP�]Ms��g���=�_�4������:��^�9�N�㘻.]�g*�;?�Z���\׻��\wwN\�ӹ����q@%�`Z�����߲Q������. �1��3$�g�Y��M�����Z!Q��Z_�E�2�''���M���{,��p�j�n�1�I�3Ȭp��#��;�l���]���=4k�	;f�
�A����O7��m]��s�T��%�)>��T�^�;��>V������Ō��d��¦Z����Ymv]�σJ:_�|�:n���~B�E\oc�c��5�5��Ġ�-��8��L���nů�v\r��/�C�;8
}�I�zg��%c����:8��(pr��%���+0�O�d�Ʃ��#�엱�VQ<�F���{�O|G棾mW�c�RO�AA�2�����uq&�@���딮?���O�:}2��vܜ�K�V��}?���-��}J.�C6�F����E��������Ӂ����ԁ��q2l��(�/h�h�_���u5Q9����S�I����+���&6m��u�`�W�"/�uܢ��^���[0�atE�P����t���|�������V �<a��W�g�p�n�0t	J��}?c^���E�
���e�{��^�:e[v~�����F9�e3������@	��������L {\f4�c�u�=mm
�IZ��2�xQRj���G�3�r���\��r�]Vv�6���\7.��532㔿���iI{k��Z��Q'��rU ���� ;:D���R�˔�7A�_>B��@J�"����/��r!�jޚ����1f蠙G<�d@�U����<1`���؀8�B��{CY��4
7�gWi��|�Z,f���Vj���~йY�K�/��<���z^#�Aj?�P>)�a���V-��WRO ��xvUd7�1V�U����h���ߢ�|�Q�:��b-�ϟmu<�40�z{pS���t�u��S��l���_����Lq��I���:�a�M��5��j�ꭣаp�0CϪ�Ʌ}~��ɽt������;�uN��"MC�%�َ��.o���9���{IN��ڏL�����`�EB"�C����1����"�?�G�A3P���!J�ۜ�p��D����f_�!�#�f��=��%�`���U�V#��'�2�4ݫ�}�f���ֳ>ܾ]n����Rg�X��жt���8�6��s8h�=x���~�
$
F/�#��aF���AFQϧ<u"��wU��NӀ2z��W��L(��љ�Q��\Kcw�w��C��:zE�C���D�,�TC�\� �I]��#�j�y��)J�coeX�#�F	��dy�����pc�0�1|`��
q@����I��z18J�����h�_�D����%��\���8y܈�9h,zz� �|�*���+]�^�c�_3y/O�
�tM��etkxz�G����K�qJ�v65�.&�9�
��;�T��`o'�hb	��p�����iC@�|���Z �2�UPJfr�j�{{�w[e�P �!1��j	��q�o���?��B��?nx�Lz��N��~��XZ�CUIK�ه�#G{��fg��% a�2�H��]�sF�]S������S���&]C��q����B������b�ٶ2�+��e���fg��U���q�����zǽz����Y�Ӎ[���xg�|��Q�"۴GO����Y�:��s�wh�yճ��Ւ<�
����l����1�>���f_e���9�8ʜʾ�	�o}�ߕ��1W���2�ƽٲ��^�IP���!���N���{�y�8��x�Q�;v���/��|�d�{0i0[,X�A��I�JШ�A�IP�Fp��a�VԨA̠�G��[C`L��K�BH�J�����IkX�~U\� �:��`�;� S�^S�f��n�8_�gB�,�J-�M��^�}���x�{Z��o
{� ����L���af�H	�d��5͇`�1B�0���a�&�B��vG"b^M�/U,ڥn@���5P�p�s*x�x��sj���c�@"���@�׏qM��J��!*j�K1�SVF[�%ꜧS� HQ�[I�)G�);��5����}��64,�5�2v���]jf��cl���G IT��1۴��$�*f��Sjg�E!�b�þ�=���uڦ�gp>%��ȱ>¼�4j�[�?����ΧujW��U�8��?�X��60�H�s'�/.�� P�|�$�9U�z����Pb��w�ȧ2XEE��g��+��w���%�$ƶ\%�xJ�I3�z,�
�"����!B�4��$є�]��U!Ɣ�tZA}KR���jE���8�%��^�J��f��!�'�/�7�C��U���ڸ9�q��x18��b�����X��
� 4�&�O��mbeC/��{q/S�h7ՊC���(QR}w�
��F>ǗH�}G٠V;4��B���խ��k������9��FxqĦ�+�(��;f��[���y���33�uǸ�=�O�q���� ���Ǔ��-Z����`��P-�	��Y�=ݝ	ֽ�z��iq�J!��	�j!��������C��c���ˑs�F�r�E�9�c�B�Q�e��{ր�Ȣ��"���jw*77=N�¹��,�����pfz�BDJ�l!��v?K�x����	cާq�/��Rk�K]؀��_�fl ����j�>2��R�b������O���(T�+R��.�ד
���@�'<x��RG>�Y�]����i�ȡ+U2�������o������0!a4���O���x��Fħ��')�N��ӭ8��v	��gFQ2����/9�mV�DY݂-���_�{��E�e�2c��|r��*R��e$)>H��~�.��Q7]D~�UH�G'H��D�si�����z���cF#���e��ɹl���� &!������1���}�U��˜"F.�IB:�3�����ғ�����TҋX�D�1?J"],eHeߕE��4K�RPD�>Rg�!e���mYm���Ց���x��jTW�JE��Z^NtR���st���s�&DJ�IЄOV��D�1�w�U(9�*1�Ŕ��3�"l#3�!Հy���$)9�Y�)f��(F�M@�~�5�`�4$����ѪN�u��p�	�h�-�0�d�e$�DQ�LXz�������޺8�X��G�׵b�v;M٩˳�y_h]0��3?�0N�w��I9v0lʢlI����)���v��������O�����������ᤑ����l�eO�ǘ��7��8��!�6���뮿�l�]��!?���!��Ft�OJ@��s�N�A��AЁ庘U�#��>W������6��:W�8ZY���@��m����2���-пI���t3W�ͩ����,����/ۓ��{�����M���|�|�t�e�� j㹹�q��qM{�p!�F����e=��`�����#���rk�D��{�w��⇸%��9m�yC�ࢁ��XU��y��o��l��z�\`��k�	��8�2��6�����5�!�[>����h)�Ȣ�c#R)2��@�̉�p�F8�M��Mc�ݣk% VB�_���}f�6�2T�6��vPàEm�L�Zx'��
��0����d{��9�a��ꟳ�ħ]!��"�*�<^K��,�fU
�pC���P�z�doq�MP�y3�%q�[��#��
�%����\rS�d¶O��r����h��j�v��Z��0��Z�Y� ��r�Q��F�Ą_w�~|��ۆ���d�O��[�d4�ҳ�I��e����قSz~�{����.b\0�\3�Ԏ�L�����LXC��RD��L��oT���%%�ӱ}���L1oGg������[)U �Hu�����_C?��MLL�x(�bͦ�zώ�GD�[�9��$�L��qf
]��$��8�B1iP$��O�Նx�I�T�W�]�@����0�[8a��韽���_ 1b�j���"��T���Jl��X`j�
8e���G��i����A�L�ls�9��,�2A{�����;��:���5]<!Ƶ2<�'F�).�A��΅BE	� ��T,@�-9�S�e�'�(U��A)®�6�z����reK�όX3R����fm��t�ܬ��~�|�2��/�z��Ty�E�����Mɗ��~-�����M�J;��vq�鉉�ղC
j�UIN\r�-�Y�~O�f��w��nl�o��=�n�+>��3qϭ���3,f�M�+'}W�k��K��:ȍm��P�c�'�ǈrCQ��u,��fC1�_P�s��-vB:r�`�zOY�c�Oִ:�h�ҝ�N�AW�|cG�
�u���2�i�vm��l�K��
����q�"̱��vԈ�>Ks8���tP ��b)��-�A�mxu(E?�bQ��Gi�Q��E2����G���p�et="�'���Aɯ��LW�q��>'`:��^�c�E��a*�H�󦈐�Q��bT�
a��J�ĽV�Tỳ+/��"CmW��GS�?�_�08q����XQ�K���t�	�)R��[���2�N���ww�*rە|�]��Ua-�]S��\b�"��l��}w��:˨6�����[p)���.�+���Xqww�@(n��P�!@��Eۢ��|����˚��Z�df���}��$���U�k�h��j�bY�����BaA �Gk�Ňo.(�C)�;��J*K� ��.I-ۦH�E}� R�*V�=��'/�.l�ª�5��@�!B�٨������«)���Q�����
�
��-T�h�m͟��JG�й��򤱅 '�p�]�/0h�%�%�Ȇ�D���g=��^ ܂G�����C�0��P�TV01�BTk������ȑqٙ	T�y����l}N��J������;�?>w���Y��s�������������`g��� ����ޮ�� �CA�g����m��}�������\��Ͷ���λ��?��R���X�ډZI�М����ɰ?����k���{T��؝���Vs+ࡅ�aF��xͷ��,�?bb˳[Z�=_�A������e޻�Xg�]Ӎ0����Z�3��ƫ��j���z�z��T��KVy�9E,\z���;����	9�n���a��G(A�1��_�[�$�ceS�зK[�4tP4��5�b�_Y��4/X��
(��e9(�6������U�x�j��A��{m����mR����4|��XL/��&�,!�MC���^L�ï�A �L׾���'�(�Ϧ
*, �6XͱE\����W¬�s�4��OX�U�8�=*�N߃�]&ez�1Q�dHM}U����b�ǏV�0e�\;�A����>u!�8�51�s�f	iH�'W�J���h
-��*��)r�����]Ԧ �@���X\�˥�ȫ���i�k� �t�Џ~R���pJ� ��ٖ/хЀ� j��%��gЖ�F��l9�̇U粁մ�T�=mJ��#��s,H��J��H�8��r|6k�w�Fj��������3g�.�#��'=���ёJ�z��E��M�18n�308h�g���"G�#G����t��VHZ4��B���C ƭE�
E�~n�oMP��i�¿��n;_'������������Ɵ����³��v�p�t���=K,�bf�j�Ǆse�=u�����E���>�Oi�x�����r��\C�/�c�����>��o�7���)(���*Ep�?I'$��T�˿�}�=���	����S��AboOt9wRau,�ZɎBUN]"g±۫HUFvN���ؘX2-\�F�r��C��vf|�t���Gԧ�:����Ric���!�E�T�VDr���m��ǿ��^�.>�Fܽ>��,�N�;�O�Ab7��>��$��
�$�F���ډ������7�Y�\
DnkI���x'_�%h�T��6; ����l!6�05C�uߧ�����q����7��Z�|;�I�9^PFNz���5I#[Z����'�+����í��l`�|���5��E^Mх���cޱ_�����%w�E,�����t�V�7J�\|^[�*%:���|[�H�}�x,}�~��Vo���a�cBs�|bW4�o]nV	����%�K���p5
��-����$e�M�#��<��'Y�@�%
9�<É �J��O)����n�;�)0ת"rgɑ����Y�C�@K6V"'#�-I��H����W�N��HJV9H�L�K�w9�e)W��`���ӯ��O'��gp>ؓ`$��=C�b����&�V��4���W�9���L  "� nY���!�SکaC [�����5��}~��\ ��w��D@��g�~���vG?8s���W�7����&A��H���(��:������ٹ��Lϟ� b�P-��(T$�c��`�Ό��N�y�b�EB��xĚ���mщ��4�L����n4����s����M�/?m.f�nz�ܾ��\>��|�38Ū2a�v?�R?=l�>mF�?^R�>mJ>|
z����Y�RIѵ���k�'~�z�w��!����_�����j�Tri����O	����f�����M�k���҃�R'ӕvۣ/ş�U��*,Ӽ�.<}u����9�a��ZC6����zu����e�"�й�Y������6L~BjY�a����2�A�����i�h���(EbT�lߞ=�7WfPQtd�� ���;ڡ��~J��ߊ^��S�N"�9��"������5�0���[�J;y�c���Aֽ*N�K�?�6�G��+jcK�|�m�'h�@���r
�ŀa��-�p%b���B	�~��r����� �|�J�{�9rC˿`b��'��}
P0��f�&8B� �}��Y���ZU���d��� ����݀(/(ȶ����%�By�QF�R�#w�3v���A�!yk}���������t�d�����M��Z�c���߻Q�����������~�21̪�~�a~�\� �������bZJ>cj/�Ĭq���8��v�p��e�g�p���o�ʣ�f����q��`i���C
�l��-�j�
�dӪ�bc2F�,v���甕�YYY_ cX���-3� j�#A��9_�ٿ���$b3���rrr

��á�_����W��x�DJ����������+&�9%:��Y�@�w����P�$�^"�.!MC�q	��p0�"j!+�*����X%;�4:�\�(4�u��a�y5�!�Y��<���� x��$ǏMP�� ��F�/��R^�2�ˠ�
���E�K+¥��>3,��>�e�63\���ʉ;ាY�j�o�(㣴�ݤÐ\,���wHD��s[-��K�X�=�5���,�՚ɯ���{�<�]�]��\�?/�>�>��m>Oܼ�<�8݅������6����E�	]M�>�k�s\�mއঌ�Ő�ߘ�5T#��AS q[��<���f3���#�k�Ƅh�
y�7�ȯ�����f���+��L��com�&��w���#�>����[�W���h�c v�^kpP��S��Tt��n�/s��*�@O��/!0��#6�oӋ�������|�/
"�)nɊ�u[��E M*�U����t�w�S�Ra�,g
�1;_����\<���)ϸ�7f�H���p���%7��܊}:��7'��a���@�+1K1AO��#����R�ҙ��l��{DM�%u	������Q�g$5���P%�^���]�2"� g���� ��6�8&
���MX��4=�"��8�J�ѭ��R��H��h#QS��SU��D��J�u��hu�����X ����?[<6vdqx
�%77��X~��p��$��E��u8����E�+���Ue_��hŲ�r��4�����3/�����j��hV�U9Ja�D��%��t�_��X2�b�y*h�*�?$��Z|1(Z�T/V}������]�7�ӒC�? ���R�>�����:�T���٣$	�C�Ơ�9�?�vY
��΀�jrJM�N����1.�㘮5��{�®톩���Q�PB�(/3Şo�}j�q�KG�8��wo�������˦D#VK�j�͘��5���m��~?
![�]^�u~\�nG��7�3"1�ϛ���3��OIϮ��L�G|�ZSk��-m���5��Ws?wy�b�͋�w��#�N��w�w��P��,����er������i����Fc���|��U��:?�.~|�����xO�U�{H��4�X�T
���+�ɧN������Fo���������ʼ��u�-�N�v'R��NZ)���':��4Ƅ�	�F3�<ʌd !1]vR4I�⹼�`��A*L����i���ב I�����N�lM�u�U'�ʹU��
Ѵ��[�z�v!k�@�'5�T �A�RW���w��|���	f Tv��%��]e[7"}Ѱ	�bU6����S��S�j �q'��q︶�����'u_K���o+T�2:@�mJ`95z�`���W/�6�f 5�Xpj�ذȮ���/0�N��Ѡ��V��ZZB2�12#=��8~����� ��i�h$W��bh.�|��;�!-&�Tq�D��j!�$d*E��0��G�����P(/�b.~��ɿ3��
s1����V��Ƨ�K�@����
��嫲�`f�2��{آfR�ɕ�m�I�.6�5X��bXbcU����2�xyy��t�Ȱ��4G��寣�������s �-,,vvw�M4�Ʒ�K��f�T*tXʋ�$���3��{x̂��]�����/��I�HI���k}��}����k����f�������J�9�a����8\�Y��ni�h4��A�@�N�0����U�}9 �,�'��/���#���\rm��R�P���A�i�P�рy܏��a���jH+qU{;��5��T>��{�v�ԭ@�?���tc�y�t�B���獿�g������{���w�}���|F< ��*3�?�ǻ j������I����a�4Dj%#Ü''"���Gr�E%*���e���=M��ܿ|ɚ�c�K��i�d��y(�1G.�=:)&�Y%u�Rg�ǸP-ג]t���7�̚��Z�^?��;֥�fhߒE��5�a{k R^�	kb��P���yx^1�(�b/�������8�ĩI68s�B����	p�y��99�`7Q��0L��V11�1,��##p�L%�-��fNE�S�Cl�7�����b�ڊ3 �>Af�Մ1���5���-��DP���+����*����l��+m�6>RX˂��x��$�r�� ]%�]���-.T<��d�t3�<:��.iy^2G6�?(f�J��d	�j�Q���~u�)�nVX�MN�q4e�LцYMdZټ���t8�����:�m���OLz�^��i�h�9�=�>5��#^�o;�h�\�o��/HFc�����g7��_�� ����3���۝F�bt��l��;��<��)�ݝ//����<8�&o�8G�t�^�w]�D��Ve_�E��-��J��t҄��ai0��P�ʖT��5e�2�G�>"�J�n�#���6�~��.$�[
��L(R�ΐ>����,R������c�2�^c��y0
�(��>��U'+����2�r�SI6��%0^T8-��!����1��G�Ã_N,��P7�����Ooq�Q��P�ȭ��?�G'����z��(�z�[sQU~-g��8��a�|��x�� ~/�cVu��{�$�D��D���w��w���7Vp�>>V���Ҹ\��>7��0鉋y��x�1]��tT��P�Eչ�}�@Ô��u�E6�����?�5�9?�|�'��ɟ{bm�����A��h����c�[���+y-5}O9�p��88iQ�2�C��&	�A2{8jd�!�|����>���������h+@�X��-bV�:���Z�-*^A�B���@����L��|N%#z�]��C�6��+A��8j��D�`E�0I��-�G��n� eQ���+,>.�Ӱ�ۭ����:�T\S%t��a�]�׼���¢>���i>�1���t�g�Q\2|";`�S�P@.i��T�B�����%�j.�K��s�<���Flf����_�)�a6�M� �8�̯M��>�i9���ܤ-8���>%g9��q^�̭��CO�cO'����/dR}��A"t��3g��6�F����G��Sk.�A���+�+���G63�������.+b���ˮ��6m^"�'��Β x�s]rQ���J^|%�TbK���7hvB
�f@R{����킖 C�8�!�Fbq���Y���=�����Flo?���S^E��<,�#�5bc�=�鱠]����,Y��җ�����n�c��
����&�|��Ŏ��-(9jw�W ������݃��1[�,��!,��&=�u����"]���y�P����i�C�L���M@@��oԊ#�@�q�1D�o�\�Wt�)R��D��`ii)�?�mnnnjjjy�4i�0F�aȌGB���靨ц��}=:87�1��1��1=�ĳ8�!��U�qi�&.�+v:p\��"���	�?�V�gh���A�|�E4'��f��<�?�����yY ��E]�_7���V�m���vȅ�D��'��r0�C:�/���m)����=G�1�_�4Xp��D�����C�D-y��%��Jd����9��Y�	�#8�0��}!�7WoY�����|B�d�Ğ���d�Ha��9���_�С�!�<��(��ǌq۟���jx�VW����Ȫ��0��Ӿ��4��è��_mM"V�7��K�,E�v�a*�@�Mڤ8RY�oM�z��??ߟ�~���i��RE�u��S*$d���&u�8[ɔ�d�qF��,�5oP�9O��I<G�0l�9�/��
M�����>��X�a���{gH���J��)Y��8�1
j��XP!p�9�}�,%'���&/$"�kO+^�f�&(sR��Ǆ�+#>sBa�<l�^we.%������5�v+�a|���+\_�/���r=�
�g�����|{�R_}��E[Eκ�KҨ��.[��g����b$UT������O�J��L�p
�R�P�M� ڭ?2_57A��X0f�i4t�SR�I����h%��^\�#�`�e���/I��G)ͥ�4�)\R�,���M�j���*�oӖ��P����VeZ��H4����x�k�I�����5���,M|�?��z��]@|�3����_��Y��r����ZMeBQ���<��7"�"i�&�4�q>�>FsY&�s���D	����W=&���>���X?�)s�./��]�H�#4���w��]���x���?P�&�<��13����R^��Z}=���n��,�+���ʒ8�����&Q�Z��ǶO��_<�a� ��	 dns�,#��&�ھ!/N�u�7(��8�6\�nP�r��K�C�bw��&�OEaG8l��F��p�XI x�mqhlC���#�o��R��8$Z.��,�v���B!:U�cw����#͑b`!�E������v*���,�z�}\*f���@$[=�����?����I�%3أw8Տ��h�`��K�ޱ�pKo��2	�B�*��1RK�D�Z��ƫsŏAtH�����2g&�ޖ�RHS����5���:���_[ �@cN:	������9���(�	x�m���%��ك�����y�����cx�@�x��z٫�%�W�����τ�����c3��4�=�D��=�J�ToW�\�=\l��ƶ_���5?Bbv/uf�M@��"d\����
7I7
6`�������!�֦KDkf��@łX'�H��8���>F�#�D�d��>�����q[���-}�q?���
��N��-ѫ��Ү_i�q�0{��`b"����4��r[�f�yw��A]tn	:
Δ�=���ճ�4.����/�Lq�|UX�1;�f�7H]j*�f�L*���"����@F��Hm`T9a����,\�B�v���H���ADǷϴ�R�$ݍ�+��жCdjI!wx`�����g_��e��/�VVv'��EP����Xj'��0}\�����	mKz'K���Lje0��z#�����5�����}��-Z�����ZD P��&����";��	�y�ep��f;Ϭ�U���v� W{��.��r{�Ϛ�,���5��������������
R���U�7s��F�su�s�b ��������~�Ӹ���!c�-��P���a�_�`��_'����U�mt?/�uV$�n�cw��/�m�c�����skl��a(��ߟ�Tx!��D�Id���Ref�IE��A��ԳH]���U��g�dD�ϙ�{YS\��kV^�Q�1^�R&��\x{��y�y��y�]�z{{X4��k�e��������1",>�B<
��X�TIH (����k++��¾>>777f<d���...���	�~Φ�H��ພv�Ѡ�n���:2��p)x�~�w��r���{��P��E82v�����������z����X'���c;�7r��n.�;�Ԥ��VȅC���,���C��>��V_Rp��oXT*�Q���|G��t�^���i�s܆���`RO�l���T�y@yM�k�}(�$7��E�g��Q~|cG�u��BŇF�f������ö(�b�F��ς�ߓ�.��>�ш�Oj>��?�x�<ݘ��*�`�;�1J��������L�%�Y����m'�j��n�eU���9�m3�ߜv��NN��=��m���a�
�ظ��-.�O�_�]�����u����m��g|G�2�n*;�8� �D	��W��V�P����!Dzl ��d�ä5v<,D9#���Q����Hq�ќqFE߇�@��Tȫ����4���"֓�4�	1�|�^�|�"oji��UC��2�ؾ����i���hs�������P>���:��J�)ޘ���F�-Z҅(��2�	'Ϡ��k*i�m,���+���*VH0��Ŀ]��֊9Kv�����oi�B��aA}��;��#	���I?�c�.��}�	FΕ�M����cg����>CI�J޹��G�|�;|���Wu�D���bW�ʭ���O�Z>!�i�cL�qSQtH�����kU}��bsi�-�_)�_vd���RT���:�PL���B�����h�E�O�[�[��J�x尘�����|�ź]��?�E�8#)�r���x�^�C)�W��6tVR4^�h�+��@1-�c��z¸ cvY��jm4C�e�:6\�.B�_]��[a�񷯽��hN��2x�x:W��	9�&?[��i�D���&��H�k��Qo���Siy��B�68̌���[��U�E#x<��|���M���"@- U;�-��l��D�Fk��	س��ANt"X���"�qG1�*o�kĳ �y3��}����]>���q�����G����3��l���<z�cx~8/�<W���Y/$4<�`.�6���~������I<�7��F��`��P��u��ᯭ�쐸���TB}'U)��F�`Rp���;�;jV�Hv=�j�
5��(*Ha�!!29��6�g\d4F���*�?��-Hs	J�rgFV^|#�Nfb�����
I+����J��H�-��`9�#X�X��O�����M�)N8�XT&4��Ԗ*���ܾ|��\�K�ɾ9Lݚ�J����*V��Q�׊P�!x�>i�N�MJY��n �T�vU���aJ=��54�p��{��ҝ���Iy�c��-7���4��#�B �*�9���A� ���l`,{�.֊��io�\M�Y���
�6_�ܦķr�V����:F1A&b��3y��tѹ���_FSI�WO�G�*��{~��Ӏ������'������e��� ���I��,�E�r�N�b�U��ӣ����Z��դ���F���2$����a�&6i8���Z0�����V��(f����\d�BN�u&.3}�-i�����6k�2��o�KH�E����|���t�m%��SS���FΖ��	Hғ[�P�m�j���bea @�_��K��X��E�ƵӔN`ޠCR�
f��4�DS�p��~��@�q��ڢ��k�9bbB|#�؈3T�y8��,�����0"�xx�jߢ����ȉ�v"��|[]]][�hoo���������|�Q�3j�=�'1qz:���o�x�\Y&��cU�eޅ��3��D���Ѱ�b�*(,�Nw���	�\7�C�����i��<7�����VX� �*^AP��4�������Y@z8�6=����Ն>�`��\����l��舄�1�T�����0S)~���~��Ԓ��R����C���B�"�6Ɇ��:q����3=�gN��%}wF^�G�EMޮ��U�NTB2�v���{o%֞{�fL�k����S�r�h"I�ľ���i������9|��Y��̅�Ij������֟���;nA�w#�KhE�'G4��e4O71����iQ5�%)⻋��	J4
*�#��;􏗋�2��n5�o�Y�.�g�g�_TU�#�� D�i?O�/���˵�B�\�OW�R�:;<`�L��-[�7���>E����\����0z���:V��BCO���SN�e��<�U��)8�tc�*�J�E�=KEۤ���(ᅯ�5�ߎ�Ӣ���ꑃD���u��H�����]�o��օ��=�N��7$�o'g>qhDDe��TZ�猪�9��b�P���,�_c���q�jrU����$"#*b;V=��e����dq��^�`EW"�����AY����<%2�ᥙ:CVZ8;f�>>`�DQ����<�4�9���H�������ݾ����x���Hx�T�>�$sQ����^�7�i<��r�.��I7���O�C�<څ���z����Xv'�PO~u@}be�qf�e��#S��@!Pm�J�]���t���!Vh��'E�0O;!�B>��6DPTZ]݁�Cev�}?��E�4������{��/��'8�b�6�9�:ޖ�F����=�����V���Ŵ�p�rg�)�Ļ�}������ٔ�k]�F2�-��d���Ӣ�m:C�d�[ɀBl 5�_ef�YAԔ!J<��n�6D���eB�d�/�0�s���c�j�+�}/V\+���[w��d�K�O�	����Vo�~l�*wW��eʰ1ɨFYT+����T���g?������~g�tnZ��$}�ޘ��w3�]�z>9=��m�W�?3RSo�$FI�$x��0��6[������(�������]g�X�OF��5��4�ZWY��RY,Y!�q)Vj��;O~�k��k�\�Vc�P~o��ʄ����Iߥ�⬝��DgG�Ң����EֳI�R���ʄB�b��v�2���s5�E?�f�C<�ʧ�˥,$�t��}�bfe����Zd?�f��{S���^G/�΍���
�Ƙ�oӍ;�;��O�! ��eۣ?�̰(���&�L�0������̬;k�7��V���kHUF���,���	^5�`�����7�6��g|^�93�?��l�S�)<��sC@�+�@��O��-YsB��Igz3�Y�?_�p(��jӤ���k?���w��<�C����$X��v��}��K������I	?�����cݹ�U���%���+��L_0y�P�׎f.��A�Gр
�t���Ҁ"3@�$��7�C�bf��Sb0r�Ģ�c��w�n�������̯�pb�O�YP�X˫�
-�ShOf4�_�K#�+O�NGx��^�k�L�>���0��$b4����B�:��iL{Os]���훨���]]]>/C���bc101���4�s�՘)�.o�B��S��,^Կnq�.��ٙ��armmm����W|Yss�O??����\�,��S�S����6��K��1Q�Q	�B"�tc#_¥�oN}��rv�R/�:[\��J��Ϸ����i��G��[c�ڰD�:C�@��/�B���3}O�P ۶�7��0���ھ͍��3p�q���E;� �>�=��1PB?��5�o���âB�r��vE��oxjexz㸸u�P�P�%hy�cg�ߓfQ�ѹ��]����^%���YW��:>�NH>���}掳��_�%���K` <ni�R�ס:�d����{���bH����������������_1jp���������o��IM��gK�����=
�-N��T����?��2j��-��"�G�
��+1Iz�0y�sd�/�#�ø���F�x�{d�n�+ݚ���I� [�3{�[�h�Ҫ�7H�u��s��ܼ�o�L�Ұ�&�MD�3~�*ʙ��I���싻��u?�u�P︰�OD�3G�!	�ىAm٘R�&���㻻$a��R~SnAK�?���M_n����k�-��uXo� VC�5�hP���Wx�|��{�pQq��P+�;@#����;��	�Cn��?0V�۱��Ȟ�Z���S�oP�~Ze5�Q0Dx< �S��ƅ�S�zb�0�lQp�C2c���x�2�e��Jnf�����b�x��D(��<0�p,
�+\|s"JM��	���7kT���t+�Ԇ.�%��Ѩv�ϼ�۷���4������l�D{5���Q����\��Ȟ7�y��ټy8��ujlҿ��Z"Ca���C�{�R�H�:��p�F��s]��Ur"�)i�{3��M��S�{!c*
HG�)�"��v�����f /��!Ј;��Xz��{8��W/S�M�0�ֲ�,�h��RJWg|m�>�a\��vRӱL9��H_���`�J6N/���f|�����75O\nG�ܸ����fHE�G��P����41�ޗ��-���9�#�|eJ��o��L�<����m�^+W��x5�b�?��[t��N�n(�e��s�im��9>3{����8W\�OL�׻Z�դE�E�HRƖ�í[�I�|@�i��n�j�Ϳ.ݸ��(����B��ꌫಊ���Fr�3�VU�h5��`c�`')ҡ���N����;�&zaniߘc���eUKZ�R�%�1h�X��˰�Ő��e�e�nd����)o�n��}=0etp�r�{7�����ό��^������Ϡ�6�Z��B	�CS1��5�����б�h5P83s���A������m��hW�d|�i>$�j{��m�E{��7�t⩙��SI��9��5��x(�TZT��y���]R1\�u�C��m�w	�C�����-*�MZ����3�$��{�Q F�=�
E�K�?U5�-w�&o�M�؟��?�Ae�?P����~��r�0��r������A<o���Q&>�G}TW�����"��~�����l��w�Qf�����JeTe�ÑO���s����L4�8�ս��֐�֞���"j�z�����r���:���vo9�8j,Sg��S��+e�;%{�3��W/�<��.�Bo�A�)��f�D@,��q�qV���`���t�B1�u��śB���C�7�y����Q��}Vbec>���;?�N��4u�������J�BYDd������\p�S�OAT��#�l}�����>)�n�LFF�c[Y���`���u���74��a�������~D��7W�ֶ��37j퀀��bR_��0�z�Fa;u�s p��XE� Pa�E�"���
C'�WI�����^ޡ���ز��+\J��Q)i�C,�+���n.���m\�i\�g��d`w{�6���	v0��R���!�oܸ�G��^�����񅡜���t~kw�B���>�����d��f��L��t����#����r/E*�g�X\����3�5W4έ�
g�_2m�o����+�����cr]7���ε�F��(\�� ���B-�Q�it
��Y��-.NnLuue��?��j�  ���U/�b����VG����=�#��s<`��c��-�#������C�U����]�LV������S��\�x�d�T:�َ,�Ƚ�z�Qa�	���luq�51��V*�4!P#@�F�Wi�5K�8\B��ݟ��9N��U�OZ�W<�����g�2lꒆ|o[��y5���R���������a!/0{(Z��8��ȏ��3�ȍ�b�7��SS�P�r]	]*2��?{q_<r����q�"�I6�[�c!����t3�T�z��!�;����j�t���d��q��
�f;�<jy��W��d�;�:�,J�`��W�
�&���o�tv�b�Td�)i8�/xB8L���U_�X��7�⮾��ІO�K�����")�-_�1�͚� ��2%��4�&��d01�� ��h�����P!ҥ��(�T��1�V�e#��Ճ*�6���v��?��0dl�_w�հ�mD����a���1x���[���t.��ŵwq~���XD�s/P��30�<f,��2����I�<[j�ɞ��G �
�*D2}�!T�6Du�?�Ȁa_�����#|�[��?���
6��c�m77޹կ��U?JkV�� ��sX�i�ԓ����W�~D�϶7�o���+�vh�x�ҒnJ�z�>�����Vt6�u�O�K�,~n)/`6bK��F�:����< V�io�ہ��Q�Lډ���P�"_�F�7�<�)Ɯ*,Y��cة�l�m��+�g��z ˆ�u(���FE)���âǬQ���k:���Ⲿs}:�w��1�M��ISe�x|C~׵ֳ~��yN���vy����)��}�BWWr66�9GC����>S��=?��<�5?_��<�%}�7>�7�n�����y:�f����}5��RW�����d�	���0�.h�tq�`~���+!� ""����ܱ��QU���w��g�.�pI��8Z[E����7m�*��xi�}�|�%ů����j�Q$�O�>�>��l�F� ,r�:,���7������� �����ShNQ�w�����^�n��'�4�&��?�W�_�p!t$���1�\��̚�	_,�9c�U� �1	���MOx������x���ȇ���nAӏ�.A�s�L`~�T~��/<f�*&���ܲ����?�GQ�*���]�*��*������ ៜr�����*�r&�ZRC=ќ�z�^#�)�'^Жp��s��1�+���_�2������Ǜw�Vs�Hg�2L�,?������S�B�sP��'�Q]�tq�r���J`���:tI���OOd.����))��д)�SRR"!!����g��1�1����W(H,vpȑ!ml����nK�o�'�C���U7:�2��qL������
��/g�0�F��j	�xU�#T.�1pͯY���;�$)%/@��νCac�+����T>�94;��������w���@͒$�t��#�B��|��0�=|c��]��J�� (�uhL�H�#�o��)���6�:9�AN�!FB1\���i�+���[�?����:[쥢s��v&vX���8ڊн�	�0>^��z]{E��C"M�飇�_�Ws:�ב> �Oq��ȅp���k)W�QliN���qi6����6�������n�|��k=�"�y@���XD��=�wY�1�þ���5�!@ fR�	��YrH}���@�{U�a1��#����*��G�-rl�-ZI=����B�	F�;l�h������:,oS���/d��+F�x������0�_��<��Z5F��;A��״��WEo-�R��I�_��"p__�`�|?��J��*��\��
�� ��xNO~�Y��K��<�a5%�xat�I�Ǫ�'���_�!�=7K�������%d�{���|�&-oHW���^�6��V�c�+e���(��`MK>��bE��ܦ�q7޺��Uņ�����??� �魶Z�g8
��LK�U�8�lO�Cʿ���ѳ�����ٜ����լ����w�&@�
6��;��_�B&�oө�Tu�@:�oU��S�Kcw�|��Ä>`,%�z��%����#��n�4�٥����kS!��n1���W���<G��,,��C�KG*�z�:ut�O%!Ĥ�6W���}֍�
��`��7,���E)��2�Q�&$kl����-lI
�쭞�D
F^�.D.�`�����(Ά�*��Og��%@��}5J���4��,��^���hl��"�{�Q/�Y$⏼�Gu��Dd�t&�*�df�մ
����;"�r��pG�{V�P����C�?sc�rU :
�o�G|�ߛZ����)+�g�h��hu��δ��(l(M�?\����p;yQ�t~E�|u���{[�������x�%g�ۃ��>-�&W�*�Q��_����s���"���j�֟̅������\���$�J�F�W�4>*ח���Բq�j�צ�GĄU\���eMb�_Y��ny�
 �hN�?���2����f �����nz��v���s�b~�Tי���;�#��������+���f���Yй�l�����`��Š���B��A��ӌ`�}\��$� �.��ݳ��׻�W�F$>\/]Y~�츾"�4�ȡf/ ?�����1�@
c#^�3��QGbgL� ���B�Eǎ�Q�SC$eػ�s�����@ /&�	��d�}��	�\P��v��Q ��.���B�ģ��'��N��*%#���pW�s�Z}�%���仼\`܊���q/��� ��ʢ σA\�޿��.��U+�r�z��K��H~�.�ewId6�fv���������]�0(G�OH�#dvҚ3������`��/gO�DvXt^[�ɞ��1+ ���o,,�]�� ���E��E�baN��������VQm�m�5Z܊�/�b�Z�8w��R��/R$�R\[��]��S������OwN2r���J�u�k>��.����d��Pt���F�' �ɋ"D?���B3�����2h�S��Y�ч�}s��O��OL�0���	%�R��LС���wyd���R=v���W�����������S�U		�v!�BU��)'E썎�R"yv�	@���
��P��SRR��̧��$ƴ�eRNb�X��ٞ�8�8y�7�y	���oz�k4R�B�{Ɂ@U��������k���~�����ލ�M�	�0u�#��7<z^n`dr���4RL�ʳm*�%~W�
m`5�;.���k}���ep/Y���j �l�:®Tȧ��[�nI���XV�����C��=	�u)$��c2�=�Q�U��L�ɲ.�NO(�\�!���!�h!�m�g�u|�v���
əE�)$`�@�H���j�}u����uW��}��_̳���[�G+�b������x���xgU�c��w�	�"��^�~�HV%Q|��}.Uzp���@�E:qI�s��C�����ӯC�<�}��؆M����?��h.]#�������H����.��f�vH� ����`΀�;�$�zM=�Xw�Xl�A&��zWC�Q��;˞eb�7�S�^��R9\"�� ��NDU�ݑ�݂��d���k��: �GDG����C�+۶�5�[CZ5���� �z#�W��}��ndD�e9�����)M!;�{��k�!�S�ItT;�[a
d	����ym��x�sҼ��_�~��YBi�CE��Xv)P��P��]�3�Ğ�6��_y*��p��ĳb�.�k���8�1�,��nJ����#6�#6�R��F��Uꛃ*~��{N�����	�/�ˏx��H0���1�� �� 
�P�]%Ғ��̯lʞ��5��#��Q*U-@9�����gw5k���s�'x�Td��rɄ�E�\7�_�[}M!^�!=.�S!�� ��.k�ϵY��S�3�T��Gr�Qk���D�JO�̓�������Z߹
����G�0�~h3#�Y���!���n�X�2#�1��=<��Z���?BU����r�-�tsEF,tn��x"���ϰ_��KW�R����Y�A�6P�6����D��ԑ��]45��=�5��׻���Y�|��æ�9���/��ZP�l:�9K�6��Z2y�I��y����d�����D�CTO[laVdo�`{�X��J�C���W6$�^��e�GȞvx���xX�7xaU�u��Ŝ5�M��幱F &���;�@�퇄���g:hJ��!Y}@C�;�W�H�� ܅�3���u�w��^��KU�bQ$I�PL��8��Th��w���Ϥ+�+�͋��c��MoY���J����rEۤ�淳I���9��+y���Ko�o�-`�%�+����'�K�PᐌW�}�g��E�ݑ�
���]�Vy��*F
��cm�0����u~_��ʥC������^l���if&�X�9����m�/r[�,}=p������Η�D��@���\8<�h&�k -��<��EFY!&_�j���E}D�x݈�ҩ���__e0�L�nă���0�T,1�=���'eӌI��Q�G!a�B�J�7dܵ��=Ϟ��v.���Fé}��.{8�x],��Li
�q��y0+ߐ$��))�g�(ۊ��0Q�+�>��tA����Tٖ�o��#;�����'.Z�jV��� �"��o�$��A��?+��jwO<�m׏y����`;�-�x�����~0�b����O�� ��� dK_�㕍�,�c�'��T3G-g��aå�^���,/I֡ �.����Ǔ�����1�ֲ��.V��F(�(Q����ן����F��Ʀ?^4�\�J��(yj�op��"�GcƩ�$Q���ƚ�4��U����O			v�������偁��d�����4	�+T�{�f�VV�����N�U_��Ϝkq�<p�At�$�\���,A`��Ř�� �y�	�	��F�P�ŭ�B�X@������@�SC'-̒\���G<(�4�b\S��ǻ��.�b���i�>������3�C��MKϭ�6�3y��V/�����)a$�����q#�I ���jw�&��ڒ���{\9�+��F����δ�x�Dˀ���jga7�ۗ8�ъ�Zs���#�	�
���^�`S�2�ُΆ~
�f'�!��U�9����G��_�՞����?%}7���Nо�h�<F)t۝�,Z��yu�,&T{�w��ԍ9f�����bp�4�^8! 9ս�����I4�c�:U0�z���b&gm�R� �c��C���E}Q���A��	��a��\6r�HO��5�#.\D zOc�O�,��RKꖳ�͑�FN<��Y�2���o�&�CL�@H��Iŧ����������k���F���m�"%i��ke�[o�����݉�3m��#���)0��ɽ�!�z��軩����漶��W^+7��+D#��X0���K$�|��wOp�\Y���+��L$���FV=ք�}*�hmU���ik0HvS���4/�t.�<���jF��R�Z�c�����RM�oi�j���"=�|�������Dqi`<��ba�3�󈼀i�[�(q�G���?e5q�H��w�j#�|��\v		W��p�[��_����k;[��4pf�8��f�h��������:k<�}$��Wе������g�W�(��|y-g�Q�U
���/�r-ŜR$C��B�*������8�5 k�n��D���������˛������2>	�[ �~a���}�G3����L�V�%� ��O�Z��xn�?*H[ꁃө}9�F������7��v���3 ���)���Ѿp�wZ��"VO�Z��,CM	f醧�7��p����$߂j����E�x�xe$��b8"���ڌ��"~�n_��AOݺX�"ѧEE��Z9�*Y��jh��xtoT�.߻�IC3I�	ƥ��� �PYZO�9�W��u�>d�N(gy�éA7G8Y�������O#�O�:��<:��(��=�s��D�����z �h����sl~��/��1�:�Zk ��IQ���P��������3`{+l�eա��Ty��������u����6㲪�m�]�_�]c�Af��r��kV���=�$�������u�7�5�Lف}��e����x<�����i�L~n��ք����jM�g�M�S������!b���;��^�"e�?�w��<K���Z/��bM�'m/�8��F/�mY%mOc3���?�m�RF�2@��W.sQcc��}Z�Ė�\��߮��K��83�A��/��\����3��+�?�Kw�5ECh� MC�l�jf]�h�\�?�+F%y#7Hu��L�؊i�*(�q�ξ��a��+I�H|L<�#���x*x�3i_ki98n!hi|a<(���(���(�܎l%_[��y��sB�H��&�-�=���dcA3>m�.Ëbf�8����c5�O5͋v9ﶮ���,H(
�1�Kf�P|�0�����3u@Ki��
]���'y�� �Ƞ�H�O�Q���>!�o㙽;���wv�ZE6"i�h�d�T+w3�]�֕
=k��2l��O�ƽ��Y�)�h�b𿅚Zm�������[�_�x,�B�a����u�I=��W>_3��y���~�ޖLp��~J�fJԔ��apz�W����(B�@�ⲯ����#`s�یmK<mN5"�ao����/M�OZ���q5u�S���!k���	fAD����;Mv,J-��ޛ-��rܸ�}?�0z�Bd���Q���X�����0ե�Z�CL��pl�r�z
�]�uA;��M�������u�~�(nG�������ś�é̂�z�~g'ā�c��*j8>M��i|����X�Q��[�5��8���lB�`���*|ȲzO�,X�"M��X=�D��P�%^V��;<�b�i���f��}H�m�qq�tv����<^G���|�c�|����Y��Gر	�������$��>�&\/y�^o=-�rP�k���CALƂ}�ю�~>�C�c��eí���0����@������)�N.��#��v���T�p�<e�`���>������>\}*�*;�~�5~�J���;�d5�g�=�Hkf��\и�~�M���`�;|��DY�\���Y��6E��G�A����s����jt�Q���_�j�%r�{4�0��B��?�D��9��G��nl�/�0��tD��7��w���[4�p�
s8k�]6&���s��}~����Y�P�l^�,��S�U������Ɲ�����o�ڭ���&c��bEۼ۝��U
�S83�Q�c���g�O��0�q�N����*Ǡ�l@�	���^_E'*,+�5�ᣏ�@5_w3����9{o�ޡ������g�V���J#�s[L����w�#�nV"hO�A6�^E0��B%��;�d�����H�i/T�9����/y�r�1�h16R�gR��Z�
�5���p>I������&I ������ܙ�əu�t�Y���2n�,�ab���ዀz
h1�{%�w&Ml&c��g�I���tΆ�D��x2%�.�\A���s��\�յ��	��1�������ՆE���x����.���Js-.�wKv:���4JX�օ��4�
�R��H>�̹�S-�U���kX�tiذ̼�~w�o|�]�XmsLZp��Ed�#�A����y�@0��-���;�հ�m{��.�8�z��p0ZF3"��Ƃ�Kx+<v�h�����c��1	��Mj8@�F��ݮ��{����״�n��8�|�G�y����Me\�=����Eќ�?�E�ʔ9�����"Cp'�F�?$8�� �d@x`����;/gKV#�7������(E�E��"�ԇH�=/��%'�y"�ID�x��hA3����K4.��5v����;��+ʜ�a7 ��.�4䣌�͙9�[�ʜ �bt��Ѯ��-3��Ƨ�z����g����v��z��LGm>���Z���"���I�H�L���Wz1�����{�[��O/�#AF�(`J�$F�Bn����U�ƫ�3��}/[N��K䷔c�<2��WTx���B �i7�' ��P喚((��� �>j�*�KP4h.�3��iut�9B���q�WTվ�	B_S~�e�̳GLf������Ǚ#�Rܻ-e���T����9���ى"�+ʧA����T���=�hy�X�}�r�����v���y�����(�Z��6|��7"j;g�F)a2f"0򻨻1�8����~{
�}�o���9�j�*fϪ	WN��b��4H��G0���$�]Sԯ:n�����h9� /
ּ�w�W�Ҍ]�_��{�o�����E�Yh�����L ��@0�A�����C�5rΔ``���oہ}�R�~�\���ld��@N�1����0*�K�ѓ�a�g�\����[ps:�2�&��JN�H)KW6[�匸�i����i�������t��qjl�n��4з��a5�Y��g�t���J�x79RMP4���Kл�~8�/��X6��x�^�!�w���"Sδ�6�>��f��eYS:��VP�_IؼM a�~��Qj���=�Wz.���S�8^�$�(��\U4�·� eb0�*�鷗ߩ+�'����pi.���`��T�×��}�� (��o�ng��Q7I�s��C�-�J�O� {D�v">��w��7W��R8*48�2[;�����[���«�	;7u����`���b�̰{��tU%Uy�~W��@�!�8l�O\�!� �����������|������%	�.�M0�-��T�b?и)��Q����TT��I��F-/�+R@�c"��OrP�[T��pE�e")�$I�d��ؔb�A3&6S��T��׷�W�U�۳Ƃ�Mu�Yu�	�m7�e7��%��G��N�������N��G㹣q�jMOq$3�������p���*{���܊3�D�~�۷:�ҡ7�#gg�f���/�#jʘI����y�p����-�bL�m]�ub�jŵ]�J��Z��1�t���Bz�B�-G+Ȏm��P�6�q+���ŞB��>�!K|�FrL]��ӽXU�!�3?����L|D�6�S�1���
�3��D�' t6)�͆ {��r;���D���yxrr��~i�l��#�ҏ����a�a�63���)T�*e�tbo�1��l��_�9k49r�	�� ��� �TS�}���=4ob4������3�%����{C��z�ݴ�����w�-e}��f*`�p;��r�{L���mPZ������]v������5�p���wy��)X�hl�:�
l٤'S��_s�ch����$C����mG�� �7�z{�������E���q�~�FyD�iO&*rR:��Vnk��ԣR���ݲ� ��a���Ѩ{���x�#�o��6�ު$O ��?�ʉED��s?�\?�~>9�i8���7�ul���!�K�*|}1��w&h�x8����Э���s6��K���t:2�|���p��f[Q��|w��8�#��w~"���᣾����L�f]Q�]i��M��e�b��9�$� ��{���p�H���]�VqF��r���a��{��[5`=;:��X�n�{�_���5��[���^��,$!�q�v�&.�-����?�9�U��T��g�3�\'�&Vw��ٜ���	��������	h�7�H����+�o��"�݆�μf}�[m'�j�p�G�xj�������yq��H�2s�}P�S>Z����]s�v�T��C�AXD����0�a�[޿��2���eY���e?���"��i���j���y��"���ucv��>����d(1S�����eAj����,���=��n^�3Fnc�.ky��7KU!���,�^qD�bِT(�)=�� ���vJ�sǥ,NB�3���_�c�#]��fd�.Pi��P���� Zȇ#	�����	�~p�8~O�:��3��8���V����e�����X�i�N�~t,�PG(��r��8S�cm�x<U% ix�c�
4H2]
)a
Ԅ�&�%���!j&U4�*�x*_Xc%U���ၵ挌_䢉M����+�|���uF�g�[��^�?���I�`�����2j�e;����42Oԋ��Rn~���O�
���]@�z���s`�9W�L1�VZo4��>�6��M����-���'�D��TT?H�(��F���Rmi%
z��	��O���� ��������RH#6��j%Esi��<R��T��O�>l�iP{��X�`6��]������m)�j�=A�L��;��-"���gM4�S���-b>Dx|b+�9~��ykAD�X��py��d<F��1nr#�w�Z���] _��Ϳq��۾�Z�|�4����צ`�=�f�NL0#��J�9I���8_��r?�pr�8l	����1?��_�X]��꘹�M����?�h6���n����,FT��`́�0~���W��d��j�k�qQ�cs;��l߻O��i~��r��hc�L�L5��~8�ΨѪ��>u��`���F��2���sr��m��xS�6���x;��)�6�޼<��{�_�Yp�w���#|3����Լ�C^X4��%������ᢐ9��BX��\{}!q-���v"h�܂YY�b�����<��!��׉�0����w ��9��R����)dpl6�7I��g|� d��{�0I������:һだXB�y��o^���/V�� �7֏��`u5�W���)#��w	�!̣�͵[7NF@@��?9A��t��!�0�Se�����L؅ק��^�^J¥��!�<��S�r;�Cy {;���t(^i����݅`d��~m��"�o�/�&B�&����-�%ӉI�S�*?�%����K�L�vmؘL�O��λ᩹u�Q�Q�ߠj�*�a6e:����1�����`^�彋_U�EMe���j*'�($�(��SҲ��UW�^�V.�Q:�dR�7W�}��5Y�jV�
8��AE������!;0|dS9�j�}�k��3�8�[����:՗�W��O\Ó���j���+���ǟE�Ib��7%�� ;���y��Z���R�I0~�7�<ӛB�bi��ǌp(�AtSL,f'9u���D�?�
CC�_��ɄK?R��
��&*����y�?��=�����7
�tg6
oә�����ǿ�D;����a�㓦��*����������.y�N�����,�����g^��G�4��!A��A����Ȍ�oc�/������ê-���Y1kɠ0ۢ�w]D�<����^�@&{V\N�"_u���1��F�d*(���LB�Ks39	����Q��Ĵ�Pb��1(k����%�eX�a��V��8¶d�z*��x>��oPX߾�����'	RԬ:�{����T������@�����SsH+��mSP�'�?��u:F�w�����o��:��2`V��!;�6���;�O1P�$�?x���-�e�nc�T�-�������{5�P�F��1U�,f����t����攷#_��Tz�Ƕ;�f	�Xf�����a�G���-�o������#��os�sK��[&���W��*=۪��JJ��^Jt*ӵ�*�C~�{J(��%��6��7L^�0(5e@�����Lk�5Ę�j�o�_�\�L	����C�z���Bd��
X[��d�ºy$?�~��m����20!E�B���>5^l)��KJH�h��l��6�\}]:vx�������:̥��۶}`�=�R���#��d��W6�z����^�x�#�j�3>����{�8p]��Sz�����>Yi[�ݴ"����:���bY���5�$eF�£-�#!��M�F��!���������P7ڏ�\ʛ�#mM��.����?�m�y�0�粑	|�\�w"#ϳ��"rb�P+^.�HJ���z&�c��L ��T�-����<VY�"�+��=K��fG��P��
q��"K�aEڊ���[��H �
�#��ygYSK}�*������� B�/Y��w/���,��toB�o7dվ6����� ��4�T�\��6*�}�E1$�Eg���UIj����*Rj�5��C�,D��NgF�TYF�<�`�&�0!k�����R*�\Cdi�{��yD� �<C �∦r V=�������d{�<{�����<� D����i�d��Se�0lM�w���;� oB��BM��*�ٞ �f�X,v���!=�'�J���A�����7�@_H�`mF��H��N��M$��%�����ӭ6��H����Iɓ�ͩ����lP�ပGp'oӍH�틫76���4'����l�̏��D.��-C��e�ƻ=�!���,Qm����>[�\R���0�g��ytf��76���ŏ�������T��TYYT��'��Yh�K׋�5 ��E����E������7�j��A�D4Z	�]���s����K#"I"�I�EZ������no'�������|_�Xa-8e*�HA��ױ�m������U"�Ͽ{��!�_������"�Ƕ�o�Cc��eXE��mp���#v����ՒV���Bh�+��{�����Ԇ*���hD~��P�|��P(F�+/K�q(}���LT�w6=�[�j�J��X@��Z�'��"Bs$��s!"����$�ԃ:�SK(������*3�{�����?���i��ɜ~nHȵ;s�Y�Ai��C�����,;	R�a0E����K�Ӡ�{/�Q2i�h@�Lb~d��T{�XM��7�cI�]�z���Z�����;1�!��@G�dW����yHEa8g!�qG$I�-�K�dHX��̦vf�+��u��3V��T7�����'`Y��^���K�W�Y��K	ax�Yq��	ˆ`�+��"Q8��Z��m����8��)eі�g����2[�r���{"m�+�>b�f|�f^�l�i�֫{���ujV*��	_������'�(x��נj�f�7V�b���G�&z:;A�S�Xt��)t���c3��R��������$58�]$ S1&��Fz�d��� �5$"������,��5D`����+���Y/��(Vi���ʏ7!k���o���U<�I�)"�
�J^_����j�bJ��E�Vz;v*�GL��ؔû��m��3C�(�\�̼�@���j�����7�Xd*`�/�wig��������:�P!۳n��q��h$Q�C�>�p	Gb������5�0�$�%����#���M�4���C���M���܈�pA�j���<�!X�2\;���K(�X\0�s2����mQt-�FV���I)�jo`ū<�	4���<��t�v��>�TE��A	����k���c8m����Ӗ����߫�~ގ3��5�3�R�*N�1%�\�ww��\�K��W�s\YlM>U1s+~%/���V���=e�vpoq��!&�0*k������aF�:��&#3�L�����������(��S���Gѐ�.�O�3�}1��@��UqE�I3�+�y���g�)������_V��ҋU4����d�C�A�ӡ
R�;%d	R�gK�o Io�鄧��)n�,��k�[��o���_��q�6m�J�7J7o:��7��O2s�~Ͻ��'=z5m~�'7�/�۫~���q)��m�Wh57�롫�/���h\
���tw+d�,��0�J��$'n�����p�"QZ		~ֽW�͐��3\�*9N�+��xSF���u0�TB�aD�.g����֜J���g� �do��%�g�s���DT��5|�����vv�8N�^�c,̒}�-,SM�i��v��dJ"�}��������v'�JtY��܏|�֥l%��)�G�#$I�{��+|��l�d�9)f���V*w0���|��Ĭl
��X�았��r���vIp��y-P9�����e3�x��88�#o��wx��oT��*S�w*9��JV�����^���2����#el���j�q�W��I��mĘt����$��%������?�)o�0���u�E�z�qȆ�uf:�{#*�*��iR��0���cߗ*�04,��}���q�����?�6e�Y޸��,�ؾd-�����v=\S��×���ƎW[��f�9�֍����{Y��|����,�ӌ+ɯs��|��I�` I�ޯ�*KR� ��N�ߴvy�h��o��v��8];Z_���>8�<9�^?�9�^۳�8t韽��L�	�8yB�;��BCh7	���3������p�K�w�_B7j�uֆ\��;�[(��g��k��\���i�a�)3fd�l�\����ی�����N&x�����S�/O��+M7-�\��Z����/绛�+_�Nm���Og�b}��n3�dN}/F����^g��C)r�Y�^|7��{�ٳ���CxIK�+�����/i��+g�9t�J�~�q&]�FՉ_M�K4+�M/Mp�]�r�e���H�����ʀz�X9��j�RqS�t�OɨG2�嗸�	�3�;�+"u �jL=�P�y�\f�'i �D����#C��B��p73��c���>L'�{��'��ȇ3fI�=��ư�?:�����d�hd����RR����܏
֔�_���J�g�{�R��r|�ru}���j�u���P��a���Z��F�Z\LƏ�2��ISm�٭��S�Ρ�ɦ��"Oб1ߧ��į��a��#���-��ɱ�I��`�i�ə��՜�7��W�U4��׈�ω[`��JX���+qU�Jo��s�yv����z��K��� �;��=�eX�p��Ƴ����Lz��*��őg"[��À9m0�&zR�F� #m���;����R����Re	�E����+ ���%�v�UA����	e!D��.73��^i/0O�R/���D��|S��o�I�E[�u��z9��yD6�SA*��������tH�4���Pf#��?�
���"�k��9δ�ę{G���hy��$���t���1Xo���t��Bd�0>jgi�K%�^������R������+xq���whWk����Ġb���Js��|��M��f�#1�����y�PO���oǅ�sIm�5��Z�+�5�O��V�Kn�7�RtW=[nZ<�^1wQ���Vs�;�SS_���q{��BӠI��ٮgl����kx;[S)�o$v&������\!0��I�2�ZI1�2��}���ͣ'7Щ��Hĸ�>��ݬw:���/�B��˂g�i��=��{�f$����ოd<[�d�r�a���$q��ݟ��Ip��<�zG�66O-7�+qv����
|Ը��X�~�\6{���ߘ7jݷ�5^?(�=��W�Aﶗ�ۚ�nǌ�n���G����*�䈻��n�T���喒�H�v%��vFhKz.%����X���(�L��I����ϤI�Dߝ���A<z��}�'�Gzk��g���
v��<]���ꚵ �_�#��tl��(A��ƶ�{�L�������J�T�Iy��C�ĕ��lh���]���msJw
{d�,H4�ŋD; D��d����0�A�+�"�n�;a�[P��!�U2�i�v$U&��I�����f�?�;	��	#��_��*T�AVgP���ʧh9������.��˲�G��f�o�<ffN�q�R�9bi�V��~�W�*�O�t�hW��m
5�#�~�oo�)V�}�t���UK5��0�p�iM�lD`+1`KEr���to�yX��{�ff�Y[WT� ��j2Х���$Z�r�F�x����`��,����i�憎����QТ�~&.�	"�c����ޔ[y����=<`-���P�������|��D�p��=n(HH�7�_�^�O��N������x�UO���9�<�/��6�45Օ��lm��6\��c���⧧RY�\U��_ɢ�[�\��55,�v��W�ռ֜����~��9��|m�BI���~�jA

[�vYm�=obp��%��?�O�țy/�3ɸ��4��X�2{ˬ���)�S�?/=��ڄc0�1S��T;t��ba��8�P�v�����J��d���+f��P��|ñ���9�d�9sq��lԨ}�X�+�����{-�d��gS���,��.+�|�!�����n?�a��>Qg*u��� X�Wq�p��b��M������L��%t-(�o0�Y�Z��G�%&��`�ck�;��#��
�ť� ��2��X�D8b
�Hr�� �\�&���$�Bu��`s۹�OfR؏6JaȜ����=5�TEs@(�ޫ��_#w"�ف9�&{�,�kh����$���mT���+aL?��z��);2o_���-g/IiJ�8s��L^�n��oUҿD��"3�]�QB��D�����b�m�	��0aݬ?��z���=#D��)}�,s�I�El��ﾗF��N��.q#�
�*Cu����`���f�B+Zo�K��.G�S�֛����ϴ��]H��*�^W{�����Y��X:��Y@��t���DN@�m �)$'_p�!���f�������d��l:���N`�T.�a��5̭!�s$�5��t\Y���yDQDe�є�WV	p:&�Q�<��0q��[jQoWW��VD"��LL�{�����+i�cn����߾���(,I��x&�xxxv�3��������G<ч���%e?ßh��(��T%��̽�.���*�s�`�E�� �6{$H�w�i��b��R�����@�[�$8�rkB�"��TVě�d��t��~k/N5X����Z��i'���G����ݓ爜�,��E��bJ4�2.�����G�_zk�	�`�UL�����0�?ߞ�ȎD�Z"P%g�ñ�;)��Z�˝��+]��2�g�+y���Gӳ+[Թ
:	��Yc���B6�9����?<���o'��wՔ��E����}�b���>����V�5x~�ݒ>�D�\�n^���ʧ�M�=L5.V7�ʡ	a,�&��M�?Ց�2I�E1ɸ��\F�1�~��l1.
�&�h�x���g.����vlsG�5�*��*����9�&�
�<�b� Y��'5��u�����ۅ�����D�)�����Q���)��[����ũ����\����덟�����Q���u����Eۓ��\����ɑ���}�oK1���ZD� �<�U�r�� �B���r�h򁹅����.Q+6�1}�)��[���{^�0�	�LQ�t��]���sI�	�9�}�^pC:\�c�#��fM�F��w���1��������vh�R�f61�g�y^����5;�6�X`M:�����F��۩ɾ���R&ʙ��c� �� GArӣ�7e��R|��ۭX
�_AX:���6���<�����1���}E�E�AY�����1cq���xQu�(r:t��ZE��xA�$J,u�J �.�A��\�85FZZ ����o(]0�P	� B��aM���šp	��Ah�Y�Y�ds�Q�.2\!�#�8)]�)f���Ш�u&�1ѹ��Տ�Wd0)�)!���?j������ɀ��3R��X�<��&�??�EJjj�叶/��A�Y����^T��>��vub�fJ�<�>�1���q4$>R�2���,P�:9�f���,�e���RxT?�cSH�������z#56}�ƌy��~�����;�s���ۛ�rlI������&K�PTV��5����뚠�hv?�_i��횝�\;::<��<��<�;�^ۇ�y�����2!�#gC�%&&G�������Z�)��d��lJu����@�����9�����L��������;緫�������p����O�i��S�S�Ys�=��E�\��\�7��~W=��׏�~�Ocm��a^�f��*}�+�ǭT?g��[��}��VEȟ�i����v����J��j;���(�V�h��{UCp�?��?q���p���\݊.�(�fb��mن�+�\�ˎ$N �jb�k����`�`�qUbK��Z*�y�^�P��,�0'��<�ك���(\DaI���:��|"�����i1xc���֛��w�3>��a9���w� ��)]Ȃ���v?nX��s��^�6��7;d��%�B	�9彟��# �G�35����� �(�ί1�I�G��{��}����)�*�s�n>'���σ8bƌ�� �r1����fV�&�R;� ��_:͡��Τ�e/����3Aw�	��cu��v��7ohs�Z`o_j���m��VbO�S�b�k���ۼ}aq�Ze#��װQ�N���X���� hA���kR����G,߉WΈ��p�bh��|�K�JYzy�H;^�4[�[���Ks�x=�D8)���F+Hǣ<�.>��K�M��ɮ��0��������,�����k�AM�L_E�o�H��ᡥ�U)e�in΅�]��U9��� 6��� �E��@ ++�*R`EEEYY�ϟ3�g�\\$'�擆vh&Kx4K�x׷�D�wnPZ�s=��l�hkh�B�W���+l����ً	��,���&:����������5��X|�����u�q�~����ғM�X�SsK��� ��ae�|����Y-�M�o�qh��߯�ca��|[�y>�+���b��K_��AR��4� ��R|!�;}`^��Y ���q�a��TY��Xc�0��o}�.���o���Is�����M�ûj~���?Ї���1�f���/�mP�+��1bQ�����F-����C=�����]��;���(����l�D/;�����V^p7�:�/���_�40�P[���	��3C�-����@�_���G�}��|�����q����r̘@,7�.������/L.��.��r|j,T�1CEAVP:9]�mg� ��\�|��-Mu�6cN�ęR���ɨfVV�(�;g9���R�
��JΚ��ݡe[v�k�7eru�������n����d˪�X�˨�k����5������|fPlI�n�gN��j��mW��ä�Oz�� ��qEs'�	:�P>�ǩ�:~F�������H�cn�ᕷZ�������Z!�;��թ�i�+
����w�S�]⤯���ɅW�P�s W�����9սyM���,U���t�eP[��S�-P$P(�]����=/��]�S��-���܋kq�����9��L���d2{�}����}��RmF���>�m!i��`u�"h��Y���Ls��k�-Dp<��jN�4T�@��E	��62C8GZ�򬚨WS!�FZcd~���r+����O�@E�����������c8q!ͱ6S-�@9Uښ����& (4� �� ���H.�4�[�����X�B��Q�_��4�g
�"|����!-$1�-ه�g��8�A��Ӯ�5uD�a5��6�ަ�v(1�{7��6R�Sqn�P��$�4�`���{��jn{�~L"]��s����_-4RC1��7E8ˌ���m0�9n�h���!y�70���P��p��Lv��2V5"a�Ӓ���W�J*�[����|�D|�H����I�x��23��wia�oq��B���G��&����~�ǋ���3���������%��r%٫�	2�G*㈟�R������3jr���SJ�
�%�����E<P�7�V�(�d^뱪�]?���j.|�2�ڶpB8<�6�ۂ+��K���D]eDբ���CmɮD������
{�C��6������\*�\c����b)|����T烼����"�q}�v{������H�~�_�9�!�BO[�^7z��ve�;��ד��?=�����O{T{���k�,�b�������w#H��S{�6���~;��Ϋ^��nN9wm��Zw���N%s(���N�1qR�Hr}Ɔ�a09.�gurkB��E�G7�៘��vf�5���G�!����F�?&�o�!
 �X���D*+3�A�*��,�N9~���?�Z����5{�S8S�|ISw�셋�������#r���E����3��3VH_����:Ԓ���jR벜\�/��/n>�ge�S���O�c�7V��S?WW{�1��d߯����؄dO�n��wE��ɒ�H#qcPr�i��)�A{��|�s��DT�X�1��2b�~<��7��m�m���_y�.g�G�T�nW�j�rV�rR���)�z����83��8�������YH�p�Ӊ9E���a�-6��L��m��\ ��'����[�Ѿ
ß�7���`�{�������aO�A\�Y։�`��[qԮ?H=D�TP���Ñ;�(����ѿ�:n��S�'R9R[g�!t�fU�R��QǞ�6�O�/��Q����:���eM�Z�Ȼ��ڥQ���h@�
�oau��sva�lN&�n�s`���� �O�"l�/�g�s�s�[R�!%���T�$��T�X��5(�� ��B�DP�&�a��/-LP%RN��Z���.����QF�ئ�Qk�W�}��'�����#�ױ���E�.1��W�%���z���]ܽ�y:@x?�� |�oi�����v/�h������"��FWʇ�� R����&Wʗ^�o��l�wF��Fj��z�۬��XZ�\N�+����īo�s<s��+��Y�8\�I�@��ş�v���ʕH�J`C6��2��:��t��f����f���)~)C��k�F�,����9Hr����k<B(�%ޚ�1w�٭���s���L@4 f|l�~�@:@W������p$�� .`��{g�헿�d��_����V��=}^M�[7;7"���o��4H	�׍ǩ����Y�6ޛ]¾'c?)t�^�֣�C�|w����si�m�gK�P;��VϭXT�����_*��Y㞾�:sN����;��v�9uq��������� ����=(�iJ2)���D�b^W"��۴�*��&PJ��\�p��~�$R��a5w8筙pQ�
n�j98��"����=���[��M7�5�=������v�H�y��t[�Bke�@�َ�Fbs�����(�%r���Đ:��q<�s�W ��5r��,MIkF�R����Rf�g�.�/�D�X:[0������d#c�r���MZ ^���ic)�@��&?4z�Y��\(�A�"Hs������f�����;�����`釗�+��CF_c�g��^���%-�>^ߵ�_�8}�dA5�Z����x�e���-����`��ѝ�]`f3j��9,��7��!7�UA�R�������f������Jq � |�z�u<��,��s�M��V��*
�3�3jG���;|;��t,|���*�pq	j~KVSY�\?u2ƚ�>�k07�����ʭ�%��*��~�@��aa���x��rT��gܲ��ۖ����W�W,���Z��W�U#��&�ҧ�����(���u���V�;��f|�KW|�
�����Yg�
�4P)�	�L��;���h��eQ5�����K7R�h&�Q������"�a��T�P#�$����,�,�s�)X|_��*��|�;�b��(|��Mw��C�� ��
�ݪ���
r�U���yA�����K6���{��{���܅~�b��$�3fG�ӡ��]�b	4]s�ߍ���*�>��N?���'م���O�^S�~�:�㸘���i���R�H�Lu]���>�n����Ck�J��e*�o� {V�|A��X�0��(��a��<���N�\�C��wG��%��4"���um�S� w��,.:�/�2S��x�\�G�@�q(���0Y ��s7��L�,��ǣd�!��0�*��*!𸤺;���W�?��4W��&z�,"v%�+�٢��?dX�╣cj�=���8�6dGj~X����o�׶�{�$�EhOg����ǻ��^x_LK���@W�Rh0]��0mZ�r����(iX˰ia>9�Y���ؘٔZ��}��ys�K�v�O��~{I5�$�r�_����������j������u�������_��W9��0Z&�!�(+(�"n������2�J���9�Di���-�<	l�m�XL*���|0����dS� >��`�@�փ����|�m�\�J��圀 ��?刨�;���(��B;�K2;6<h�=�Z���Z��r��%�PF�����A�R�L�4ߘ�X!�'ں+!��ƭ�ZJ%�Ȳ��ޤCQM$�����m�rJL�)��&������3��9��Q�����{>�{xPF�	��������>��p�
!��~��梕��+M&�3y��!����$e�Էo��ڑ�T��?����R��#�D��oE0#D	������bŭSt���SW�V/Õ�4�	����C��2����`�y��oc�FD�V��'ʳ���K)���I:��!K�#˒cj�l�0�ع/-�d3��SFt�V��e�l����e�g�Z��U����e���;����B���E����,G`���[���?��,��~:���Y��������c�M�@e��F:��(:�Ȥ�f���٘��s����6�).1����"d���Vw��՝�P�V��P����R�/o�`�:��������8��Z��$��ڲ�צ�Ҧ������`x,��ͻ�w�o�z�w�߾�E�rq��G��,�w޲�mε�L�W��f�{��a����E����1d.,k�
ԩ�߫��b�����t]�w.%�������t�]DM29x�0�r���Մ�d�O��G����[�$��$(Y&(�2T�ܿz���WM~�$����Ӛ[0��W���h{�My���/9�i�^�判aS�T��)YT��J�N�R�EeVb��ȹ��)��K���jcM՜�M%�A��%?ҏ�|L��#}Y���hֿ��������u�V����6[y�_���`�V�=�1�]Ʊ���R�����di�P�A����iEn���f^c�O��e#�
p!B���q!s�-I�`�U��Ŏ�%�kr8xoS�����㾡������wJ�{�`��(�D����rqx<���N}�N�e������	���R�W{;���,�~e�`7�Rސ��pf��R�����9'zU̾�+^�S��;�p9O�P����j�7�Z��܁#3�pF�7�6!bv"���(�f�Yb�ׇ�H-�/�e����ž�NĲ~!id����'^.(�a^?j�R�(b=�Ċ�>�_u��w���_���v������/�s�`���PD��9n��O���IrN�-5���',���'�x��i��,���<�,�+����:�r���1b�TE��׏��:, �$�5��\��l/
n+9d%I��Sf�x�x��N,p	9!#��ǺNs*ML^�\�z� ��~�B�BT�uݺ,���)Bv�h�Ht d��q;��ib��[�"%�)��w?��S����S,e�a���̦��	����د��T��B�)���V�[����A
{�B�w^0	a�K������0���6�4j���L��Un>���B�(@�ݙi�<;A	��(�m���oQ�V�&L}"��K ����R&=��\��'��?5gz�./,�E_q)	>mᏟ,Z9M�u/����
^}iD�=�K���r�v��us�A�{���r�������t�ϥ����fE�TD1T��VB!Wjߋ!�ZJ���>��y�r*���'�t�;x�,ڡ±���?��������è��d��b=쩾�=���e��L��)����e	�:���섍���)�a���׏���Ɣ��LR�W$����Vs��8h>��9����<�����tFAQq��U�1k�e�&k�b�!yS��~��"z�#	���J;��V��BM?�"G��/��@�l�k�M�9[������x/��V�k���b�P
�P��\�&� �Xi`�z�0��,����Ej�9�,��s��H�AA���Vr�0Z�pF1����c5�t��/?�bt �%��nvW1���w���T�� ���\v.����(�IBZS��wAB��*4��x��ԩ�}$�3Ng����X#!vU0��Q��]F4��T(������^�BTAx[BCn�:1W&�H�`�HU�1��r��3fޑ!�l	rӢ�6d6�I�#�6�ctC�W����C^e�E���%�aD�S¸�&�*3�{/��d{��t ��Wewn���z8(�Uӧ��#�fA��n
N���f?�Á�D�Ӭ3&?
�t�=ZhmJ�T���ˤ�K�%j���8RE�h��Xm��[2�,ҽt����:���'h�����`�Qs����J'>w��>����wi��O�v>����Z}�.��'�v�;[�N��ɻu�|L;*x
C<��hxё{sh5i�\��Q�6.p���W��V}�5@S)L��{֫��	se��9b�G˕4��> �k�P42N�S?$���ͬv<����ȴ�=�� 알�r�����r���7��&4��^x�+gϫ%�F��ʠ�	�`�8��)���?^�o`����l	?�8�{I�4�0f�2?�4D���榾�N�y��e1��������u������վ�U4 �R^��Mu�� ����N����h�EN��s%=�iy���W� �;�C�T"|���vDcgu�H����*��+��	8�v�7���" ^�u�\�^7�7�/�bi�T����Q�V��\z���N��6�|�oia�8�j��qP�v0Pʬj�TӬ.<�!Ľ2��=[ɣ!����/��I�ިu�(�� l��M�y�{�Czx��fջ�x�jL�mգu�6�]������+B�^���N�հV���t���B���Ԟ�Ɣ������F�����kKW	�Z�dhh���=��#7�',j(�ԿI���[�xb�co��0��rJ�� �Gw";e���!��^B��PЫ�u\�N4��Tf )}�jA'/�uN��-T�����/��x��մ����ѣ��ӳ��������θ�	W�ks��w�xC�4�]�8e�'{�o�ڥ��� ���	xW�����w�����o������#�(D���l���z�daN�cER[2�/2b��/�2�oO�>=x���!�1�͍�w��V�5�c��>�W�z�N�J�LOWui�F��@���+�\���l����x׺>�fV7�����%�N��2��FR�^��槅�`���ِ����PYT��S|�#�:��}�JW�^��|�;[���2f��7���t�	�$"e\f�v,}4�Bf2��w���up:j�yk;E��ĸ~�a@ �}S�����h���SA8�&`l87�`��鵜)��K�*�C�K�FK>���'H�t���p���l�R�M^�e���p4���L������<�՝Nq�{��P��	EDU�{
$f�ӝFp�"�W�3֋�J�-�6�mI-��I9��h�L:^H,aY)L3�ls̐�q{����(Z��31�o�g/��n���L���9 p���1=2����a�.�g���>[�����p��j(�/r���xW���*�VF�D��BD܌m��[�6�PZ��v]%6�
U�V��Q!�x�ǃ���������@���ja��G[��[W-}���U�~�\M�f�x�%J٧y����P�u��tTo�{n�����:ߣ������RQ�K�Q�0�?�Ĭիa'��U��f�8��o`:��O*:��3�'�L���	W�+6�֋��w��0e�PL>.,����T������]���4��έ�7T��Z�}eД������ϙ�����y�9;f�s���M���5\�ӊY�|.����]f���i������of�_�J}��o��ݲ���s!\V��խv��MwbL��zڎ�F���ߒ�4t����9��kI�F��Mv�:�ǆF,����EL�׬F]F�����#g��S&��w�rdf{�j�rF$���;�͏��N�Ɗn�*x喳��?�҂ө��^��O �.c$�=d^���P4s3S�a��(C�c�w�Q0�J@��XK\�'����a�Y�͍��ƣ\�k�4���eN%{>� ��g4n[�ݵ��m�'`(^�#6��S�\�W��e#�9�S/��ӧUuB˹`R�pB��hG����VF��Ѕbձ��Vj3���~1j�т�]<F��ƨa�f4��)����t���f��v�����]r8�-R74���Ajf0�d�}`��im1��mZ_֦[�'8��Q���R^ﵸ�]L*.Tp��/��y_��	���.�}�a�=�X��z���a���IK�Q� ��83/<�{�a�D�p�m���ٺ��&E����M�3l��˾�6�s�(�`<�pP>��C(�N���Lx�(;�(5q�c�.��N�,�Ce�?������G�r�|�&��̘�d������{��dށ����M�q�J0t��^���@[@aF�6�$㌔2�������L�)�{F�?q�nlc��~}N��a���A�r� "�7�z���Pژ���7�#���pp�/)g���$����纺�܏UUUQh��
�tb��M_�d���8�V�V
���Ʒw(���"&����p�=_�
.�&��G�@���0%vb���S��}���o/��,�����Ŀ�(�M�Q�hY*�̚���j��-�N�����wO�M�w���W�R� A�@B8n���χ���;�Sw�y���l�h��]�/�[�u'd�	��S�SU���M(l���g�����bO�\O��׏w_�#[��0q�`M� �ZE�*�	��v�3I������jǬ��Ʋ`>5&.��ՍN\���ՠo�XN\0���a��l�^mmZ}�W�*M�)I��a�ڤ^��Fq0-u��\���ȁ-<Yr��{�x�x�'��.H+KL1:-U���U���r�`�\x�*h��q��P�8��� )�u,����ZT���'�"��A0�A�i	�M�68�
��5)��T����Y���m���1�Ԋc��)&Y�Y�������!�Y�}k��!T1��e���&�4"�n��"�BU+����	��'\w��W��(2Nڜr�k�ݒ��R�~�@�f�KϪx�H�p�_�ś��.|�<�"�^ ����H�)�ٗ|����1��oE���RK=]���>�_��U&��y�7m�|=x��x�aсKD����:U������X�@��C����$�Z��E���ɢ
8�(�����-�O�w�.��"h��?*��ؿ���a����6��W
1s���}��OX �@�@������i[�%�0�$'��_<��E��Q�XT��
����e�Gm�"�\(=���mZ��-*m���JB��e!'e$#/�Q�T�k-^��t��)4(` �����C!Qw5�RV�N{��9Y�k3���
���� dsT�Wj7]gC9:1O 9s��7���(X^B�m}���F?w��%+q��B7=�C��ll�5���:vm6[�yZ�-��B���TM{=C�b(��d#x�y������w㥊r���8�g$�<2!���l�N�|5���B�Z������(�	�M�@��ʛC�5SԮ��,BAx���|��R�3��/�Y��/tJ��7�J:�c�_�6ƙ�]�P����G;�f<~�s�r��y����/~m����{�)y��tqB#�H�ᐯ�Q���4=Wt���_����B�9=�MŒTU�FӚ�_1�;��օ�2	))}^s6_66�ِ���z-�W�BAVP`_�J�"��M��Em�s��'���-���F����Į��Q�/���L}������Yz8�y��X�7��c�Q���X���HSE6)��S�㶒p�ۿ'ߗ����e���ϓiR�m�\_S����}��_�)���������>�G&�\yPG�Yv���=���}F׏jC���"'p���U���2�?��i�R 6�A��[ �$����_bOK�j�n4�v`��cƞ,Q�!�Ő��q~f�o��⳸`����8��:H��\�7,�nw,�#~cI���Xu�V��n]c�(G-:�t�*	�˫�'�����f&�1�3%���RL�=[Rޠ$7vf���K�x�"n�q�gx{ci7n)�O+}�}��{<[� t��߈R2[�C �@�5N���hda��aݭ	��r�#Kʿg�Ǚ���j㨤G�'{��[�nUI�*�s{U��&Ǫn��(��G�+��8��!_вq�A7�qY�b^[hM�)�����ɰ�4�����{��o1<hF��� Z����_���?�����M��x�z-h��zV�]s?���
+q�$�t!)h���Oz�*F��ܨ���YY���������MRwT�JT`u���A��o�:^_��fۃ�;M�b�bB H���t�k䕓�ְ^5�Dc=m ���L�2���xSCb=���o�d�mz9��Kvm�=^=���u��)iD2�O�2jp�� #�������K8 ����t���fG�2���
H�7�7���	�d�9��X�iv�:T�I>�'!�}����qlzU���YWW�B�?�/�Rw�Ǌ����m�@�k[��Wt�W�t�w+_�?�_Ko5�� ���+Լ)��p��N�͘��o@ +�_$gs�?��Φ�|>��oN��B`aى;)��~N������r���X��9��0�����Vg��]�^m�����{�ן������(���7��kב�a��a" ]�hX4�Ty���H-�Jz��e	5���(s�'	M$��Q���h�Ks��b3�F���ˮ��3���@K��I�����s��|��&���c��"��R⇋�U|Ys��Z��Z�WΘ��ĕiȊ�Uሊ�>ܒ#tA�X�Zը�V2.��x�(�^[��k��Uճa���64g��K))ë~C �K�pf�Q�T$g��m�lvmLpP�����S��ղE|�+[`�Kbʢ�~\k�e'�+yK݋��i�'�/�Iu��1C�x�R-Q���'�zc� �!%�}����\�]�v�,`�și�#<�}5'h��d_���?@��s���ޑ	1Ӈ�l��U1���l�b�	3�o=NHo���E�b;��a���F���M���`0�hL���Km����V\=��R�m@籣s>C�L�С��3�j�id���@����T�;=tAƫtit���6�O)�7��.d�>���Rr �iĜ@����\�
���%�0Ď
 ���Z6갎�0|�]�mbD^�*�F�E�2�.�r���; I�=�ڬȏ�8Y;�W����!@��X,�kY.*ppƌ.'-�.VQ�#�[v���:����^�"	�+L� �wl9԰�v9���@r,fff�\\�
6�����]]o��GF��M��5��-�(����z���GED%�k�d=�"���כdC^��lO;�Gx
�vZV�>:��;�=�o,�"
�³�':�PN�&�FS��!�NTv�>_��K��}#6�߻ػ���7{���mI	��F2\���D
�jҴ
�V�&(��EF��G��Յ�lg���d�O�f>)�G��J�Odj�&��}¿DL8�Ā�` d�������-e}F4�(�Û���$D����1Ŗ�rni*�J������J@g޴��^�ك��S\�1Q�s!�8�u�S����	AS��"�)�xiQv�ҽ.��_��~���[�_i��z�m�QX�IŹ �Z�����R�O�!6�����3Y{�� [,�&����]����F��O\F��j\�*��k�`+©�y��,=:/�O�Ea'�1;�8�3����<�Ƞ<�I�6�v�"z`�g�쪉��j��]�ס�#�:����zۄ�u�cp綜�.�Nf��������S8U����:�7/g��/'�l/�Y�//�O���^/wo�)���d�-�'��)Z�/$�{�zӬ��.�����/P��Q/aK*#'W�`�)cUW�&�r�I �ۢ�ϓ�C��������������]�!��Z�wЌ�g8�N^A�i�2�9���9�F20�"c�U=#}�μ�	� �'�V��'�'�T���0ՙ雷��P[TFub�v{Jp���Ui���di�X��"����x�
���̹xV��^6X]�# �.���T�(�[��K���!dثU1�p���e���W��B�<V�˙Pg8)��h�4��zgUݹi�L�y�I���e�4��J&�o-��Š?[4ۊM��S�׽ݯ;�aEO������l���n�H�Z�K��=PF�#�ӝ{��S�#:��s��s�Z����S��.9�i��������Ķ�{�\�#��t9�K�p�۸y%�46�v�e�q<!xٹ��	i;�j����Y�GG�]�Sk�	]�u[ �ύBX#_�7��L|���4l���U:���tv���ۭ��ػ�9�2�_��	V�uu	b����D�� ϟ�s��Ɏ��ِ`N���<�� *I7lġ���ق<aw�"m�d
 ��O�i�SK6��DGI���+�����g� �`�"z Ka���'��wA{rttt:::�=��nͭ���;�%u�|d.�_z�9��xFy�y�M,B���P�?�q6�r4Z�����P�M&�	�d��(���;�{���b��Ǫi�Y��`���BIL��7P)�R�0��������$��q��1^�4����쟉����OY q¦
����w2���h�%�`� iY�y>����喢Q[��1�� �R0��O�u��ԩ�B�^��Zd��Y���8��J�$<���N���o$�� m������+�d#��s��r;8��7��oۍ���I~�P�^�����N�3!H�=C����0(p�;��R���ƙ�A�!�h  @ �U�e�<�UM�U�8����#��`w�f�Ea�W��|�T	G��];��+��0�Y09t��M�Gq�f3�ld�H20��%����y��쳚��bWE�@�QN�q����}[��Z��:��R�^r�U�l���J�{���]��%'�?��ր��+^>a��(�����8ȱWj�l)Q"O�ښ|-��� |���Y@����5�-�	V3�L��1���L��,|�D���y2xp�Q�!Q��z<�t��yE��E��Y�,hJ��>���tV�u/�A�о��l�}�o���7��|�7�Q��Me ��:@m!�m"�%��$�4lc��i,*�D��a)��B~Y�����!��Ai-�TE�9��D���"�]��̅bC"��7���w�Aq�O|͋��'�����[��K�. ��Xթ��dz'6{���.�}�`���`��
>��6�)\��zC-m����O\�tC}:��qU�Ė>�E�ʱ�Ӻ��)�N���evae�*,a�n�hl.�v�2����x5�Q�}];t�4�*L��ʋ{5�M�o��YM�P՜�-����@���X����c����P�� f>�n6��9�z��>)�������N�@g����"%�F3Qز�>p|8���.�̘Zט'��z������xw}W�ŎN�Q)��K�В��I.�q�vu��Y��&����k�y?0٩ߎP~%�z�O��Z���\��0ڲ��c�LPq�m�ARP�F�3I����ǭ ���Jl`"�I1�}��^y�;q���񿎚ӎ�-������α��������oL�iB��Փ�Ԏ��������HQLM����*)/��i{�m�y�f{�n�h~�xq��T�}�=.ڟ4��٭
?�)z?�o3��9��-8<�v7����-�N�s�ѱ�����u��%ae������1-�]�;�;�bCy���AV��W���$f��vo��]���$tE���0��'��|')�y� q����ã�at��N$}��Y���Q��g5���F��0����s���HUW1Rrtጶĵn-�7O-��7m��a }SY����m���*��{9���Q��IB����ڱ�~OS���+��f�an�M��24M�Сl.W�c�����0g���=iRvc�R���R<Vȭ�y�$�ȨQV$E�nJ�/��ͩ?S��?�*q�^���+kx�����_�G�ے����4���m�4m牏tI��'���͟Xƿa���u��Y�[8*�z�o���y��]�8�z˚�D����=�W>�}�0H��y,~4����g�����(������fA��¿Zm�#�)Q�j�4	$��q�V#���QKj�;���WO�'��Q�%עa�ݤ|�� g��[}py5��
��zqd&'��)-N����&�p��J�6<�������q:�H&�b�-H�Ω�/]�#���9�.O��|�z$���� D�F'%G���~h��g��SMk0�u��lk�b�b}�!y�7������u�§в9��B@�g������stK�YYZ�` L�1)���p�������cV8 @ v�� ��iX�����8����~���q��&B�?D�X��y����i�����b�u��{)\�h��oߒ�����њ+���wq��V|���Wq.��Q�u)�j%a��yvM��)2��-Ԥ���Hӻ�f���=�Q�5J���j9E��9x��w�Mp7zɪ��߅z�#�D6.>�ZG>�����"�a��n��o)>�0��sx���������ٚk{		��'�2��>2*�[ʖڅ�_�.^Uv����;�Y\v��e�np�g���fĵa�}l2Ft�j�$����j��O��(����`��ʦ������a��c+-�X���%��16J�b��5��/����x����52���h�UL	���b����y*;l}Sj�x��í�I3�����m���x����sf���n���`ogS��$n�m�]�i�)�:�@�0���IRE�G�Ӈ	~y�ĝ0s�JGZ*e:9쫑�ײ�����.[��~@�H�\�U��=2���,�S}(�r�T�u�z:T�K��ǣ�/M�&OI��� ,=y�M�B������ŕ����� n���a$��\�`}.�Ly7�Y?$�C�D��ªW@E�xG�Y�1�gEKq��B U5�l�*7��`#��������}��Ve��FJ�;-�L������:l��.�t��N[��uا�!4mR��\�?����Y��d[�wj�~͘믫����!L�+T�k�A �y��㞳�-U�m)�� ��-��Gؘj��qO���v�))Nr����95Կ$�@���.�H<?8��)`}u1��V�A9sD"����<��M�������v#�ۋߟS��m
�CBv����C"��)2c1��trq�	������qQE#l�
٩$ �ޞƀ���{ n�3/��%�Ѝ����S�u$��ܽASW�c��e��)/p�4�|ug�m�,�+�ޣw���?�\nZ�� �2��3�su�E�8���2���T�Ԏ�tC7X�>�+M�]r8~�]�|4�mE�a�5q։��6]ʓ��	���!��/Q���Y���=�}QN#�S�0����$�������羿 Ԧ�nh��e'ib��9V5��4��7�*���s6y�U��͵v�d�~���F�"0�a��)��-�aq֒�E��1�� z�Ӎ��e����˶�����M�~xӯ��s4�s))��/�f;r;ɲ���PZ.�����8���f�E���i/��{�����~)&��E�8L����99H�[�;������C��	�d��8�&
.	����pg3�u]:,��D�k�/���������+'KV��ծ��l)g*J�O����~� i_'����{�x'��5�Ί�BT25��,���Z��Z#�������BQ̓Z��V-���{5�'f5G�\~I�P�%�l9MQ�t�{X0�4;��0nq��F��*�P�[�|p��hF��C�0�]�qx�}bi�R�[��F�	Ҩ���+��CuA��pȇ���n����#[>�2�����־"7�b[�����?��Y�[��疚�{X5xyd;y�����v�z �U��&�?��f�^�S�w�	y���/�L ��dO&m_AkOI�\^�BqQ镗�6��syь���6%{}&l�2��Lo�B�X��2��9�*�H���W�u�G��^`)�\�]:<���f��7���K̞	�h� c���(0B�n���cD
$T�Q��C�۟әus�ă��9������N�f�a�#��@&b2�:�a& U?��0\�Q6�d�?4�1y��͍.V�7�oP3R�c� �'vJZ�t���ϴN�q�����"�	$.w���g���#F��������_�e�@q=[w�_AN��*�[����3�G�"Vm���R���%���zE��s��@�ȕ�S>09ى�Ij����	�i�!q����>-�z�}����S½��]+��W=�J��J�D�v.��Q�ӏ�f��H+���P��k�_֖�Ge1DZ�E���,���� �ϟ� !�|_"{���x�n��@?��oh�K�`|I��$*�~�:�L����/f������������ܧ�^K�u��%�G_������wg�J�|{h�t�h�)iYBi7�O�]uo�O�4*�ԯ�J����/�9�.\����x\%��߃��R�V�Ad��B8��b�{Y�}�oM��) �i��(44ǥ�8d��od4G7i��%�K�|p�`��k�/ҕ�x��~�M.�]^=�y�Pl���vP�V&t(�5�}����/?�]���a�E6C����}0�ϱ2y������H��M����ձ�V9�d%��?p�mȧgo�)Q���E�Jp��g���hR�[��|m��-�GO�+!m�&V�~l��B���#�X���>o�70tY���?��S���԰�w���G�{��9�lU�=<��|���[r[��}�Y�3g��U{>���2�dZ�K�Zܐ��i-�rqj�����]�;����x��W4��GA2&!�"vM
� ��d��y+�;m[�0h2�vL)-��K������dcM�;#���͘-���i>�C�+� ��4��HR
wd�W�7~m��
o"dQu֍��M�F��m��Y5�隂�/��3�ƘM�~���@2š�1�mr�Z�����3-������S �(�5g;���",Q���;��\���%)��Ă�ok!�[�ߩ�*����G���?&�K!^UT�g�]�?=nRul�T{���u�@��8���a�" ��h�n�G^C�n9��CE{D�����4	Tc��~'��:R}��� �҇��-�i��t3kq���,��Z�*�Ag)f�
�DP��`���z����@�Hh^��=��,$�xH�������R1��A�v��2�y��hm�f�J� � C=���S�9�ﭑ��v�]=�y"[�����@d��E���6/׿��������	�-N��0�k�	�������Npw�A��wgp	��{.�9��Z��UWw��Ou�z���y��	��?kn.�i���������x/�<�>+Ũ�~����m7~[xmV�*�5x���؄D���.xO�j��I��|�z��+�mªI�!,1��Q�p!2�@�84UL��(��o��CH���ޞ4��8��LQ����y ��X *�1�1�-���-ڣ�=�I��f�I��,!�9�w���~,�-��⁎l�@'�t]}B)9��f�������O��A�6וϪ�cH�QPB^QZhgZ��&\Q�P^�BG� L��C���)X\B����B�u%�r}�0�E<u�p�H�D��L��sl�Мϧ�zV@q����0:��0���hw'��M�(�^��!+��F�pX�^l13��(�@#d&>�K�k�0��XX���X��~�Rv��$��Gw�����s�F�k��ۤ@�S�"�z�8��4ܨw;j�͂n��^���y�� 
^�����ƽƥ%C�2��D�ω�܉�ܛ����܅��ѧ8<D���IGc���V�+�QˏI��v�`-���`�zG��;��h�Y�έ\Jn�w�]LSO�z(�n)��|�e&�/�eV��%�Ŭ��X����i`�u�M#���ؿ��	>����{<}�Κ 8�!;��<��9UԿ��?W�ᤩ�=��Ft@Uo����l�%���v�gܛ��m�%�*M�G�V��G����j�gv���V�Q����j��3H&C~Gq�u�n��m����/�ZA[вR�_�Z!�
ں�7YS� �@�uV~�
����cd�I�軂��2����[	��M�63u���(΅�Mc\_BܣF�% Ȅ��_�C��e���R�1ǂ��ϖ+���Z�o91��T�N�25U���9娑����D8��T��rd�
ܢ��}ߜc̜/���]
���U0s�&�k�J�#��\Z�[���Z�L��&"�ue%�����2�gU�A�9'hP�h���W`Y��f�G�4�}��3l���\̮�+��23ƉNuP���\��A��^�U1q���-VG�ϵ��u�Y��7�#�UU�4�C<��Ta8��B��t)ʄ?^ό�5���&zL(@������C�&O=^�
�<�E�VV Y���)y���U�T��WR�|�Q��7x����R����ݻ�{Di�;����vP��=�V�����t�����:/�Z;Ϫq:�ʚ���*I��.jjFFv�7���J9/��Hya�^J������*-�Z��kJ����E�#�5̈e�_�8�o~�Hs�ml�¬4	��ӬQ�Y� ��;�v������,tHk���.���
�P��XL�dbn���aF���'����+�"@��!Y7h�&�P4}�tּ\���7�ąJ��cOީ���ֱ�zI��B���@�Rr��09!�iY�9R�iׇ4�MSa!*�q%UdJ�Pj�T��ݎ#��!J��#
|mzIͼ$xAMљ����ݮ
)���{b�%)�4���%���R�R�zRp�(i#�M�Y��u|��}𳩔���H|W���Zt�IF,�AP���i�A��`Z�oȵ��͜~�&p�:g�aW3��@�p?DD��Fͼ}f"��A�jx��/�J3g�)��i4��d^��Zed�1����@�ۄ�wAb����b���S(Z1�EѼ����
G6ҫ|��f��4���%�nHۆde-��J�t!�D�	J�w���+/���%e��q�U
��f�^�/���s��WC��)�z������ �1�ͱC�E?2�	*	?ѷ
��AjAL���A�+����Cz�}���J��ZZ ��(vc�w¸�wgͪcVc�ॳ�j�ߵ��ꂪH n���tR�eP�%}ԋ�6���3�D�R��4s�G?��!8R��\H�����F���9����7+��a~��g'��Ur3�h5���YiJ8X �j���
D���@D~���8($C�?�z��jH"��Kaοʸ�2�J��V���~%�a�~5uY�[תM��;ߤ��Ъ5�>f�0�'��iM�fK�ğ(pz>�����Q�6U��(���* ��ɽe`�	�j���y��9MH6ӛ��"�)Sz,�r0�����N�Ȝ�Y�埜�����ό���[=q��=��{4����"��L���T0�rB��Ei��~�%B�|�:��+���Wf��w��犪�?)��b���c�\Q���� ��єR�]~<�����?B'�g�M<��v�V��R���P9��i��^<u�!ii�s�3a���d����3���U�����8Q[�}Z,����K������sO�h��fi��5t�����5᫠B:~���!�|��Ї��P�<ddg�9���z�a�{cd��޹w,hvg��{F>F�g=� �z1,�54�*@$  �u�z`W�%/��� <w6�Smyg� ��T4"�7���>
#՛t�3Ih���,�i�����	�1���%��W��ҵ�Ը�Ɯ���� �L1=Zlm� �b3���K���3�����FW�zW�i��"R���0xin޽c�w�\w8�";}��\�x>%b'~;a�A��9��-��i��1��X�x����g��M(6��:.G?�ê�f�t0&��]�UH��R�/�"#񐑹	}9�R���!I�x\�7��q�\hZZm[[���]/ ��ڀ�L��+a��|��&n��\���f� ���D���^"X�6==��n���%��m��ڷK�B���6T��'�Y#�B�F�`��i�Ph����7|�Z�N�w�_�˚4p�k6�岱�v��r,���V�:a��mկ��J	C*�E���̓�%2�"Y��8eWp]vqA�WG�j�*�f�ق�U�V�O� #T�:��H�*`@�����5PXXdӫ>1�HS4%�M�X�x`Q��cxA����� vRN����҈���������<!Z�e'uU��"ˬ��������AG��I
���.U��4�R�C��40,Ѳ�j�����=��������Ɯ��DEE)?���Th�GP�E[pd�UhT-�݈ƪ���;�Xx�+��=r�pm�1�(Q�ʘ3���A�3��m���H'
���|N&�L�ATUT�2ilZ�Uk�L�����"�2�8���E�b��,�W>�^A���0���v�ٙt]0+*�t���̜����t4���ɫ�5�.�Y�%L�k)�k��{�k�o�y5��α�[�vN�-ý�b������l%�ͯ�������d[�z��RJy���0<�s&PM�뢸��u�|�"h3��uE���`M�&ZA�?/@��oϝ�¦x��jD���a�ƺ�6�#�`>���p3w̠
	px�ZCE����0f������Љ3Dg1S�ȑ�zuP�ա���W�V]U�,(5�Y�^���@3Y�
">������0���|�7
36�V*�{i�3��U�F���֭Kc�޹{�����7��if���ަ���t��r���a�6ɹQKs����-b����:�U33���6x�6�A���^�[&#���!���h��hEp�w�A�l�\:xb�=`����"�IEq�V�DDk%�D����֦11�?S�NG.xUzG14�I��(X�ഀ�Ҙ�z���Gm=��֞c�c��C��m���8i�P�S� %8iF�1�G�K�I
G��y�2t�^�R���FKA��m�s;��/�Uja����`�T�q�d��̳K̪䈉�9dєl�j�'B�����F��Sk]_c�&#�#�� �r�1ֽqx��@�=Nh5�6I�4��}6�kx��S�1�j��%3��C����M�{jm��	դ=����2k�/��_а��BF��ձj��R���&�-<�7�a�
�\��6:�l�[ٗF��W��TT��3BΞ�u��b��P��9?oEF�5�~Z�R�o�p'=X��}E�;�h�,y(S�{��	����T�<�Vp)`�7Q mA/��[����M�`��<k���l'J�S�V�@&��l���XB�:z�b�L���}���|�<gY�Kf��\Ē�<����懺-ۓ}���3p_�t��4 ^�P�w�v�[\G����[=n����P��N���n�/�Tf�dStF[cN��1�'���ҿ 5��Q�����m�@�-�l�H�3��o-B�Z'�F���`��kʑ��]ؕ
��3���Zل?k&QG�K���ĩٷ�Z��=j���������F�����p�1��p[���V�,VF	X�A�`:��aUFh�!X/��^2p����s��>�Q�ĳ�4ҩ��aA�O�N]Q����D|Y��
8µ	�裓q�9�4�b�����=v��6x����~��Y�T���<x��G|y���4Np2�O���~cC��+�˗l����R���x'�V�&��@��Px2Ǘ������B�}���&9��J.�m��I76�#���TƻO�`�@�=��BkN�=/��W��lUl&)#��Q�9�C��I�F_*RE���	�WA]5f�:���L�����k|�LBM] |�<��*�ldC�c�\d�L���H��Рc I�������14�~���4��@�����6c�gH���{`	W�V2u�O0�ĉm\��Y�a�S�/�[����
�j�H��+�j~��lӣw�t��B�\��:I 0�A^
�7{��.���i�Uȣ���(Vd���C)b�Y��<oq82�N�T�	�V�FV���	�;#T���
T5b�4��t�lf%�k)C�f`��QZ��7�+b�+�/� �k��0C�'R�'��+�Tŀ4o��̓��3��`V�XW��u����Se��|F��j�y�do���z�24��Sl�8�QV�Eh�;�����bcAnG��8&&@����9g{it �>��1�� d
��1�9~�8a����RD��g�|����u|����J�E���Y�sZ�fֽA���C��L����j9V���d�(��U���t)$i�wJ����(]9���O����~`��M;>l�MO�}/����Z��5�M����cjc���Yb1X�PYb0&��fb�)2� ������h#���e#�����od=.n{?�O˴֬w֔o�d��dOC�!�(�h5h�����S�p���;��������vÛ��֋��w����b�M |gv1C6�߂��K_�Y�3��5��U2wo�W�c���K�K-���\�#�AHA�N;��54��}��,j���4����wG4P|�2HLҨ��N{>���u�9�s���Z��̜�¨ޞ��(s���M��8�h�U	T�����>��G�p}�Y����ڿ�W_O�~F���
�����"E"!!EF�~���)T��a�J���IP&ʕrd�BB�{owo�H1��YY�QƷ%i���pH���
+�F(T6���Q��Ʀ���?���9#f�����l"/`Yf&�z��|���Ա�+���?�G��0��KRɍ�3�V��6����!��J3�G��Q�?���Rߦ���ߖ�D����N���4����	8���qK#N��g��j� R�޻���D}[O�8��2�=�Hl�f�i�pQ�%{�ܘ���c�~P��ϘT道h����F���N�{���^�^a_��z�Nr�z�x�Oǁ�b؁�cŐ�ܮ�Y��M�3�\b��=��/.�˛�Q���U�xD|���{���Xо3��C� �-��(�6I�Z'��n�qoǅ�@W��V���@;�c&id�Xs��S�>k.l�sV򀿶�7ʃr�1��;5�!���3f������~i�_�?|�ߞ&����="�wXf�mAgE�N��8����������O�����I�x���N�f,�yX�f��^w�1uX���1��z����i�q1���7�L��M�/�nj����`��c�r�j��,���
��EirA�U��}$�Ri��M��� �y��_���B
���_]���$����3�N2�wI�0�~b�	q�U)f�TǵK :���A#�Os�H�'͐ڙe�?G�"<��U�װ�߷�O���`FbmKh�݊�VV/���4c�`y4�Ykb����vm���Z̥�;�b���+v�Pm���t�i$-b���9�\���������������J�g P������
���H%N�����*�K�/���\.�냆J�^9g�W�x���+�ܐ���/��bv;�E�v+n@���!���y�U����Eo���q��@��>��R�AҪ�DM�8,��\Pـc#487�:��(�.�u}t󛦿����� ��"ae\d�
_�=����ޫ��N҆�w�$i�+�J#�j�ie���[�;����m�Ob��� ����vj�ҟ��5��(	E��/n�2*�g𺈶���?4���1[��Kx5��F
HX����<��	��*ݱ�-�<H�D6�Ȝ���s�1��אQ)��O�՟]4�\`ן��M�Ő��~}׺�@��!�T�I�x�<YW��|l�����,`P��9w]���A&�%K�������9�=��RX���uj)���ݍ�R �v9�yRv��O%���Z4Fͪ�p���/>�Uq� ˶���F�V�B$*ˍ�*}MA��i��3�:xɀ�|�4���Q�T0Z���t����Q-���A�^�����Kp���/�����r��S7s	��ׁl�ebhy��\,��"���t�?�[̃<�n�Q:�="W����٣�� �+��"zO�Q�H@��b�����F�D)��:N���ؐEQ'0�)�_N-:��t-c��S��
,aU_�/%�����y��z}�5	���@9��Ic@Ƕ�*NedV�a�z@��΃�M�:��|/�@��Z��˼�[�N��&__��2�rc:����h�0�Fg޵����",]�����@ͬ��/��0ѝ��&uU:�x����)��<Mǻ��V���@K>@��If�G��c��s�[ߔId��	rl�����S��5Z�gЈAj��1�J��M9>7.�'+��Wã�7Đ�Kt��C5�ӧ�8uX����U�L��~��{?���� ��K��N������ڞ`v�)��A&��@�1h4�-��*�����=���ꢊ�]�xfzc���l��ȯ�9�w�ӑ��SD������z��m��'�cd��`������q�@"݋XM�Z�2�x���!��-)̜(:����)Tdp����	�8�9��4+r}�A��� CK~<4��"|��B:��L*���&l�1s��<� ;P�>J�7 �Mi�&�BL0_��RI�|�A��Q��� ����By}�B�X(Z�h��I52�X[C#Ű�l��S������ ό'O�E�8p�,*�=�� LE�ٜ�6�[��@�Tn�+R�';I`�1�	on�[#-4���:A�U��+��fژ��`έj�=��>&@���X�TTD� Q����m�X�TP��QH5�y�_#g�j�Z�*�Ks������'�9����]Kɂ�̻Vkb�2�y��(cxK�eD�7�e�� ѷ����=�����5�O�5���<F&56���\���u�L/�ʩ�������1���Ԛ۸6@��#�}�'���I��/L�'��&���':��s�.���}3�o����=V���1�o�`�2�0B�߫)1��l�'��#-d�	зշSмY8p߶���A�!�7�&�甓����ST]�j.3>�L�h�QC�v{�6��a���7Mp,r��J��&�t���]�����x�D�M��y"iC��މ��ߍ��U/[�&3�Z�:$���gs��]��1�2&���Hz��X@�O0��,����Hg��~&��eofR��ݦ�Ի`׷$��&���R!�h�eUʣ�=U��!)Ҙ�z�aFP�^��hU�Wec�J��v64U9MJ�0�?vU������Jr`s�A��'�FP�F���KL$!��
L�%?��{A[j�jWd8�%��� 7S�2��gF�g�iH��[IF���Fx���0!&9����Ω�G)��傉6K�8֡;�f-�a1��.J�$�[r�N�As����b�de�SHA���?����/�H���}�� �߸��%F^���!뢵�(���SF�
h�¯�"�ծw�	j@H�(���,b���.{@�&d��$m���̡zίR���`�E�B5�#]��p<fBcg�峂U������}�)plj���]���b�Y��  t)h�E��)�����rL�,bp�����u /<kzh�X�5���狺+�/�}���'�|Q�cQ~���ç�*�G���)즼��njk���X)f�4�j��ͥ��*�P�!�ì������J�=��	%m2q#�(�\����`�ݬ�S�"��:����+�z�����KK��n&J�l� {/�4�̴�A�)����q/JCv����Zs�/��8=m^����B�֝�����J���)��E�^�3]`�F.�<r&2Xm����,1	>��V84�E���s�rW?x���G
.S>;H�o _vbnx�j7l�
��W#��q62��\.�_�$����l�!�/��� ](��AF}^F�z���^� ��a��l�W��ZR����_+>��<����V���u�6>���Ĭ����7���Cz�zT!v��������T��0/�yPu{B�jQ��}���1IXY�l���EP�$���x ZU'3M�����������v|&٤G�IB9(OI�j���q��ָNVP�+*a���xZ$6Y��jQKIP" ������Bw�'�i@��:�B��"�X��d�*8����a˄�l��57yǷܴӺ��X�G�'�O�8�'��h��+5U���`6�6��\��Pi����I�>6�yk�tW6JCv7_��uA��Ml�7r�i�t�u�q���+�O@��"�05'`�4=�?'��f>>�5��ٷd�1���'8�y@y7R��>M��r{�.#Z�R��B5��������`�g��ԗ�-�Ұ�����|n��f�e^�^6�m�\���c,k�dOB�ҊS�F�A�UO'��Yͫ�y`�����k���5��5�~J��to1��~��%J��b�*�� ���R������:�?��f.Y�.�n�z^���\��7�~��~��؝z��6��K�z/��j�'�r�_EU�"�~��Ed[g'�2���q%E����4�(%���l$�6ga��(�,P�3"'�Ԏñ�v^�:فٴ���v�=�γ	N�+�Em};�f:�L4������rɼ���.Kz��	ED�
�)��+�*�vv�%�yKIH�>=���{��UUU�$���ܮ�LB����8��7=f�qEc�|��>d*j$^��'Λ{�DE�N���D���7Fxi��j�G�qa�g
��J+��3Pǝ��w}��,1#�D2ܺo
�np��@ǟ�<�f��@ɥ��`��~�)KVI���n�$m���O�|�����wuΛ�cÖ�
�=,��{�<72����>?4g���ɂa����!p}׳][:ܼ���\[���{�&���N_ �\�@Z����3��U��l�������_��-L�Ԥ�`44{ �,�9���w�&��Ia�g��#��v�?_�-�ŅxhC��7MA��*.���� �1>��Ū���7�����M�3j�7[��Nq��Rv7�$�`��1R��ZR��DM@����5�l�D.z�V��BW�F�.,���25}O7a"�;���`pwMF��g ��؆��`�uD���ct�}��n�`��׹�^,�w������tSE%�V��l2�/hn�(�EY`�`-B��(�Wj����+W�8`����.�Xzo~Ǚ�(�@a��Hq:,�w�Wl������71�����%�(ғP�ΐ�P?�+հ$��*P# �R�&�?��I���b�$��Q�	�u��2�Վ����5p��=F�ʧM���F�y�/��]�����"����	�rCb6h��@%0����: /-�͑f�g��n���c{��2=�7v��������0
�1U+os�|�%nf�[˒pP6i.s�W`rl.�ѱ@���8��kFa�~�y�`Y-�R���ҷ�f;���^��>�
�}�7M����H��(C��7��a���0�VHIR����-To)��P�G�L���ԫi��)ݑw�em�Wt�� � �����5��I$m"_��ͣ�hb���Ͷ��Y�V��؃�aXA'���H�Ց�8|u�+�VR[5*��	y����>Oj���(������.�H�4��+� ?��~j?�+�(m�M���Z�C�*XY�EBݭ�C�ͭ���fsc���`=ڪ�"�s�Ї�N�/$V�O.��W}���@ѷZ0����g�ef9���UQg��������wԓİ���P�8��oֆo:�9���ז��ZM���nd�������� *P�1�/�L����N������]ϓ�4Dd���}_~�'(z�/�ɝϟ��.���y��/MU�W�����)kC����pu:�j~�N?�`�P5gA)�J�M.U��
��s/	&����-�0��[�/��e,�=&��~8||���Ë���>��p�4D��@,��{�Ϗ��X����w��K���-X����0��^8UL��ɟR4Td��,�w?���KA9*�i�ǌ��ԟJyz>��tr�N�v����)�?�(yb!(��&���K璠�4}����_1h-
�r̼�}'��"z��.SP/K'rky�3����Ʀ�<��������:����\*��9{~���.����}�]|i593K������uшƤ�,�Db*6���\)3��77|p�7s�A�׀�W����KT�v�n�� ��x!��˸3����s��Gy�Wi�/�K
/aHlV�Om�@��Y����Y���P�A��J��I�����E�$��W�M]��~["���&g�rxq��a����4���%����ep�Ǣ�H�h]���Y�t���/�}(����	�_L7z}���{74p�b����~�=���W����Wq�'��w�ͩJ�oǓ@����zv�n^�F!��y2�o�u��� ���u��#d5�7������i����xF���j6I�$��s�p��P`c��W��w���"+R��)M��gH�̈́LEG���	D�t���D�G�@�L�c���(��1a����
�a&|;AbC*A0*���az�P=���ʘ�� c�*�8v������r잟��64(��z�e<R��48�#�H���1��>��`hFAA���������>܀�����z�ca���3^�4��mќ�-�-��&#�5C�\a�I��.>q�5@]-��,�ù����S�
w (������h�������қ�M� 9�WT��Ъؿ�S��h�� ^ǲi*z�!�f�:(iB����Uw��38a-�Ik~^�	�v�^�'$����T����U���Aj��ö��
g�b�z+�<@�,�h��N@�e	��M��2ʶh-2&H`U&Kh�X^`��s�ǐ'<�=�x�}af��P�|=h͔��9Ĳ�O�juKHKD�$����_����7Ts��߼͞�.}�r�FP�E. ���Y�vȭO�`���C}��ƥ��z����'�MG(��3���ZO��YI:��T�� +.5_?BQ��mc�1T���Ԁ�
��ȑ��̯�}�=�B��%<�	��?�,8~�Qȑ�^�O%������p.%�38.���$���� i�o��%�҉�G�З��S�������x�̏��S�}��_L��#�S�x�p���} �G$*��XM�8�J��8�;M.�gj86X.ꟳ�4Զ4v?5B�c�$�~�
�r�1� a��O��%t��vC�A���|�l��؇���޶�ބ�t&�H�|l�?�d�.S1/SO���#�XT�����C�Fwp\"vUf�,q�a���QE�u��#�@���uũLu���sG��&
h��1�d�e�/���p#�a����pZ~̥dO:�
/��i)�����!x��D;˱���xv�ի�֤fB�c�=Q[	}�ot?z���;W�N㴓
o3���a_u�jh�f7��h,d,?�S��ݬ�T*�J��%d� ��
�TXZ�T�a���
 x�MkX�m�[{(���G�`D`=���z���/��"+V�`<������;:�u��6���pDP��*=���9К�x�q�(~h��`�ǌ�"k�w�L�fh�CHE9���h�#EEdS+�(��RRɱ�WO?˒�ϗ#�8�����=^����V[�w�+^ʞ�"D�0Q�l���6�!Pz�
~'�����wuh��P�缕`T'Z��$��p.��m0�'G�x�!w��٬9�ɰB�o��o�a�]�ۦZqd,g��C�
أ��֢g�!ԼH"!|~W<��H3�F|�t�nu�̂��N�S���K�/[�7sm���*w7�J˄����w�|ŏ`�����i0�-�3�9��>2���$	Q@��ѥ�OܢIk\U�jJI�k|B���ȏ`�jjx��>=�Axg;�۲W�w���S�.��s���[�ʧ�����_v��jυ���0�ө�k�k$�c%����	6T���?3��rA��aα{I&�[<���(���R�7�	����U�D<��@�*�H����<�r2��ه�8"�%�Iy������/�n))���A�+�=]��&�u�^C�@j�X�\�Xx�M]>j�)%0�I�q��1���a�P�Ҙ�Z)j~�m
�^�<���H�R������zO�1ii �~��:�\lY�9
������7gGlp�q��Ŷ��^�;���l��Z�j<{�ב[n�Y
���0�D	����N<e�R@���?0��8��0�8�8>8��S,TR����gN��ޮ�����%,KPf0�f<(1�&;>��wn�|��q���'9Y;��!:�'��G|�G|�5�#a(Q(:������-�z��������Ûo��[��.��{�g�"KvF'���ʯj�g�g ����~KR%�I{���ɂ�8}��/JI��x�������T����.��QL�=
q�C��M@G���Z��������������v��b�q��U��ni�ZD��݇��	�� s�Yt`)`N-�&�a˴؞J��Q��U}�
�Rv�����c��m90�|�Ň;k���˜3/�*�g��ؿ22}�ee�/&����BEE���9��l�ufj*V��������/�c\�X�*M�T�x��j��Oa�+�:ۺ��qX��D	JL_+N]�"{8:jY��>�KceǺ�d}��]` c$��]�<��A�Y�%a��ҾO�� $�TP]�jV`1{���j+_P)<2B���3��l$�7�'UʨZ�t���W�84w_��$��g��?��>ē<����8_��>;%[�"���(����Ώ`^�:�U)���g��_�`deS;gM�Y�š�<����|2�}JT/����\�_/����)�9>j�"Ƨ���������p� �1�9�5�o���������$�l�څ�?���a���Ow_�����w����7��yvªN��������Wkw��*L�/R~�8��g�.��<�S��bi�∀���S{e���e��xZj���..��|���	���Џ��:��;��'k�Cϗsx~@�n����.��i����Tnu���k�]�'Yk��n����0`n��T��4�J*��r�T^�}MG/؁�u�@����i`H�y`!Aqp"#qm���_��N��N饌��v��_�t��t��;S�u�� �M{"��y��sJ�I^�� ���"�N�ۨ���7�L�]|7/���#����.�s��~ڟ,p�7��=4�y��gu*����$�8�?ȹ��b�,�&�mvW?�v�����b�sֳ�U�N^~��Td�ig:c�t�f8"�b����كq����7����/ai�ֲ�-�H�6��O\�(�F��I���aƞFa���x�!��3?�
D��G��� [�pj@��U2~[�0��Ί"��V���$��<	��J?����j�j�Bc[͐�炃��f�s�7>�;df����5ٮh?"�5k�� ,�rHAĘ��\����pGD~?y��pBP�[;�۫���SԶPZ��h�E1�)"����̋:�;�Y��%����Z�l�*C���ǥW� 睭��x��.?��~�s�o���f-V�Q`F��b0�S9B/�j-��5F�&<B`{��XR��Dｴ��*lVV?5��j��=/_Uys9cE	EOUK�p�=�O?`����������U�'�t�2��,+엯"А#C2�X6�6!�{�Bi�z����a�n*�1��.�ɕ��2H�E�z�����w��\gI�s������n�n�k��3�V2J��O�&V�, Ϡ��h�gs��~��`\#x��!"���'�?���x{�/��^4:5�P%눅���3ltۗt���3��D�X�[0Ɨ����@&c�}8Xt�rɑ�1ᤣĨ,��$��*)(T���0�p��Q�D�d�|�tɩ�>�(xHcMg��&<�u`[
G_k��JD%��$a�.f�u��a ���ւ�C}��_L16,wUu!�����֢�Ņ4`�Qc�#̪ə�L�T��O�����Db/�y�eo|ג~Գ�8�y��]��>V�|��W?1���z����^�G8�~$�scn���1�ź}�"���^��P\�&�V�u8\�xq��-#�@��Y+��*K��6�$y,�q�3�ؖ^��S��J��dVz���r��ְ0}��n��g%���<&q�2��_�:������;�|���e'�7fd��ߜ:��z������,�q����<�������ø�r��ǭ����6�YyRΡ�fK}���&Rb�SVPO��p�'����c�������_~@�K~�+ߗ5��5�I[(.�(\�}�]���>-v��A�� 7q�"v�֟ιD��|&����^!O]h�hD^�Ɍ�q-l!Y|!�r�!��d�����?�|�&f�-(��xAҽ�b�^�/>�PG�9A����ZG񻡤q��p�=�����k�kW���,���R����x�XN���	//��R`Z��2(N5�X��	�Տcm͔�����-Q����	�����ۙD�CX��qj�����9rh>� ��W,6�ϟD<��s�é����P��m/��V��ԋK�|�>��Jʨ�qBj�����U��B4`0m����������t�;��K0�><m����@!��_�3F�k��4��a��w��y�GN��|�~������Aٵ�Iږ}u�q��]���U{=�/�~A%��J�ɐ'|�9Gڲ�ٳ�ǧ_t6��S��,�.���+X���{�����E�[���{lX�HP����ޕ6�6z�tIRo�D+G
#����a��9�&s$�f}3O��44��� ��wLI�� T���/�/Y?��J Xi�Q9c�l�"��'b႙�b�Ε����\:^#w��������x��7K���:���e����L#
�{	s�E���}�s|��?��fGN��O�]�����N�L>G�Dm�!�c��DS���x���3U4|"J5��2ڌ�F��(U��?������	��0�ܷ=7 ��EQ�����Ì���L�L��Ȃ �&v!.a\Q&�9k^e��rj�0�`%�`j�A��+���������a� �朙1d�� �Xt���F��lp���F�CJ�G�:�V/�"�g8]��x�Lj0�~M�3=��2#��C�1$E��fLA�ɦ[|��M烼�*K���Ґ'��4���z
�MU�ӗ��g�C��
��Jr0-�+�c`��U�qg5��ݴq�bl�1��8,��蘄`�s��#�+���N_�_�T�a�@����9T����H���1΂z��o�@���wv��GQ�e�U��+��;(O����?���(m'����ȴ���ZPh�PwW~&Fu�TǙS�=���ʑA��d�\u(ޟ�
�R}M���� B�O��M4��5��"3HН����1$7��=l���K�n������
k���t��8��K�B�w�C��A���R<+%��[�Kp/�����]39�Y�ޝ�~���ۙ�
���)s�V.{3�/����X�f�%���eOFnf�=6�z��3�x��5Y2h��]7���#�"��w��PZY��Ƒ5���i��k�t���H�(�35~����'��2Ny��F��D�ˢ�m��7�I�2�5ߵv5�B��~ԕ��8�Y������p3�cWq��}*4�=̹��[b�c.PM��h	䨰{��Uh!�o<@����ux�I��#�W��Z/�e��3�IZM"n{�|,����,n���+�D�񓎹�a.�G��q��/MVv�!��xS��N�W �1r�4��0����-���cS����PO��5*�������V��O�`���!�>MOҕ���	�%37x�R��|܄����$"�1���hSWG�W+�)�'�Q՛���khT�5	�yC	��Ǖ�o��7�}�]Ė]0�#Ir��`B+h��Kl}yV<��
�[�x7�/fr�ݙe�$ ΢p���A99��Eb&������
x���ks��~NXC�j�Lg�O�n2�{&Z����O���/��8�$k��z�+�؆�7���7uV�Ga�yd׼��N�����yS��+��*���ys��3	�AM-���ڵ�����Ay ���l$�Pt����x�$h�
]|#&�g��h���:j1����z�)[��#%��4��rF{��oʼ���o^����U�N/9u���T��l{�T�~�zn�zb�~n���_�N1۟��{���:o�;�6V'�c��vxl�|�Q�q�z���׃�����_���^�j�_ma,���I�R�����e���$����@]����D���m���c������RPk&�׳�r��T�: �h�7e�g�K�`��AB!�IO�T�
�LL"u,���}�����S�U��R�%�{��lؾh��/��fH���͝����|��W��A��j���l�K}V�B^�|f�	Y ^�� ��+YFP%��U�(��	��&\�&��D>�n�;84448-W���4����"D���-at��������z���y������v�֡�⠣���5V�i;O�:�J3��*���R�L�����o[�$��[���"���{#��?�k�D|��m����վ&^�aRSQa$� DWx����?@:<嶯C$��%�í|��z�`l�ۖ&�,�[��ۍ���&��ܝ�&�<SPFF�섌��|�!VbF�C��I�j�_�2�.��BM��M�:�n�E+����)�Jov���s�7����~�i҂m��*�>8,��7P��o:�|����R��|����C�X�?�tF��S�Y@Ye��k2��"mF?�O�u�i���*"�G�N_R*�Q=�d�x���L���ol�<��f:w�<_V��g��> ��/���C��i��Q8��i�;�\w6�V۴���5�hW5|{�VY���M����_l�����o"-b�m��&�rnn�A�w���������s�9�����k�9d�	;E��f]�h2P�%�=e'�A��OR��IN��{��F�~,�v��2��ޞ>�Ipο���q$�f�dS-O���iD��	"�MU� #աד>�1~�_~����D���Lx,;.���UOk,-��`݁�I�CF�����#��	(`����PIH�.��/ϭz�,�k�T��p!��.KMV⦫���`�w��2�RX��w�nnn}��J_���c8RY �/N����S4�|�o�B��i��h��J��n��D^F������Cx/"���Sp�qnye!�6�.���@"xA��<h=�@���mmA��0��8��n
�
	��	81��_Ә#<8��ę�:��x�ӹ��Wؙ���/9*�K���\����$��	�j�e;��RȨ������/��4�Ơฌ�~ol�(~�����#@;?{�Α���WrTV7���9dZ_�d7��E���)w�鮼�B����j�7�yհ��ϡ�˳�mY%G��I����Q�EL�d^���x*���9U�%�)H+֩i�**jj�z�{��:�����1�7��P=��{����<�2WS1��a+���G/��u�F����)��]�W �O���y!F���T�Ē���<ٻ٬x��ڨ[$��d�(��ݲ@����D�ӄW���L��9S�n谮���8�қN�0fC5�i>�\���D��x����h�d&bkk����@��?�1���e���QYib���KN�k~���*���[�}��(ne���o��3�Q���hjѤ����¡�R߅��Ɇql�Q5DO�8UK]�����tHR�Ft���Z4�?\|�ը��e��0�2��7�Mm̻m0ʜ�~q��ƈ}f�L��g%�|��;�w���K-ʂ��B�l���^$g���Gj|Aڝ�ŋq�����>4u9��f[�J�Cx ��H��@� 2w�4=u�ؒ�V�~��:x�׹c�%m�{RR����J,����G�mH��������3]��a�3�</�v�NhmR1��ֺ�'�B�G���R0�.��ʮ���s�C�=���L��)����v!&�g����Z�/�/*.8��/=�.���/8�*p.�$�1`[鹁�6�(y�H�ם��d�/��p���o0˥�;���3�M1 =P���}oDe�����7�rS��r���;��+޸ր�X/� ���G�jχ��A.7a����ѱ��a�}9�����Ǌ^�xL�	�nɃ��{���=��nZs��v���~l+� &JF�}w����K�sw���9�z>R5��H�i��e&�Df�!��I�+�m޽ѩ �粗��H���VҰ!B䯞�MB�;�y��Q�6��&1�|.mLYz��/��>|G�yB�)V5���۷Cǃr�E�w���������Q􍭭��=,,S�58t|{xӵ`rg{{{sͳ[CXXX^^�"!?G��v�����#��+�BMK]�������쩤.�S<Ob2F:����D��5"�&b&����6U�rT#`�)Liy{S�2��v�tV�O��|�w!�Ӟ�f�!¯�M�� 	e��j&���é���(�l���c��ǣ���#��{�N?�մԿ�cXf����X|��]0����-L������|�c�y��R�\z1��$�G�����xv6��+�"�c�E�\��������>��c\�%����+m�V�H#nȜ�p6k08߆ǹ�F�9��7HX5{5�<����mz}��.�DKy�@�lrO~������H<��i69����S%Rn�=��I%!�:j��y.͡��.E�{B���6�����z^�g�m���D���Ġ���'���~�X8?�Ϧm[}���Op�-�l��5�\��t���&��Vv��g�L���ϲ�J��дۿ�w��^���kө�\)��)���_/Њ�޷��ya�������I����j��3~�JI�@��y`����#-z3�Byb9(��~-������l^Q�юww���\,����Uh�sЈ(Ӷ�8�����3$D�J�6ː�Rv#c/
��޺�?�����E�3�������k&ir�a~�ˤ���$5���53���X�	�47�gw7��=
��`�%|�-�s�,Ý�dM��ove����AL���e��N�=R��m�r�p�dQsY6fގ���ׄ�z�8}����K�$���a����w]�d=��	qFz����>���8ٳ`�UVQ",eCz��yT�\i���%�kRp056����O#��T5<[+C����5t�Qt�i�Cޓ ���;�kn���c�R��O�űv�P$-Z4���K2iр�l�v�y���ݯ� �a�C�x0k�;l�(� s�I\�曹Y/�Xkֵ/�]�^�pRlӍî��zp��##��|^�<n��XT���
�� �}&�΃Iz�w-��m�)]���T[ �ȿ]�z���04�S:�e�}��u�pOpz�[>|�F�7'>1���ZK����ร��ttp��0�oy�.�G��j�,h�-�8�F�������xTs% �T�G1�Bi�k��ْv�.���q`S֜��X�*&�.����X�B�ӏ�n�M��v��U��Γ���Ӧ�A���+Mz���||����χz��~~U�7���}bjY㯦��5I�j��O~�G�Q7aͤ�����{(�]"h�;��A�rA������v�X�TW�{���	3���*7u����Mz�y�ЂK��W:�EA8?O����{�}
�d���X��?&?C~�~�R�a2p�$v��X�0��63�gN��<�Ts䎾�b˗͡�Z�����1Z���\ί�e?c�_l2u��V?�e�2��odp��&\0��;]��S賕��s�s�[Z_46��n��r]oO��-�+<�g��'[��.��s����!�QI�����x���i}�b���4�35B����v�U�6C��dI���Oq��:�#%�
{�hHƂ\�u'Ø���Y�K���/��F�0Ay	0c���3������L�cU��#�nWO� (�z���i ;���bhB՚r�VT���N�E�WQ5Y���_������?�]>��y�^�f��t��*3���:I~�rӵ����q���>�tg=U���H$�����7s
���:db=�3�yW-�F\��$2j��F̬� D�T�dyj$��*�b���5g��ǳ�
r�l�aF��~��,ԃJ*�Лؼ޷�צP�K3���j���5�NN�D&��LB�32�_T�]�y;U~���?D����J�_�~�U�)gj��|�}>�|�;�ܴ1	8�j�7�W�Y�ɡ`�F=���
݋3�S�;T�[F�tg@�3Q�7�������Հ���EJ�U�m��;��R^s'�Ɵ������:S{�K$mԨz�X �>|��I�Q�Z2�b�`dS��|��'���؅�<�w,Dv������_pT-hjq&P���W��n�E7�Z=��_�O�-���9n{�X�f7Ew���Sq�f�_�7��p�A�(}C���! �h �kjDe���!aMr��{fplf�ofr�U(wFX�\A��C�^٤m[[���*2���]���]վ,D�������%T��׷29:69=�}[�i)s<��z	+lԕV�?�`�IJ*h���&�(��7�n���>tw��$���_>�@�3G��%QU*:�mz&R�=�|=���
}Դ��[�o����ڃn��~��l�ݡ�Tp��k�5�Q�1�ky�(�y5|g�������5����52~�(�A^T������R*�$�b����7ex1�ρ�!�M������m�D�FaB�(�	c�ܺbԀ��,D�~�>��������5�_eڑ�vb�H{�ښ��v�KD�,>bQwP�E�<����.'qi>�Z�:0�s����W��L��S�c8+"�'':���~⾈����Հ�E|@}����R'�gۺ��2��Ik�C?`[�ՙ6�������;w��z��bp��u��=ԭ?gm�+��?�x$x��ъ?\a46�O�wZZ�S�&��KS��\�HϘ������f��G,q���eDBB���+�hMىA��d�������ڲ��Gǅ~���@����a���{R�ҭ�m�O��:;�5"m)��2�Ǯ1=S��9�	a�;��f���n��?��^�6�W�j��'x�����K��,�FS���%vM8��$1E+d�5�y���'�X��?���R�d˰��*8�����c���}z�L����8?|�`����V�8�l���� @ ��DW[Ͽ��σ�y���\��D�[$�἟���ԯּaOp�j�|���-�<(:�>s`Q.E04R�'6C�#�o�gڑ綄Q_�z]��5.�E`Od�/�5V��b�p^�2�f�
A��؎�6n���^�śٰ�9δ{�l��9MV2.�n�G�n��U�E5��8*�X�f���d�.{Z[���qko�Vr�eT,��%�r��O
�@ *%0�[O�TZ�Vt{��a��D^��Q��m��*򍦴�z��ߨ���u)Z�ǀ����r����F��KJ�s��p圾>uC�{��X����}U��x	��,�TBQ��Q~��W���B58jI��j�i��Zf��������O��(v��|mR|oһ�E������أ��~`aK��4A	��� �uq<����1ػ��1��1O�f�qy%��u%.厒��}��?C���3++��~ٴ�ca~���M�O����s+���߬>@�j�abO�{�E����΢T��݈���%�f����M�KLq�H&ϐ����gF��W9�h,����7<�n���C!Ew���dF�2�	bj�����_M��(ZT�rf������5�.Jl0_FA�:i�^ֱ�J��Ъ�ky�8�8b�ʇ#��7���T=�k#A2�:4:�$%�����e]p�s��Cm�/)��*nJ\�\����jɃ,.M*qoL�I�B���<\>��x!��t�L-��Zڨ�9n�M�.΄�s�B;y[.;�R�"������(�cA��G؋��#�h�7s)5�k~m�4u�ZxAuV�d�_V�gg�t���k||�Lu`B+��j���=^Vv�n��>͚�o�{U:	�|��>�98�ڴ����q���Y7�T��U5W�1Խq����v�0?j�_Yp-�r���|�����W4������];(*T��z`�lK�g�`K��\�s�/e�f�A��a�v������yI�P���ьm�Y�|d4o('"���TYE-��o��`����q?����M|6]B�w�bɃ0�z�� ����u�ӊ1�8��Q��$#�����^4,�MhO��r��܌�6{��v��h���������+��u׮F^Hv|ym�h_�
��ņ�MT��o���Ɗ��zz�b\��
Z��M8��`s������vT$(�?}"��I)���n�D-�b`h�(�#�o����J��"�Šf�ǩڂ� ��Z29v�ڶ��
>�u	�?��G�MΦO��'dLjZ�G�6����b�]	TQg�d�Nеe.uW�PI��+~��=��yv肿���Z�Y�L|9�e� K�e��S�*��2S/V�	pf.���<�2֚���D�)�[ 6(T�����$���`x�����K��=IVF!���)`��|�G��$g�&�����,��;�2��tvKI�B���^�:�(�����u6B�iBcm�BA ؝L*��
��F�~���&ܝ��{3��/���[2R��Y�i�*2z���h޽��z,Vx<��@�f�iӉ�P�鲑ك�]QG�������۩��[L�M�0�6�<��nk&�俅V�H��N�T��Ec��63�|R(z¯�H������<�2��v�B�W}yQ��;u?U��V������u1�=QP���m�הЍES��a{	�!og�'Q�R�Zy��S'�4ؘ�]�a����,c&��Q+�\�:S��P�=���e7���J���ڽ��en���@�V��59�j� jAd�kIF��4�5�E�.��OT�2��OF nS$��$������ד7��KvWa��:Oe��������Ч����Zݤ�6�d��0��27�V�����j�N���o�G;�����u���?/0
�8�>kpG��ϋO1����`UQh�Ηa�TQ����=[�KC��++�������,�X;���2ܤ����1����Ȯ�I=ȱ���zv_W���ͯ4����������r�將����e&1N}h���E��p�y�]`<$]�9�c�h&a�	8�dͻ��:(iWW�(�I�4�Gd�YaJjzW�8�4?d���gp�2*�<����{�o��RfT��9|ڸKI�8����O��!�4�@A'��F0g_���OuLT�?�&����pl0ޓ��#�A�MI��1�e����y��1�_���*�1Gױ���c����R��Z�o���%���ϺNq͟1���>ے(�c�{����R'?~d�P�U�j����w3h�:bDS�%�Z�L�(,)G\�E����w���|$�.ϭ�+R�}
nV��Qn#�yq�-�~���lx��>=����������Mv]��N������;�vx4�_M���~��qi�z'�u棅2�D9�KP��+_��?|�`�72���㘄ۨX�j_b\4��y���B��k�q��� ���˜��%D�ՠ8�0�v8�aCf�?%��^������0�wڛ4�ҏG5)�y����s=5	u����1�Vt*��zK��f��̐jhV�F�E>�K6�I6�i3Qp^R0\V���y���s��x��<J���9
{��.��{�~��u [U2 V��?H`r*��h���P�p��^n�%5��E�1*!���Y[��i� u�b�!��&�v.6+�F�.�*�s��;VF�:F����l!�������۳Z���է�E��U�ONn;��ʗ=
4#�ڥ�&�/QPhj�	-:0?��bh�i�*x���o��y=���v�ëp{�a��f�6���`�߆��V_�Ô"Y��"q�Gގs��a�:�$)`%���#3�y�!S��`� e'�Im<���!f��w,��H��UA��$�}ğ�� ����5,�y�[���/�@6"�?����S~5e#��+�z͞���Eu@봙�4�x�//9L�A��%����x^p���U�FN�2��0���E2cY�H�.}�U���e�4(ú���H������fffVVV1�2C��I����ݫj��<��� ��s�f�3B~�W�q���=���K)f��Ʉ�/�C��(V����3t�z3��)� l�,\a0E����yV�.�\���⾚�S����-��)���5
�c��Of�S��5Sx|����$�@�t�Ss��{=F�*����QWj�����$��6X��=�����M��JP]�%�&_hL�Bc�H������.���@��%�b+��b!];�Ȧ��[�k�f¤����qN���
ʑҋ�IP?nH$]+Xy;{h٫,M؎���7rǭ��{�;L�z4r�tz�N�v����%�w;��5��JYmG�\.g�����`�yޮ��$��D}�n����m��s��?���R��ӓ�r��e)�|���i|�,4�6aL�����j�r�X��֋�D�ٮ{雺����G� �A1L��@E>��R¯y+�1��٦��@�s	+\�bJj���)ܦse]o5�ėo�{5�p^Ч��Q��&� VG�TW��-aο����^
�<I��	a�\�{��tقW�Z�^���K�T_�����X5�h.��E��S�9��n��bP�)��{z+y邐�آ��zx^�8��RrgXDFh���b���q�R���v���}�ye���)Je�r���_� ���P `�M���\e�I�0����ۑ��3�����\�1-�oj4�ɡ<���-y,�UcMV�ڋ�cG}�g���_>�3�.��WG=�{�_���w��9�& �.|���8#��qSy0���c������i�@t	��dbO0�thJ�U;U��53\��Us;�����_��՚���\�]`�2�5���+���52pljӺ�j����Y֫0�Q�(���<����)�o����F���c�B��'>����Ns�k6)^o��p%�R0���-:�TVэᇾ�ك���������"G�̝��٫�����t�#�K��������	ʫ�o��M�	���#�ʈR㬐���#�Y�=�4~9�����YVk���م���M��y|G�I82�펰��8M���0���=���yQ�T"������Ě��@��|��I�w˕|Hbg��cV�OD����bdɎ��o�1�n�����M�з�(��X{RУyo����j���ӭ����X�'��La�b�['c�b��3q{@������dÕ���n5����;�wx�^�mnr�vz�z#�� \�8�ۍ�k�F>����W���[�NM?�=��R���w����R��
ɳ����y�ù�T�츤P4DT>�
���ˬ��aO����$�S��HH�ܕ�N ?}�lǶ�h�����]>ΣB���)�e7��&�#��ʻ(����{�ܶf.>LJ�3L�C��Or]$+Z�ǐ/DL��A��4=w�k!��
�ֲ�g�����݌y�2���I�p�A�	N 7ɰ3>s������

���t��z�p�u��8ԇ
sF"�o��[���,f�bU�ԗ쟌}��CB�$�g��6x�$a�A�Ve.\*~��X�oY��62e��k��U��v��vĹ(ǽ*�U�5y|!��S�j��n��Cw9�H]���il�+ak��p슑����6���{Z�J��#���Z��=r�3B�1�Ch['������x��8v��o��$�Q����b_��
�N�L�_�B ��8%�[�Q�~�sJsYi�Ҙ�)�������9���E
7�#�1* `T�J�#�<Ș��(UH��H ���}q�)�3)��H����|���=�lo��K���]�,o'���[�&t)�u� �� �<����#V$���+�b�f��ফ@V|�F>������P_�fEFF�֊��Pb�3IF��
O��[�B�3�,�K�]r��sgA-؈?>�� �W`B�KL(����th�Ul'A�J���i���/L*jD�Ȳ���Nè�C�ռ����c�����u o*���3���xv���	��6�����^J�;T)�~'��k�҂+h�2�����*�Ϸ�Gd]Vg�LU�LX �7s�w|$,�Z���27��MT%���E�����h)�F����x8�����BK�7�$��Z3��vyp$���籡�-��SRLjlr�`Z���ظ��M;pSk���J�K{�#�<ӯ���h����
���Z��1RcQ����i*���X����߾������^:_���y"%�Re�O���a�=~���H�?��_���?�O��K�𦣾���Qgq]#;k��l��>�g��r����z.��zD��ˑ�$W�-��ɑ�TG�B����H�5u!�o����B������I���X����GoW��+S���M�fm]ip������F�L�l'n�D��2e��T���C�T�_��z��$��B6�H?�[j��p���$]7&?r1������|y��aN�R������"�/�1V.&Ǵ��A|¥�^�N�5��'R��=n�$�Ks����b�B	4���7Q�݈
�/s ¤Λ��C<�g 3����<�"�J(�>Y�A֘L���p9�x�p�Z���f�N��0�D�Эc�bK�}4a;#�QO��v�/������D��#�8x
�К���R�$dJV��Z] GJ݂�w�%A�{�+mC�i_�o8�p�ɮo��t�?o�2t}??��oݎ�ݯi�c��x��Ƕ�	�ĝ�1~7���/���Ւ~C�,燮�H��-�� /������Q�����}�Ӽ��� S����!�b�I#�+>/ ����Z�JI����.Iޔ���k?����8׍���|=,!_�j��˴�s.����&���t���rb�,�-��#<OԲ7������3:�S@3eCy�:b9$ /O�Z4���: �ŕ���������M0�#Û#w�D"�������)i�兲�'��Fr�G�����r\N�}��D)��\F�����o=���̈́}JΎ�0� �>�Gˑ���˫�/Z d%[����o���d���ϡ���y�.��a�N���a�b����s����m[P��Bx��vIe�x}��;g7��=�iާD9J�c���ϕ�u%@:MJ�nm��CΗ��0�[���O�y�,��䌬�R0���$B[HBo��ʷF{�k0J����R��/����pl��$�Z��5��v߰��/$/$_֬24h�p|�F^ �ly]1����9�5T��uk���$�T"�x�[}�>�1d��G�sH����4'���B���*��*ۍ:Kf�����l��Bt�hJP��e��WWi��h
>���kIT?�����<qy����ڛqv�u��;0�Ŀ辝c#��,uɓ �L6�zi���3ݶ:��V�k|��	��>�pqYq}]�w�T�}(5	�ݍ�}x�5yu����G)��J�L$��1~�\q�R���u�'� Dì�����0�βơ�z� s���\��U���pn��ɞl"mp9���[6��!��zQB���I�UwBTsE���� [�>D�QTs�<ނ�LJ����9��:�Zk�T_y�!uݧѵ�
К���o�FDK=��;�P�3�����(iۄc���w���*��h�J�Xb�p��q�w Y�ZLJR�S���Mϻ�}l[Z^f#�
�.	������7{���+~U,\��T��illlh�(��ή��s���-dB�RG��3��D ��ոfP�gʈf��~-;48y�r5��ϸ��Dc��ݹ�w���ɇ!�3GA�yR�!@�D<�f��a[��?���cJ��zyXd��E�7z�k�2EM��a-����>&��R<Xۘ$��)�(��UA���}�up�Y�S6��3!����8䞖���}�h���G�gf�"#�����Y����~`t���4%SI��� p�^|��F�����HB#$>�������X���ݚ���5d$`T"��O>���v���ݹ�}k���t�6nzZ)we��;������z�#� �ʣ�E/���v��c����T�J�?����;[�UA��V~t5�'<�!��u*h2��7��(���}��hԮx�;��6oC�9;K�e�6�Vc#G��o�@NC��E0a��y3�ځ�#v�b��Pe�H��	h��c�$�S_�s<�="R��G$�$�JW�f��V������C�ԯ���0���ʣZ���ǖ��.џ�~T"J�'6�`\�q����	��F���G��%�g-���L�f*���^(Y�����X���իSC�h������#��ѪNU�˒���?�a�k��~Ś~��Ȭ�(�O��F,����������ʻG�e����yɾ%����B�U�҄��XY�!C_��jAUO�fH+]�HG��Oٙ�穄L�L(G�{Zޥo"N���]@t�-V7�h��&�!�w���wF�{(�Z��8�'��}�@��\l1�|�1�Q���^ʥ\So �o�[�]x���;�ܘ�"��\�V���|$�.@�u;��6�a+f�(aOh��u��`�����s��(�D�>��e��_l}6�����ʚ!x�>��o_�֘��n�@�zK�Y�tr:Z�Y9�?��giXK�=�]�������1��-�>�<6�dN�ހv�6{���[��-��$�)$,
�yT������Eh�<�
g�-9�Ј�ci�fe{34�s�s����£^n�y��<��rZ����٩r�=ܯ�����?��,����$�V)�n6|�[i�##D?����$ܼ]�vg��EF��mpp��1��уk�9���0�;���pw<�aG^1�oU�S.P&4׊��|�k�#���-q�м^�b�8R�z�C�
]��evj`�>Z�O{���}�F��W��q�mC�̀S��B7}��٢��[2C��vd�6F�_�64g.c��c�F�}/�^o��]zC�Ui���?ت��k�[mY=�9L�_�����-tC�n��fiM�sez���O=s+���I[�I_�3�Z���܆�1�`�D��%P��by�Ծ1�b�nb�Ġ$���sMk��c��Uƥ���e3w��+}"�N:��!���3�����yQgwq�:Jhz���b~ݗu�4�V����/U�mjF�ܼ��x�\wz�$�+�e���m��������1No,���A%�oI���Z����RE���:m7Y[t��/�r궚�������@�����(���ɰ�fR���=FϭN@�)����χ5ֿ�G���W��^،�\[��M�����ȧخ��Q�#e7�u���N}M�oC�k��k��j�k�x����۵��ǽZ����l��w���0_��f<�v><�w0`�w��5���C��r���n�ޖ�5��������J����=/ZQ/��ޠ��rk�Tj����f��)��*?_#�V��y1�W�U"��?}W�f���}���?�:��Spi$����z���#���z�%h�hjQt�)�G�g䙮�������v�T�v3�>���Tg1��$���.�ó��+���k3�h|nnngggbbb�)Al��#���o��Tb�	�7	��W�򬯥{'���˕Y���>6*�U��QAgiW��q䅼�V�J��*��y[��b����׎�1m�4ϖ	���~^p�f�F�V�F[�Y�%,?����5G�f^����"��x��-�^�>x�a��ɴ��(Ϛ��>`�:Kz�Fo��Ldj02�(�4��u��NC�� �Zoe����-O�u	��.-��Pϡw�'�2�=QN�U�o? �pNr�� ���֨%�O�??��l�����iN���C.��-R�DT�B:�\m6?\�,�.N�����fWĂVR�"�4+�AE[c�^΂b-�Oԟ��;�o�f�h�[���c�-Yd{��>�+K���A��?��u�fs�5���.3�o)m�U7�����:�2y�y���"0V�7c���t<bco�}L��+b&[>s�j��/����C?���T��C<GX�����bƕ���Em�A��㝳PA�cwiB�S����6R��#B�Zez�W�5�1}�$��?]�f�g���@-چKR�K�k+ZL�2�ɵ��R?��6S�ǫ����/�:@�ބ�a9!��<ړ�@c������V[3[�B{���Et�,B��s�G�JkFd���� m>%�(8�<�b"����!��c����rdnma}������:���z�fk2��aY)�a�im��z���8��f��v� �l�ô�W��A5�}@@ 	E��6th��R�>T�3�@fҙbk���2��^����u�
%�ϫ�}���.K�����������(�@P�����{9�v����R�m OX��y9˴�0oL`Jf�:7ez$���\?���a���ͫ�/�F�,
��ozE��DO��!?��؅�ߎXM7º6��W��N�Se�%���vR1�Iⶍ�B�ܐJOޢݸ)�.��D��ݤ>	�q��sM��es��Hb�W>c>m��y�!o��c�K&�,���w�茥ݐ�va��O]ߩ>�?%�h��	�L�S�a���65��}���}�"A |d�TH!���%=��gB?�װJ�mj�fSݥ=��I�2������If�}�kcx�������9+����	��_�'��=��a�\�)
��&f�d���-�J�1H��u4���F&}��pҮ2S4ڷ��	_�O�ł�(i���Ƴ��6���7KJ�!ɏ�s��c�DCNߡU<X�3���&�$-��6]��j�Y����+�����~�I�)���)�&���xwg�$e[�B�Ư���*��s�Z��O����bUv���U�k^n�׍5�+�s(�n<ݦ���b�t>;.:O�=�NE{^��WvR�n�2t޺���V|��gkk�nm�bm�Kml��.���^��f���:��B�Z�)���m�By{M�^�W_��̾�	�i���ݒ�mR��`�\r���i z[@�
b:["� HA�j�J�K��p� �[�m���"���_�@���c�	8�xNu뗨AΩ�+k_�~82�Eʮl�s�P��(3��t�N��j�3�Y�\��d�Z>���($��cw�;�\,
�_� ;��}v�E�O�)���Q���p����<Tk-ň���������|~������8e�V�m���ԉi���Ӵ�[i��JPa��E8[f�n�Yl�	��M���������M��+5�D&����j*Q��j6������al�M���l��DTY�nFo�.ϭ�� �H�@p���gǛP�x��}�&�t|��~�_�����w�M�t���ܯ�}�G�V8ߺ_AC���@I�����(�Fw`s�0��^q!���	X@Sj`�V�3��@�i��<*�S�ALxLzT����5������*�Se:p9V�tc��!�/��>]�+H21Lb���3	R6S�e��\1�e�g7(�J�� $\0�J�B.4㰙<���% �lK��\j���s�.g2X&%Z�BBA=�D������O�e��� X�J<G�H"�������߉�'N��<~{�%П�P1�&>FD��S�������H��Є+!���#(�Ԫhzu�&�	��c�ų�	�Z@"�(SӞ">�.�>P��)0��&�t�E���إ���lm�Kޟ���e)�2�#��*�Jc�B�a�\��:\�����f�ӕ��2�D�r�r`�B	��TLU�f�Y|�P��9��g�F��ʽ�ū�'���fp()<w�m@c�z��A�.� �����Gnj��6��'�«�N���Y��>�L���LTj�05���'���x�9[�m)�w5'�.�M]�\|ko���#���{�V�{wz����7�^��p�r�[7 o���y��+M�/6�<�pm����k{Ww߹��էK�2��]�nw_}u���F�����כ.]��;_��\��X83��ۑ�V�ZS��hNIp�g��g9ti���XAf� �]na��y��x���&��9�Ԡ9�h<g���+!���B5`�H�5�0\�)u���XV�TE��B9 �JT#e��r-X�x�Df&�D�REƩ�1��!���U&��i�:�lIXZ�΍3��T<���52�N���3�xi�\�(�*�L�P��5 bj�B:�K&IX��w'k�D�aP��� 6�$�4r�A�4��F�J�V�E�P�?��è�Q�&��4Ȥ�,�J15� �t������u�Ru����Ta���9)�����l�ffjθ���8�_��x}�~���L8j[��Ҧf��4���h ^�e�='7jjP/�P��(�*ЧvQ��p#冿���� ��A�q�� ԇ�W�<�%�%hj@��
- �*�]��/��t<;��jw��l"k�K�}%��lY}��=[��܊�smΝ���������%}�����l�p]�@exm��9C2�s&Ou6W����@q6[Қ&<��U�����������i�'�듷����~m��0QX���I7[5�9q5�	Q*6���%�~������SϿ|�S����sϜ��'���'_�}�e����z9 �d�1�i<Ð��z�*�-7�*?
?�)�k#B��"]U���t'��(Ϝ�={��i�1_�>�N����:���/?�ı�=�w�y.X�gX��$��j�l���Г:<��AL�[ӸMM��e5q�Cf/$Q�o?[��ԓ�ҟ�:躸��4��\ͼ���2 ���lw�&����;7��{���w�?z����K^��s�b�k��n_/�y��;��h��/����W����o+n]��Y-���wn���fɥݼ�����ҵ��鞂�����E�Ee�	IfW�<5\�%)���H
"��ܲ(^U��6Q�`�5��V	��.49D�f��%Y���3.��9�3Uѕ���g�s��&$G��Gf}z�L��M�P��g�G�4 �O 9ƅ�լ��4�j�f)L���l(9畼5a�Nئ�1����K|�U熈��B��Z�N��J�:_t�L�®��o����\�_
�_��^����͓�:�><�����bW|0���� T֠���U`)`�������4x�*�tP���f��in6;4�8�]�n��زk�+ƨ�zG2���������94t��B�n������������������Ǿ�����|��o���w�������/������o~��o]����.Z�(ژ,ؙ�ߙ�ڜH�M�qm�&o��C�����~�j_�Jo�Ro�bO�T{�Xs�;5�������d��j��n.�/�	�lԂ��@�zo�R�i�+� ]�г���!i�g���U3G5��܇�d�����>����;z1��	>AM��*�'������� ����h9�{0�������������%E9�#qk��rY\&��f���J.���tldX�Ӗ��^��]��U��	�9��i�N�-1l5�j�FfJvZ�
sr��$K\tTXh���e2�d:���� X@F�!b� L�`����)��'|O�t��c��=���s/ß|��w�xJE��b�
R�����f��3U���"�)#��������A�����>�S���Ob�YXPn��Z��6�v�����Bb5�85��|�P�T�ь�G
T���^7]�w��n~�� ��r$���LW� 3U�w��.A���{��-�����>�9
�o��� �B=,��w����զ(k`h��B�QCqT=�� h��kwhd�����Q�z_?h��GXm:|H��� ���|���r�.A��@MM y
*�72C��P�4�}����@���4d�:f��5�W86V�?��>�^��T9�[�<Ѽ��~~�����7^�����woܹ�}c,'߾}���k�n��|�Z��������8r�b��ƍ����q�ak�ry�zy�vy�za�jv�p�;��9��:���^�tE��Ԇ�#Q���ȵ)�,��Xvn�8�Z�@��'��kݲ�&��8�$���Y��,4P�4g҅^�Ho���=	 ��n��-3�����p��P��9�`�j�Z3P��+ST�F�C�"�J��%�1�$�8B-2�$j�\%� �"�2^��O
�j�B�U� �̬VFt�Z�N&�r��O�"P)<
�K&rH6�"�,�A��"�BQJEj�D��@�� 2Z�'�fЩt:I���g��P(x&(�@�1)1���	��/O�IF�IА��)��dy�cv	���6��No�3[�;���i��Ϥ�Φp�ܳ>�e�Ёi�{��
ej ��Zp͟�4�U��\��*�- j�� P�����(5!(��A��ڢx5��&o���im<�j�6=T��k�a/q��u��0Q���=� Cg^�h*m��{h@`�Ct�*��4(���������6�=|I �z���5��w}^��������	�5�V���: ԭ�f�s�'P�E��>P��(�����P�W���W�gI��h͐��Qv�kS��HR4�/у%2S�㩷@ٓ����)�:s���-	ܙ��\ř9x�m�2�R[�%uN�����s �6v��[�V��*S�������e̶��1��t��g��'�=�̳O<���^x�g/���x:��$?� K��bE����s�Ǟ����)�(�$����r�}������x�]M�������/��ذ��j�RT�S��
���K��c���S��N{�姟y�ɟ�=�4�������2l:Az�47Z�³ihIj�UC�jHH�'-%YKu��V%Ţ�'x�ᒰpi�ݜT���_k�w Q�gӯ������,&�-�/m��<�{�r��׊^�^����7nܹ�~eǹ�b�ZJ9��}u������[ٗϵ~��з_�泉�}��_����^�Ur~7gc5oc-k5{m1kq����i�������:2��,y�����������Uj�$+R�%*����J�b����Qm��>I�5R@�"v����8E�NIG�ʚ�TEw��'C�3Bs�@�P�d!S;���s4nG5͡��y�A����"R&S����35c��td,M3�jXp��TKQ���N�'��6I�s�e:�*�q�Ÿ�a���ɔo
ķ��$�<�2�tC8�����/v��;m��|Z?;:�U�e��5+���~A�5���  �d������Ò;b3*���tЂf) �D@z?=3A���� �|0qC�c(�l�_qN��)�����|16���������վ��z~�oodx��{uxxyxxidxyt�oj`��ۯ��������~����՗���O߻qichq�fq�du15�3;3�[㩛�)ۣ�[�Nhj6���Y���:}m}������{o�k͟�j=7����r&d�ݴ�ʻ�;�1�|�u�< hP����ǩ�+�����fj���A�s�!�)�K�iV�=�݅����Ɯ��Xq�����<�F��H�
1�\,PH�����u*y�Abt$%�:m9���9��y`���V3S�3R�i��d��n�O��I����� d���ʊ9�`_�)&"ԨU���,�a��g�)�k�a
����{*������N������/aN�D�9�8�:�$����l2b�����fh���>9Z�b��L(!��������jU$RE��f�Ų����@��{��K8QwO�
�8N42��h7�<Q��*5Δ�'J�L�A��t �V n��|oa/A�]�A�^�����CS���ep.tG��	��{
�CA< ^��@�r?Sc�z�CuM�w2S�}E���,����)���h��:�hYHo���4|�=mu�fc�kmcxi{���/�w��'o�����^��sm��^���+[��s��c-K�`ٴ0 �������ڵ5{f}j�����u��n��i���<�;x�������������������8�En�Y�EV`��[�y���(rI4�2�\�ojj��5	4��X�5f���ejPA�i`����=`�
j�@e�
>�a$�+3 ܆k���'0��bj��5��*uO9bjFkB�"zJ"J��Y1r�Y�dR�T�ke�55Z�J�RT�LnV+��Z/S#d�a�G�p($6��" \�1�B�]� `[4Ź?��Ѧ�O��i$�����B6�F�cO��v�Į�KELM�C�`�6&1[m�V;��h�����PS�i��O����f�X�)k��x�Oks�Uy ���(^;��djAՌ��9
TӌW� gj�]��'��gP�
`�>�T�< �,����Cm`{�#|�p� ��������
 V!���@���� ��9LӠt���3��)\@k�L��td��fKz��Ïvm;��Ƚ��#m����(۳䨩�O�jjJl��daY���!+r��R�YV�=V����>���c/�a�}	�_Ƽx,�����cԗ}��8�?A{
�|9P�b��&��PBOL�Sh.�
�'(�A"���$�;�:s�]����VknKLJ�24�.���ɏ�	N�O��02Nz�$����_|慗�|�﹧�~�U��!9Y����G�2Cæ�ٵL��nӒZ�SC�k�V5բfZ���Pi\�>.%*�6'g�9m�#q�ݱ9�wg�r~�vy-��V��M��U��eץ������ߩ}�N�T�u��իe�\.�}���լ��/�߾Zz�r��%�.�]�Xz�|��˕�.������//���ol��l�n-��g����5杩�k�+��v�B6�3V�dF�D�q��xYU��&N\/�K7X��I�&�� ܎��u8$g�ҳɲN��+Eѓ��MW�s����`�0���gj�u�wG��.�AL ���65cnG3�����N�k �i�4`2E3��_��c�+�-�dO-� �^�0����d�5��q�ɼ�a��^����`	o��W���A�����=?�Q�gzBe�1kw����Ɠ�ӈ����4�XO;�=��_ܦ/,���Gl�]�Gs:h�g��,?��	"�"������,�2��n�;<ɮP�#�m��[�E���9�Jf�����zwd�Vύ��+���#+##ˣ�PFz?A`��~����w��7�������ߺr~cpy�~y�by�p}�`{�`w6gg:ss"mk,u{<ekԁ����$hj `,��¯-���/��߬�w�vg�:\-�k�mtGl�E��zW�Vo��`�����9�-hP~T��T�>X ���ދ�t�U3^��F^��ȇKd���bu_����Кk��4f�I������0�
�A)�)�:�ԠQ��
�Vf��D�&�F%�� �]��gV� 
)�ӚhK�sٓ `5�i�m2S������즺����������'*�Nn��m:�Y��0��0�t2�������~� _@�ω ߓ��x��D�S4�S��S��2�I3�7I�M�ҵA��L�o����L�}25�3i�n��O`	}���}s���B-45Ȭ[n#s�����=��Q���A~#Я�C�*	/����Aۀ����nZ�Ss ������
z�B5��!��n��45�%�����BSWQ�D[��H��T��|�����ю����ަ��*Ke�1�.H��*Dqv��j�|��(��T�ITR���9�����;�+�ڢ
SSZ�[�S;��z;�Gz���*ϖu7�6�g�$��Yr��m!��!VkѸ���I�\�8�"̏cDS���e1��x��L�fj,��$z���45��b�h`泥L�
>+(k����5v��A�4(�ڡj�`�z�Z�_��Ԏք�TE��DT8�y�
{��mj$*�L.Rʄ
�X�;y�ij4
%�i4Z�N�W�C���.L�1(��E,��A�����.�̡�XT�ȣÜI\��ρ����â�4
v����g0��	
����H�'!W)�Hy!�"�a�Ĵ(N�K]���O���uVvM"�j7w35�&;�Å��T�:���
���jPYs���vP�7��|����:�u�cU ��-�W3�r�C�Z:
O;�W3��/����5@PG3V�<l��S�	�aw�&�l�a�Qx�A@O
�<*�W@�W� =ԡx������ujd �Jţ�܊�{�f�x�L�'_љ#mK4�p�\��T^G��@#�Zz��-25G��Cd��W��*v�K�B�����w��,K�6D+gѨ�A��@��'	�N�}�y�D�c��u,H�c(lyT�*�B].�*�DU�-!����� ar���0f蓫�2�xa�$�U�X�R/
˒�f��v� �"����� ��'?�<y��K�'�:q��	Բ�Q��(̎��G+2C.=+Y�8�t��d��}S��a%��0Yl�:�bN,t��)Oi��7;��3���\�,�s��ͫ`�~i͵��y~���v��B��|��\��l��c~<ir0n����Fӛ7;�}��������/��b���Zo^�y���Ŋ�լɱ����ђ�������֬������3U���Č�X�91Ig�W:����)��VYdUq�75�v��f(��i�3�n4}�J4��AW��45�����x�n*G35^ɚ�TͼS�h�,D�WB$zю�NȾ���#�P(����L������ߦ��`)�����l��e/v��pNn(k<4��X9�̚������l��	�~�_ܪ�'t4�~�%_̼o0d���hS��"@M3��4�9�B�l�[<	`�#le*�\D������?�}ct����ɱ݉������ѕ17�C���淿��������ͷ���������_�pq}p}�is�fi$}"w�`o.w:{k2}{<mg,m{$y{d_�xv��i�m06es��������Θ�<�p�|�͸;{n(~�'r��X�[9r��h��*Ss�#���� �L�Q�jƋ�R�h�b�H9T�.3����̵��x���S2CT�p�4ܠ
5h�M��0sd�	,c�\��t�#�au$%X⢓�c�	���8�%�8���6K�Ӗ�l�2S���Sr2R����������LkScmUYQ~V��b��Tr�F!��&�����t88$��d��)���ߗ�C8�8��Y�;a��Yĸ45!S�����h����*Sӑ*9�.�45}�pA��z�/F4�E�}SSf�.7B��_��x5��AM͏��:  ��IDAT/S����Y�������<�a{x4��SX
�����2��15&�g9O�� c-�4 xB��A�<�& �mj��4��GdjBfk�K#��b���ݵ��RKy���6')=Μ&URT\��(�������z���	~,r��ǎ�����#��k���>̠�q��c�3q9V�A�Q�4ۇO�0�/D!׸J3��	���y�̲ԴB����MITd%Hr�y���xva�8�X�?*SS�Ą�<��>�.��x:��L��x���vx�~�^ #�Vk�MM�z�R?V
MM]��Т��J#TB�L�����/�����%J�L�T4Z��j4���Q&CL�)�l�i�r�B��pX1���a��l:��ՀK=
�h����hj���wM�J%��AA~�)��˔�x2>S̡Iy%���eDʓ50S����8���+��� �LM������eG2猋�9T������^��PSs���/k�U��@S�v4���^���KРx5���L�g�:��J�a35��Cw��A5����sӡ���Ú����V�r <8t�_�a�P)�ޘ�Au���^N�{�z/�Ԍ��o��=$p[��5�ߞ!<�-�ʕ��4 �4 K�ɀ%�4�55�LM�K�ʚZʚj���)w
���87I�eQ�b�Qf%�I9y��g�?���?=���q�I�ҏnd����rqL	/����-d�Ǘ�w�|0t����K�c2{G�2�'�0ErcBŰ�aڔ�.�T�f�	��`�d3MY$e2^f��RX���č��
?,����C��4�������iv�$��uj����&z��Q`����)�)%�ygk
��d�tg-�nM6�~���[��i{�v��Wjo^��y���e@õ�5�vj/�6\9Wy�jw�h}�2�m�s�d�O�޼<��'�BƧ[����������ݼѶ�ݰ�Ҽ�޹�ݽ�ڱ:�8;\;�Uz�.�,3!%:*NkI�:թ���hqv�(?F\� �JT<�L������ @}w��;M֓.��P@_�������<=`<W?�k�B�5�و�A
��Ը��6�R�j1\�bmj;2�9�<�z�D�J�ޤ3n1�7�̛l�m>�5��:��q1���_�(S���n��5��f����	?�40S���OGs?S�� ��Y�á�f5 ���]�� �DS���A4���,`M3��-��+4�K Xa񗙼U�`A V+��[u���t�9<xkx������������������������s�?~����w���o�����9washs�us�n~8we<wk&o.ww&kk2}k,uk̵=��q �X�5�jf;"�M�|e.k�7��\6�n^=���݇���5�����9
ϧ��/��9
T�x1U�-S�(F���U���a���J�����~�I����F��Ó�cc�,q�Nk"�/�N�f����H-�ˮ()�./)�͂��e��f��M��)Yi.P[ۛ:Z��+K�@��562,̤7��!- '	����K�B�}���~=����445$��T��4ߗ>Ǥ�h�&C������U��L�R�]��r5�ڡ|�pޑ����`�l? ��S���Ԭ���2� �b�g�2⮏�S�=�1������x�`�+S�u�BA}���A��{��R�h)X�����WČW'��غK
����Y�2��N����'��??��?���Ϟ�����|6��O�b�2SF%�T� ����%�|)�y���Q2R
�-�鱎<�1)\��*��|r0�H�8��$�DBOj���	f@x�1&V�/K��g&�s��	��8zI4�8sT��6�Vo�� �'��<X���f��[Р���'c��J�p�z�J�W��ЎՄW"���2MEIj�Y��e"�D���<��{?�45&�>���a��F#ዸ,�����<&�ˠr舩�tT�@;V����^�t*���3X`�t��h4"�	�=E!`��T��p�bM!d��X==�[b�W'���-)����a�7[鈩�3[�V\�[��v���� upa��O���n��ej<�
������L�#05�p�=� V�j�� �X����p@x
�,P:
l��@%� <��A�Nw�{>h^@��Ԡ�/5�Ńgj�[K�F:s�g�%H:&O�2�_	7u��`%XK�䮩��ej\�Cd��[�֦I*]�B�8�"M�Wƅˍ:�X*!2x��֝�j_����>�<�bʗ�[�9�Nn|-��]ň�+{e���q��g���c�������1����w����7[6����W�����ݏ�_��ݍ.�9�,��Ob�9��)D�#����OsO�Sq8��#0)�qzE�Z�4�S����P�j�]EI��,*�EK�i�6-bj�Z��$����l.W\J�+��0����Uc�K�i�n�k�17V��+B*͵���|y~��4_]����2�G�T$�4Xۚ�R����N�"/�\Vd*)�(Ih���KikM���).�+-�UU;k�\�59����Ҝ�lgBZ�%5ё�L�t&ғ��I��DeN�4/ZT'.O�<�L�AG6��)�R��i2/Y@�6^�h��5#9� 5H�|�x� V�|M�~"� �����L�x�zޢ\��/�ū:����-f�i{T2jj�35,�M.���ƺN�_"�����a�e���۾+k�>P /G���{�7h3�	jjP}��v a;��@X�GL"k�3=��	ˁxD�`qZ�f>�52B�
�����E2s��^�q�K��7g���Dng��n�{s�����������񱍉����1��x���R���?|����w���~�ه��9wysx{�mg�~�?ky${{*ow6oם�AL�H��X��("k����hg;"A*�o2�d��Ά�+���f�7j�;b��t��v�����G���O/�|��'���O�^��35�A� ��>�4�Y)Cn��*�5�#UQg
�j��ى��(iR����F���ᶄ�d+�c`X&�aMw9Ғ�.{��3S���K
r�ʊj*[j��k*J+K�J�
s�r3�`������ʲ��z@cmh����ب�pp�o����C#<`B�:�F�������`|�!����C�;E�=A�}�����x:�ǩ���t���65��ԜI��M�����,�}���|�P�z(Wy(�Ԍ頦���25G����� �Vx.��W�����o��y@O����(��9���1�j���]����ךf����U��� ��ctcej�¦�쓵��t�=�m���,�t���S��O�A41�!%��x2?�-"�e4�����yR*��!�K�YLa��������֮���� O���h>�S�1�^��ߧ��~�ٗ~v���@�I�������K'��1��f�-Z�䂇��x^��W��*���'SSga�%�<;@�X���~�v����sT��-¼-�V���Ȉ��	
�T��+�{�C[���V��$�T�Bdb2߶\�Gt�}��F�R��Qa᱑Q���ĘHH|Txd�ѠV��"!�)`3PM�8*���N&0A�F�R � OS��&&��D�~:�Ԑp�\E�a��T)����C��X=5�[�$����2��O�6'�ɂ� 2`��j������NvG2�3VM����/YsS���v���	�7S�z?��� ��9�P ��<�{փU(e	kj`c����
T���VQ%qh.e�3����J�Z�޻�:�=��Ԍަ��L��
P�@Q�Y�;�	r����25�)B/Y}Mc��!]V�"-�K�,RW�:6\��*�!�|M(SEV&���@y�q��P0��R��Q��/ m���o#��/����t�7��j��M����v��~������3�~=�ƿo������3����[��]�0{�Fb�Zx��!D���Jh`DUЌa�q��X ��b2�j�<L-�V	�:�C˱��6%١&۔�iP����۴��ݦ�i9�����kv^jzI��,7�,'�$�\�S[j.�Sg���Ru��t/1�b�&���C�T��\�S$�c����:����?�$?A'���(�FJ��O*��J�Ň�~��}���1<��Q�m���lknnE[[CoW�`okϙ��ڢҜ��ؘH�#N�a��YI�Xin�� F�t�zD�(h<��;U	�IS��ˡ�����d(3U�LO�ȴPP� s4����|�D�q"�0���TO�����P�^���nH��|���K"@Ss�F�Ig\�ӯ17X��\�M
��v!����4��OAs����)h�*������m�V0�*/A��?n�X��Q6���F0	N�j��K�� A����/�5�"�4��5�D�<�9Oe-�9�L�����f�ܪ�zo������##�Fw'Ʒ''�&&�'F7ƆS545���������_������W�_��Y�؜���M_�\��ٙɆ��l��և;�ɻc�;�ߏ+e�޸��k4��@�o$η���MHϦ��Ș�w�yZl3��K�>��}��~.ۣ@�H��Kgj�G /F�T�2U�.���]�xM�peD{��2E�cQ��HQJG�19!<���g��08��l�:m� 4��d�8s3�J
r��Kk�Zjۚ���k+�*J
���ܬ����"P	�6�T�T���}aB')>�t,q�	1����0@txH��`�(���ޝF�R���� R���0NrOh��� ���a g�Y��l����~�O��~��|Mo�z _3��-h �9
hj�@ � u(��Ǘ����\�� �t�h�'���=A< ^���R�P~4�p�D��9J� �s ^�Pe3U�̒{���Q�f�$j���W�%���#44��D!��NP�<)Y�aIul��.T��r�Z���8#�h(U�dp��)�/���/9��76ǗW��K��2j0���C�R9ADF@�O�S~�cO �0'O����O���S
F��Y�x�pFr$#;�[�į�r+�i�Ѹ�255j��X�g��Q�u�x�oA���h ��)UV����%��R�p�q�<���ܒm.IR��;D.4)d�L.K��C���ԄM1�������P�^� Wo���2p�x:� �qPրz�c`|�O�8�l�L���C��ID<��C�2�x.�"bS��N.ӈ���(N�E\f�ւ[�ik����j�P��h����6��퀩���D�5��xu���v�ej<G��zTР,��F��Ԡx�k ���@	�� P �p�'P@�(����(��<����.h{XW�}���A�B+q(����}�������P5M���i�s�W-@�̡x��љ�׌�#Tր%(�R��D+�Y��1E�)k�����TI�KZ��ZUi]|��h6�`I��4�1��v%�"�v%k����Z����+�ș�0w��/�v�*]��j����1��Ҧ�/��*w�9?o��/�[�.P��Y��?t��������/jw>����v�W�����,c�NH�<k@�������G�LP���T�D*V��(�آ�t��q��)Zj���(��ƪ!AS8͢�peunrMqVEEA^q�=��f�9�I1�0#ݤ%k$������'��g	�Ǟ|��'�'{���^|�����Ӊ����Ǟz��ˁ����29m��Xu\Q(x���{���~��c���??�d ��*�ⲳR�2�ҭ)��	!W�";A���ȊgE���q�G�����SӀ�])r��5��/M>����f�ᝧ���h��t��B�d�q"G?���NV/GI7��u5C���v9�*i��?Ot�SC��R�Wh�k�m6��zC�������b`��Xͮ?v7�sW�l����P��f/�p.���!��H;X"�K֠�/V}���W�qkxD��6�I��&�����bIh�fCX�>��`H��Y�� :`��Ț)eO��0��5�p�/�
�5V�^�,��獁��CC7��/�O�MNlO�o�{���~�%45�|��7�BL���?|��'�z�����R��\�DW��@��x��L��d��x��p���sw,�PS
sg�Vz�V�����͵�Vφn�F�Aj�u��6�B�� ��/;�ɏ*S���Z��D���*S3R�<��2�0�Ŗ'*ьW�UD��ʜ��$eZ�29F�JIM�J�ƥ9�9�.GR42�
�����@��0������������������������
�W��T�U��V�A��\_�PS	6�J�I
ڟ�d;8]�{�bhj �^ߤS+�"������L
��&��qj8�>B���-�'��9FZ������=���O��#Uc5`	�MO�{��#25�Ԡc	S�e(e�}����w��55G�����<�'h��kwT�ʏ���i �s��dj<�N�1��T�<��	��	ajBǫ,���m9qJ���g��4l��<>^ !��4����b_N���-[�f�5��
)U,���t;8<BA��*�LK��h����牴S4�?[��K<�+�sx����^~�'Ox|*��DЩgB8V3=915�VA��W��(�&���M�45�3G��}����|Jt��pT��=�7#e���@���y�A&�ϖ���|Ck��آ��92F�\��"C̈D��P<M�^�	3��@M\|BLt\T8�n�eD�Q��K�<T����F�S�8

p�?hj`K�Π��.�3��L�/>8�J���D!����
Q�F��͈X��I�j��)Y���7&1i���ʄ��"��;��N�AS
h���x�4V�'�O;�im<�ʃ�%hP��}�?h��s+*k�<\�f��4|�ԀJ(kP�
`fm	���ex������#(�UP	��A��8��4Po�O*OSM���A5MW�n=*e������W�. (_ໃv��~���e��5���z;�>YX�,)��
�,{�-1"42���*J(>k���X�����k�K��L��>��k�ä��Rf>*���t�ی�_����]��:�1����g�}\���ҍ�j����·��kˌ�w��>H�z's��_Vl���s䵤�K�u���3}�/+4�����r�ƤRD�d�Į�;4�d-=�@K�m��D9&A��25�pe�N���	7juJ&�D%�?��ĩ�O��<����ߓ�O���{��Ǟ{�?ߗqX?
şJ=��|��4{��}*��� _�I�0ػu��������ܠ��`�x=��3�>x�ɧ{��gO=��O>q�Xd�Z�0�X�j�{_�%ώ�fE
��y�тG��9L� f�Ёi����xџ��K�@a C	��� 3v��PS3]h��7Mg������Z�dG+�V��=�l����ǝ#��~�PW(��T*2�0�}G�H��	�<�}:h��eg�8�����@Y�l�"�ǐ.`�q��8�.�}�5�35�����dO~ص �FqC��R�q�-���,b��	ڟ��4nS��G4�1��NbɀY2c������D��bB.[��|��콎3��w\��}uz���������񭉱}S��w_��/��ï���W������4.OVL�����.�flNf��d!Lf�L����
�2�=�K�q�]� PX�MX�lZV�#׻��$ܫgC����ft���	u7��g�Rf�#d�L(
�Yn5�VPXl�{��k`{�
ZB�bj ;N�Q�g�?��:�l�}������At����:V�-S�(��倱�H�|�L5R�,3���u�)p��NҤ'R-a��,�%3Ŗ�ڏ�@@9�=�SvzJANf~vFanVEIaS]u����������������ڪ����ƺ��P m��Kښ�����t���8?N�{H��.{�40Vn�CZ�J�c�{w>��cR9"��������@99(����Su��PFA9?�g
���؄/1��$rm�+�>		׀r�����C��d�zs�}���<u�| ���Tp8�B-� ����5�3A̟�T�0]���x�����<��x}M9����^�^���5/����_��9�7/��(�p�á��q�#9J+�E� 0M3YipO׍�~/���<Vj-1��.�[�)�.M��b4�XO��c^�~�) h�bC�L"��|%�#�C%&7�0iH�,4B��ED����r@Ml�>2F��qy""��ϑ���Hgrx������L����Ǟ{���O��~���s�>/3p>
�x1%��Æ#
F��b�5��P�N�T'ҪU4�UX[]���w'��"����]��/Pܛ�/V�H��[�B�8mq�C�s�Ur����5��ͬ�eME�M6{d�Z�w�����(��&�3P�c��R�0pX	�"6U���z��<��L��d�Mĭ�Mh�$�K�9��H�L�e�>��s��t��ǒ���=��(A$A�B	� �DA�m������������؊<�F�Č� `��q�i�D1�uf$����]����#���a
A5b�w��n��׏�O:���ԩ}Z	B���������V��7f����Ӂ#� P`ǧ nЋϬ4I4�ih��~����Q#���I%��i�E����"E^�x�g��9��1�{��Dq�CAhv
?H+��������E�p�38����N��Y��(N"�D]Y���Q�q���6,��@`I��O�b�%��\��ꃉ��ńY)�� � �0��Tē�(j�L���Diq��Z�]�G4	q- )��N�4B�,�N�!��Q �)�k��ake����=Sț�^V|F�z0��jv�>+��d�` ]f�D�Z}�5�q�_\
\5�԰����>�Y�p���~h7
��	;��oO�s�P�c��(�o@�9�(��y��Ͷ(xM�>��t�G�U��#/�;�4)V���y��M��s�e�[��~����5l���������ouK�(+�G�z�Y'�vׇ��\-�V�<s�(���vB_������{UY�<3`�~lj�%�,8^��lr���8��}E�]��wԂ+�թ�s>M��M���-ɠ���Ԣ����ǇG�~ �?5�\i�m�mv0F��:�]��g[QA�mC��U�~�6>l7�d�v&��MN�O��t�Y�u���5Q�����OF��9�{�W��8<���eN�{��i`n,��,��jr2��~�
�U0"�N"6@��}�� gVf�'(g�)�[��?�� i-�XhT��M� ����lЂPO�������i��q_ͷe��E��E;g��Eb�n,�V�*��}�7a�Y��
'�a���q�k�eo�ӹ��k�}��v9Z���)[����V�W�E8Qh���1R�L$"�C�/-ѿ ^��4Ul֯�o�P9iy9�27���٪�t��{�|f�$�D�tg��ぜ�Bg*���"S����n@�5��̽�Ӧ�K ,+.<Q��6�/�F���2��9�����(p�4�s�;�B��R�M�s��NÉ�7}�'����7�]^]�7�����-��Z* [�P�BŬ�ݷ����V�ϛזo���ޞ�]{X�QY湛�s(j�R���_.�|s���S�*j��'v�6K`(��A�]E&�؉��KBW�<�T�9@'5ڳ�﵊޹I�axR�Z�� 9��];𤀔n�����򆻮턚@L]�k���P������[gk� e[sǡa�?7FQ�I�_�˜��?�r�|��w� ?8D�F	���b�<Ӣ��<�<�<=��~�X{p�[��ш� B3��01�� h[��aj���$f#I��]=	HV�OU�k_,�1��@¶	����H�_��ԂQ��h��eT�	�Z��'ڸ<h�=vg�$Z�ޓ4��c���弾q���l�X�;���I3�dR�����������5�'15���+�=qߡ�3��"=��	gV�MzeU.��(x!&/�;�������15d%�W#�>��7dc�A_"��+V­yKR��ynDZ��� ���7��S�dd�,�`�J}:G��'�&��Dl6��-�"7E��,��{�UѺ�Ь3�3Yb�p$z09�/��݇?������2�b�����^��?b��?�h3�п�˕zywD`�i�3/���e��P@�B(�]�,�#D��.�*:0�"��f[��0a��&5gh夡k���x�@1��M���:0D�)�o "N�Lhr�X&Z����G��ϼ#K�f�_"ڠ���+������O��C���QPn�o�p0.��my|y#��1��*b�H P����
�n`�[��+�=�g�=�_�7�J<R9#V���32�����+r�}>'�Rfr��Hi��	��x�F		��oŎ�𰣖\�U��Ľ�=[qR��~��<�M�Q/�ZP[�S��0��o�c!�|U��s�[ ��x�S>R��=%ŨARZ�H�1�l(�q��qq�h�S" p��_K_"�����jռbV|�B��I��S�Ȃ��,��?c�>/��><��H�6�f���Y`�u�f�T����>O��9���!w�%��������S�t���#�����- �{����VEo�6r�Ǿ��<r���m/��f�b^S��?���<6���t��l�u��4��ڥh���>h[��jh�b����β�+c9��Ąg��I�>H�,��?(W ����hR����O)ʛ�F�Xݷ�P�AÍ�r��� `��bD�g���wC "��¡%������r�G���K�?�d
��F��y���DRF`rV�-��mYz$�u�)Իǹ�{�{�/�}�uS�Td����I�2(1P��kWp���3�K�l�d���J3�L�?��N���#���n�e��D�s��Z��#��3W��`<�
����>ul���E���M�=�0���8|���_��p�	[�L�8_���S���"�l��8����#A��J��9#7�:6���ٷ0��-B,{l=�ix�h�t쿂
���`��08�?�����AS�ž6��>?�F��OpA�RF�{��>�P���v��������.�G�*8�#^|O�@�3�:�4�2�_�j$0F:>�m��%�����=������߁ȧՍ�ㆍ���>>�4��iQ������(���tP��q7��`�W���Ƈp=�i�ZR��
��\��v���Sk�mA�8����߲+��)���i5��<�9{&�l->$�-_�ŠJ��x?Y�'�&?3���^���sUgW{I���o������Xyz8*:��*���X��!Z�bo�E�Ab+kHl��Ms�ŰH�%����<86�2���m^�O5*����2�>���gĨhM��0�e)F@��x�oY��ŕ�������-�I����d�k@i�d��14�0 ���4lw�\�+��9�vh���@j��G����D��~^�X���to��B6V���7Bث�t����Z��;��Z)}�uz#�)�� >YlƛX����-x��9�$�[�M�+G�8�)�>R�M1#���O1�:!��Go�tŎ�l���7%�7C'zD��:|t�y`}=�m]���{�!5Q�A�JS��1?i�P磱qC�G9we�RF��N�,%���E��>��҂�N~l=>\g0�"j�8o�0�\a$����>�[,��AHĚ�cZ��wQ9Y���ՉH�8a�F����=B�Mw�X${�br)ҥa���@/K@`{���ɲKNՌ�P�c4���n�� �E��q@l6��;�PLKx�����:TQ�q�Ə7'i�E�0���H_��DKUo��S�������� ���.�s��A�¬�#@�>����ꝃGD�W��j%WRgW��W�EZ�F��?�?E��_��#�aZ�zK�#&���,�ꉜmu�D�Qjӈ���ǽ.MM�K�i��lԥ�e׺`(94�����Z��W����Wb�[��ɹ���P���

{ت:��s�ʊu��N-�}�9}�E�VD�h%t���o��/�ڑ}Q�����?o�q�t�k8�����?#��ggm�m,�)q��v�?�8��@����,���,�S�$���i�m��=��Ff~�fS��B������V3[�!�W]gE{O��r?S<��>�/�v�ꦘ,14c�s��B���Ո���9SQ:�)s��f�oZ��9�L��q��2 ���]�ރ���d1��6\�B?R�.j�1|�f;�W��@��$<cz�
�6O�Į択�Gʋ���į��R��W4%�৙�<By�ۘ=�z��&-�9*2
=���K5VԇB��?�����M�V��Q۫�L������L#Ic�I��'ן������Yt%��1�9U���IPz�-ڛEB �5Ƨw�|�N��W�z,�S���B� fE�PnKC�Vl�2�7�ٚM���#��ɷ5�gm��6�|���)� �{K��)�&'e7��e��%Wl��5G<��/|�_\�s���.x�[q������f=/��;;�FV�3��|����9y�r&�\-y35#���C��ڷ^�K>&7*��f�Φ8Q�~b���O��Jc:�ܑb����&�|{JI�b~���L�$NG�-V�0#Beì��������/���D�:�x�h��H�|ķ�͗�o�Jm^XaJ�jL6jN=bA3��].�QZ#We�m�-��r�6�PE�B�J
G�e-a�H�0iЄ��M�xE���rbƙ�	�����H ;IS�͎寑��3O�����g�UW2ťu�}��"��z�}�q9�N�~�������,һ02SI���O�?ůo�e&�$O>n;R�p��[ ���������G�P'N�n-�g�)��۠�+0W~`�J$dTfN(�`��kx5H+U��3T���0/zq�	�0F���D0p���&�%�@�J�Zٹ��?xA����� ��@��.b�
���c�9H���P��c�2i;��p��?G�;p�V��L���T*�3�����j�u��7)�L��$��R^��S/�y��O��Ԧ�yKi�ޭSXk�'�V"�N�P���XYh�Xm�q������ڡ��Su}+��iFR��oU�鿐e����Tv@�zW����DB��_F�g����9�^�K���;Tt�>���}�H"�f}�軚z0��h���F6ӛ1�t�	m��ӵ�~�o��f��E���/_YP��XEu���gv��@��ӽ�GS��I:`��|�������������o��*2%W\�6��S���L�,r�S�h��㱔�`DD�D�{;�v{��99�9Y$D$;�;��eL�9��ڌ���l�d�Eju�H1?�x��H� R���ҧ+q�`��������G��vx=��Ϣ���yl�|��԰�j�Wֱ'��O�D9P�W�M,��|���	$�wыX�J��wJcG���P�J.,}>���}�֭jwBK���C:DR}>r��K�Ω��f��]��n5���w!g�$C��΋�o	�t����#r���4bҵ1{��\����/�B�C�AV{�o"%fn����ȣ�D�#�����F�jW�z��ϧ�$�,�.��n$ ��h�&��\�ꋗ-a���(9Z�����I�f�R�4�Ö�U2٧��
[L[P�|�Es[F��Ӵ�mI�C��MGJµLB���qc��J��ӖNmO�g�^�]��z8$u�=��?���>7�<��Ʀ����<��{
~��
gz�p�j}��^�Mu��=4���J��JO��I���˒����=�W�fF�	u^W���ʾ,��~����nM��(D��(�8R@����������a���87e�~{����Ź��ɹ�	#�zxw�࣑�X=�G��b:njx�D�74A�r�1r1T���Y���&0���]�$�@����B���i�� 7ٟ=���u4!z�7����E��B�G�m�S�F�p�]\"�ǲ��Y!e��m{���zQ�5�ntRO��	h�
�����o͠5M���Ø��_�ԙg6I��ț�ц�cw&OJO�2Dg�!ÇBϥ�p���&���ku#�P���Q1�C�抵��B뼑(���!��v�����N�^~Z
a+���9sݦ�m�Y�j�e�Bd{l��")�+!،���F��)� =F�*�A�����F���R��JAl.�,KD�[�0�y͝U<@͝�k���>�!>�>��}j���&h�ow;�ñ�*o_�Hn�B.�ᮢj� ����"�O������i.�i�uH7e�e"n�/��
�п|� U4��!���"���`@��H(�Tm�l��q4�PO�N �cg���N]d=a�د�a��@з���S�"�Ȇ�N/&�\];9�:W�y�G�š�H�����l[�{o?FW	<��ce��b!�<I�^��:X���R���v��vx�j2mY��˜*����!i���yј�]E�j�R��u3Q�`1�z�*�z��f~]���d��/?n�3���C��7/��W�b�-^=&���f.��m5��"yЩyq�ms��r0���/��f� 5�s~�qmqU�I9�T���}t����h��H-Q�H�� ��i���u~�c4�`�"��ҷn��}J�ʶ�.�����|���n�}��b��V9qO�Q�iU�.`/sZ�[�T��Z��~e1`˪�*���y;��0��a�n��D�w0%�j�2�䬹mɿ3⮛� JI2(Po��*����{E��bH�d���a���X��=Ic|}�%K�h$[>5kC�{BY��`�x��$o��)�F "i�@(���X�S���P*é�1��ߑo�����5���߾Z��o�����B�!�*���K����u�HV:1d��l�t�~T� K =>�+�H-��;�v3��(}�L�Ҍ~,�BYfgd�WC�i�f�I9�����T9l������
5�8Ltx ��2F�	3�I�����]��� ���|��,,�%�����_ojuB���`(_�R@6������2�߿�z�(�.�Z��J	���g��̭�T-K_�x}!��>ʼ8��ѢO�-yf��i��)%��"����g�ʫ`rnc���+q\V�^���z\����B�����ٵ��s��\�!��N`��G��W�������߀����]�����1.��%jUp�{7�/�����"����O2�~�|J���s)�/���x�e�_��Y�U���o�o.�O~��|m�>�-w<�<߮%��?.O�|��Z�St,�\~;�ꯆ�	�Ź��}���پ|����mg��z�<��w�����Yy���u�cUEL%�pZ�HĤ��㽅mV��bc�/�-�r���t,�k'-|����:j(�C)��;��c� Uz���?H��N��'Ts���W1�R��Ea�6AZ�����L�P�zR9����u�iɷD�j����f���!�9V2��H��0�]��[���#_IEgS�^D�6��G,��X���bY��.�+���G��3;`0f�I-YXȯ�[ߪ��2sM������9��M<U{�'����Y�|�����_��I�ؙ�k����?���c������� ���Z*\�,���bF7�P�'M��<��3�a���I@n��*>On� �pb��_�o�����
%�]��n�+�Fу� �Y���xC���ϋ+�}Ǡ���c��a��&�������{�G{��\z+B>$<�0�<Yq��0���8;����?O��M�y��,����\А=r7��ќ��<U;�R[yT��wM-wK��Ĕ�s��KS�`B���G��n��h<��S�*x�gK�oRՒ��&�����ٕ^�oy� ���|�@X��p�XL��u��b��\s�i#S����o�GZ���	m�PS�h[6
�5��h��L�'��a��ÿSb}���N�I(f�i���!H�V�4-�" !�d�X��H��M[�u�F�mQ.4ǭx�Ą��y�l��h��&@o.�|`
���6���H�����S����9�;׋;+�����p~Lũ����5�Xg��CJ��k��P�Hˮ�h�Rۏ�uy��wڧ�Ңj 1z��*�;���I�b��!�[��#�6>��y~>y��#�#ИŪ����XN���ż\Yծ-^.�t�����z��SS�_�:Ҝ<�6�|{��Λ辛��]�E�m���y-��b���ۃ����Ї���uW��ʯ��Ȃ�'F4���޿����W�)dd_��� 
�O�-4�'���(B(#���7a�F��BrCS|��f�,̍.�(���c1��E�.{0�z��ED�	�����41>P��.�.��K�UGjAD�ԏ�}�,C�:GG˧@a���EM�n�w1@bl�i���%F�6yֳ`�FׅH�R�q����Hf�=�	��8W��7�̎���ve�VQ�HT=;?k����3��s� ��*�/��fb�5�7��p�~�!�lF]j7��"�Baa���a�c|q0����*�&�96Ƭ���9IC��B��%���V$��lKAz�d��z�,UjB1�o3���`����"@)C .XἎ��t�^��WT�R�Н��߾TJ�`:�sp���|Y�B�N��D_ f���K��6�Z7����6-<�U�X�Xp��Qh��\q��!�w����.=��H͓���A�'u� +b�(ؠO&�gu�;)T�wo
�#�:[>�(�}��{L���ܵ��F���&�NËQ��v�]����o'׏#�u׉���Y6��w�I ~��zJ{��Y�	j��dd�k�˷��:	n�0̚%L³�W6/�Rjx��d��l~~mzV��Q=Yb����	�rؽ���뱧ѥ����x�|��H�;ܨ9�[�S���@��(����-�t��۽�!񼢖���O�~|�<�Π�#w�E��?��']�_�?DQG��P�U'�Vb�8���:~0�.�]�n@<�z����(�؁�ת���	t��$V��ENO�.נ	�[b.�Kp�|�߳�)w,�$Q���}T���=�tI��)F�A5�Ζ�$� ��S��zB�������|
Ν�dwrSs����Q��m�&�s�afΔ��2��rCPga�"�H��a�W,O7��#b���dj�����ʃ>�y���WA�2���}��/�q�u�zT[���`?��/�I�����=��v�v�Al�6��߾S�B���V�Q^���Zs�G��΅^��Ҫ�6x���swŭ��Ā�^#l,��f@�Մ��OZ2�w�7ί�ם�������$����۴\��)��9V�Ǽ,x�;��N��x�`�|{����B��r4��Ȗ��:;¶��L2�B�O'R�r�v\߅���o�ke���?�X{<\{�)h�|(�������!��dPE�aT �)X~���0�	2϶͵�����c����=�_�2��cW�WJ�O,/=B
�@k/"�������8�e;�`��H���vTM ���h`�2r�T�8QGEñ.|�{��W|��օ@s[c�|�s�>�[�X_���=+�?.�W�����*F��v�$�����
R�U���l6�b��YG�J쀬�L���3=p�pzs�� ?�N�A��AZk ?h�j�����Q����S��	�R�t��9��0��W��H�Og0϶���CR(Pn�s8+�����<8&c]�P���idـ</�jRiF�����K�¶N��CK����c�p�ˍ�aݳ�������j�պ`�~^X�Dt���l6u��|^�x/�z�:��h���Ԣk�i���{�Q0n-(�v����`�������s]P{p��f�}��/CIv�˺.O}�I��w��.c��w��b�Hc��$f�ӠuX{���YPD1a�R�S�0�lW�e����"cħSr ��w��:�ҭ+�p�i��2[��_���@���:�IU�C#�:$�������#/^���eju*��Ӟ��
!�J�K���G������F5��9F��y��s:f�Ś�	X<N�:��y
l�A��l���,�G��z��~�[�Y%If��C��;B�ޜ�� O%� ؛�A�"
U@�}�fӝ+LJz���}t�D����T��C�,.Z�M�x6��Iϧ6��*���ň��E�	���([V������,�R|�+H��f�����_�k�1�Ĺ	kD��2A��Q(�@�s���	�(���@8-@�� µk"���{-c��֞��&4WO��*��:)F�������S��o��7�z�;	d}��{t���
�����$!�� ���9�zÿ�D,ш��y��&p��HG�rKs��k���w�@��^��ta�h����Z��%��r0�I�g�;�r���+���vB�픮�;����X�:���s�G��Kvf ��G���ɇ������)ԅ�3�
��\ݼE7?��Cg��)9 �ï]~��"���>%)ͽ�ZF+���S~��وq����
ѲF�a�ԕU��ܚ��x#!G�e�lG��ۯ�\vp�l!tE����I�ցt�6��T�y7`sW����������V�$�]���pk�]+099�sp~R�U�T�k7F�)��T��N�`Κ��`p ���^w�� �6��ƒ>�f����D9L��F�aP�K^�/Px�����	G����jju
�K\�u�qKGor:i��������S$�'��霡>lW��������l�oҴ��u�h�w�HPձ�]�+������5���P��ۉԾ&�Y�� �����@�9)���NnRM��Xzo,Q"��5zTM���P6��#�v���~�a��+6���};�RA3�����Jw�ה0i~����i�`@��.Fr��uι�s��	�O�,�rLM�Yn,���Gߕ��YAԻ��K3��5
�2�~x������u�͵G�����ݵo�G��?�
�F��?��kP���џ�r���[���J0�}@v���/���|�ex����p�)x����E^-}�4O��A��p�pv�sܴ��j�O��ņ?ʿ~b]?��K4�o_��C��˒�9Հ����=�,P�8|��"ke���Û7�]#��%x���:	���ү`���9@�Y����C�đyh!��ı|6X>�����h�Z�a�ؕ�)��+߸��rn�ʫ��������)#�J�ǩ���QƼLRp-amcD6%���?�Bd�[鬼)��Z�"���* �xhۦ3�☗Jqxc(����,���ɂ�MN�/Ex��Fק.�f�48H-�5��C�k����J�	 �p0��>N��������F��w��Q���S-�m����C�Z�Z�k�k�U:Y������4�<Fqy�7&A����M/W�߷�X~�=?�̡�s��7�&/�
R����jlQ����Uw�k�ݫ<�Bu��m�����
#����ٹL�7��_k[�<݊��|hRg.�^��coRkJ[��"!�{����;=_Z��C�M��e�����11s=f��N�'h��K�T:�+�޽�3�h�Υ3E�P�4~� ��V"B�?�_�i�5���6t�� �_�$-pp*hp�c�C�=��Br����ޓ�˩�i��d���W��5�e~u�%iC���q����_G�IP�7�g���g�;�;\�����wڛ&�:�*��Y�Y�!��_F��8q�\"�_�k��7�!Lc����14����0ڍ*�*�t�u�ҕ�0b�A�/D��21o̸2#qqh�t}�F����1hQ��%��`4���q}V#��)��/F�4�VP�%ط��6����sC~X���H(ʎ6x]���d������롋�9�1�ءֵ`�A���%7c�ԂZ\��i��*���J��o-9 #s^�G.`��f��*.�<A"�����3x+Է�B6=F�<ϯE8�
�"��x�42Ǌ���·�R��Ձ�W�2���R��aX�(K"�a
�ӵa�����߮DbZD8��>uI�z��E,�P�F��7o��n�BTWO�*�#b]�"��qPhpy�$]m��JF֭�y'�\zڦ�n��]�BYNs�<�C˸C����e� WY��}@>�A��D`i�o����'vb�\^��\�o�c"� ,`��]D޾ ���س�1b����m_�p�Yw�+�T�t���W��|��/��e�&������*�j^��&s=�	�V�~��xL��U�k�U�Uug�W8�He���>	��3���W��mK}��~8�J-�u����#"�us����9���L^̜vB�?��C��$4-�C�
Z��,����?fO���Yv���������fꆩ�6)�Yot�+�GŖ��8�>�r�$\�t��sLC�B�%�a)���Ty�s�88��sX�>2�h�
%����&"����rq
l��*j�EhP���z�&BT����{�f�@��g�<!�0���,��r6�`;������d���5���[ʋ+�]�H�O=��Q %���T�/�Z���k__�߫�t.Ļ�H��G�è���`W�'�׺A�Fy�l���kt0�
+�!��a��T��$�q"锠f�]$�q���e�"�XO���_!�%�A��D%�E���$����
9d���L�W���Ǝg��y�����g�.�E��6�sbf�lx�7�o���N..WɎ���x��
i|nX{�]\{{9`X�|6f����r�ۿ����۵o�{��ǚk��n!+6C��O�r��z'j3'�O'rW'��#��|�J4�Y�<�V>�A.�A>�8F4j+d�GX��(������9�H^��@~9$!8�#�Ì�v����Y��=X+{k�{�i;.]t�~ =��Ž.��x-�+jYځ���b�h�D�RQl�DP����!��E#+�d��~Io��"����������Q��R�"Z�� +tH�T����tW�T�f�{E��ļ�jxLmbB�ut���Ź��ݣ�����,�󗞾���錖��I������2� ���JH�# i�1���X��l���W�e���4�m������fx����R�����I��ܿ�28�������s?�e�~L�L�˴y�\�+�&ciG�)�ɫ��F͍%�C'��b�V�j�J���rR��z��EAh��I1�׺|�)@m�"�L5�qR��Zí�jJ��zx�v�i��dqɿ�0��F�Z��O�q�u�QhE�[^������������<�3�7����=ҡs������@����+���eL'��v1L�-�h��޶i'DH.T���|pԚ/Qq�&�So�ᔱ�*"��R8bcA�d�D9��^b��n�a�\^@[V	
�������]6ߦ��v�>W�C�%0t
����*������
k־������tJn>�v�^�Y�y���֪/rZv������c�ԙq|��s��+�S���`�tO���yu�bo�Ü�#�:+��I��h��8�$tf����b��� <?k�8j�x$�m��m��#���LMs���F�k����"��Q0�o�+�4��m�U���2/ DN�ũh�L��a2G��Ӓȣ��i����	L���Z�,��44���	�e���$�I�Q}�v�839��X5R?��s�CY����1cu$,�e���&�y�)IH�;��K�r�&��M���Gl��12����2jV�o~���8T_З`���A�R�1b	�؈�vt�se�^%�����)�9ų��S�L�dcTj�Z5(�����%�ﱮ���0�y�8j\i�/����B�%D{=����C�6�а���Z��b��p�R:+�ȗ�m�u����i0q����>�"�Y����f�,=���Ҽ�׽�΀�-�/e8T9Ȩ3�ʻ��-�G`��f����4�q8���'%�>�ܟ���uL���I��(�d��uK(8�0��X��Z
��,�k�!�l3I��⑷��ǁ�_�����Fڏ��O�ۦ��v3�V�����q��:�%��h6�u�����E�n�;"� ��G�X�}T�O����u����Y$��:��E'��%�E�ݢ1���H�.������;o�/� +���H�E�6}� ���^�ֳ�9{���4�	&�Oe�������z̎�|`���[�>?�D�����D?b²��vg*�wY1�m�2��A��~��wzS[W{;c���,w�2a^s��Ӳ���z!ec��L�]��lA�y}?���I�ZǨmƙ%��{,��RШ\���Nc�	~�j�*�[�ybS%�)[hF�;&�����y�i���i���K)��%|�E���{�	�%E25���e3�pz��q����t�u��mvs�8������O�_�e�ɦnuk�]>][�����.GPK�t���^��P�:�)c�������9f�����\*�T����;��1��U�2\��q���C��7;����*�Դ�*R��m��V�4��Z��-=�'P`V�1ߋ�@�W�A��ݒOŤE���6����k��x-v:��Ɠ��eWu�هWy�Q��(���Y���N��y	ט��7Ƅw��q��� ��~��I��&M�ƨ]������s�N&V�(��,!M��,T�/�+�WZ̅��t�̬/���.�����5��Ь@�Y�?#�����1�����]���w�7F�8h+�X��8��0L.�M/N�1�Lp1,p����}��i���E�c��]�A�Z�}h�է�4���C�|9G$��}k�w˹�7�D��9�1tS��s�d ��-��x����"L�)V���n%���"Z�%�@��Z,�[eϽ1օr��Wz]Ϊ˽�#~зY�M������q!�O�{��!��˝����S�w�OOc�O��ϋkaW#A��_[xBݻþ2�}��������pt���;��%�p�C�<S+��c�?\�rbT� �(�J0x]�x�(SW|R��L�,!H�L�M�Y��Zo�<xC
��<�K9+�+oC���%�=ۮ�	����S�$��ɊA��#�C&x�OiX��#�I��f��<��������������u��u¯�T������CLmum�M5����p�pK��sW��

�`�׹�/F5^^	33��ڧ��Z�d��x���:��J¾�q�mZ���`�M�>�ET K��Ja��-�o4y�t]�f_n!���Lֲ��)�$@��5Ř(�˸����AlGk�M&ǟ��b(���E��[Cý ��䗴�*�Yw}A�zy��8��Q	B�w쿸�
Q��BJ;�$��T�,3͑Dj���� �����؂�.����1&B�>��Z�x��Td�ˠ&��%~I���_:?����:O���Uuux�v�LZl��azXruUn/�U��s��ݻ��*��4Dx��鳻���xW���-���*�הah�a��a `gqJ������������рk��՜��D�w�w���g�|�3kGvڛ%����M���2���ԶI���ȈO�k��Տq!@�� |@=��,RP���ʟ�,���%o��ǘ�J�v�����~g[~�����dD�T�M�N5�/|-�\��R�D�&��*�����"n����*�
�/����bޤy�6�%0=z�t��)�o3ƦĈ1#�4������N�
���DA�m	��b�f��Mc�+�'6�x��~ooV ���'�����d��I��G)jx�p~Q�ZS�&�+�-�}WL�R0|Ս�8ﲛ�^㾙���[x ���&�SD�Gi�h�g�	�Σ$�i8G�|�o���Y�Ts�{3'��JM������	���fMz0�&Z!t��E�^����u4�>rŕ�C��N�-#���^;�WY�c�a�Yn�c4aW9�D/�PG��k���e�Jy B�VN��M���w_Q?Ӧ�C��=��P R�s�NS����r�UnG��<�:y���Y�
�6�-�:N����*��*|���l�g`L�C^���+Sw��j����y�+�T��d2��4$t~r�cq�Ы�L�bF%Q����B_��c�	SҐ�gzf�l�:3�(Ԃx�8$$'u<�[�cb:���te���l��:m½M�+�M�9���R�$�i��<^*��M��t�n%f��Ge!��f��b�,��f��+G�?D��ڏw.�������C4���OS��[����~SI�a�s���k���mwy���Ƿ�����6�>
�8Y�	����Y�ѽp�px�>��0w<�m&�ii�hlnS�$ �ʷDD���9���5��ޖ�)b=��,H>�#��	���:�;}��)[p��) 4΅0u�ix�݄�
La&/i:��̓K�HVc��L�+FBP�5�W=�=?Y3� �-�(t��	�y� x�9�}g��~;��������`B�a ?�a�V�4�e�4y��[��L^�	��	q��$�a�;�?�[�y�1T����<��=A��ɛ��i�u�V�J�3��%u
6��I�������~��X11�����kWxW��I鉮Y$�ߪ�?4�ePo߶����^�;�h�܋(^ܵ@q^�w�"E��wkq����Γɷ����u��5�節s��I�Ф��$C��b�H�Ǯ������k�?��++�>E�%���z/��=�����r���g`z�#1ä8�a�ֿ��Yޞ�ݴ�]���"���f^����YGw�R�yr���;�u�S���yӇ��<����G�v�=��>4K==�6���X}ػtK���&1`���d�n*�jbqk�kV����*�d��$ �d����{2)Z6�����x�{�>>���
TN����8�p�F�ٍ�c�a(���3��ݨK&����À$g��̖�����?�V9U�;8�:B+��R�P8�;�}�G��������אX��ĥص.�*).^:�
C-���b-��o�8J	2X̧��ʾ�|�Q�"���0�^�T߀��	�-��z�l��i#}�rk)2*Dff��8u��9dZ��	x+�-��,�ˀU��2"���ӵ�7+�?ڽ'(}��_5��z��Ob���&�?��AQ�Hscuq'�m��S 4mK�l��Ja���忕�3���׷���mnK(@cN��b=�,�ύv�Ʈ���Y>9�
O�g���	���j��B�Ģ-&l=��Ԛqc*qu*�SL�Xۚr-X�MN.�[u���Z5�O����ߑ^c9�N ��>Y�,�dW.sB�|�u�ΪI����wdz�����Ǻ�6W��515�g[X����nb�md�
����9���[F�SG�6��q���~Tm>�?^��*�agS#H3h!&���6��MC= �ĳC6A����H�@	pl;��R"q׌�����l�>_%L��
�p���i�fʏ�F{;��L�GfR`�C���?�0��Pe��_���8u�)�sȧ�xU��so�P�"$���?�'4�Ҍ;Jߑ᪬�_R�2M*�@��d�ꤷ�k�ȡqC�(v��xrC�S�~��l�ɴ����������?}k�TZ�$kY{VL]��o%?Vc�g���q�L���a����@���dz<�6�ퟰF�����Alw��7�7�)�����s�kl�Ę��58�Ǯ�_~����7��:�Ѓy;�蘆�X����r�����,kQ|��>�!�� }�����Y��j����K��P���ܨ�$�𼴯�� ⮞�T���f� ���Ȕ4[��ȯ|
��8��f��3��s3A���Vv���-�}�B�F<ǢX�M��"�_)����U3$�u3�E����G�"J��sG3�-<Y�$	��R�=}�$Fq��h�$K���d�^~��d/���\\�Ny��Z�>��(��w�p]v�T��Zɡ��_Ro���%'$OΏ �C�Co��΄�'�Q}glu`�d��&L`�����`�:�pY�t���2�x-�vʧ�}/��7r,}����\��Ƕ���Ivu�G��\e����� K��s�~�u��_�i�'Ū���g����N3]�w���N�^ϱ�yݿ/�sҮM���!�<M>�<��gy�|���M��z�?���|�Y�5�h6=n�;[�7n��92x�1"o��=7�m+�"����_zV��bA5}J��(�A�|8<j�[q1��޶��O�P���$��i���[B���+,����]�@��Վ�^y�-��p+���S>�\|GxI���.Y`$IנN��b&�< Sg@�� X����U
G5����YW�}�ќ��\u�X��z�xl9y��h���~�Ns;OKٲ`��0�V��%+�Ç���j����W|x>���R����=�?V�c�L�5�w�X?���=�C�b/��G�G��p�#�k��i/�_�P:c�fM�.�%�������{w�缒@��e:P.F=�R�Q��%��P��	/�����Z����m��4�9}��QB�ܼ���fW�� ;d�pw���#�t%�t"r�Hbf���b�/w�a��XV�ə�������n4kܹpr���{Em�|n�v7���.\KD�W2^۫�
�G|gyo�dQ�}�?�DD9#����-F(W�4�Va)M�!/���G��n���:�U�WT�9�P����w�'п��h(���=�w��3N����] $p8=�kR*�-�2h5bH.2`��"��D�r�}k�c�|��G�}�A')��\���cЕ�c��� j�ǯ�:f�(�2zvyhF����	���i�IC���|%೹����D��^9.K���p�[����t�6����U>DG���${�����)ҵ�v~74��i2)�O,�f�;Up)�VF��p�#�����k��ו�8q��6*b�K���>�$�gM%�\6�+��u���܇�LN:;�}�w��&�wL$ҽ?q���}�n-��z�y{��y����Aw�}V�s�Fw��ҧ�H�IH�tӱ����vK�K��U������aX��ǋ��x�eJ����p�������2Ee���PK~����c��� Y�mA6���1K�5�+*�_L�6�B���s;ئ�)�].y��/ӌ
웈3�JY��J���L�� ?��T�����z�6x�p(b�3'+��h�k�j,��0'#'�P'�M��OTr��U������u���Ən!�K��j�1j�+���GD*D�!�E�?�k��s�q�[ /,���/��C�o�ҿ��l�}� ���
~f��x_�3�1� J�x0ΎrA��VbE��$E���=Z7ؤ��-I-�X��e4P�1M?P,�.�s�b���MԱ9��9��s ����ƌ�7�l�y��a���\X�n��B�)~B/=«�5��] 9u͝.��'���ќbL"K��������/'��� �OR�Q��� Ol�GD��Yjt�c{����&�������}�რ�:��o�ki]��4��l
3���w*D�g�H�ъ�s�����˂)��DN�)yM�<ҟfy�#~�4s�f,Y(��ޯ�Tb$J�#�?��p(�Ώ����ͼ�-��[h�.�)+C����9b�_�|v�	�"J(rI&�������@U���H{7��5��x+e�����6�W����$w��(+l¡E�{%y#ņ�l�]��:�]����K�s�&�~lϩ���:MN�(_���a���jҕ6����Ae�N:]�g�g��G��;�ko�k�^H��j����qn�)��p6�z���Q/�Ԑ-���$�|�����ݴ�W[�\{�pc�d��֦���vɮ���-h���2B9�p;�v����k��{�(wYd��|I�����L��#]Xgk3�LW�L
I�LU'�fO�蠗q�,ۖ5I�`��4�������ʰ��	QmտL��#J�����̦>f�Й<����"���_9*U� �|͖!� ����׽�²��G.��j�Z��z՝9���+��5*`�k9@66�	�z3Jb���}����pVp���K����-��Z���6�����������<�˷���q���4y,I���D��hs��CK$����Ӝ�m$Jg��N�KkJ�u�(自�%��o;��n�++�D'��:JI-5;A�n/wMO��<��]�>_eU�Ǽ�z0t��'ռ� �/Y}�p�������w_�9R��t(�`�����o��������9��ަ��=��F��;�]�.��Xk����0Nl��=��o�4���ek�:���`��]	̝�tj��L�S �:�+��M��rN��[z�;K���N
��]��e�]�|U�5���E�Q��S�q�u�[l�*F��R2��A!�t�Ԥ�v3��X�m���Xw�KИ�c�"�"1�6�pL�5H�ͷmJ64�_��yIV�"�	��k[c����O����7���B�V�d�*�	]j�o\��9@[�O��Ǐ&� ��t�h_K0��ΓB��d���z��v�I/@��.g��?��'�ڔ�U�A\R���`f�Hx�CQ���ӆ�ۯ1���&M����,G!''!R"�<�HyxS:��[R]���]m��x�+���7��щk1�i����mUQkJ�����҆�܁�Ո�β�m`�Ɖ����'G{�����k@��0a���a#�����V��8F�R���K��> ���òmfho��$����4ݽ���7.�k�N�N�n8�|��6�#APB9��Ue=eDW�r����\<�2MT̮�'��IM�Z([��Q0\��-�4@u�0�Xo"�V*���>�<Zہ_5�4\Y9� _�u�&�a��i� WθM�� z��"��)W��yힻh�*�i}�J�RT�����S���@Z�R3�Z��`��fԀl�"-���j�Vy�oU����z�ߕ�1�e��♾'
�{�H��G�����'[��p���km��!A������	���O�+�e�A�w�OkZ���~~*��0��/�P�����P�n�YM��~Yh�b�SAdU���� X�"bWpPɚ��:m2n� �l��p��1l��]c_�� `�T���i�����h�&�����ƴ����Ĵ%w�ì#Σ�1�Sئ�1zI��#Q��.P�P��^�
6�4��efU1&���)�h��Q߀u�P~ׇ!L>�Nq�'��G��qsD�O�S��>��ȷqD��M2���;�j1�����pF�
��Ʀ����xs�dJ��$ٙ��pD
͓�hcΚ�j����"H��	���Ay��H 3���_I��O�=>L�����8P�ؚ�E�����p[�x�y�	��ⴥ�}��vQv�~xyUVd_���6m��;�§�TW�:D3xן�h�L%�]�#.�u�������Ϟ�Dz�S/W�Lg�R�2eo�.�9i�C:�k\��Vy�^wY?+4Znox��j7�S�������n��s-������D�k�����QR<�օV����޸����Q�ޜ� I*i���&��?"��U�V�z�2¢K.�dù��|���0�R;�i&�8�Uy6�"l2�<$h�U�=�#GÊ?���U�M�������o�f���w)mUl-�V*�W �C�<��mjr�E���@���Lԯb�0R�d4�~i#���QN�B�J�X�)Um�8L;������������r���ID{qF{�Ex	����t��`����x0�_)ʏM}�Q;S�;GKKD�H뜦@�v,ݏl��<���r�%E?oM!λ3�������@���>�k|����]$����!vqf��<��9T7	Y�
�|x0�2�F8<�0O��B�6Z��^�豳TEU���w{����J��=��W������{��/
_\�^������V�t_�(��!�hX�K��+>�1X2�\��*�G��;�!�?
����w�H�A�>� �+�?n:wgh������}_�ɟYI���Pd=�=7j�j�Z���a�cD�l����ŖE�<��৐ZΦ�̧��]6��_�;���.�����9�D�R�vl�̥���TU���b\(w�Sg,X8�p��X�7��������G�\|��\��$���$?��P�H��I"��$�SfI���f�	���*���US(����	S�(�?yʡ��Bb]�����D��`p�K�~{�����������Lز�y'u�Pk�8�w��oC�q��FPC�2c�	������@�Pp�-о���ê�M�.�W�E�`muߜ�:{��݁�l�w��j��I-_����n���m��ڮ��*�7��iw"-W��]����d��j/�4n�������D�������d�@^[C������@6��~�5i���J��i6��WD�8;�֟�m�S��v,ӘJ��gG��>�pg��o�,��go�A�_��.�n]��Z(�e��L|�~�>�>XdT���deM�o�F���BD��|�X���fd��~�g�B�3(����xZ�H֢�6ss�J4X'g�h�2�mbRJ��H�|ب%��S�_c��K}o�#�LB��!����Ҧc�B���+������+��l�[9�%�����O����F#�d������5)]��ܸr�3����dV��lH�_��V��fx�i>�ˤ ]ON���7�t�"�� @�X��Q������G�{�=��, �~�1L �!�! ZscJ�$2�c�,����`��cr��8¥����K�$��+�U������.;�lPS�?*�/����Z�|\a�Ҡ5���<(d�Ӛw�P� ʀzV�0!\�?�"������Rk���]X�r��HkȠP���Y�_`���8>��fs�N����������5jQת�:�j"\��Q��-��/l�6}�ӵ4�ę#UW���眢*
*)xͷ���)�'k~����{q��r�2������aeu���
��p6P��O���׊�ti�`��ZO°)T�\K�ɤw_UѦ����Zv�2
zK�O_�������g@����[��t��<�@���6�E�0���u�Sv��7zzHe"��Յ��Qy�c��:-����f�}����g;}Jvz/�|�+�Z�./6�f"��m�h��/��Y�P�������k��%<���;�]O,�L�M��re�o�^1��3��_5;�;��+ع�Rv�fIm�l��n�2�yGi��Ή��r}���Qdh���S�a	2ꬥp��@�(V��^���)�����I�/-yU'T>��RGKO��3>ڢ�����3�!^�[$�M�`�Q�	�u�t�3�3�J�F��� 7'u�Y@cr9I���*�b��E>��V鎖#���ړm�zml�m4���0�;p$L$��)����
o@�1�ߛ�9����N9����dH P��&�L�̨!�����i���ݛS9*�\��m�����(]�g(鄜�^G�⎢b�Q/��8G50�����PF�
�Sl�9.1L\�Z4�VG�����
���M�����|0�1]�jL]\$u�~�(����Y�zx��{�z��x�g�����o�����s�`pI�;���ʞ?ކH�Y�C�_%n�~6�9~k�'9%^V��L���[N��I1c)\J�(S"jysWe�H��U� ��Pd�"�}�V򠍊���[��i�M�]]�Em����ͅUe5��:Dd4+���᣻�,
ׯ���`4bm���Y=�_#̈́�(ȵ@;ҽ%��F��Wd�,k��VAA\:�UYR�w�g����ٯwer��?��z�� � Ǐ:�����Pe9��N���B�� ��K6rߛf	�� ��|Z���z
C��
15@�k@�M��!R5� ú4���^����t�Ό�y��&�����e���Զ�;�EU�����*�NY/��'ȍ#@�U%*��,nX�!��0܁]rΝ�Dd"n�n�^o�>ܲ��(����!T+W��˱��Xk<j3sT�W2�+�-�-�	��bM�ݡs��U븓	��S�����}�j�;�B��SH�����>Ý��1&�j$'�.��p�R�`U�z:�A{phj�:��ijy�f����_G�%&:�ڲqa��{ ɜ���h|�� �.�s�R�4\�=J^6ڻ�LtD�� �2�qѣ��'�2���ZM�U���o.�\��|7����Z���f�p(n��ZLYB������ ?XJ��B�=4��1i��Z3b�|�d��%Z"`߶����х� ���c1�Y
�Ԥ��W��1Q��`��3�!@QX�'��Dߟ���9�
e�TP��p�
��=f]=ٰL�iٚ�L{� K~1���A9�ɢ
�$_�I_�A�)*�/ӆ�¢(��Hs"E��;U�5���R��ZA���f����t��kT � D2�:=��b�XV�1[����Zo�f.�������炙��#�T�5L��K�R� �5�����?^p���$�|9CJ��Z9w~&!�c�׫�1݀�
س	b&��5������op�Ί���ӜX����o��K�Tp���*c��&W��,l���/�M2u;���FW�3j�u��68�;�o��������6-
k�-h�m�,��§��|�( ��V@��@���[g�T(�Q�e<D(Q��h3�"��3(�"��UE�<l> .H���������Դr�8Ԃ�"�a�U���g�L���n��ǝ���&�P��q{��m���˺{!��
���4|%��hp(��Ҵ[�|�ำ���\�i���`��}��i��U/e����쪟���f�_��{����W�F�c�߭�ovuը�Rm�>^U��+'O+ȧO*`���GO�zc�U�ۇ�m�͒
���)3팗jsBgs`����u�j������g�|�QH1Q��SZ�?;��󭓢
e��H�0L^E��d�h2R���Fs`�s�,��ގwߖ��	�NS>������n��/� �tS2�bD�:>�L`�R��7>@��*���`�5D�5�P↩.#G �O�H��O�z� ���-�cř�J�����W3��i���Nӻ�~�9����b7�}�M�����y��v�r�bkbu���LS��Qa�Rw#P�gI��x�����Çw&����h@7�P�Ur�η�X�<$�@�Y������~-D�ۯ�a^��8����#$Ի�q�E
hu2�\�k�̕�+����p����g ���i�oF_�L��޼^yZ�^�
��~H�/�c0Fj��^/s;߶�Q�PM��z�Z�q��1{�\�4��t̂�N}��xg��ĺ�$���sr�`-T�4�QbH+Ϛ��+{I��k҆m�9ՆE����p�{�eI�u���Pan	6���L�k�;�X�p	�x���v%�h@�>,�7T�>��]I!�x�$r%�q�n{��mjTB@!`ޘm�Sin�tB�"�r��/GϑGm���&B�$t(�'���	j�2�Փ�Ŷ�Z?���R"��},5b�O�*��̰#%/wG�ψ�)���e����/�Df�\��|�'�Ч�/�9�5{�	k^��Ju� ��(���l��<�*����΀�)�UK����C����q�X���������N�AJRtX<B�z���#-G�דeo8Hz}���t"�XT�e��v�<�t���k���ߙ��F�;�l��1�����k?׏
UІH��6��視E��[���6_�TWsgW?̤�BR�vf��W/'�'F�̭���_#�ې�Fa�
(��S�?�R��G�B����mS�;^�PG�Ueh�B��m�����q�aw;�T���2�Z�?�'�>��/���Go�gxl(��t��Tx�|��zi��}H��Z�/��~�,
�L���Ry`Θ��{�0����(�ʗ?ศ���|���;��t]Y)�����e�a2i���ԛk]���d�~�Y���:T,��cb����A�Q'�����`#�x@���n������;�7��M���٭�2��<���5B����{�t~D@���|���� d˭��i�B+�d�2}��H����@� �*�7'����Mn`�-����q����#�$�fxpd�b�L4B�<�I,|>F�Hg��E�
���q̀MA߸ӯ��j�z�C�Uy��}�� �6�'VH���m�=�k���,o�{a:Rݜ� $(����G�Y4���P1��/oh���_�A���)=_�b�����)��j�n�S�2W�ӼR���\�jt1uJ}��W!Me��\�:�e������P�n�,��~@D���ʙǺ��J�����[��
�l�w���VW�(-E">��O}Ԁ$W�n��!���^�g��S.�t슻��j����/k[�6ϋJ�+��}��/�@ҏ���^��t.C�b�W�~gy"UV�:\�lv�ml�Y��~�:�S����Oa5�i�пڄ��p�La�ܧ�k� 3�<h�P�n=b�޾D����'�(7�0�ծMۣ����Q�p'I���r���Ѯ���B"��V��g��I�>c�Y�Kl�)���b}Cj�������=-���N�z�c�W(��QgA�]*������|x�����P(E��9�!�-r+t(����� �7(��A� ɔכ4>�4��\-�T�.��}�����/5s|�:ys�p�q*osRkA,�8�������_��W���^���I��R^������S��#����no ������Y\<�m�����=:S�Bf6������x�"Ƒ9�km~��������{+�t�QE]�PKR����n]E��O�.--���s��ջ���P~���H)��' ������{���WS�ʲ#?�1�5���W�?�Z���3Z��\���N���0׫�uX�7��7�A��i����q�\U���)�4^"��yi+���:���/�M| :G44]����h�_惬���F����Pվ��-�@��:�D��?�( �(z�bd���x>��1���9��Z�M�S�w��*�&��!$jo)���w���S�C�^/�۩%Kc�t�B�7�5i��'�twu���YLe8/��ν9����~x�+�3㎏C3,�B�����AH��q��P�2��	$e�`*��G�H��٫:���LDh���	٨.%NOLNN�����oQ4g0���Z��kM���p40��1�>l����u������.�Ѵ�.}�{|zِ� ?���?a�i��c��cj��B�ē(�6���Ht]��M��8E�i
��B��:Xd�o��%��֑>��^)�´Y��f�#��<b�����J ް��JC�����H��������XF8�`%�"�a��� `�)���z��W�yC-O��t������4(	x�Ϊ�V�5+B����}@����d��~
�>{v�M�j�_�_��kFi��%@�O�t냻fVo�4,>�i�GH�j��jN�w	�D�.]]�W?�� n��i,��������8��D�;���u�~PN
�2�h���8(�ৼ�ו�	|�Zj�a�p`�ё�T�lG�vv��Y���(��k����ˌ�Y��D��(��E����	��.�>����\����T�5!b냘�Y�\��Ă��w��l���� L�q�ǚu�+�(��kMJ+�Rd�����*�QGS�#<�Ԅ�����Z�	phB����4ܱfdIw���v>��}ފ=I1f�5��yzQ�6rZ��E�??�T�g[��^��VU�d�B��l��Ah����z�=>&G�{z~VK�(E� 2u�M2-��"s*L9fyH/�9%)
~B�+��h��-gz���ͱ�Q��G�~ؔ˷��k�:Vf�����BRM���A�EJ}ݼ;[��W.�/�+xz�*�UA�N�ʩbB�B������d}��z-���j�aOpd��p��/�@�_S�'�O��dF��R��J� F��s��#`�"�(p��L��ļ!��뷃hX��g�C�,�.-��ԑ��q��Mâ�z��lS1dĵ�PTg�]��6���%UՂ~��s��䭾$[�[��y�3镯�ޭ�*d��[�H��0�]�n�'̽J=���NĒ@mZ��p�F��nBʏ=.�����:�K�_����z��"	�*�G��X&1�d|@t��s�Q>"؜��[JU�!7�	�N`�B2�@�����G	A��%��M���;�R�����t_���huF�����L�jۇ��w�'0)�5*jo֨-�^�a9I�41�X��ϖ�;��B�F����z)��	�J��7j�|_�����$�D�^�>q�5�/#g*�:��D�9�zl{�uA�+{��3S�U+	uC���zˎe��D���W��Ξ�~Y�{��\��m��1���fY�'�w�v�õ�1odc�3N-Xx��·3��hX�ա�>P�G^Qh�u�HbЉ����Z�B%C�x�lw�n+P�_f�k^ �O%л��s�C��`��!�rY{`�Պ�}�g5��������ν.��qiW���S�'���\Vm܇k�&�՟�|ѻ��vמ��[T����\�|�*A�Cϙ2G�HW%���V��K�����e����\1���F�[w�Y��.l�}H�h풀�����{����P|����H��/ ̯�ƺ�'�ݻTA��&�����Tm�.sR4:3���ZȪe����yK�����(t�&a:a�����`�K=Ŋ����b2�@r4�����k9"����X03 }�C���j�!����Z�c_���ŏI��|)2�+1�b4]Rjk�򃲸؉��|�42;c�;��j\/_���h�w;�W�<�|/as�Ⱥ���	�x-����ȋ�X�|a��K�0WO�d��-?��*5�� �9AF����KR.qJ�rNl_l�H+�ǋ;�����9_6�[��B�j�c�l�nd�ܳ��m�l|Q�azKu���2�S�b�1b\]�1;��T�<>v3�VETK>���|�Z����*�΃�����z�2;[�������K���`��%��jc[��!u@^3_�9trJ����?�Dw(�a�ǌ�1�yխZ�^a�l3�O��b������"��ILx[7��}fU9�Ę(L;�asA�|������*����B��?�:��SwU���wJڱ��i?�qB�ԧUDxUX>���ᅊ;͘U+��4?��K�ؿ^4m��o�+~3�����|��$�!�P�@���alc�|��E�|�V�9��R)z�u�݋����(�%�ۙ�"$�W$G%G��Q������o�`Qҳ{���@� �FP)<�GN~Epq���dF5���G��t���|�u�.�wZ�	�
��-��z�!����˄Ir+,%T�i�?�%��k�V�w�P�aD�&���a�a��,@4�ߔ�������9Uq�����[������̝gP�>�*��+�a�eR-���`�Ȅ���qu)[^1�pR�rt� �� wפ��8�\C*	������ۋ0�B�8�}�w��N��!iYUNy�G�����]k�!�kS�G��طAm���\y���:;�'#��v�3^WwػKզ�-^]7S}�w�,X�bw��-U���OThV(�N4ҥ�S��y�;g ��}���wMh׊�l�1�,�n��v��:B��s9��swb�AA%�0�O�o-���G����-i�1��a3�Sę(Na%�_}砠�ĸK��S��Tw^�蟩�u��±Bb��GH��z��脅z�i��a/dIj�|�/�|Q�==�̞o�8|Y2���ii�g�0�Oc�DD�on0ie�Tx1�1�aJ�u�p
��m����<?1V5>tg�~��+�;�X�d�t��ߟ[!�_����;Y���P��'v��� ��]Q�[��{���g���VMy�A,˄rB�=�o$gx��1����x_4&ߏYc:,6�B}�cc�V�<<�jm��ά�v�p)�շyS͋�(�*�.NTf �������T-��n �5#�.`/ICP��d�Yer0Аm��ʥ��\�U�TuB�],�X�^�Sa4�c�PހLs ,���7�c�&�&@�#���I�5��ν���ʑc�m�^��0B�űҹ^�B�I��	��g�x���C�T�����~�s��XG���G/7��`�Y�����ay	��8��br��������&oY��{�h���q��/(��BC+@�U:%�M��%��J���	�l�.;��d/(hY��+���#"��R�(�m�}S��ۊ�N�������s	�����?Ie�~�d���4P��^�~��&��!�Ձ�0���n�Hq`�`����{/[��g).�7��� ���ɩ\���,�ʦ_u�x�Q<��D�=;d��S���q�Pr�n\�g�Ϲ��dv�0��:��ۣ����$�l�K�Hr�ǿ�p�6�}��O�B}@��K���Y�������틞K7t����eߝ��!�7�z&���Rb+|���n��������萾�>��6�y{�n|�OаX��K�ЬN8|<%��E���QD(ͻ� @b�VD�ή���إ�}\ʴ\l�*�Q��C\��	0ю�a����E����k�|�L���u�z,RkP�� ���q����_'�y�~m�b��b
���=y�z�8��q�vr�F}��C���5��O���R��T�o�;i��:�q�3Z� �g+?,���θ9����M1�*O�6<�QZ�buG��R8�5DZB�ܤ�u��!5��Cb:�������Z�Bݭ�\!���U۸��4N�2�j%�����`�drƃ��p$�~Ş�K~T-�/:U��gYLҮr��β�I#��_�-�j^>s�uu�wt%��g�=ܤK=�N�<���]�ݾ;h�&,!+�&�ס�c3D3}������ؾ����9�������߁VH(N�R���vj��ʬe1\x�4zj�z�F�5\t�Qi)�����������#�-ν��ȑ
�3D%�H���vC!���e�� R����d���XT��������,Y���5�&y�2"���0Ώ�m[����d�+5ٯ�_J=^N<�K=�I�zl�FkL��E�W���?qӳ��Opp���7��ċ�#G�5����f���'�R߿�s�.a�/ ��+¼���\��7C�.�������
��uٛ�b�A��oI�|�X�f���sp�$,���i�Pn]U�����5p��5n�p/P��%� u��B� ���fd�x����fm�d�r�t"��cYC�@͂M$B�:~So��>㉀�����qH�bp��*s��9Ȥ�Ώ�G7�	=^9�ׇl6>�I���xd���R���8���{ ?�$]�2�5�2��VEM���g���;�ow~�.���\i���l}���MsU�I�����Jp��v�I��[�����e9��1M���g�ݱƟ��3���i����~�B�w?���S�-�vlï�s�����ca��j��o�*��0��uP�(_CT�
@l��rgtl/��;�u~o����䅬+|��b��tgLG�4�YLr(5x��b�eP�;��~�*L.��?��YIb�%=�X�����7wk�{�jN��IBc�z��j�ؑT �d$��f�p*X��&��x,�
�;~%^zv�ޑRaP�%Ѥ�����L���V��R�=Q<5��v�?��w��Q��<*������Ej6�����0��ϯ}F��;��V�R;3Y\8�z�k���k���F�
�M̄�
]:�Ky8)�2Ri���]P���qs__��c����3
e2ʄ-'e��6AsS��V}���$��Y2SK����W����# �[�����kh#��A]���dj����:��T�������ү��Y��kş���m���U�w��	�O%3�FF���ɪFE h�Ri� F�Ȓ� #��1@p��	�<��'(���P杒S��S0��t~PZ>�6�s�)��h=��_؞݇ې%��Ե҄�|&Ԧ`ЄT��숆���w�	y	H��VK�LP��H�H��V��Ϭ:��ҙ�y������*[e�FJ���9T��z�\mT��.�����fS�`e�P��2w�B��Yر#�a��s���r���d?�;�%�l7���+��\K�G���#�q�D�+�Z�x:�Z��0�=�>P��!J�d��R�(��7���>}��d �����������p������fگ;K:/s-�yRQ�������4��wӳ��m�:�|�U�/��)����2�T�^sU��/� �������3t�+p�_�����\t���U��uyx�՞���3\&��N��t��f)3<�̂�ۏ���a�kb�(��5u0��|�������Qf"�\��`��!�G�WW��{�86����4��n �֥L�?�b�Uf���t"vF�0��,�7JԎq
�а�s�9�̵8=g���?7;�6���i4���f|Q�>qܾ�BrƖk-��8ـ�/��A�(,w(�}d�Y��S
3�0��s��	ŹʵF0�~��`%݄�n��0�Zd�׎1�6�h>r�ڞ�����n���Q���
U�ir����:S�ܢ���3��*���S�؛��؀�/��`֦���v��m�zeIE8��\�C��8��������Z8ӓ5Z�*��ퟅp�>M�[�4 CpV C~G�8�|C�9{DA����~�]�<�l����u�4Vt����CdV��C5~\�O�=l�<=���{)v�]�,,ῳ�������tK�2�=l� Bȧ���+ɀ��?��*(��׃K� 	�.!dp'�}p�@�<h�6����ap���.��T��������^���zm�A+�� ������kH���U����c�@\U�;ɢ���EN�CB�9�4��G�������Z��]V(�����S��(V_�T�>�"����9�Ѥ�^��g�+vsi���U{`���3k�%�]=0��b�1Ț�CΦ�Aؗ��Z��)���$A�,�[����^��T�����O�Vf�Za+��Ҁ��~aវ���,NB:��~o�mv&Fo�
��	��Q?[���$���B���cd�V�B֋L�5��L�T�
��14	y��6L�K p�\��^D0�����P�
YDn�U@��T?�RW0~�L��{�� תS�]m�Y�%&٣:\�#Ձ�1���?;�bzqr_T�w�vL��V��Z~hU�]���7!���F2p|ڮd�)��q'(T��$÷b�k|��@1�| -�����HdY�������/�)Y����.SGL�7�c�i���d�c�m�s����?���ն���c+������!e�D���|Yb3^O��Ks���Ѣ-ܗ}�>�*Ǎ�%O#9f.
��yᛵhLC��!Mon���w���ѷ���臝�1����k�+iR��}@��4 ��вFO� ��TM
ĭUJ�g2R������F}�5|(�`�Bw%��F����0��`N(	=%����{�4E�Xtr�Ph��)E�`E����CP�uT*�Rz�$��o�������J��a��<Z.1� ��Y�Yp%���sb9wFU륷x?��Ĳ@	���u�7�"�oװ<��,AѱѢ�Y�{%Q_ۦl�<���C�3������ �ն�+��<�x:!�vf3�&�@?I%��P���5&�O4�>��A��~o	�>�V�/����s���kP�H�A5�W+��[�pG���-�Z j��J ��g_�[���֘u���I��~-+�2�����qmT�^���� F�lt�[�b����L�6|o��c0�7�8��M�>Bb��� ������F���/�z�q�1���$OȑXM�k��ٔ`�"�q)�O�% Sw�
�Ľ�l��G" ��Z�#�.��#�ΝBJq ��K�|7�Zː9��wahz����)����P�p/��G8Dc-�Ê<(@�|{�V8\b�����G�f|ڑ�9����]�_ܓ\\hU.�.���2.����
V�C;�v��&�qԝ���^�����p�Z?S�|*��(6�(��������J(@\$���"a��In��a������<����癔��-߂�	(��<�>}���sEVab*攆���1�pp��Ȝ^���/��b'?�Q��5��=�j�N���i�`"�H�>]��+�B�ooR��t9Us���{'�����Y+����ƏU�����der�t�T�j�Z7�=��=��*���m4-�t����8�fR�w�k��Ȫ(��C�i~A���?��d�-��JX��L�}��i�;:���A��PRa�������y���q��2��?�`߈���ê /��v:Ba\L#t��3��U�!=���ۄ��"��,�9{&��q -���Q���&���S��:���\Ŗ��
V�{��g�����f�.j	តbc��W�Bѫ�K/O��Ѣw�_�+k�)2Z����K�43�a�iM�'䤺0$��Vt0&�.*O��4Nn���J����_�����V5��m������:��Lm$>̿���͒����	qU�jI��iq�w%68x$2�f�7r����x�	3hQm������tU�k���V!��Yd�2T�/�bO��?�&�~�����>n�_�r�xBo��T��K����Y��X�@�nuw#�0����L	s���.��0	��ڬWx"�?�MN 2R �4��m�+�w��J��!X*,~lz����L8��a�3�v����D�WMchV5P"��Z�;7��	'��g��G�aTN&skW`4�1�[�2|�5���~�O'�Y}���]�>�������b┌2U*��P 2�&$a�Tt.������E5����U��XY�� hT�,l�liA۪�ޤZ�������$���o�'��*���mJ����9���W��9���u�8S�.y=�qze�����o�X��YE�*'
��@���@��h��PL��f��UU��vB���,wB�%sQ"��ߧN������0���~ަCJ�o���[K�U/��jo�i:i�nu0l�ܮ^�����m#�/t0�vp+s2���I������rP48�?.O�L�4�g�鉵��4�ܲ�x����~�h$P��y��UÏ��gϗ�C��X��8������ǋT}m����jQ�ۇ�ۤU�y��ݣ����k�D���B���2���(���9|8��X��%���kt����[7u罅�ݽ�Iu
�N(���tGa���]BR�������������g0��I��g8e ���I��m;�4Uy$���KY<�n��6Drc�� 5Q*��Zs?>GEuV�8u|Q\70�wc}��g��ٛ�/ tS�7�>��6�ns*�1:��ӹ)�Zw��k���\u��r������k1}�����6������ҽЌG��r��c�MSu���Q����%(/�W.�i^8s�$�VL� ���л ��[~‐(�*����l?��/H�4���A1�"���#Ԋ|)��%ܑe��c��.5C�ƹb��+�E$e�~k��!.�o$e�QӋn�\9���Ѩ�_H��W���������o���!��؟��`0���\s�E��q%��/�n�T<��1$RL�����oF�2�5�xQ�q���~�k�kt"��ܜ�F���'qOߡ��6�y5�"�>d Kvg�4!V�>cd�D�#����.�b��7\@�:	�5%��l�L��Q�����z��
u� �Fv͝�D��h�@�`��?�������l����+��g���ǣ���9�Myϋ��Mt����}�;�K������#���7֙^�g6��]�"hT�������s?���fc&���j�&����qC>֢ڶu'}�i�6m�0��+7�����8��^*����&"b��x]�H4�9���p�e���J��ʸ��gaݙ�Dl�ER�[�ۙ1���8��
v֭�u�;�0[��[4�gu�p-�ƺ���;��@O��Y�Y��ݺŭ�C-y����a�1��o�9��d'�oh��*n9I������L�v!+�0|Ⴔ�7�y\�s�x/�(�2@��>l�O��
��mT����p�����u��N����qeg��Qp"��(�n���;��i-3���°��O������LT�\~q���%+��M �8gvN=���3�Mx��3Y�K1X��՜����}�N�����ÙØ�#
3�z&�L�muF׉eߟ��߆hS��u��y����y?��������*B�ej�2�S:�]e���d�<۶������ �B[�v�	��O��V�;�vl����/y/�Q�{eꗀ���V8��"�oȄ�9��!8U@��Kct�,��azs�4+��O;=�:�=�K�EP�K���G�v�l]�-���{}.�󿖴�N���7��|�*Y�{pA57����A3��`�m5J�΅ʘ�n��3��t�Bx�M��#|@EaMy�q�
]��'	Q�p2�ź�v���a.�`|��I%]p�u���^��ݰ�=�'�jg���(�}��ub��a��-�|6��8�&��d��q�;�J�|����͙�2H8�!&��"��h?DAe��ݝ�U��
�M$��2��>�-(�U%^��?�g��d�Z:��@1O���7�5��ޖ�����'�����7�YfG�Z9�Lۡ٤��3ë��a�`ƻ@����5=E�˾�T�� >"n�����*ƙc�g���U:��)d����uV�Xv�w �����
i� �l��}��g�<R{����d�����V5�@G�jG� �W�����D�8��Y�̊~uU��$���j�Ϩt�;�2�{���9a�*�
Me�z�OS/�d��i������G�B�4"��h�=!ޖ�߽��'�V��u<wO���[�6/O���G���^��k�]���=�E��+�zx=�
�8�Eiw�r<�@�*_%o���x���G�s0>i��]h7�y�Q�6�7	/9�B�Y�x}?�,�	��t���|���ſ��8i%���*�+�=Kh���X���p�t����I�N�l���2\'�>_�O�?ԲF�[FQ���a��\h./�����5�� e+�˙@u<~�e���~u^POv�8���:��?j�d%V,� [U��n9b,^AR v��l�(��ܦ��8h�#7�W��c�΅��4�ĪC�2��k�n*c�_Yx���D��̂f��1m �gl��{[����cLG/g��F;s�u��U��6��~�4OZ��d��x4�D5���̻L�@�U>��`��J�|E ?t�U �ѯg�3��(��Y�=��A�K&�X���v�d��l�����|�v��6����[U7v6�IȈ��S��!�@�mg��2���wKT��Aa1�a�'����(�"�&uDu�WEN\�Q�gBFP�*D������a�u��u�[�xi��xHZ�U)�K�"�� ������%Tʲ�B�B�m��;C�@�z)�L��k&X�h����M����
+�2 �(H�������(c�ߤ�����d�ă�<F0p�N	<��3l� =��-6���H���]�y���B����~6���d}z�6-��7����+CB@��ł��CB���3?����}�e�D�6�nKZ���=�ZM�Lgւ�ڪ�3�u�ߴ���f�W�;À�&2���՛w��㶖5���$��V�{����_Sq-zq*2����9���.��Jf&��W�mh�VS�����X!�uV�V:�R<�=	���N8(���[A�%'��B̆R���]�KjƀX�5��7��C�V����K���'��x�/���J��@��D��Z�wM͂�{_ꅤ���j�0���W�:����c%��?ܙn��O���������a$*ڊ�������v0�&��{,��n̋
 __gD�f�Ċ�C��jis9����9az�#{W,~�I4�����)n�Qiv7�?��Tֿ�݌�vΡb�]l#n� ��l��-�@!��`����y�х��f%���&��Njlf3;�ý�ѫ/�yY�W{�?���ڽ��_����l���=p����(�
���GD*��'QM*���&��E�q��kÛy����bBEa�<�|]s���pZ_�\�5xՁ/S�y��*,w^�<�|\�d�� �h��i�v������/T��mM�_�M�E��2�neq�6,Nxx��v6�{_��\��m��|�{�'�����ۖo���\����hW��D�f�����Vv�l�����\��������U��=����-�#�~�t�������&�����D��Mn��$"ZV�_XW�l�8�z�n�u���:�\5�6�r?���XxI�`�G��4��Q�3�K��y$�ò��I,`Z߫�2���/���?fI�﮹���ٙ�3اi)r�S�������R�W
�c�͠k>�Y �~e�����#��*����ȼ�زW��3@)�H�N�K�E즇F��0�/JJU	��Cl�zL��������P��ɅE��`I|�ͷ��d:)��|�|��Z��h�����=������,�dmTp�'��y;Bhv����W���1�/fH7�x�<��EW��C)�;��_�xM��; �<y|��{F������ͱ�R�7�Y��S�`�du�Nj��ۭ�n[�S�G�_ɫ@�r�ww��������2���"�'�ۇX�l���{�.�2o���������A�՟�J��Ju���=g�
o���8�w��Na�e�o(����?��o2uSm!ªm�����|�0�Hj�=�9�9=K�$2�t��6����0�T��o��5�T�`�ĵ�_������%���ݷT��ծV�t_+ԫE�҅��g�+:��h�j0l4`�d��޻��)�q��&J��I�U-T�LXˊ���"�U�c����!�a�Q�����2.��4BhZ`k�CU�#F%�]�7��W���j4WLN�Q�T��iOM��Jrw�d�Bmo �,�}�}_���W�J|>~8�~<�}�<��s�[��m�mwg�^nK����@�1��8�ra<�v�6�L��{e�V�L�f�`ǘWOu��D80�x��~���~�Y �4ϰ�lԘ�������KѬ�5ЧnPdj�����-��P�����D�ˤ�|�Ţ�d*n<�΂�c�7g#a&H5�M���S�0�s�w�h�Z$��o3�l����F��I=?ݡ�>�MR����(	~[�e�0r�o�(��'#1�$���d|�u�����,Ä+�m|@<�لNU��߄�}'�w>�7�?��B�ٜ�ˍٌ�gųc1��R*�P�y\?�	��4��� $�)�Q
ĭs���W��]�E�p�
��#�5��:e^ ����@��22uS�A�qj������ާ�a��3݇3�?�e�w���QT������$�!�ɵ�b�g�f�F����B$
��o[�Z���;�-�sۼ�!��mv��Qf�����x<���i��ↄ���r����9��jK��fԛ����,y�� $�;0=�@�k
����cw06��!G���G��d�q5��ؾ	��j�4��J�>ŷ��6�Y��Z��%Ą�L��d�^l"��$��=���?�G���ͷ����K9Fff�q�,̘ɰI�����W/s4_��� d�Z�������l���Ivą�s�3�ߣQ��;��B�_�f��ݣ�'Ђ�78\{{c�a��^�uW��y���T�/�p����7~M�=<��'֋b���(�O �#b!�O�aY_�&�������Ҥ�-���D�������|z��ꡦ�!B蹟x{t!���[�V�讀o�|��s��<��?���jKj߆�t=1w2#� �6e�6�w7��6�muf9�lC2��I����OE��O�E�~z_��\�������qhm�-���"E$���5+��$Z��^E%�gY��V�C�`yK���WO�22Z�+mO{C�?E=��;~�g�����=��|_w��X7���7�O7FHvJ��#*m�`�¸�rap��/���N�^W��j��	ħ~�i���1�:�Ν��ji5��{5��я+�"��.E"O{փC�'B�s���v�FG�#�� %�r��R�Vz樨:'��O�Ȕe�xRʃm����fRŻ�h�I��X� �d!X{��F8�l���x��._�]��,�<����^��G��z�Ol;8>[x�Y�E���صDo�ٟ�2$U΍۞�l����{���E�Gߛ��q/��l*�;J�˲@�^��f����՚��$�H�����n���OGC��m�qlU�f���f4��R-XA�����X���n����hQ2<��B�.*BM�e��e���Z��RfD�K�f�;0dC�O��<�U���[	�ٛ�CX��E!tZA J^�~O���!pq����ٳ�{���y�O���a����ӛBt<Lf���rx %���׀hI1�ţ��,(�U�6��'<��Ю�ܮ�n1����y�����ѩhX���\dm_洱��Z�RF!��t6�ۻ�]�9��d
j4��{w��5+sg�j�:� �j�����KA��w��:j%�����dÈrJ�+�(�KU^���QC�*��<]<��ԿV����eT�T� 7�n�TșO�ڲrر�ز���,���Ks=�8�?�3C�?0>�zja]�͜�3G���$>�w�����}����B���+�3?�j�T��:��F�0l��&�{���FyD�XG�;BM{.�i�N^��,�ܳ@yDsޔPS<��7l]}P3�K�= 0��I�)ޚ�0�d��(��{f.�=y�#ț����\U4J��e�s�d	!B�|�֐z� #"5{kќ<9�T�M\ya�IB̲�z$��kWw�@�����;W5M"Ҫ��K�@���C��C������O��v���cB1�hWۘh���,	o�y3�-sHҕ��G�3��@HYgiU3�T3��W��l+J'�OFG{Hp��\�_��F�cw(Y�X���>;� �����qO�d�;*�1(�6��R,�`y��/��Z�M~�n�5w`J�Ƹk���0��꼥@u���x�v�\gu��6B���;lJ����2S�&�t  �9@a�P!�_X�=B�����7�������o[t@��>A�df���E��RL �x%]6j'��rH�+?�뙕=:�������M1��C��g��?����	��x\dz� ���c?��8��~�1A�<s�a���Xw#IQB�}9�cj��|W�+�LU��[�B݊@��X��x$ \���(9�����F��G���x@5���Q>��Y=�2��	�@��G�`��[���o������Ø=X���`
m7����� �7��l<���c�}���)H�տ�YH�:~y4��dp��8����`�rv�]��J�;��j�z�Z"倒�:"���v���qL슽%��.�j=�����<���p_�/������G��C��"�띡FrT�TM�bn���[��^y��7�Cv�%.�qa�z��,jL�<r���$0(�X� �N<$`pSX�ʌa�Z,�c�ɞ�FWJn�sr$��Pp��B��2>�)?Vǽ*F2��E�7S��������d� 4�ƪ���9c�ջшZ���42�ar��1���6~����8Br�x���``Doo_�tO�̺S��D�x�zO��E�[��X�X������i�"ǋ�|�}��<p{��%H���Ώ��Z��q�FA�J?�:��I�Q1���r�'iTUN��P�R��sm,_K�'x�H����V<��E��/yo�^���D'N�)%!X��X7��8`p���r�atǍu������#��^gD���-�����E`����a��Ұ��y�Tx��K���K2?/�ȼ�i��>��zڒ���7q�����(0�+�zh���g9g�ǌ3�]e��D]�ٛ�J[�u���?��g�_�'je�z�Nx�>��G�N�i�������vb}�}4RE8��I@���թb�i�i�GR�Y�_��&}��A���f�3N���}zz�U�B^7�Y)��"S o���&x��_dļ_�O�o�������WoWۮ�j/Cn�(a�\U���u��T!mgϲ�-������j?n�h%���͢��Ֆ��T����oG��j���D��8�**�����G6�</�]+F�m
@%��$�y�
�T4-2r�״v�jE����ҩ�^�qi"��:L��XQ����H�ljI�J����@�	n��-@�P2��<�7�vV�a�IHi����<���ˁ��8��Wr��u챑z챇mq�i���̽"RqZǊ/�	�3F����2b`;��>���M8�}�@���ub ��:췤�L�O|�V<�4|��O��!`$F�I�$4�Q��ya���b����$f2�T�
����\��4?=t�b��3��by�V�,�sd��)��)[��������Yɟ���^��[��܇o!��pqOߜe�w5���h�"� �����EXMc� ��M�;��,#	&J��������"�L�� PD/R���BJ�^6���Y/���O�5�����t�ٻ�����%�F�R�&��Y���azʢ��%����P�9��5�׃ȯ�v���6�y7������O����ҳ�����*]b/.x�hd8Wiq�������#�ѕ���K�Ն	Ζ����U�#�B�B�A)�x���}K�}vV�m�C�C[\оk����"��9�afJ�7(&R')x����G�B'��>C��Kd�
�2�4̫b�����F|C
�g�Ak�w�		uZ|	ZD�5�w	Ѹ��Ran�s����a��q5]t�����F���+��*_i�L��Th�r8S�!�#��$����9P�+y��Z��k`��Δ�g��e�:JJɄ���RO�� a��?�QId�ť������'��E��x�H/XW�j{<IX�3�E��r�9c���O�t����=Nhc ;�n}�������d���@��_�JT=��Ň`f*��E�Vp����I|�����N���oҒ��@���K�l����7�Vp��N=!_�#��B����vb�Zɣ�`v���Ę�E����xܘ���=6��\�p��.�/��ދJ��>y�u?A���BAW�lbS�8�8�'�վ��ٿN�����E�����`zpZk2�J�ǎЀ ERAC#��'hp� ۳��<#�=��:ZF�
�)��x���4$�zB�(Ҫ��Q";��E�h8΄�F��I>�� R��L�K��TZWS�C�~��Ư@J�+�1)��fz���&�9�V�u�5B��'�}<�ǘ��#���gh��帎&G>���ACNcK�Z*R��b��lmB̪[v���pi���^]�DŹ�|�F@���z��\�
�\��m�n�GѪx�4�.��Z�*�U��ï��j9�P�E��O5;��z.�����J^C�xh��Z�ƃ3��(�M`	 ���B�t)]7.�債1MUA�9�g�dHMI>��:���?�m:�S���J/����.ҫ2W���s����Jg��_O�_Y�(cS��_Lg�Ǒ���[�Wħ«E��y���+�ْ{���A�o�HE��=�4���ĀC��';b��5=I�i��m�\3fJ���Y��
kY!��"�����~�t�9c����De�yچ�q]���<�_��δ��Wi�{%˵II�ιn3/�����ѬB��aN��/��$�"���#�-��ǘ�����H����5I`2R�aj|}5�O���,/���T�~��:۝�����Ҽ᜗P����^Ӎ�4@���hj�J���ΪR�O��c�Ã�������7�[�_'�X�r��?��7m
6fr�Z��0x�Y�݈�K��}�9(r����PJ	�>E��E�����,8��Ȣ�tV<�d&�1���{��D�'G7�T��1,�Qw��hv�p�`j��]��N,G��h�ϐ[݋��4�ޙı�nN��;�
'���6U�!S"Vg�w)��0��Q��� oK2�c
����F7e��!�������M���2J� �o��j�[�����O�e�ԙ��p�6�ʳ��h>�̈�BWs��L,NZ[.�5ǜ�JL7���'�hș�C>�i^�7����Wn7BGQ��5����(���h*"�~�5�eb�tb�/�e��D���W���9�nƬM��+������{%��߄�q���e�q�v���oڛbP�q������W�X
�#1���#V���.�ߘ3s<�:�ֹܺ�q*p�v�j�YN��n�dr�1d����G������X���ը�kv�k�i��3�w7q����G�ⱝ���w��9��*�B�W�׆�\�Ҝ�i�� �y1��a$*f=�z,��fߞE��z��'�M�껫�鴞���y��HI��g���<H�k9��_�o<��Ih9+.Q-iJAG�C�į�-�(H:=�<L��D9L��ʨc!��l�Aq_-�[3ɱo�9%ӫ�m���/��l!��8�6K�_g���j�ϛnc����*�Ѽ�bk�`%�)%f�J��ddq�ԫF�@�ﭬތ�	�3Ÿ3~X>��8�b���L��z��$�ŻL��2F��#L�S��gڏoW�4z�K�S��C`|8�T8��b��歕�y����3扞R�)�����7����6����jc7Dx�}Fv�Į�L��h�C��?�ո֓�h�gf���3���{��<�5S��^pp���� ��\�Ԏ�$��I���J��<�V�Í������w��/Ghb�kK��mn֖5����S�6ܲ���l#��=�vv�ܾDDT�����6��sOp�utl޾"~��r3�~�3"]�w �#}��5+�A��o^����!S6B�³�����e�*k��t�X��wg7��8t�r��'(p5�IB��8/�����(W������|.'��I*����R�a�`7 �('��&�-���"!��_���9�gS(&[2YG������7�uݹ-�>}�gRd��;;�X_\�ԯ� �?Z�H�Λ&����}vGO:?�@a��f�s�$-�@�|kJ'��o5���Nn~~�h��w��J��֍�Bv��u���6�r�b�`w+ykgۊ��%��<��>�}P>� (j��Gk}{.�b��2���G�㑶b����n���1���?�*jJ*b#3NU�������_�c����u.i�����W��@^��!HSK������ʮ��ÖM�������R���gK�wAv,��q����	&m�	�:-��T$~�7EU�ۭ� �]K�~��ðA%�fpȗ�:�% ���I{O�� ŏK@̕V���FY)�_�r��(٦�Cb/0H�]����g��tZ�J�B��~��u�z�{�]qk�tc��v�l|��U���ٛG����@��߼�����==�ܟ�B�y���º�[���ih�#;��mg�Yݗ�� k���LE�
��c�*T@X�Eo
Dkɮ��Ӕ9�"��������p�4ͪeT`��I?2�r��P���;֘I�]���t؊DԒ\���)��\pd�V\�G�(PK<��d�6)R�8@	�!��O*lR~`��&�(Y����.��b1�t�I9��c�'l[�r�5J�4y�"�¡����ֱM�8Ŝ�1�3�^
�M���180��c[PM�SͰ���|D�%�kR���Hٶr��9���f���!�x� ��ա��H�V�P�]�UR|)�;�Z�X��I�o� ���U7~�p�o��x��K͕Ո����QW&�i�+�Ŵ�c>������?^��A9@B� l��ц���`�qL P�k��1��Z�Ҭ���lS��%��.D�:��W��i�|G"X��TԬ��]�/:�s��ݲ�|Sӊ�pb�}�s&V$O�]P4<	�򜿼|���o�-����e�I^�H?��J3N�eK�����sñ?��:+���_�"���ẘ�~,�ԍ���rX(�������v:�,t�0��闱�[1YR�w���I2��2��ƤI�Q}�},WzwVx����k5�#y�05L%�&HLN�y��?H�GF)��oV�0HzY�՞�V�"V�>�Չ)���N���s.��a�4���b�<��|m���vڴh�؞b̞9m����~$�T�|���`��'}\,�H��iY�;f�d�X�D�_XO�D�hͪ>3t�>�Y�)z��K���h�S��[�-�9s�Y��vvڹU-�߭�ldj`̻yg�o�CǛE�ɗC�O���b�/z�R�;L�`~%����+4_�R�z���!Z	�O$&M�$��.�2tBf�a���������f��8���@
���<�8�)k�١Ŭ�F��C�;zGf $���{b�J�D3������#�p�5����=�����@M����V�e���2�mE�sX����e.�����>��h����ϻ"Ro����*�a&Qvy�Q�YQ&��rbb�9�ߐ��}����oe����k�b����H�ɾ�9��SM�C�)5V)A����(3��5X��@$��%bThtI�L�mň�
��6�Rv���إ��?��=yy:W+�w������[�xn�E�a�zY#{~�<^��Z.��덚+�M��|�_�.��L'PW��%��2�q<(��il�yͱM� &��L{pv���
�|�SKB����iD�>~ER�[/e�h�==�'��z���Y�!�*��j���-{rR;u����o��z����wW<�Åy�qG��-X�o��V�u!J��F��iX��U�A}���|~T����bOk+2/�T�sb/7|�w��W���q��yA%R��,���I^��(�gd�s��1!l�@��b^������5�B'�lN �}�B�KIʹ��^�%Y�oI��y��p�4��%�7{�@��X$�� �2_��Vo0�#!P޵km���k��Dh�6��u���B~iKZd(9�Њ')���˕��Qԏ%^��+|g~L�M4$ ڇ�
�y���{�����=���k�LF���P(��;��Ƞ�{W��º<�eօ�*�����A�sٙ����������ۣ���~lN�cq��y�m�3�Θ[�˯���*s�`�NMgL�Q<Vu�6��Ӗ3o��f�Wm��d�"$�>�oSAm��{�Zq5wj��]u�a�xA��`���9� W\�P9^��Ȃ~�{�_A�IU=�m�E�W�����{��q%<��c9na��J�ɤ�#0�Y�c��� 4�a���q��vY�,����y�]���m��Y$[ݪ���5>t�[+ímZ���l��+�������-\d��5�H���eVC*���M΁w@�������hJ�_��ɾDM@jA[1���n��(�6��O�C�|A�Ra�+@�5B)�Ӡ$��xw�;IH>�x�iS�L\չ�VKP��� 
�4$n_�3�F1:n#a�#^LIi�7n��̔G:�:]�Au��G�x��A�d�Ym;�����nΓ�H�?f6��y8\��$,�!Z.5t���{F;�1�;v������g[I@�8�p!�[ ݅'���%�w� 0-*H7`�������^+ݵ�=/TE��C���W4�[��s!�J������㞽oٷ�&x� Eozdk�h�ݸ�ܔP��Jay��݌�����7ݞ�Fn^�[�?��5oF�㑝����h6�\�9|252��'��E��"j�Y�? ������Yh�	�� ��A�?����1&�G�=����hHb�v>��>F�bx�C�����\rG@��r0�a�ф��Es�T�� 6wL�U�����%��ef���*KՕ�Ji��J���"�� }#I�6���|����L�9+)���H-CEc}[� �V�;K�V��q[K��D2�4��A� -s���y�Q�F�:�$P�&����������[�˟�-�h��u&�ª�DH�,X�P�k�YUC�g9�ֽ���V��c��H�!~sԼ������M���9Vy��}S!%?� #%}��?�����J�A�6r6*  ����ݦ�WP�cTlsh _���ϡ��\�_��Vk���.��J3����Y�x!lq��KQ+|��O�;���&e�0Z;����#/�a����0A���j�����𻃨��U��͛�a9�k���!��\)���]L.{ȼ�%��m=W�Wq�]��F�Aa �YY6��a�K�A{۸�܂l�iV6�ň�+���5�m�ݯN3�0�76���a��d�ϊ�t�a�
ty�L�¡�2�*��o̉Xjo/S�-�%�w��\���>��Բ��~k:�,���<Q���t���� �nt;?��Ɍ�>�2
�y�>��|��}��-��נ��5+�Zu3�'��������|kIg�#�#7���$��^�Y�O���wl�& ?(��H��H���LgT��5����������M>��%Y ���P�~ט���j�����_߫ì+Y��|���^�oO��.BO�~VC3�qz���{��u��K�}M��,.K�L?�o�*9�o=�.9p\ίx���CgJ�����-���Z���}�qI�l3a�7vl	��J�R�����,;�׮�R� �l�!A���^���s����.�E�����g��%�=<����|<]�=~8ߜ:��z����f�&��-ȧ�l�=���弲y���Gj����ת:�_��}��9|b5��_�HI'��.&� �VRtk��l hf`�p�uż��X^��6ӦBe�)j�!j����������W|���a'GD-7H�.9W��y�*�R�q'��su|�}��1��`��y+-�Fx��I�V�l\z��U�Ӛ��v���C��i��E���]s��3�����?!Q*X'0��7$�4���>�*�K�ҡ���K�]���ue����}I�a�%��fދ%�
�m]�?D�eP��w����������kp�-!,n!��g���!���ߺu��j��̇9�����ӧb��n�-Z���i��1��C|�h�qQ+�ŞP��c��f!I�Xc%��2� J�oR,o<�SF6J@��G4ځuw����w*�(�|�sIw��	�`p]��\�����QE� T�]X��T�d������.���)h_�O�	-Z9��TH������z־7�Ή��:�i0\ʗ��,(�����%�E�b���*�IW�h��t+��>��c�l<���Ă[�y����zϚ���Pmt.VȐۈ���ǱHg��ц�8��:Ê*4��>%d���ʏ=�T�R�#�����N�?J�����c�Y�L��c�y�c���+5�<q }�>j.���9"���sҩ����m	�g��ۭ��?�Utz���B->�����lK.^�1��& 2�P�gO
~�6�j�S����~KCW�b^!����W�U�;��L+��a�b��u�u����T�]��
�Z�h�m;9�8%�O?��(��0|�ƭ��-�i�$;Ժ�ںC�ĵ����nc���i�*�0J���kXD��XxMǙe�ó���dK⏿m�m��"�0����J����o�Z]��Ђ��z�`��1&i� .���X�`ٻQH������t�%�����L�.u��
 T��|b��oҨ"���0�����T��%F��Ia ��Q�wK��U���r�ud�Vh@ ����1�����Ǯ�,f��\���{i����-Rd1E%U�b���2ٷ�ѳ�e���p S~}%��#u�|q8r��^w�M��;q��#k �873��4[9�H�Ӝ�h�qK7��7��,ng�9�Δ��A8h�E������yQ.�7��+Q�����j  ���x=\���Jj��g�k������1������}���-���7 ׵-��h$z��_1Ǚ`�Z4>�3fh��#BaeX�"h��B�Ү�)m�c��XT��e@k�tm��P8�t���ܕ�(��d� �,�.�ʢ��]�G �Tv%�� �����?_DB����o�aUU�#�[#�1�FE�4��sA�!GaK^ihϦ�?і֮g2[ȫ8�wK.o�K`���������v<T>�u����I�{&�e�{�o#6�eU�mV��7�K���e���%,PrfGL#b\�8��;�x�J�pղ)OF ��h��b"0S������-��~n}�܊ˢ1Ж���^��(�?�hX�E�Y�:'#��3���^Xl]:�>��������+���W�Gõ�3����!���u���D�!�lovG:ѐV����P��x3�/b��Z��?��XL���������x[�B���9��ح�������1b�jn��[�'�}�����d���]t$uFV$��o �o�Z~_���Jkk��r��-��_�wH�` ɧ��F����Ȥ�i�$j�B2�k�1�?�1G���%Px{hр�ǂbA�8�2���(��M�,-��(]�#��zaQ�2��py�I�	LR
�� ��ˏ�����}�z|�Z�ԼkZ��5����f�n�?�.�L��U.�	��W���"�����<������ǒΗ���`��^o��	�YƑ��s�����3��P�L0�a��*y�?bb�0��k��ǢƯެq�K�B�F&���?u�|�	�gM,)��u�$��-���{��]� �sm��^1���L\�D5�6Ku�U�/o���/���P��%t]��_�=�<S��ܭ5ߎ>L��Sb�����VWK��g��FtJ�c�&	�`� ��Qp��Q6�G�H��@���������Ip���|�&���ҵ�R�X������,=�v|���"#����^gy���a+��i:-�:aFI��cWv~�`�"=����ϋz��
�YFU^��|�	�r�l/OW%_p	���o��H����s�����o������&��;Π���� ��j��@BLb�8�:�VU���>A"�e� ��Y�AǨ0�Q�:�<�vS��6�Jy��YK��G���)�u�l';�L-Ӫ_��9UG7��2���V��Ҳ�I$��GLħ��^�φ�qO#7&:bAxTC*��"�ݶQZy�������M��:�������t��/���m�1��T8��eT�6�;_1Y2i�>9�k4��'1"F^F���./ӼH�O�>�NW�hnn��E�c��Q��
v:���9�Bcv���l�X}in���m�(l�|絅�љA��Q��?|�9��Wc���;×~�<�/V�aC���a�t��@+����� ��8�t-Q/bF'r� �H�=�4�V��[C�*�l=�l�r7p�, �@v�ê��,�z<�d!�&��dB���c3�F6�}�����"���6y����N�$?o��w�����bl� �E�h�A?�=����JY�D���?;⩂K4^������d���Yi�*Z�r�<���x���J�8T�Æft�f]ae2��pPT� 0JvԨ�҉G}/�ۛT�a���H��1�R��~&O]����5�P=贓�J�dcZ����'i��,=�?�c����c��Qd@��Ͻ��Lw���g޿�}�#>)�B}��k1�������j��9����ف$1)��Xz���[������@ ���	AS@�ʛ��t�	$g:퍐&�y���|sS��0�-m��b���1f��f���*����@E�d7���L���*���r�"��D,~h=v�_��F��<��:�<�*R���@G��8X�:�@�@��w<��B?t���u���{3O=¤��5���s.iW8�á�֩3�+���v��W���%}5�+ ^1�_�Y�ד=WZ)q�������I�1�w<�K���, \�_��_��_"��]9Ϲ9��9G��	~d~J;tr))9di�7�k��R�r�H��a�H[a�=Iv:�Z���w���hD\�C��O0���?�/�=�u�P=��#���@��Dvk#I���s��F�kǽ�c�{����h�WX�u�T���x�����q8�$� |1qr'�sJ�\
�4�d�.��F-�ՋAuM9�}?�9��K�~�����5��L讳~�q��Ll�P��ـ�㐍_�+���[��6�z�AP�D�d9囕�/Á_��е���a����R�����\RYI�y���*^
r�z�y#3��p�X���l����w�r�W 
4�V�%���h�6���3���{9�U��ܺA(��QN���Ï�L��XK���=l�)7�W�̉�{���@U���"ƴ��k�a�Q��E�;W�	s8�PY�����P֜�|UΧ}���/T�
?!����/���*s_ݘU���߶E�!���i<0�ځ�.����3�t�gP�g�H�����׌�kJ�zD9�T�mV��T8�� Q���(�I~�bY�i�s?b2)�KJ���37q_�EoX�=��;ȃi��.*��pMS���2��_�N�$�^���Φ�8�ۯfE2_���7��(��o_|��	������nv8�L`�"em�L^��f�Y�B�N�=~�v��ת`?x������5B�D��)ݲ1 �����D�5bx(�C�������A�Q���xl�Y�'�D��'[N���j���fޞ��	�?�{�*�~}��x�������ա5I��I��=��ӎ�EY��,W�ޘ������2!�t���NĻQ������$��x���~lV�%J��{%�a�+�����͏��J����QI^����
���X�7�a����d�ٻ�h�\.��'�^1j\��1"�51�b�c��_�c�h̛�g̢)�>sƘU�I3˱z��#mO��׊�����������u��_l��wQ�bs�����z2�|���NA�'s�ΐ0�͐�G�B������֎r��/�1R���~�Ҏ���l��f�"K[f�N�j;s�<C���v�o��8������N�<+#������@�BdO��ߒ����A�9|k��ۇ4 �<�d)����[�BL\��oz�pF x�#����Mk]�FUF��~�~ǅ�z����". @�����A-*'Y�o��u.�Ec��#�t� �1��h�V�J�Ui�f��k��za���j���&d#⺇����&��H0,�e���*[?�ˁ��J�t���G[R�jք<^t�6ĝ};�
*�/3v�-�X�n=&�n>L�q��4I��М��l��=p#Y�ge	D���
�G��{{5H�i��Tv���)ih��g�{XX��Nefv����[imҴ���@��'CSыRa�xIg�X~��#9���|�6ß`�2
�@�y���,�I9���E�h�r�K巘r����c��oO!�b��/^4U�)4'ږ�C��E�X���޸>͖�_���A��K��Q�s��1�o�Uߐߤ�{	R}����X�4�:iijbZz����Z��x2��Ң/�.��z������]��2t�X�>����*�Ji�K�PW�C�HY2��ih���՝*���f�7�_�[Lt�'�b)]*�+��%�
�=\���	�R���.�]R�&��rM9��h����<�_����y��p~)��"��=������b5���]k�z�Ł��Uy{·*bW��$�ԋa:"�?���<��R���̑��P�J#��S+�/%$�A�	q�|M�K �c�eG���1�YQ$)m�F4Ўz���Y|���3T�7S��İ����Ƽ�a������L��ﱎO���:q���9_�aʯ��	)89@i�����I0��-� J
x8�R8�m���e��e�dN���t�/�A����O�5�Oz�����H��58�/��k~~�!�-��a{�è���pK��S��Hj��AV
j��Ԭ���� N?���=��Łx�õ�W"`����5���ˠkm�� f��O�JVj!P�|5�=[k+��?X{��Ֆ{��h��Y(NFQԋ�u�`��)^W�-���3�X-R��S��1Q��:
\)\��^��.BĈ�ȶw���r��C��]��M��u��M��G��a"
R2.=o�Ka�Vd0T�I���#�*�%�:@֔�İ[2 �������ہ�c�I�Az\�Z�YqIC�˸7X�Q��R��P�4#�K�
��q��ռ����Օ�n^?��;7�-N6#Sٞ8�M�V�Ϳ<�U�	09�w�t�/&?�]�v���1l`1����|oX5�y�{­�����b�8̀����y�,Oˠ�7ޤ���¥�o0��[��}f.�=���>_��*2�!;�yo�����@תA��a�BG]�a�F�+OA#�i�ٕ�}�^�9,+Р��%=�T{�,Uɔ8�tcm�r���Y!�).s)�%�}�� �8yy��e,"�6J�y��ኯ�&1~�S�q��͕i��i�'(aB�7��*+���a���kOQ׿�i��k�������t������Λ��丑lw�%̯}��?���DZR�@(�c����D�8��\���vs�U/��υ9n����&�����L���/�L�vdv��M�!�_��2kt�� ����]����Z)����=Xo;eЏ�d����\�)���	��]�濢��ۋǮ繤���&�����{�
����+,�J���j�K)r������0{�8��\#�'ν��S�rɦ��k'm��5�p�C]�]�s�b�%�!�����@|*�#��k˄��+�{���"��N�ߙ����ŻT��v6BRxv�U͌��)�[BF@���3_�Ӓ[#����}N�^O&ͺ��_�̞�<��Y��EQ����sR��F���XG#����ә�TU-B���3�����x7��y	�=g[��e���>�F��l��>��iI�*��Ɲ�rÉ��$T2,���
����у�V�����8E�hEh@%pO Kn 2�Mx����6�Au^����4����O{���V]5��S�@�ڲЛ�	8��7�Yd׃���K�7뫤�e�λg�$��Y ���x���x�	f��{�1>�1���#�=�븄���5L�H+g<�X�x��b��'��}�U�i�!R����^O>��S����d�)�~���W4��l�^�ln�8�/p�z/��u�INlh��ޚS�V�꯬p��yR�Mr,̳�)�g��(P�3���m���XL�M�B�J�����J>��c����o�Ec��v����/�-����I#\�)�'�=�T������T��_�܆�'c� o�j�345�x5-���������)���}�g��1 *.��5j�}僷��2��C�U�Jg�3�������Tr�n�BA.�<���	�vC��Z���8�����n��iY� �7���9L�(�+�a��r+�8��� =�_R�
��i�p��]�W
e��4�F�/��K�X�p
{���?Q�j�����xZ]��6�e�uo��KCKBI��h��ob��+n� ��?��!����|��i!��iP_h�-_rX1��H��Tn�ώ���DMv������� Б������w�m��*����c2�͵�8�����}N��j��<~�(��"ܸ�i���$C���b`�%k��D2"�qn�~8G����Ӛ0؄�s]J��eh5�."��w��u�����M.�|U�0d Q �@���X�ǲ�=/�����?�����C{Y
,⤸5��U�y��G�D�����j�E[غ"
 �뵢����p��1��1?��M�%H ��)������m�x��)<��K��[ ��C{��D��|�sOˈ���U��;ع�#�[���scW���qc�P�ӧ�ۚd�Nɤ ������Ʃ��/p/�&�ɍ]��R���G�)��N8lZ���#N�Ń�4����\�
&a� >�(�E(�	���k��w8��$���p0��n�0�`trd���;��/92yI�6h5���sy�����<X�J�鴅��^r��˚�ŉ����!������S+7���9w�趷q� >J5í��J�t�]X�]e�����2O�u�E�.e
�k {��?�%�*��^��0?�X�"��8(a!����t
��T��5$���}��Z�X�$��-����̗����'{二;�/J�?�/*��9G��'~u�+_S����M�&T;nF�ݽ[�?ߘ_$�1rq��v2�G��~qX(`&��0d��x%;|�����wc��;�Q���L��L(*�����V�`����(��#X*���-z1���L�sf��>����Ep�w�>a�[�(��Ⱦ�"�S�(ǟl�ġ�H�r�G���SE��qz��5*���ҕ�&��*�'��zFb��ߛ��7	>-GY=����%�+��3��t�ߝ[��!8n,�B�ȡo]��]��t!x�#?6�x�o��T �Iw���ނC�J� ��S����� ݚ&��~��Jzٳ}��n
�:}~=ˋz����t:ɫ�O����'U'P��R5[U�� �܏��f��hXퟣ�Ph����-tw:�lψ3'�|B�
������"q�d���WCc���L2�[��4�fAo�~l��c�sǕ��&B;M�z�Ċ�}p�y�\� 49K�.��Zx�~j��{�]�x>@9[k��z��R�՚���G�&,d����;h�##W�������ٓ�7�煷d����^�U��
��}^>�H���B��C6��l�G��������:f}�kXf2���fa�Z�&��Fv!���	�Gl05�S��N����q�:��F3+�{��u���&vSwJD	�5)�$�j��δ�e2�f6'3Q⡩��f��X�a�������6U���DX�M8��tycxO�R�Ub��^��\�,�,~���܍v%�)������x#�������e�x�(2�����7Fi���_�����0T�$R��;=�\2�Z/;��`��L�i����x�z�\���1�GW��������{�O����&��?R|��nMy�)��H�:�]sS�MW��5L�P��RR>R�YV�;�Lp -�I��,2]%,����qK	&����k_�Xc]S�h_="�]|� ��Rd�,��uS&Y�/Xv�A�Q������ΦoF-@�	E�Yd�lHwm��M0.��[���zF���2��M��FV�	A�����$���ǜ���0_�f��
K��ݞ��6��������f�O�]On77(�mG�G��Mz�"?·χ�"�b�%���&?g7E���ε�;V�p�����೵��SF�(�Bw�1GZ�h7p��x)F�s�ū�}8u_����`2S�4k�6���w���f� �:��P���?�<7p
��9� ye��Dhi]c���Ȭf&��=T�S�9��)�FQ��0�Đl�h����ݟr��V��>�!�!���qv�����@�o������\[���x[��9��*�]�
�x-�Ǡ�a[l�n
�����������9���;X|��������������������V+I��l�>���O|�j����µu3�U�ԫ���МΖ�����c��!�y��p�
?��Y�|�NG*�|o����E��I�p��m���f*X�64��{|��W��@��Cg��^#�TN�)�%h�a��5�#�ܯ�TJ��*w���64��5-MK��mA��%�ո_寅$ߧ���T�+a�	"$&�
iR�6�mI9G��O
�׭���h�l�3D?A+p�@�U�|]'<!c6��o�|�1�L)u>x�(�T�"SJ#�Ty��3!�R+�9}�;�"f��>�*���Bm}</f��>��m!���O C��q���#���d	����,9B�]��I"����rh�4�o���X������t�@������v��m��3�c��v�3�����7�Q3�{-��?i�N��v�JR��?��F���T��{)E�F�'߷�^������G�/���)�]P�1�<��� ��Y��=h�#�K_j��Y�U^���ԟ�%)����q��1u�2���,���/,3��9̹�:Y����r~�f�lt>��W���ݜ�Ax]���]�0'����zw���&�p'E:�ܵU�O�^η���~��~ը������$e�]�R0���jK�'�e�P���x���i�^��_�4%4"�#�6`�ià[էU2�E� ;��[5#��u��E����?t�Vb���P�tR�~����-+���u����K�ϗ����q��Q����|=�R��%Ӛ�F#�_z��'��ކg+�_��v��`C'��{����[�'˼Nk�~Gk3�	E����n"�͓������.�R��p����el2��T	��&FD-,c�{U��$׳��<�ff�)�tD���c�ET�
{�*�IkQ,�u�h��z��p� �[63� F��ٚ��l�[�����
�~��s�S��U��\�N����E�z�n��Lc�s� �<J�W98����b|s�[�V!\I����I���\��؝"%;#��P���~ll�	P�<�G���GI�J��o�I܍���?�>�d|Vh��M���X��>�&�R��}\��m�6�~׾��=�l�HOZ�e�'���<���kC��^
�S���Y��Y[ �}��B��BF�U>�Vd�+�����g�6�d�z4Q]da5��4�vn���"�M�N?�<��Sw\�s~#��~G,`�w����x��~�:v����3�GRq��%,dt.�@��GU����!U����č�~x���Ԙ�T@(���/�� ���ok����N'�Q�#s�_��[�w����ոfR.zÈ	��J������$xc_PD�ֲ`��5�����ւRq���~=�;�T��k>
hl,�88���o	�·N��r��m�c8�}�@�t�B w���o��x2q�������.w߭5�4u�&db���Q?]I<��n;�?�3�P~Q�J|�r+0g�=ۗ`CM\MC+q4
ߴ}KQ"�$�Ȅ��:���K����t
mv�Eh?����K��@F��f%V��8=��!��g�Fc��
�=d(t%I�|�,nð�/a�(�s��Yn�����i�%H9�L���,�'��4��Cg���3əXE��zDQ�d'w���O�aVՑ�Fǖ�
�是���&H
a�  ���v3
v�0r'`�GIgW_�un�7��3��i0��4+�=Gv��m�s�9S���4S(PN��)j��u�%#d��p��OȯqT�ù����J� �Lr�L�!e���ƣ������DO����*A�<��Mh�X�x�.ґ^��Y>� �,os����N?zs�{�Ͱ�=:�����|�ȹ�<0{�z��{�9���3����K��t��,{���Y;�lkBv^���ߟ�{�h�^0�d<���� �2�K������n���=~�Y��[t���[J��D�Hx�j�'*S�X�w_��ǘm��G����f.]�X��H!��/��|�C�9����S
��j�� {�epb�JX����|lA�<m��_�)�}aѲ��5���rC��	�?C�}�48�tT5k��PXϴtT�c���1<� 7"FB�֟�UB����F3kZ)R��H+`�ߞ�C9����M|��(�Ԭ��U�$&�R��g8���M���f{���;�c
9�P3��_�	>�����\ޓJ��R}C����<%v��W���.{һ�u5-���9t����:PUѶ2|��`0}2�q9���'",䈿�[�Q������(�\�����tQ�\۽xv��A����@����K
	χ�B�{xW��م����%̗�E]f�ͭA(Xfߥ�E){�}S��"�A�V�F�C�P����䑲� |�!���LB�������mc�]�n���E���r3����PBP����mȲ�jr}�a(�=/W�Jdo<0����-ς�Z7�i�=�r��:�o�[/�o�@n}:��*؃.[�2�*�1G�6L8�#�6�,{bH�V�P����:�D����=Υ��s�G�A��t����0�+��.��>$F)�&o�}����:�s�' G���l%���c�#;c�������2�!=��hdt���J�NM�'�=�S-ax����[���|�=�_����Ιxf��ݭs[iW3���S��-��T��A��VY�/ߕU��U�+9�t�9�?j �%�S���x�d�`�f��Lۿ�a�&��nT2%w
�qF��1m���0x�êB� A+��^E7L��[𱌟jDW;����%[4�_����zo�&G��@��7ÔOw�h�w&{���U�`�a����]#��.�u�
<#�!�x]XO]S���m����A��X��)�m�9 g�{�f����Np6����L?ep�f���%xu&T�sœ�}}:�h���ѧ�T����Q5G��~�$��3�^�ȳ�$z5g��~�o�
\!�$Ud�v`p��(�ru��t����j��l��\��]pZ������7���0�^��<.�9�������@ׄ�݈~�{רt����T���(��/�����/���O��������u�Iw��;m�``0�!G��p5\9lDl`YhUl��s���$+��ڋ'�T��4��w���k2`g��A�=�G��K~x���7�/��҈��������T���-5���d��f'�����¿���D>z��1�^-<y
���v1�"���$��(��0���d�3���ӂ��t(خC����.Ҏ�gp���yN!���g\�e�I��$��%�R��Iղ��Sk�=ZmqP5����}T�_!�lr�kO+x�lsx|�K��p�I|&��U��t��|������S���37%�����K����2K��N���^�"m�x'-�?�pf^C���[�S���D���T�9qI����}V�<���C�:�OG�M:L�A0/7�2룭sJo�o��Gfb�[qeE	�o��w�u� 3�F{.�H���d�2���d��h��b�6J�ğ�;&%^6��ş���_�����`,,�ۢx�61�U�b,�V�������!��D��lG5 �&в�l� J�5(R(��(IM��H�ѕ�4$�{�w| ��v5gv��"sP@ � ħ��(��0�X~�[B>�}�9�=�e]������J�g|���-���Z-���4��k[zPS鏬����ٙ����
|������&3��εǨ��볠��ם�wfm���[�l+~r��~?a±��?k����3Kr�_Y����W�y�� �b�/��UV��j��t�J��3��|RP,���m�E]��Z�r�%m�s|.3�ƫh��=$�d�����������'p��[+C�Έ�W"�d�֌��"柹&���N�d�+m�\���r}La�*TwW�P$�%��;���� ��x�	�\o<�Jĉ0�qͨ}������I\5�/?$	�.X�,�ݘ�l���4`&f���㰊Rg��n|�����f���5?d����2�D�����C�ZL��II^�yF}c�L���9{�$����<��=լ8�y�|�Knn���W���w��g'�^�+�^v{l�j�w3ϰW���g_n�s:��K<����Z�n8msVk67x�#Mu
�x����OH�M0���ЮH�~�.��J���}��{��l;A=}���� "4��I�̜�-M!��7R�Ռj�"v#��A�̧�pc���}F�ڜ�`���-��D,����o����"�ȳ�"���C#��Oh彨��!\#9�U��֔0��P�����,�dr>��#���Ś���|Թ{���3R��+���Y;D�+�N|mG�8D��"��	{�����ԍ��Ϣ��<�Bq[њ��У�&D��D���;!��R��*�u52 �I��Y�m8` )Gmđ�!�����-؞��x\����K���!}��,���ŔI�l���oWv�t(���u���L�`ׅ�%'�v�D��y!���k\.��Un)���ж�j�*��.#�1H�aR��3(2�n��6��zA�T��l���	��#ZM�]�w�U��J�f+V0���s�	�-��zV�����ڥi��K�1`ݻ�tϜ��2#*��7w�:�t/YF��L�@y|1��S�|t�aL����"[��Z��C�.k(�O"b��9��Z�-�b>F���\�n-b@��a;-z:8�nK8
��~
��fB�D��p�J��Fᷘ7]�����L�NDx�����ȵ�A ���/7����Z2  ��&�8��r,4d����S�=��t�-��T��̵R�8_��M��S�pPsqRJ�=�#�\�"�y�ÿ��yIm�9�nåk��i@ �����GYH��*d_? X
�둟�/l��J~TQՎE��`Ӵ�:Ļ�u��d��*��h�ډo��m]�]�.���Ԧ�0��\E)4y4_E�T�+�z�G�����N�C���vd4�@� 	��Et �&�/�L���wa���;O�]�Jn��|'�N�οC��2�N�m���]yi<Y�W�������ᆦ�~'P�Z�\�T�vt�yX���?�+֯���ǜ��iZ"~�5RI�)_j�I���_Q}���	�Q�*�3;�S�*jS�x��h��yǱr��d|�Pf�`��5��%���z�\��vd�On��#Ԗ�Җ�+��LΐC���P�?O�v�遉��l�sJl�mE�6�PFd��������]�C�
H����C�X9�c:�e(f8����x�.C���w�e�'UU���LkGL'�D���/Tc�Ć9�+,��.�2?Ϻ���������Z�|b�\N�h�k9�`m� \MV:Uf���Frż������jfy��!��� ���eRVX{M|����A�������b�m~��D� ���
�U��Y�MT��@_��H_����~��{�_R���~oo�=o5�Me���}c�x�s��qȸ��3��Z�K�2��k�ޖ�~�3�q�ġ�T��9���>��tU��=�F+��֟�#�v[]_�������l���������;�Bī���'b���iY�z��A��6-m�#̘R� ���ߓ�O��wA�oTq���]}ʁu2��%q!�:~WR� Qe*��X��Cm
%�x�C�XI�ږ�gh���,�fBʯ�Ȭ9�I���T��̴+1�Z�ѿ�֞��rZ�і�k��6[$�<�W�����r�s??Xv��;}:�<����=�d�<�{O�����t�0n{��yEl�������ts�t���+�����WC=O�B.�q�'���T0��Ic�	����6/&�P��}�l[�O$.�j���IHy�܇��Rʪ�Eɀ$p�����\��Z�8V�^�>�6���J 0;�[j��]z��W�
A�ۢe��'۝���8���J���m�"j�v�zK�=B?LŠ����T���A��-��'ɵ��HAu\?�.}R���B�ħ٥E_D�`!��y���S5�7B�\��r�������<��鉉�Y�� 5f׍�zN�Ί(�ÿ�==��N#,ε��z�@���ۗiu��f/W��2^6�N_�8��_�L��|���>�����v��Zl2I8��׀��O�G��ɚ��}��]��M[W;�L��,�?x�*ʚ��K��ف�US-G�J�/�د�؏�:�wy��a|�f�`�&fc�	N�}��������+d�o�#��(*�� ��4�_��Q`!O~�.�hgr1U��>FA@��=��N8�8|���M���|`0VDu�<\+���=�J�^v���P*��"aDx��7����ȕL�Tݞ��N��%�<G��=h  �-^�u �8��[@䁹V�:��=p2S�`�mO7�h�*-֯��V����:��"v?^�C%f	�a����.�_�x��	�k����4E8oj�X��{a�e>6��5�Sjp��*�آpI������H��� b�7��e�"b�Q--�c�[���7R�U��¥�Dgv1\h� ̀?x���F_�ݗ77�I��Vl`���3�D���^5Z��W���J\��2�}�]�C�	�B!U�At��_�hN�;@��3���+(��=ׁGrܚZ��O��=�eER�3G}� $*�A��Mح0��-r)h|(���M��N�F������z�qj�HP��l�Y�m�J*�&K)voJI0+"�e�����;_R!JW�{��x���g>��NGǥ�Ȥ :���b8)D�ˣ������w��i� ��W�8�w�����4�V~��Gu�ve��vq)Cbβ��O�l[���<v�Ĩ9 8囯�2��E��%�D����@ʑn�S���dYX��=�V7 ק�JdE֕�j�ڕ��' �{	��!�I���(��� �Z.89�Ը���OK�.��M5dÚ�UIE�)���Z	ܘ6�� �!6��	������{��� ��>�g2o�li�$:ag���ē.b��sS�Y��.W�)`�5ۯ@�����V���F��j��rG*=kk�p�ȩ��f,�Hm��a�328�{
�>�º��~W� c��������-�`�X|�`C̮��1N���0��4���a��dq��3��S��c=�d?���ʱ��	F'��JN*���?���f&��f��F�F&̆��Y��8
rK�݊��"G��9M+��E���`Ӱ-3p^^~�a���Wu!�Գ�~V��w����s����@FŦ��j���C�4/�#�ӝ��fqah��B�ot�m
��1����i�K���2OO���	c'�zzt���o��8Ǘ8�S�}$�#�Wr��Ȣ��){��-��p�"b�0�Q� 
x�PY!�o�Q��@��8�~<݉?���n�k���_�;���֬���xg����|g��'^a�xs��m_��J���!���t�R���xh�����8�����5��h����ϲI���~�`�'����H���Y��Z\���8_�ȗl Pn>��n����W���8�����xi�4��A)����dn��KyAU��1�1U]"����u�������vA���x�u��^��<�Ӥ��qu������#y�6<�mo�l4�m���x����5�m��$��x�w����|���:�}�����)�	�i�I�@{۴Q�_� Xp�.i�>a�!�O������P̀���������s�(>�����x�W�L���7�Zk�x���!0�AT�~����� ʨP��~�"��V�U�m³����ԋC�6��t���ل]�ܟO��ׁ7��zݎь�������}#�Q���"�q��qF�;��;���B�z
�ޏ��g_�/���g�U�ڰL��4�������F���`���䔐�R.G��E"��P�-<�w�o�WT��A�:D�I����Pt��3�ι��T�H����w�#y�v�e�&w7�!XjW��&7�Y�A�T��ar)AqJ�x���*�lp���;W���U�����ć��Ǽ��,�hzS�}M=�M���.EZ�F��=����O��d��� ℺�UDM���{��M4�����$���K��ʯ��|�o��~s�ג�lv���h�]�����
8�w�8��L���kl�����ay�-L�}j��(�2`0=��n|��r8�mt�y��]۳�wp�����8[��Ͻ~�u����תߪ}�K���?�8��.{��	��?�9i��[��Ab����"�g;!Z셺�k��Q������a%�u��{@/-�HE�F2�
��b�sp�#�N�Ŵ���#v�{�SАߢ0�@'	�:ZUھ��c\_�����|��*��Y��,<̅���J��=�^d�ӞσQ����Q�ȅR��)*�`���-�]x\4���s������G"�'Q �s��ʑ�V$dm%�Xڸ��V�Gg���D�	��C�aI�a��&������#�Y���U(C�T����%�C,+�W��md�����W	ݥUZӀ���$�i0�7�,��J�� �8b:zy���~�SYx�E�C���!�k� &%�)5Ӈ�[k�1M�qӷZ��(�k3&X�v��[��r�UV�H�m�,5����N�ٖFx|�0�GD��A|f"͑��˞��ˮoܚ�jw�c�GP�O&0狞�PDɚ0O:億� ,�"�*J���N� ��;��S����qb4�'�ɨ@���4'`���~>Q �1U��D�0L��ʆ�"%�LĠi�7�Eu\�!�j ��8DH�h������O/�/�kf�B�7��ς-��g�_�䦕�S�#��0�s���z��u�nc�� ����J���N:�q�Z�Z̡���O�T�1e�ǆ��D>!i�ue��gՊ`G�k-�6�ԃ����U�ĸ B���
����:���bv�D���r̔���4�K�<��|�E<YLM;�/��%�����E��N��Q��a�C/�v{�Rc�Fg�Bk�z ��V�f�z��D�F���Fm�D�=��#u+����ru���0��:H� ��l��d�<x�n􌵫t�����Q;E�k��d��I�˳ڔ��[H�`�t/�69�	|�=�|N��sY�_A��2�~N��z��Z���4W'.;!�;ש����۶��̃����`hY������Ҁ�Ä�ū����£�ƫ���������ٞ�Ȼ����R�F�d{���L�Q,*N2*Z*�^P���έͥa~\L%7�Mw���B Ģ�uG�$�+k��Ȃ����ND\Zj
T,ġ�uͪ/��6u,�,����Ů��;VW�hZ�Ζ������M��4�E�tpٵ�/P��'��k&�Z-�:1o�L��MO+)N� ������v������ "eɗ��kXe!����v������2�ZI���ޅ��G!��''������=�7���N�&�����G����u�<@�{�{������F|��VU|x3Ii��G��3B��s�kI�j�P��4���ޕ�W�a�
��\�����ŀ�:`��3�Է�� ��K����gZʂ�g�ٗS&�V�ݹ(,����mj�ʛ}�{�2�_ދ��㘬���S����t�d��C%��kCz8�.��9�7�)�FO�قq�V>�^>�-j�7����X�Z|�a]V��*U�R�_(�X �v�����l;�����%�O�r7�}FM�_ϊ�"�_l�W�1���<#�<�+)q�+�k�����x�^#z?v�?_Cf��>�;[�,r�$�2��ni��0�\XrVWWU�v1���������z(,9���`����q���+4�����W�&1S=�@�Cv*�^Ɂ�U�T|՚h����/��ma2;p��ڨ A��,:��t�6&R�N�@�i{ݬ�u�w�Sƛq\`ve��0u#,\E�Gſ7f�:�9ڊJ�����|�����f����&"����_�ֿ�%���_��y� �E��ų�*w-���{����n������y|%N����j���\��__��j�k�mf�����N����F��3������Ǿ���Qm��g��Q��a�@N5�̽��������f�0���"�������Q{�]���󥺨�(���	�������TI��$s�"L7�7^��#���Z�9JU��e����bu@�lܾI$�pWy1ޒo+���χ��f����2r�=ӊ��^��"
6��krs�&+�.���^;�����-��]�i��Ow�S�;��v��R���t�j�03����n# �7&l�b_�4n���#rJ��N�b%x"�\���2���L�7���Wnm�n۫�CD�M?�� ,\�^'gc0�O�¾ �V�V�0� �;����
��|r
�x�#��q�%)��[�\��b�;X��&$��O���[��4$�,���5Fq�lN�ޞ���9+ǎjy�E�й��0+�u#�y�w��D�� ��WJn�]ð�&�8�弊��<	���#�&����l�\ XAD[¹��*��,�=��Ŝj�o6�R��#��ծ��)�sF�K���徆�{c�8uǏ���^��=pں�LJ��ܷ�cb\X;9y�x]M�7Κe�����f ���=f�`��"H�抌�" q�h���!%!��F*�tqg��v��`I��p.#���6�Ku�حӁ����
�9�?�M�<jz�F̂S�A�A�:栂,P�Ғ)��vn3������#d"E��"7e剡��?9�J��f�W�A0�8˛�K�v�a�}������)%��p��F��uޝ%ʹ��K%��D0a7�)��vh�jSU���ĆTiJ�\O;F��7����=����w	-��/���(�8����B�߆���GTϺN�Zf�Jb���NR�6i�&F�.N�z�&�ќ#˩l�L5�\%�L5�-H�.[��3[Ǎ��Q�v��r�]��`mG�pL�2�;|2�1}�Q����`�<��qڌī8vIDm�=��E��Wt�J_:�:�Ȋ�6Ɏ�Z3'~�>N������M"��R�[���V2H��z䏛�Kg=��*9�QF޷;|���4�D ���H��������������������?ڏ�G�2��ic��$����J!n�]��T��!�Ӌ�F�'�o�8��eG���f����eM���p��8S{
���@'(�ʤ��\��ܬ��N���,isz[��QO�E�?�P��s۷
��T�;�@x��4�y���h��l���i�����y���VbgF��e���+1�~1���8�NC	Dh~�h��fL�fjk�'g|i|ol�`d�dlvcv%M�x�i��a h\��'�ƿc���S�v,���8Jzn�� I���9�9{��V�	�>�=na�)1r����!�v�����@uD�����%���Op�m�X1s�9�&�W����)��-��pp˞L�onݞH�pH�?*���N?�Vy��oܐN�@&���.rȀ����oSH�'<f4>� ;��U.
D�&��9%R�L�u�j��j�9��`���G�--��z�K����^.���¯w�hB���y~#�N�ݍ�B[�z=sy�1 �臈���+J�
����2k|\�f���?p*��٣;]L;f�R��[8	 ��U@���O��aPE²�/ruM�j_m#��ȑ}̗v 4���ۇU](!�)y>}w%��xL독]ǂ�>�����,0VK��z�w&�^�ҟ�����ɧ�G<�ϻ�_=����ߧ��;}��>Ά�K�3�3Q1-?2�
�R�1��vSaݢ��Rw�T�M�{�v��C��gT���J8�H*-�B��)�PTF�U͠�ԋ�x����� �f�6v�C|��L/��C�.vVh9{Hw�u�3AN�o���F���y7{p�"\�'��K�yUOͰ�?*`�zW���ם��_�G���gB��8�0�~ө��:���51v��Y�m���r���[[��������C.����rr�C�B�$��R7z�ΕN���G#��k[	}>wG|~$G�	�=�}�X�t{�����Z��Ϝ����u��Xy�u�����$������\o���eC�/s���W���|~=�=��ri1<��Z�F��r3ͮ(1]��9�)2MD*Ƣ��geC�gOs��u<-X�2�fT��%E�2���%#j�R�~��r��4��c��Qΰ�Dt�J���@�@�8��1��["�̨��Ri�d\�R1�6���B�f�n?S��$,���7�a����!�M�'�3���s=�S��*v���/���i_zLL��W8R<����6�r�{�7�Z	�Ax$�gw�^�%���h+�b!�l%�
ν����:$��T�bN V�Ĭk���Q�f"��������_ �̊�"��5PU�ԁ����A]�"���{t#l�CD�W-�o׼�����;�ԉ�`Ϋ�mP޽G	���E�=4u6����FG{Ɍ��#�Q��"O�>�U1q�� j�X�nu�B���ǖ�ZR���k��m�����z·�	�{l��������q��s3�'Td֗7�Sw=j��э)���<pon��V�u�^��A�<�7:�"%	���@
�!Dkw�ԑ"Q�31>�j�dyp���&2b�,�?ƟX?ۇ���(v~��������F�P��䠳��8������k�p1���
\9��_R��g��$�N��l�هG��`p#1Ѝ��҈�x��6ۭ�?��g��y�(K9��|�|�>�>�f?B�7��g	��E��Ό0Uq����&���A �Ft h���J�ū�N�2J�G�����ˍ�=�DԞ��kJ]�(^�����Q=���s���35�2�Ss2RH1�-�d�؎3M���{�_�e%1��T�_#anu=�˗�]�}�u�y7ğe�}bs��p����5�0`�ǧ]d��#��B-�L������������<$4��}�l�9�y�yLl�����|��-C�J������o`�`�����e����9�T��fQ��|Y!����ՑzH�oɃˏ�;��z�nfp��,{��z����̬����S�-m���;X^�^xO�y?�,-Q9NQ;��N��p�Ԇ�1�.��|+Ŕ�*v�f,��-�8�[�U�6�V�v���UR�#��g����8�K%�L*g:���ʺu�и$�3������ɓ�L\��Ǯ��7��*3VY��o��K!-3������_���>-L����|�^��y�p�f�>�H��(x@�9@�y��;��?W�g伂¼
FUD��"TN'>H�~���
<r�z�E�z̜����K���g�����_�SF��%�SNVG��#�������4����a��Z�]�4�Ll6��uɯ�c�d[���\�g�7����P�,$�([B��N�P@�s���L�sx�8��- ������Z%�<� )}�N2�/���x��癩�����<�=���Fh��Nҽ����_E\��K�>^u���3�ED��~S�>�^?{y8�_*���/����4�I��:�:9�VYLS�7����5;%�,Y҉N[�_ՃE^/��q��R�}$�2�mn���?�uZ��}j���p�u��^T�&�qW�ϔ\�U.6��/g�����TR�G�G�q�X�[ζ�8;�^���n��y���
�;�j���6�5�{��:�w�bflhd(�RR!�B�M���|�B�pIȋ`=��G��a��K�Q�K%_:c�� �ɖ�����m$n��,��b�d0c~!��-ǟSz0,g�9ɚ���
Ȳ
�f��J��	�lz|�v�Fɾ�a�R�W��� yL� z��}f���(���sL��,l���n ]=GĔ�p�j�KMz��5�Gih#j���M�������r�ƮF�f����7_��'r�γ��[���z�;/��q#:m�t������9m��TޝH�]د�-<�]w��~�.�cy��Ms��{m��7��ؐ��9ٛ�C˩M��I����6��6�@�q��Lm�j���e#~-8m1x�-��lw�6w������A�dYhn�`z'w��5��=:�(�X�AW4o�!�K%>�2L#$a~��sv��F�E�6�z�)L�N������j��-�(�sh T���hG�E9�`��o8J\s�ጵز+���V����{Ty�2~u�:��x��	77�ɴ<����"��A�+73_'J���y$��E+I7n�L�4�]�%�.k$ _vF�H��Di�T�)�w\���t��t��f��vuq*ia2¤HFgal��ڰ�#���tzXT�w�7�)��I�f�k���hi��	e��f$*P��G�(]1�v<]1!���Qr�:^�;�oz��"�%X��B�����As"�,B���M������`��ǏB4�~ZEiPUKO�̸�YV.j��p�r�E+��m���g�i����&���N�L��[��'�4O�k�zz����c�Ǫ]�k�y��v�O.��=>p��e	@)�lI�#�c=�
�#��b�h�r[g'=�WbP}�/) �ƵN8ĥa���GC�|����+�a���>-t�� ���ƋH���3��JU��ɐ.��V�F�Ef��I�YS����0�R�^ (yB��N���W�l�����z�%���pb��!ɗ"�0!���!RaZ��L��Ρ�`�dǉ��`��tQ���w?z��
���pz��]���}����x�2~綶}^�j�4M�� ��"�f��d�O������L�8�(���ߕ�Xp0��w'ʥ��ۀ���	 �5��VQ�Au�)�����^ha�a0�NI�cjÑ&�2��O���4�,,�A������:U9��͠�1�{6Cr����������	&��DU;	 B�$jH����������
��o�12B��0c��)7��.�	�.����	3�q��	rM�f~�O��OFs�����_T1��{
 ��b�t�	�S�^�~������~���}�����M�պ��Hl��"�Hz[���������5�;�Ƙ8�K�<W��ۋ�ۮ��^��<��>n��Q�Q4 �~�{c�|`�}`]a�Lao�|�?�ӗ���tb)�xR<s��
Ջ��������U�	�e�v8d92J%54M+�\����R�A�E77�^Y5�5�s�.F�Z����	��7��г�r3u�H�!9a=,T��'"���e�������)�gȊY_�^k��ڶehC�Ze��eg'��,�-�@�T,|D�p����a=8���ɯ��}u޹p��/�rjv뽜��t|���y��}�FH܆P�3җ+&a�f��W�c�>�z���4S5k�E��:��Zb�!�.�&�4�V��D��(�r���9?�S�V�R�l�d�3i��~"�1�d�G:���sR�r��K�*��k!��t,�L�(�v��v����n�o�~��9�!ۣ=���ȵZ\��o\F?�w�==Y��,͢b3?���3�YTřWŁ�c��q4��T3(�U:��^��c���PF$L�n-M?l�,ԋ�_��a�1.����w;A�l3��/o&y��(8�GV�b�˘��-y�6z��~[ל���;s��0��n��}_�<:�S�����;@C���m��:�0�Z�}�Sck��a���������_�~�[J����[K�jݕ�����ՠ�D|���8R,�����)��(��J2a� �<��e5$��@,ь�� �H$�X���/�f+\�G(f�{ė��A������\A����fG_1D�s���n���uj�{j���/yc[�{��A(lGc�>��'	��֬]K�a�t�C�gVA�Sq���B�s}@�-Ť���S�Q'�N�.R�ˇM�ÜE"�=�{�|:k;n�x�֑��8L��&r�J��_�����q=��-���*�]���%�:�y��j%�j85���;���5'���v0�I���/��ǂ�5�F��Ǳ�������6hy<x�ր�t�ݖ���mi��i��������	����̼�n����˘����Čܙ�Ǖ���울���⮔���9Vq�b!9,��lL���崗'ۘ0RbQC2:�*\g^���J�@�~?�A%:;��a�Q��>��4���L�dӘ�:V���s|�����*��)��c���eBN�|�e�n�_(���`m!YU�pa��KZ���X?�����;�
�]��G��z��~<��Ӯ16�j�W\̨�Q~,�u��r+�u.W��U���w�Y����2OuI��q���/t�����N��v,t���cQ����:��DHf�ɬ1�u�RHύ�Fr-��T�^�T��C�;z�H�7�"�j%�f/�3xd�͙�P=�)Q˱Mg�$�NcR���ZpkX'
*n��vD�Ú�=_�#���B|N���2�޴�`V���3�y�"���l�_�δچ4d����-x�|j��L��b��`a�W�p`�G�����:�6՝��y~M�%�;�6_"M!#��d��Z��^e��<}�;�����B�
 v���^�,�k���IS혈�(�=?1�3��Y�?��Caٿ3'�I��(ɞt;B2��^�����O�[�1쳄�U�H�>������KE��@���Q� (=�D�yK�Y�+y;ǡJ0���-�H0$��'�r2ɖ V�	ㇱo���t d� !"P��`��O%�y ����R���Ʋ�F��F�c���L��S����ę��_�a��r�S��yg��� �/R�&�Q:��uUL#�!�7�2j�Q��.�*����	1�ŇC�/�l�jR�LBߴJ�_�E�@��!UOTg��,�=�NF�#��>��a�1��
e�{ƉI%]|R�����0���k����j������O������߿O�/I�.l��4��)
GI�L��J����p���m�Q*r�t:�0һSZ7�a�?��,\k �'t���
e�������	.�q�w���8L�e���Q�k��*�F���p��(>ɞ�m$�#2�>��J�~PϘ8~!n����wǌ\�
3|r��x���?�w�͐%p�'� L��,Lmc��5���E�������!qC���o�pEV#��_������,D�އ����t{0;r���r�S;83مs���-^M���%����P�F���Z����<�yr�j�HY���FD��JH�d�wO�T�-��&G�'�A)>����ND���P�R���5���yU������i��ʿ�OR�
Ӭ.v���ǳ�B�:�q��Rt��A�j1cj,���j�Z���)v��;��|�J�O�	� ��2��eڭ伊�:��dI3$A~i�Bp�L�^�U� �� ��KwǕ�����u��O�&�:���܉O�x�L�"�����D����,(`��z$q1�X�+�/c|�9�UE�O[3�'s�>�U��%�ZU}�k���k�)�^�»��?�o�r�[��V�O<�mj����=�7�����"��k��7����*��l�-�L���-�J3ܸ�%�hfAXG�h���^�:��_;���އG��w��<���n8��	mqmer�dsn��$�p��]ج��>��.�P����5w�M� �$�;�����|}��_�S!�(>�7x;崇F��SLk��8V�gy�A	�AŒa՜�����P)��	fW��u��B���O"f�y��D��}����[���<�ky(W.�"6��d>�u�V!�1a^��n�`�&.��\�Ǒ9L�n��	=���~�|~-�� c��X<OGG%R�XG�?S�KZT��/>��6g袆mm,���|)O:�*y_�p&�P� mV�w�_eH�ɣ�~y�rE��;ܺ��Q���U�Ha!�c����yc�o�����<H�u[���n�FS�ES3����9dGّk�5�T	��視�J}ł��C$�����Ú��'�"xP��0�qOL�[�yN�Z�� V��0{<*E��.Up}����_�Y�O��'�[&�A�XmW/3M����\o�-��M�J\��5z4`P�9�b���[�5�V=�M�{H��v��S��=	����>���A���\���u8�t���R���'b�.UC��0��c�cfMKU�Uc<�ս"����Zv56Ӷ$Nd�Y�]�F�f����B��E9Ov�d�7�����]���v}�D��´�Gl���8}~,>�/��^�W�Y<]Q;8�8\S]^�\_�\]�^�oO����洷&7�f�ץ�;'4w�77'�{pX9Pz���Θ��������i�H�+ۑQW)caKG�V�|�A��������VYԐ�e(z	����od�aH2,i��V�$�L��x����P��,�W'�w�i'�he�����v�x�-	��*/�]/�=�f�߃�f[$j�����!jP���V"���'�|�P���,�ܥ��FJrk\������!e怘I�F�����<�N:[�����Re����EXI�a��I.Hu��������qBh�;���$�&>�ȾO�T�Qsʜ��&>�A���yb��Jl4��ng U��G�CbBJ:(��jT'$���@ ��,��t]m�@�n!�z|�݌��(��Yj8��O>��t`����!��EnH�T�H$D��@�*�	���9�|?`6�+� +� n!Մ�$�l���ه���7�q' �|�ȅ�0N��7F9�P/�E�_������+�O��fgT#��!-�=�q��vt>�lb,�J�����㠘CJ!��\י�͡&���H���I�����dP�ҭ�N�ת������{?^��丸7y��:;�56�G�%�K`F5V�H|�)��L5c;%�J��h�6-Р���BG�
I
XC��g^s�Q��[@t��b#�?u�!��4( �pF���g�>�I�Ds�C�EKv:�th%���叛��`W�|qws���pS��>D̔@��GU���F�}�<1��[�0�Yͬ
�]�Y8Io~Dl�}���Y%�p��`pL��b��%�V�:1�a�����:4��溷ۣ��l��X��4�:�a;	R��RLX�'R�&G�zd�ǲ���� ��7��F�2��&_# pV�F{��\�kq�m�"9\L=^L�yz{X�]1�N�`k�d�K�zd7-0���jK�3�a/[j*�h��4�����*�����܍)�h3XDIrB�`����n�2/�����R�LmS��q��P�P��I��k��A�eN��\���Vw���-W�9	Ė�x�!n��$�g�ҋS�$4z�vv� ,F_����)�ѧ�u��Rcp	�®9
��T��UGZX[�@H�^W
*]��4�;����M����Y%���	ۻS�߅��3~[4+X4�Ɓ7`�Uj�0*���"��OT��b����1*!랠SI{A��q��)�L��p<rD{o9��G��0��D��	Fy(~�(�h�ylk�Y��B ��
�D]���趇�8D��M��&]���I�������+��C+�G0@���Z
G��U`�
���������K�s�^�c�n`S�=�_�A
?,����v;�:�c	���N1�������hO/�7]~��a�i�4UB���S���kC_P���n`ޠJ�Ana��S}�e�W�zO3�h�xm���V��7��N�=z:0g& R�3�z�sh�i�+��j_0�'��OH�ls����dv�w⋿^��Sw-�?�Rkf�z3��3dBy��KҾ@�~��8$�������|��<���x�:x"9�6�㪟Ba2��|�?fk�mol{i�����t˰��dB���WpR$)�!4��-]4��� 3���c��'S�cgƉ|�ZX���h� ��^e����q�b��IL�@zg�뫽هQ�ӘM3eO��U�^_��	�/���G��\Y]�||�y��l�_g�0tm$�-�(*>.#��5���3�i�=�i�7�@ۦ��尃�}գ��t\?`�H��E�^<�RB�~��P�pȶ�cX�R�
(�l���-;q̯����D���v�C���g30�`����鸂wJ<V�<Q1����:���Ϳ�9�����}2��O�������pO��������ffO{��VRۺĵ V�P�&�X%9��� k�q7��i���'b�7�
q������p�����C:�}(P�7W�����@]�+����0zܤ��_�Vb�!Ft����{N"-C�Y���i�GC�J@e8=�:�J���K��
��Y��EhK����n��X(��=�ƻo������K�,�o &��[��Rs������}������Ȣ�D6|eY �:T��
�3s�ƙG��i�����_��Q��s��=�HӶ����k���5ȵ�r�N��٧]�͏#����;G�v�7��2�;��ôƻ�z5>��ǡ.jiqh��������
�}���
e�n�l�	�b7�ew5f55f���7��u&x:g8g�8'�wf6vfv����wv�56�w7'w��t6���esy�t�w2:�}-*�S}���`�Yg�]�`���9LûTC�g��N�BL,W�*z4lA k��&k1�ٗ����\WE0�(�{[ܘ4&R��� m�sNX�鸙��hY�2���V��Z4���K�	���:�U�+
)�)7���x!cV �}>!v�y��%jHl�Ҩ�5iTZJdD��o�Ĭm��%�����
�r������۩�>Lf��3�S�Djv�D�jnX�Y�t����(����rƌ� U���90�ɷ^��q�d��)�cO��_����0��8�� ���9,gB�+Y�s&�ƙ��L�b�U�jc�تqU+�(uPf)�fk+bca�Nˮb
��JͅD�s*�M)+����⠜]���c���1q���ڙ�B6�*k���Wc?�B���$3L)��� ��g�}�����'�e�cg�N�/G�E`;Z+;������(�$�0�9�aȏ0����`�E�޽�^�-Q;u��7a�d�{��Ї�5�94&�C��o>�0�C�R�� �}&�<e��<7R��������Nr�}Y?�%���B��	鏇��<<<;;��+T�+V+W�Æ���v�(���P9�UCT�U�p�DRea=�i��L.H�g���.gs���g?�a�)y��+�h�'�&L+�L�4�+��	��B�]���y��,��u�S� ��2�}�pՓkl&EzNZa�Ҿk�����0�#�}3�vQ�����
������<���p��/�K�=c0L��4�����V�iD��T0&U��T/�rO�1u��s#�B��/uī�5ս'�����1��:��R^��F�@�V�b�!R�He�����K!B�F0���f���C�y,�?�c�쐡dl:��� 	¤8t /�ǔB[b�'� D���~�d
�ngM��"R[�hB�T�Y�
��;ScS��Ej��r���|���	~��8LW�yy��H O�7�O8��=�����χB���>�-��ꡋ
�j��*��:��
��p�4�۞��B�w��c)5[ތ�H���ƿ�Կ�@PP���2ӣd~-2a�ߥ ѥ���D��ɠN�^$�R���҇�اۛ/�4��B��M����
FLl�V!�$�Ӫ�UY���%���E6.(�9~w�m��p{�g��x爙�m���g����Z=kb��+lcq�Q_P�3�`�h�^x�Z���ƅ��\	�X�����f��y��b�Sl��������`���#��B[�!�&�u�7�[�CV�/	�߃�[�u�����ܜA�d�+�~_d����g���M��R �e�ǹ�7��2����*R;���/|�T�����g��@<���灇��&�������~E��L��,�/�y�_�Ŏ.�-����I2� X��'0;$DP(�n�x��3�)����=?ȕvz؁���}�L.�9�f�Z0,��)s��xmĽ��-)I�j�s�=����Mm�^v�m{��'6��w;���}k���|3+��(�q��� ]������4��������>�`��0�<�J�k�%��(��aj[Ս�#�������*����QA����qK���/����OMͦ�_�O�T�s��{_^�?Gk�������g|k7�o�nP��=m|+�*:�����+*�,��]g��ۊY�h*P��ԡ�m �lb�@G;���� �����9�n`��o/;�
�9��CEEzL����ֻ�J� <��:gb�~��V!�9�:K�wd�%��E������ъö��v�8�ju7=�L�E��c�d��y���<��lǻ\��,�?y6�}b�s��7b�c�s�f;�ݟ��0*�&���i/*7�	���B;c�[��� �&�ؒ{s�{8V�J:�7y�ΞO�*�	p}��)��8Qm�����uc)ƃZԢ�%������2�e
)	6�.������XGO������H�EH�F�߻߭\����g�[��w�W��D����H^�S�Ѫnё��U�D����V�����NP�^�^�\���ݴW�pqY��N�e��'ɮ��������o���%C�f�k�WÖ�
ede��� ���1 �\��)H�^�ϟSN��3X�}�� _�v�@+�Y��/dPER��s�^�D��1��$]�>��H�m����x�8�A��Q!i�.c�
!��Fq+���Ɣ�0�^FwN"i��F~go-2<�Tq,-r:፭hv���c5��m��mYe�(_�HE���/D���ci)���~_����)�*�+>��hn0 +Sݭd���<&�\z�@���@>��Z� �q�D��i��@hZs��d�m�T),�9��4`�@�&��> �u�yi�IwV��Rz-�δ�����E�Ώ��ӳ8dE����&ٵ�e.nE���
����Cb��Y�*gG��%
[x�y��YXD!����g��[\�����B/=� %/5"!�������`՞+Qfh��[�49\�T�\3�{��I��9*tx���ubֻ�,^K��?�>~\9�P�����H{�_��%��n�,rzCz{Q-�R��-��\���h_�����?N��"%%eH�+�3.R��C;��@����^E;c�T�B�����q�a����\��I��e�:*.��c �\�#�q%��� [#� ��qK����!�M�4R:X�?��9�u�P��E��_M�m�DL�yU��V-?�:]c�!Gaz?�piR�VQ.jjۅ��|��h�}��P ��KjV/0U�$j��1���&9�-gs,��&��[��"��3��DC��b�CR�&��@=3��z����s$L�7PC_W����#ơ�?��w�4j�WA��4���h�hEn� ����@�c�a
(�³"S*�H$��tŜ�����X�E�3�H� 2�P�DP�w�[����=~> +#D�Ƞ~G�e��-WĿP�k��fMnlJhgO��ja��1̃-�R]���t��r�jn?�q�,;�Yϥ��Q�������pf?|䷼���5<�Ւ��\�Q3�5S�S�տ�W�U�?�~T1T3��qZ�ц���*4A+4��],{+�����Z87�>$�	*/G��*�_�����Y���u ׈�'s���W�z��F�.�S�zIq*V����90�r��{�"�2�t5��^�d�:��g��[K�hc���k�G}��ί��/��]�����D��jk����b��>������!�S%3E��E�Ӏ2C(��/��G�Y��E{;8('H)w	�-�݋܊S��	.�[���	�Ž�^��͝��3s���9���^{�n5��,���z��FĦ߲Bo�m=7�e�¾hu̖𓹪F��m�wk������_���^̶��?�m5���NJ�Rh�Ii�)8�LGF@�2_@D���9��K�Ck ��>ypC��E��(||���^�bT`ȉʎ6�&Y�R�6�|�vw�ogH��&�һ�,��t�]��|����>u����wP��I�T�ᥢ�AH�r���:`�1�A�nv�q�S�.����|+�.������:�Z��x�<5��TeC������
�, 4�����5tL�R.p.[�����{^_y�0��=R���ү�o���X}G1~�-�K'g�[�OU+	7��aI5|�rl��*0X
w�/s�M��������J�`���R}�T1���-�[���Er܈Gr�S�� �h�Y��W���t�{%�?��{��?����(���[B���.l	 �D��A��Ցb�Q�(��L%�&%�К�x��7/Ƞ�r�o�B�A��'�n�����l�C7[����`�����0��83p�vnj�� �kI����x$�k�>m�`�F3�����&���0P2T�	#es�`�W����-���f��p4i����x�n>u�r�F��н߁ߵ��7�?O_^~�-ɠ=.Ԥ��fut�k�n�_�����{1=�Q~3���]9ˊx��+���{����i[��6�}�צ��������=��R��.���ռe���I���@�7�1ї�d3E�.�Q�QԴ�Ԓ������R��< X��B&��-���l�"b�~e�/��۝X�l��v��~�M1]!��z��z�x��;Z�s��L��ɪ��D��;5�=����~T����ۙ�����d����@��B�2�FlK�J}��\�*z�W���>��g�.��1�y.��3�!���,��u�[�^�����v#(��\���[���6��{W���V��{�c74�Ţ��Q����J�'�Onxʊ���8{o�5Tn#�am �}Xl�}�5�(��P�,��5��3�x	2�������uQ۲p\͘.��R�%ʲt42�� �C�	{Wݷ������"Uy	q"�{�<\W�:g�Wy'�d�9��]�	xx��Q:����saL� �Cq�j��agP�ĄK��(�%�4�b�Zv����Ŷ�e�K,���o��)���9j�y�鐾�EИpA��v(�!Y �?o-�/���)�9M��k,W�AX��aw�TT0�P��� {��Ua?(�:���=���`�L�$��q	���!*��|���L�_�ݦ�����Dv5�8Hl��AQ���!WK&��hO�"Q����u]� ���%?hװ��*�fq�.�0��k�& ��,��+��`���T� �\R¤��>�q�ne��QՐҖn��qB\TB�`���,+I�1�d���+�Jl����՞�,���4���eܺI���]6��SR��^���O��G����tVr��V�?L�K$WĲ	��7G�_�\j
�tT�t\"�US�9���(����J�HF���Q9�<v����E����֬B�C���p���ʔ���{7S_��䳗�����������^�cfv�� ��,����:�!��l�3�5�Y8��]% >r�{4�i�Lm��wn��vni��dm/-go����y6g�Y�Ͷc��~��=(�'
�g���&�r��t��4ΨZwYPǉp��$��K>� |�S���1
��R��ʨ��d�$,�M��0�����P<Bj[���GA�
:�t9��ʔ�T�eAh�����a�n����l�N
��a�bj}����*-��MmZ��)��ʦK�g���94�C������-��1���������t�h�л�1�������A��^��q�PY�Lq�*���+�ٻ����Bj�"X+�-6�]�o����^�{Yxңo���nE���,���`��J��*�U�+���E�F�MKu�W�Z��o��P���Q#q���o���2�K�5^c��g^8���]�z�~I]�~:�6�=9�iy�i9m�j�,6&v��U1/�Ĉ�����x����(��v�>t��t��p�{�0�4��!�h�O��َ������ò�T�k�S{���[���:��Ba�6)�j�����Y�N�g�S��?���&��/w���=�f_>b��:[��}=8�<��kkk �Y��;G�%eZ���u��QG������:�|�I�z��6�	=r�*���յsg|�o�6F����k� *(N|����t�#!��s�Yd�����׸���Q�V���v^E�-���Ĵ8�wD6c�	�G��Pޮ�?Ժ!V���dϸ'�;�:����^�W�$��~< /�j#_�6�M(���p�ǿ�g =��@�1D�f����(�B��{5���ݫ����j��䤍0m���Qh��gE M����P+_�����ίU�OU3+�W��Ii�Zj�i����u�V�2����ʎ�����҅8@D����������1�&S��\J���\�������o2a�h����^f���E�&4�C��K�q?{f���$�W�p��J'��/��!���3�?���[�e�Y�sv�d�*	��>xB�{WN��5:�\�:�LSC�:oXvѮv"6K޴��Nڰj�~��J��F*�o-�AT���$yf=wq|uf��ž���`��!dp�"@cssG�6�֢��|_��_*��I�/�tD]Wf�<����;�ܲJ�%�d���Ի׼-ܒ.�{����v=�WΤ6��S�a�L�M_�	A�-m.̀t�J%�N>����5����N�=q�q��q@��M�5������3Nc�t���p�!D&J��,���bU Жyx8�4�����?ٖ�(D�+DՃ�`�3���j��|�(y6_k�wk�'s����c1{�2m�c5E���K{hH�8�X��T��o"���&f�؟��ڮ8���O�*�dǻ�Ռޞ� ��T�rsskl~��� �7��JguY����BZ}o��wQ�{k�� ���<*K�����l�۫��U���S��xv("�k=�x�4@�q�0V:x�������wǺ9��?�Ñ�Q�br�Hm3m_�|��)�_u��4(ʼ�f2��q���U�f�P#�SU�x��J뽣a���Q���D,�K��S���b���a6g��� $%���6�����C:�}��#}�z��M�8���WAl�X�џM�Pƾ,L.�����ZU)�XGJ���Y]5Bx=�l�i!��!�[H}r��廋S��ŏ	0�%�z�L:]�����l�L�5�$�C�y`J�W��.9�3B�;��D�ƖL��	Quˈ�~���Դy�/��!=�R��(��Nы�
�+�Vr�u5�S�Lbs���F��?��wh�U�[{����_񮸶^H�����O8W���Ev�	[�S���6#��L-�j\b�M�*-<Y�BFM�����u��?�;@�m���m��}I�Ec�����>����ɪ��I��d���������r���Q]ɒB��6��MØ���{�uߜڼ��M\�_J[����ٴ�y�O���R���ھ�Uz C�Ū�a�"���T ���`8i:H��>V�o�jqis�l���uA���Ǜx?~�?�<�F��#5�r���Ӑ��U��e #���w\��Y��I��AK����R`�ѧ��a�7fy�e
��;���>�Ur x;�Q�ߢfn�[#iߛ�!��C�_�l�G	�C��b�S� "5���~�F�Y(/5��R�(uXT�������N($9˒Kö�\P�;��
63�PJ�O�1��)N|���\�kF�Ս�$�G��:ݳ�����\o��'*�S�]�B@��Jkc�]ӫ^>N�OËg�u�,���]������F����9�vuW���sv�:YZ0:�����ۋ��GT�cI��_��Rg��F��"c�o��I/Ŕ���_΀� m�:P�@�q -� ���a
�|�j�.8���{*�hZW`6եv�Nt�ipm��C����Y�o��'y�����;o��nΑ�U+����{�CFΙb��?�_��˧��)ò�5�B���+}��v�8���=��\V"07�������xo�L[�/6wJ�.,SI1qf��]�d�=�z������B��,������I�E�B�
�x6vAv��)���yߵ����/:]�;nEn���;gӞ{�A���=�xS�b�֜�x�� �X�`�x7�E�x2SZ.�+u��z��o���]N�Q�c.�m.��]i��&w�=�/H�E�2a�D+���i��������~ӔЙ}sw�;���<�K�]�1����Oy]?g�����3�u�\k7�:�.J��vz��ߟHt~>���|��6���y���v�������請�b͍IX�9���2�T�����8oᒡ<j��w�&^��v)�2r�fH�6��Iz����d,�% ���}(L���)*R���Bi7+���Ay?�ُM�̋��Y��m�����-�y�/�����<�5��U��~tʰ�Y�q��4j1"���zED��a��|>d�͘?�|���O��"��(k���GwFQ��'(!q�18��y�~V
��_�m!^F�`���״O�!C���i
 j�������1��+O�*��G�x������WϮ�)�`ť�V�H�����\�u�R���o[�����ۨn�N��W��4��R��o�����=�m��Le�W�iH����%vR~!��D��v���������S�����ͨ�r�⩫'d��?�l���&��A�.[z�$�5�"�x��3u�	�J8u�tqĴ�ŠZ�!E��&����g*�
�^��1f��USV;�%�H	�FK���M�q�ژF�[�}p�K�'�/䳗�tc¿Tb��3P��������� ���O[�72�dpeeecC���������������~�S�ͥ��E�*�/Ш}�f�%����7�Aof���(8Uz������sK#�'�w���?��ĥb���bƱG���~I�fQ�n��Q<����SNƶ/���BbR��gBs�Sä)A�����j���~������������)
���:I'��*\�-q�7�F�1qa�0:�_Ä���t��ì:�X��!�)_�M:�� ��7©q5\>���~"�)ԚZ���c|Fk�+Jo��1/�b�*����@ި�I��:�i�� ȋ%������j�i�$ZP�F�����5��jq{�3��ʦ�\�U&#��o��'�G�&� fmA��ӈ�`^��a�z��G���2��T��4�g�t��Ժ<����-��.�ݎ�,+�.K^?��j��+����#Ϸ�@�K|�9��M��]A��`�$��͖x����A��ј�\'�p)�KPݹ�»�ͻ��%�������������������gY	�h-�����콩,�x��w��LǮn�AQ唂�.���bl,��B��}̯�!X@��E�
�	x�u~�,~�Ͽl��R*�,�C���]�E�ؑfe�N�����M�[Sߝ��v��];�Fx|�G�tZ�pY�)���)0����y�ߛ&ŗjŧ\����H�KJ�g��id8�]¢C�`�;�,XO �C��l��՞D,�v��S���J��\������}N@�ә�Mk�b�?���1� "�m��]{,+�Z��u2�"?J��QU��eR�X�`�j/��x�I*��%��cq��c]��^��K���E�Ƌ�J��������inf�y�̑T������<r`L���u�l��ղZ�+K��[�ڑ��k����i����-�x�6��}W�w
�\�w�$?|}�k��o��VXi�(�4��J���w"���}d2?�X�g�|�o���+ο���O���N'���Fk:}����^���s) �U����n��Z�趟��ĥt�� ����C��HH���@��1�����T�UKֿ:�7�/��?/�7yeb��`޶o�� �>�Z/�n�T_�N[~��{�W�0�ͯ��o�)X�������@�����d�������N�/�>�2��|i��🕍2}���K����
�n"�����>��q�T�E�ё��aL��~~�
u^��A�0��FG�S��yy�T�Kf�߾����d5ZgĎ����B>�|���N.8�=���q�\H߽�����;t���4��z��{v]��uj�Hl�귆/D����π�����A�	����F��G�k��7�Z~�u��~�����f���%���
�b��e��&F����Z��	��*�ogK$�f�Ef>�	|�O��kHE��f ?�m���	�������^��3e>P���@ȏ$q��0 &�́'�f��mT�k�̓`�F���䊨�1���@y��*�X�?]�]k����b`ueG��(ҁYT�_�C�K���șUV����_o�a�U�=�P!��m}Zsz�ff��:��jVj����FS�������ֳ�7�!�%����9�jS�}�?�� �b�b�� ~�q=I~�m�û>��ϡ��&�	5�7GO.?����q�̳�2Ky5�l�y�����?U��I9�����S��3�� ���f���Q�'�i�̬L(��Q��Ȼͨ�:2-J
e#P\�P�b+����Ͻ�M�B�V�A��~�y����+
Vǣ�y褉����L��L��h%�z�E	�]���D��'P������.�bU�ǠE_���E��-?yܯOOO=���u�䑅b �ETC����IkhhHJJf����IOv�,��5��Xg�+�n�-���J�o����.B���O�E6�p0�z�v�����7��QPDS�*PD�"%�d���t�䧊�*�szL..yQ�����(�X���%V���B������}{�_��V_����r�{U,�p���~���%�����&�ֵ�9�a�R�Y�e�\��nGD�r�d�q ���͢� �������\0��5�%�z����41��.d�d�ޑ#�������G�ꬁ��y]���?@O؇/�iH����z��Q��L}�tr�[#Ϗ��p|Bd�_���dt IH�'����Mq��������$S�������#�1���X�N���!^�^���xE%l�2�\�m,�|�@T:�T"_�A�LC�8	qS����`\C�j�<�J��v��R��[閛�9bJs��y/��u/���`�w���gP�������0[.X>��M��K�X��y������e�w|�Q�{m�cƮEl��)M�y]�N$5xҚ~ޒaִf�j�P;�<�6�r\֖}줆�RNyb�GJiD�����e[��P�U�VXZP�*� (����������������u"�������}q��:�c�wO�R2]T�8�$GbϨ�ߧ�֐c���3��� �G��E�_�KKA���Qm��2�O��@ڡ y���S�SrV���y^�dm^)~J鿒��ׅ<�I0������q�e1�]��>��a��9��2��.����2�a��Q�/�_���3쎖<��:z������t4��N|T���-���,���G���DT~*���SD+�_aO�h��u�6c��>�a�6z6@2u���q���omim�"a�t3���QͲΥ�B��G��-w@aԓ���Op���9Z�����/�U�w>�!��������_�����@ (��sO��Ӏ����N���uϭ�PCV��s�?MSH'����S�}����W���!%��.�⫻��W��y����}����������m���"ʘ�cZ���zɿ#W3t:W=�/����{���{~*u��V#�����QY�{o-����(����2��q,V�/-\�<%���{ 
���E}1I��]��.ܶw�6Q���<���`�#JLe ��j* h��0��x�������Y� 6�b!��%��ě��C�8�P�M�L��"��*��n�#���;�g+�F�Y'`^�H±���a�����mMK�,	8��7��o�sd!)y�}��,�.�&�����q��ї+�X֮������+u@)��|Mx���w�N���nO��4���=5QA��*���#������|���.����@�������'����N�����n�~x�>��|�����Hh�ӟ��P0���Y��3��3������5ǟegY��(*g��������c����$l��g�g��')�|�A+uXoz�4}<��+�R9zj@J�����~�����H�w���*��~��؂c�	?:�N���d@g4Ӝ�\z�H��;s�dx³�M��@�%J��dlk%8ZOU@�����|��餏R�,�����iYR@��]�~�*!�m%�9���aY<��9őto-@O6�ɏU(�5��pr�[�-�Q��)���6�J���uΜ��K�P�Z�UT*>���}��R�}Dao:P1�6�e�~q��#t�+75Ѭu0��kiX��^R2_b����.�l,m�P�s����=д��� A!,�'�p8�5���`�4��,K�q�s�����&���^�Q!68s�2�v,��)���<|<��<
(����kh<��r����5��p5i&h�����/Y6�q���A�Tybb�D�~����n�I� �������8�"R�����u#]]�����$(���,�7���d�f���DNJHHDI
$z������c�o�DPg��6���J�V�?�C�=P���D�[�+P)[8ABB������S{{����G<�ŏ���r��=�Vu:�Ox����k����j�7M��;z֖��w0�ؒQD�R@�!}Iq�o�F�<��z��ͨgP����2�c��G��X$�fu!�<���$BN�n֦A��
��K���qשP/��:�/�5�%�SJ'�47Z�-�TG�M��EL9��x8�DB�5�ǽR߹�e,<�9�U�����v0Kf�CN8;��w��Y!�yƨ���)��OZ}���%�T�Oy��C�����s������?c�2�����LQB�J��G5�;�2"w�z���3�W�I��T9Kc���cZ��|\Oj5Bg#����"�bJ�:��sy3f�H���Ï��Ǵ��
�/��*�b4XW���!��/n	?����9dy�IZ+���F�K+j�U}Ax��l��z��r��zƼFڴJ��~�F*�q��\<�|,�b��8L�����Q��y�������!Q1W7�������FnJ��n:sů�^Z6���2�`�����F�BBBBOZ�-I 7�%Rb��آ��6��z�j]��-̰�l�O�?�_��2�������OW+��)f،���k���=�X�LKC���Nknv8suy�b^�Sg�r�;or��W݉6<7���d���"p��,�$�3\��}��1��Ѵ�L��L�bNZ�e*��N/�s�"Z�;5�MmK�c�>���B�K�\h�S�d�`����5Ǻ�d�~����iܞ�u6��b/�W�J?����N�هS�J	���Nsa΢��KJ֒}I���"u�k*m�v�D�A)��r�C�l���O�����Z��]�)h/<˞	�8*�������~u><����"�?;�Sl�1�<V�,U��Vpk��05����S����ʁ�!A��Ml)3�D5�9�&���V�p��7ݱVɥ�UB�Cl�y�³(\vᵺX��7� �&��>��[����B�M�P�b�]�x��Bg�qC�0+��jn�5CkEW�I#�H��y������п�ӭ/s}�n_���$�۵�q��<f��*���&u�艑ܠ*U��*�v�<_
�dC��rQ&�%kʊlx�M���I�]�OK;���@}�D���6ST��[l���o[U�v�h(�dN�/��U�of��Sc� ����&֍Ʊz�&�x*�_�_�b��1f��RL�4*������;$��m��ۀ�\q����L�Kckl@ �	~e�C#�n�"�z�+���e�VI� n�4q�a�ݏE�V8e�껆�\�H(+�=��M�z�ډ�.�%�9�9 ��qSlȁV{%9?���ī�'��EE��$��ŏgd�J]�$��"��?U�Az�d�SX�e	R��'��dz̾vZi�z�:ZhlX��N�m�V�����9q�v>����%�Ǉ����Xht]HqcUyCxxY`T�]�ŭ�|轒�K����ߏ���\�}o�2�e�w���Ռ���-��#<���=u�5��q�0T PhcieJG�=Tӟ�>��0�7$ֶ:��9��W�"��� �#��-���.���A;��nJ� KMdڼt��� ��ZZ�+�#қ���嫊l��[J��~O�U�� ܾS�L���֫�̊ul���أ2�yq�S	7Ys-G��b��6.�ʅ`��c�q9��;���4^&�kLh��Β�'Wa��[�w���:����̦n�R;1���6��}��T^�?no�����=;�#q1��i������B����Ӣo�{]=E�y��rz˴DO�n@���s���\� ���ÅAK ���n̑/J���-����:s���}�l�/�@+�\+��w)��P|}0۽�a9��x��A��H���ʹ[���&+�/8B�7&靟U�r���0�(\��nY�p�	8�w��d���r�g�8z�����Aә�]nt^Q�����G�v �Dѧ��S�0�";�v��\�3OD�;�����X*H�S�8�9֥*ڟ򢠎�B$�����*�N��̥����E��ih�i��A�B�B��ӻ��HQQ��)(��0�g�#�����\�=�����Sz������o�yxxDDD89�y���H�;�ۅEE444��^���c�X���Q��C�R2�2����f��.\\��y���l���>��%�p�0!��9�׵���JF�9t��?��E���eI�111���PTT������T�S ��Jv����OռIx�^�&!@�"����_�I�.���//���6G�7'l|�W��yG۰6mGw_��:h����U
W��T��\K���t��tFe�k�|�@��g�m~q��r� 0�`�y196P�qx�\�zkG�+(�D"�>b�J2OY����\Y�W�+����OZ5~G8˜�W�O9���@W�;�����LW9�0S.坳�O�C�o$Y�t���'W�^,� ?��w�Q����
c��#����9@�q98�SgtV-x�5������5�ش�$��%UDc^�Ϸ�yU�us~��)d���s��@P�4{��3M��K�5�1�����
�
���\�������e�Z���ʠ�L{�F0$�#�nC�o�X535QT��3Gta^�����^62�^0z�M:��7+ MByLVx>Da�f��u�A�	��+9
�����3�Ũ��{m�X
�_�"o���1�ȏƲ���e��,iSS����S�h-3��?�9UۈV��GiTQIL�`��
�2�o^�g�����Z�;;�,"�����]� ~��tF��5O/So<#�yV��U���>6�\��!��}=��|k�+�d��I�a�b�U��@�E���,�O4���� 胏>K�$Mw��M���T\Kvb�o�-ޥ�$�{~��T�ubѴ1��d~$Q��u��b�u˫��/M�\�2�3~�s��3�����f�x�?n�&�ϼ��`�le��'=ms�{�?�@�w�.Ĳ�Zrm����Y
�@����G�I�š�Mh� M�:(#T.&k�G2�)�ǻ`�'�Y�$�Sٿ�{	c�@6½���TAa4:[o�{��ƈ�륆2w"J3�0��oB�3���;����O�@���c�����sl�߷���Ƥ@rҌ�gydg��A����}y~�G��n�p6�<Ti��Bc/'{�;��dJ,�y\�@������:R]d� x�#鵗���cx���QȘ��WI�F���
j�*�x�]V�Ǻ�L���|n���<r�^iH��nR��{[<<���H�s��w.�����Q�?ߞo���������xy�h6Z�Ƞ\�g��P���f��֭%� ����<��ዂ�!�=*̠g+NP�P��7Ȅ���L\�I�q��V�����ݕ�cp�/.L� f��v��tө�a"�s�b���<M6�*�>�y&�'��Y�Bj���?|A���������W$����$�]/�[��d�-�+@�<A�?����ƿ�P���̏7�N4�R���C��D1.h�,��KP��ь�*����S���Em �Q<E�/,��quU�Ut���V���&��>E�����?!�u�f�&f��jL��9�Sy�sX�M����ݎ��;��uݻ��&~��h~J�]\_�1���}�_�z��p�v��cf����Kӝ�>�8�u�Ԓi�jo���s��HN���2���W7#5IissS�O1Vz!��pV�~���*n	C�|pض�;�4��Y�B��<�}y�&)�L�����F`��ݣ|	��jI����d[y�M?|h�#�6�CQ�V��?��u�y�~.��s��9��	e� ��+�S*���{��iH�B��3�g˹Q�آo	8�����	O����2i��dO�h�q�������^��n*���Dn�߲�I����»9eG+�LuD��I0�YU[��)8@{d��>�"44��ŗs��fyҠ&0)���߼��_��L��cy홯�+_��l����J)A���r��$}�������B�o����CQjA��?���*����O�~�m瓙��os�IX�$�𨃇��]'ёew�]'�����&Z~m�ޱ��/?��u�_t=u���{��,T� 3}���M8��ҭ��Cgb�������p �K,�C(]/�X)�%�Z1�1G���2��#����X�3˦
�f�:�F��^�#��e����ĸ���F�X����v䇖(�������҆�Y9��5�+��bwz��/#b�#7Ð�C�#M!�f-*S��R�2��H\\�jj�݂"4��QX��h���3Gn`0������Z���pBmyyyddd^������SmpppGGGt4�0666ƛ7��&6-�v�
:�e��5�C+��C|�b  �Z�RA�D`�?���bR��t�J����Bis��d"Q�B�t2{�����d����[['m v����͇��/�<p8��0�%���r��b�F:��!��ˍ�L ��HM�U�J�9+2���s���)^q��q�_#&��௹�2�U:���{��������HWJ����4� �Ŧ�H�`Z'���@�h�^H�e��x ׽p� ���b��1
��R�?���0�w�o	�����󼳠B2Ϊ�ɏ��M��#3�c�-�!,@����B������`������G����������O_��pvY6:0�2�9�>�/�T�V�厎�oK�x{�eW�����;*A ���#�p����m�y�6�������4�h��`�Y�<$�do�%pv�"\�fx�ٖW�L����Ǝ\6�c�`����e�:4�5��r�ʎ�������Ag��bmȣS�׼`�"���bg&C�5�W8�6�/�XhD�0����gJ�L�M��X��>�M����bt�;���?���q�_XB�S]��V�ݪ���a�wap8Fl
��;	���b�Ȁ��<��6�jgKN5�&�1t�!⓭J0OO�q����o��;�Z�ʯQ5�T�Zs��c�Υ��U��s��9�<�
ta�`��
�	j i���:� �5�����lOJWg�:>OwTU��W�Q	ӢPl ���JqD����MrA�������z^
r2�~���Aoe����%�!��tB����|n���(��:*�ƫ
����r?�"��Ȭ�$⏲�@��&[��K��l�ݘ#<a0�)<p;v�uq�%���ֽ��HP����á���-w���8��Jd�!E�SC���z�b�b��w����݆��ʅ�y�k�\�M��_p0��r��m�*��N]���g.�D��E����-j�=��l��G����}�F��F��[l;lJ�r?�G����m~�c�<<���"J�w�;�Z�%6���t[83�c��>�%��ܽX����s�sf�����<���6Z.��?�#����DeP�#��8�����"�`RG2�����Q� ~����>��{جj��U��8�p��(2f����K��&�!=�O�!`	!�#��OW����v�)T��������íGȳB �B�1l^�m�����
1�;Lܖ��Y�Θn�o�|n	�����܉�W�s��)ߐ#�*��W.dˢ��ಿ��&+ʇ��H("�2��<�����֐���`�PL��Ϻi��eu�Ֆ�7~
��p�����f��c�ɞ��g �2���bs��3�#�F�J�a��J㡱�(�1(��!�_Rl,���}D�-c�Ժ4����f��]뮣;��D����u�����g�u7�aշ�����^V߽餼%QZ�ۄ���X���
�>��n٭14)1Ӯ'�����\<�9����]��w��O��w��D@u���	�������OMkݍ�Hm1�WSę:��e6��Ԙ+���|(���q_�m�VD�2@lu���o3��(���2�c�Wi<���w�1����@c��܌�#��$�B�m��D����iq�����";P�u��y��E����?��>��P�{@ݹ+c_�'�Vg^Gkp�ٌ����(+��1���h��� �h�Hzɭt	}�0���`n��Y)����N�=E����@(��b?�ᓝs��'4�↯�m�Q8�)#o-�Q������`=1�N'ٲm�>����{C��!u *U�j�a���uP�Ƕ`S���ܓg�]�tv�ː���`�S\_�]�ۻ�[K���٥�}���j%-;��d־������K���۠�t<,<<$�S�`���� �<q�(0��������(Z�@�J�$J@`�W[[[���)*,���USS353+**235W�����˫������4 N���|

�
j�P��.1��y�C������{\<\��L�Hµ���D`��D���0�����	H�IAA�Ü\\�����D�Www�\��\��ԣD�YT�o����c��V���L/��m�[f�0�$���1U�d��K�أմgh
�U�,?VG�F���OJ�6��7p� ��,��
� 2Ƒ������c9��C��'�_l�����tam
�L܈
Q_ERB��"��$�6(F���"P�a0�ط�"��Q�$�h�ؒNl������:�F�dP�}v�#����I(�Sa �i� ~~Z���q���'��^i�y��We��ߊ��$��<�l6�׌�w�l5�b�r/;E/�ZB����K8��@��m"���޶U�U��ݪV��T?!ڪ�9�6��?��B�O���F�'Pޮ�ahD��4� iz{���L���	�搳j�4�&�� Dy]̪�@U����`}Ջ�'~��d��%�s;9g�ʛ��,a���q�b�e���x"�Q:s;�o�����[,��(�h�1A��ȟG2��u�X⢂��E��!/©lb.���)�a��0�p�u`�����KW�'YI<���c﵇�MSx���ګJ�`L����=e*M<�|?E��~���Om驶`� � � ��ƶ�ߑ�M���	W����ʋB�V�]&�PN=qUfZ�t�Tygy_V��Q��Օ�dGx�g�m��}����֘k
̀gF�HFo�(FJ�N�R�_i��|����#p ��6o��|�B{�MZ:>6��P���P��p�|�`*W��"�[� �lg
�L4\�v���s_-4<�` �'!��ѕ(��QH[y�A�4Rs���U5l�`oڵ������A���E�����L���\T
����1�V&�s�)�g����R�p5OE��SF���>GB��v�S�§�����-�z2���1Nq��A<˨њ%![	G�TU�m(j��z��3/��5m-Z�J��SX Bq��
_>!r�����COQ[3�j���U+�ռү[�ה[�ҿ��p����w��w�o�u?�#����8k�#`���ET`Ɨ
S �R� }@��\̿`j��. �̋Gs4{>k�x�K~����r���F�qu�Q���_|��������O���O\;�4�U5�]�S�U�X��$@S��&�i纋� ���Fb 5���H;��O�����A~Q����Z�S#�*@�o"����ӗk��bj���&�& r�J\;
]��];�����Ѻ���������䥮���������������ж���R�>�ϐ `H��S��Y���s�,t�,dw�\�x���ǞW�25��u���M�|)��yR�XK
�#Q$k@�Rlj�_�ӦX�Z��6���ZR���k������FN/�NV�7l.֜^.Y_̘O��J���������������N\X��^�	����_�\^]X��_Z_X��-rg"��A������QNg������im�4�pj�}*j|��y��DϘ0���������$��<�՘�B�r֋c��J���I� 
8:��<�|j��~���.
�-	�BSǣ9
����fKT��8��eM����dQ3p��b�MZ����Vs�mg��P)g�&x�!0[:\�2k��h8�qq�0�RFE�$R��UFFJ܀q�'�h ���nKX�.��U15�� ^T젖�3����qI�ˑ#����Լ��*���J4*�MSo)��)�
Pc)���EX �	:�kY���e�2˒�  �i 2s#l YaV��h��x�86 ?�)+�6%��m�e���Tf�	S���ݲ�E�%�c�1���c$ۤ��%�؂��4�m���b`��R��Y���S��_�9ؘ�U�Z�����%�&z';���:�9����G{['�z�{80Y&N֦Nvts��03�e�E5~�� �DN�1܈�p�<�J�j$	��
KJ���9��looo�E"�TUU��PWW��DAA�B1����ਨ���� P���FWWWSSSNN�z�7���ɓ'����Ǐ;���o�̷�|KIN^���Sǎ+��a4Q�z���3�������������������̘�M �=�4?i񢢢�JJJ`H�{�����}���lmmutt�h4r H�����a�m�X��>.�N6��g����D&bqP�0X8DIAQSU��V�bU�i��E�#�^'뢗�a��1$q��<�=t�ݵ��ȩ��L*1Y���y!\D:� �T�"�7���{a�eHw����9
/��tYMH�M��S���飗�m��a�b��2�[�u�8��Z�#�t�X}{,͍^�[����+�L�^H�]JnX������(�u��d�6g�n����{�r�J���v�>�,wMi������`�添O���m=+��I��O��K���+������w-�����y���$s;����b��e������Q��P�S&����6�$'2ې�fDp���:6�$Kޔ�E�V'`��N�+�yJ�-�2j�'Td�V�9�&���Р�qTV���Z�(Yl��H -�vJ���S�L'�1ӈaoa�26cRm�,\�lٞ6�;��v470%��*
j���r$=-}`@#�	D-e��V�YM��%G�țclɪ��@3|�.���c���q�_Ss��䲞��2+b�Ti��0�RԄDeA���&�*��ʔ��8�f㉷�N�95��p�D�Lտ�K�H���ko�0�D�,�0Nď���Շ�TF��fP��:���s^�|��D$<15}fn�@�zW[��� ����a@��$P��*Z�р%�s
����_ʎ�ꎂڮ���2jO}VV�����T%n�jo��mi���Tu�epo�����L�i��<M�i�*bT�S2"N>�5S�T�UGO���R�ˈ� �D�*�(j@�4�4�Q�*"50C��A-������V���	�K�k�0�~�6���]G&uZ3�ݜ����s���j+*��j*��DtՖ���ܻy���sWϮn��Mv��V&u	�~��������D�[<<]��Ř5�	R��jLDJּ�W���8S���~�l^^�A�A<3kI$�ccZc(3J��m��E�M5}����� |t��_��ƹ�ɞ�����L~�Oa�[�59Ta΄lWr�%�Sh��z�r��b�?�d�ar=p�� x>d�?��E��Q����G�4���S�g���w�?���?1/����&�L)M�'v�U�*S�+��f��="�h/�j�y5{�T��6��u�o�,T�/ٞ�N��MW�LVl�V���{�f[&j"F*��k� C��}��}�^"�<{K=zJܻ�.��bvw�ӯ45��&�Q3R�j�UH�c�Դ'1@%��ԘU��Ղ�'ִ1ʬ!Ҭ:¢�k��e��|:�Ӌ�3�fv��G[G���V�
gF�Vfr�Sf'�&F�� c1S1���K)�[��ɛ�q�����9���ť��٠���蹥����^����vϖNK�ws�wc+��٧�ο�ʿ��?/�7)��	m7w���I��I��Q��~��^�+%�M;�];�C�h
=IrG��[/�W?߇
�G{?ASS�b.')�t���Od��3�	5#�+cj��h���� ��k`��D
���If4�Y��8�{��i����z�ī3Ϲ>Ū2�\mR&65A:�\�y9���A�:FR���h���p4Fp�AQ���⌠�����>�旛��{������M� ���%LLKQ�h^+��~��Pq4Mm�uE��k�3凙�CM���M�������p�ڂ���Ė�X�h&��e�4�5f���&��2��<��,��(�&/�"+X�P�����Lm-�o�E�D���遼d��^Z ?3D���d��UF�儃tMq\_S��P��d3�����;�`�5���a�^�1>�IA	!����^�&�,#7+C��i�+���������؎A�a��z4C�����I������IL��CCb�"�c��i�9�`������p��}����+`�B���ԈD���]pppXX������7�FEEEV<u7X��P����0p*�((({�������o<.�68-�����cY;�����KdjHdxpBp`���Ȅ�`SKKKGG������/:::***((������V[[֒7�JEI\v������pq�25x4$H8<��RUVA�)�4��(E�!>��,֓�6�q�ƻ&z&z%x�yĹSA���BNt�N����6��5�O�� d�@f���$9��� @^�) ?�&� 25Ge@J�<G܏�U�g�.�4��XЀL# /�Z��B�֑05�Lj��A�+5ƞ�$�X��d��lD�;�{Ep��3�z�*'#�渵ˑ��m;��g��ϧ]��ً���g���guŷo_��e�څGU������y��Ъ��Mg>�<����o{.��t�n|�������s��kٽY=��g���b���e���)n�{|�Sx	�+C���礬E;�H8uJ]E^���2!l��l#c2�D��\��B��G%��N�Վ�)�� ��'�(������*JY���U� ��T��U�L�@%buq$C��B6�PLtM��pzx]S=c&�ٛ���	oj�oni��j�	����q�s��[�t��h��ZAYSV^����	e�S8-%�������'��y�����_ԛ���_�/c�7lq���T��4���qV�D1��/��������1�EL|�P� V�b+�5d!A	P��YIP�˕+���y��ԉ~�Scrrs
��)�.Rt.��\�RvȸU2v���c�Q}j������,j�$M�<񇖌,��)��O���w���X]��:���&N �TQ�0T0����(IY#ig$ّSۖW�QP�U��U��� �A�A�o�S65�74VU��)Sr�Iy�)�:�p�d�E4X�PՉ��X8`ʹ�h���S"Y3sB}��`�����権�U�S��i��� �J"G3����5��Rǈ����Ԉ�>�4���PG�т�hU�jS��5���;p�Zr��� �m<*|��`��j������U+�-<75/���d^=�vnc{�����<����{�� 	�i`ק��� ����i�6��-��z�"ig��� �"�����_05e��p�'�Vm^i�����V�-��}������?���z��ߟ~����Vf���y����\;J�39�M�u�)��+�� �$��ԀD���C.�Ն�s��	C����A�v4/��S��MȄ���H}��)м�PF�3a���L�oS�@�p��D��T��D��`MXWExOU�hs�|o��x����ۻ�7Nw����[=�7��m�^[�8=X�ܞ<�5�=�;�9^"&h�:p��o�§_��[�&�5�65�f� v�L�H��M��^X�
�z�EL�9�g��6�&�1m���hfI�i׬"˥�:��!jitT;�K�K��˓�ū�Y�	�#���qcc��S	3sQS�	�ki�;)[;�+�s�3����������ɰ	��4!C�M��JϦv��ͫ�ɫ��[P�W"�+��f�{�Fz��x��8�y����\M�\@#!�U/�U7�]'[��"
8�BoJ��>��נ��
G��#�5?D���4�15��y���R� ���aS�ɛS� IM��}~��N�Ob6��Z��{ync�~�5�3�!`=����g7�Y�?�h����0jQ���k��I�Blʎ�@/�Pm�<Ku,���U�ݖ����5�f���A*y�(|Qc�hj ϝȋ|�y���� 7 ���/����P�\� �c�ED�5	6�(ˢZa�QQ�	4SCLr�ӂY91�¬���ئ����ā�ܹ����型�g�6'�VFj*gzs���]�me�-%��v�Lw�|_��l��`=�l�Mv7�[�����pz������ՙ�������Զڂ��:AFG=oz��[�]Y�j_��\��Y��f��+�R�S�2cs�#�#"�����\m9�,G�����݈n�g@!�S�&FzTo�{\|�H�$'��%�g���f�rr3����y���<@EeYyEi}Cu]}U1� �IKO���
���B�P�N�RPP@�X������777uuu�`TTD�xC	P��Eliċ���)��o�=qRUQ	���x4���؊n�`c�l� �cY�mQ]di�5X0�4��H$KKKpo������~~~^^^���
�������9q츦�˒����rswur�w�BƩ!`�����ã�XMuFS��BԐ�2 :�rٴ$oz��Y��Q��A��u�	�'��"��N�$7�TO�4/�dwJ<�r���] ���!b,ǟ&�i�� ?4?!�������%�xܙ�:=�^nj��@=75�.�1�z֔ �1�ԂNw�v��N	M���w�7-���ǷoG�����7��������:�w��~Žuæ|�2���Z:�z���á�ES�+W���]����q��U�}V��$}�V�����1=��[5�U+a[q�g:�c��Ĵ�ŵ�I�8)�/�K�p+�9�c�\�P�2�XM5�6�`��mg��bL�0&{Ӵ��)�4��A@��P����%��(��EMMF%�¨�ph�VK�#��tH�d�>A�F1��`:Y��-�LOG�!�t�uM�J��o�o�&Fػ�Y٘��[x��D��#���<�\Xnގ�.V�6&F�����hɡ0J(�S��h�cX�c$�c$�7I���x��ѓ�]�6Q�[W9�H#��K�&%Z����L�H�X�
�bN@Ǘ��*��B����$�*���I�X�
�*�Su2��O��?ur��̲��}ûƴ��}�C�3�:7��a���T{��T�F�զ5��556��3D�ym�y�"KW�CK�WN�O�L��7�15����#_��"�朢45��9P҂�v�z��9�]y�]�e�Yu�}��>�he��E[U5;N���F��U�=m�G����9��=n����i˚�9%�h�����ќ=�1sB}����X֌�R�Q��Ȋ�D^�h�!E�h�U�FT�#j�Qu�&n��45`=������j`�Ԥ$ܦ�nW�t�ǩ�E�:��#�^g��@�Ʉ�R�r]�pUiOuY{���VMM_��#
߽y�ƅ;����e�-E��wL�h��Ҽ���U15��)���5��i�2��0���\�K�r4�V����Q�&�$��15`��������U����x��?Ӣ���+���"�����~�� �2Տ�P&�	^���W��O?~��w������_^i^jh�'��e��G;QS��Y.�<J!G�ȇ���/����z��~�����O|
�$@WL�3����"ig ��H	���ύ��E$`&���G�k�OA�̫ e$Mr����}mJ�15P���C|��*����ƀ�Ɛ�����t�l��x��|���{�G]�zxi����&�����zz��f����ݡ���d�Jg�R{�Bk`�%r�9b�1t�6p�ҷ_��S��Sn���V15��K��W!U�I��T��W���ߗ�Xz{�5ֺ<�^j�e^��",K����_��[;��wf�����������e��I�O�L&LNELLGM/�.�D/���������̅Nυ�O��tx�t�7���u��v�6wz׷yUֻ�U��x��<3�<<���A_� �`�m�'��j�j��n��n��lwQ 45E�Bo�B]�/��� */�R��p~nhd*ēm15�Ⱊ��		^�i��������iL�DL�i`+�E�3j��SD��%Ӯ��e��{�*p�:�K�@NS����J�!?ܠ8L_�<F
D�H#n`�� )h��	�-�'�>�b�g��{�"kSS-�+U�C$����?�G��7"k@� �����H1��O05�/���55/�>�9�Ś�Tm&�2-�0@M�㫟�G��J�%a��P���������򙁪��������z�r�`���y�8�ҷ���gW��F�����Z���N��^:=uk����� ��0?Ը4ڲ<�6=�<?ѱ�4t����k�O���9��007�>1��;kc��.��gzZK{�ʆ{j&�����A����ɞ��֡���֚ޖj�J]���K�ˈ��t�v�6�a�jL�u��Z�<Âf͢����&������K��r򞫙b~AI)O �W�VV	����-��m��}��]� (-+븸''',+##MX�p�R�l6���?<<<222((���U[[�á�hp2pX@&X�/ES]CMIYSU/�[IN^Y^�Ң�����@_� _w��9��ŉ<����;�R�BI��	2��d2���r�����0�Fw����s�ZYY��Ǐc���Ҟ�n>�^^n�n⹟̌iz�:�"�Ipo����c08��T%j�3�x_;� {�(7�1	[R�5A�-�#����Z~�Y��q��n<��L|�� � ��l^b����C{�� )A�ьf/�H��6řFE\^�~a�����	�d��܁�&�A?ƞjo��������\�V�������l��i��h�e7�:6�84�94�qhٵo�v�9c[�bS�`���T6�~�p��g�>�~$��$���e�086a���m�y۟�-<.�����Q����Ӟ5�%���s.e��˜�5�W�w�Rp�r�p!�?���!4eǓinh��6�fD1bR���zΆڮOC�������)���P��7�?�+�������j���h�Q��Oҡ���Z��6�h��oa0b����'d'��R2{Z����WF&�Rcm\m����<��C�Sb�"����"<�َn�6NL+{�����J6 �u1d
Z�������d��l�Q6�(���Lԏ��;S�-6QΓ"`�E�$���AS�g�����1��X�)F`�)�+/D�`�P�U�
��'�j=�v��o������=��#s�k�zW���i����d�݇��PV�TT�UVQS��P�UW��ᶱ�2	��D$\�យ[��ne���)�5��&�t���朢�Y��F�@Q�@�W�D8+�~��Qߖ�ܑE��c���g�(Z��X�MU������b<�q�8ycu͜��%�]w�����ں�W�tf�#�ȡD�M����>�:v깦9jj��D�fXA��aeu���&�4�j�1ܸ&~L�0�&�p#Z�jD]�P�^t��V��H��Cۮ�ALM/�4���i���c>Sܠٴ��r�b]�H�����������i$g�~����{�ܼx�`kga`���^�T�
S��� �j��O���&��5����Ԉ��8J{6�(�BLl-i�J��M�oSi�.Bd�����ך�Vi\� ��;;P�8Ҵ"�*3ȸ�8�"/ti��ˏ�����w���O�����e�:��T��m�h�����Ŧ�GWlj�ҦF�i ޢ��h 0��2�X��H�RM����F15�3s@l��65�Q���MF�+��+r��ezy���M�k��֨������ oe�tk���bõӽΏ?�<�Ε�'��\��}v��f��������m�&J�z�W���z3W{җ�RWzR��;�g[#��CG��Q7�"���������l bcݞ�|)��y)���S��_�T=֒BoO���T�,�|D��X��X˶��X��3J�%�rtレ���Jy1�M�C�C�݃k�ӗ�D��_�(_��L�-Ng�L&M�Ǎ��,,��.DL̈́ON�N�AS05�71:���:>���qoj������h���k��<x|��,��NR'*�;����)��>�c����G���]t](�n�tw�Lr�h\-bjx>:�����|�E~�����@�"��TFЪ"M^Ou�im�y}�!�R4{Q�ج�E����~��hc��Sę6$��6|S�9ٲ5�ْ"���A��m�`� k{�lHUӚaם�.�L��OV @����%ݶ:�Ba\n(�+�2�A��0\PΥ`fe�!�?�x��	��c��  >"�YI~\�?��%�;XÊ *v�j~Xi�-����Ԉ8ba~��DK��k.�+�RjD�=�W�&{�R'���OElڥ�~�i^��A����H{^�CSq\Ge�x�`e�ew�������������+���ܽ�~��X�{��G/~p����;�7g�憶F��.=�u��wo�w����g�^<}����kg w.l]�[�yq�ƥ���O�]�8�]�Z[��?{zvu~pf�cn�ksytos�����Mo-��^��^���Z�xf��������`�PwswKM}UYEiayi�ۆmK��6�c��QHxM�.������5>.*==5;;��RX�P�/-I�L+(�)��痔��%�U���ڊ��2�n�hnim(-+��͆����LOOO�{?ihh�������155������MJJ�r�nnnT*�ǃ2��`0�`ynX�[т�&JY^AQVN]Y �8-����˚���M�����cif��`�I���S��5���'���wpp w�����p<<<,--uuu�M����[ �Aܭ���71�9;:�q�}<���L:�]�6O ��&apd,^,k�x,����PjE�����ۆ�ais�/:�������;F��b\�2��K�q΅��龦I��p,�To �� �~fفt@N�% 7���,�H��Hb�`����������󾛾��iG���� x��%�f�Hs~�@4�(�槹���u����>��^F	.�����F\g� N�_hzXbiDf�z�kj�K^�g��K�s͆Cöc�CˮM�6�a�Y�aӼ�غͨZ��^��3��j/}������Ô�{e;_�L?t�\��<����;uϻ��W�w�FP�E��9+��w���K^��N�N�ev���pŚ7c�9b�3�?�[4P0�Ims��#��]iF,�1ݚFs0�:R�����'C��L�:���ge�SQ����1eŷde�PQ�UR�SUWB�t)�tc�������3�́�jo��2�2c��e����gF{&��ϝ^���v~wxe&� �3< >316)&)=15+%.5.:)�����	�v�vqtw��80��xQ�H�dD�P�z(e}ME=uY]�����b�����+Y�KW��P9�B+�
{?%Ya�YX@�5.�I��2�LGb�X�d;�2��Gǔ�a4t��z)Q�#'В+��>�Ȕ*�,�9V}��7����?u��O;Z�'f��Z2n��ޠ��66���s����h���u(�w���))��)�k�N��l�h�Y�!�"�xVS�3��p�7�neٽkl�@�ஶ�m�(��:�p������(���W=PT������>/�q^^�
rNF��ɨ�R?#�qFN�"q_�r�2��YL�"oY�-|�M�����Vk�K̐��,�;��7��t-V5)J�y�D�3r�iY���S�'�掫͞P�<�2&��Q9�@SjD�FI�i��1#*�Qu��&qL�4�&�c��5	#(�0��"����nL�& ���u���ӏ"�h�&~jW�uj{p�m�^ڰ+{,,p*>j&;}��l��r��j����Z�Z#�������s����W/ݸr$޽�����}��᝛W�ݽ��8�67T�O�tW����E�q�D�f��;�>��ʘ��*w@�+��¹��	�_��*S�|Zn���,` :�-]��H����X��"�bd:m)�D�T1	��� �h���h�5�@C��`3�a�鹿��ꃉ�t��4�T��S H� R �9{.Y$�M��HC m-�o�RBLͫ�M0Ad ��	_�ő��sdD��QX� FDY,�$ڜǥ儚��D�R�OϷ�٭���;<���o�>���ÛۻK=#-�U��L��&�Y7�M�`c�\�9��<O�} �v�P��y�����q�B<ϗ (�#��I� 2D��R���+©�J��*����hگ��55M	f/�>��Z&��`�9Ѽ%	��[H����X��ԟ�,	��݀Mhs��y�0<J��79�߅� ��1��\��� y6I���MXX�`^H�YD���_ �]���)z���Y �izy��E�EN�|׆��\���Е���ބ�����e[5g��.7�Y����r��гksO/;we��Յ'�g��O^�:��;��
�LV,��td.tf/��,ue�w$/v�̵'N��L6F�ׇW�
8�|�A��@�c_�=bj������WԀ]��b���4��%E�k@uT*�d�:Pψ���$�M Mq�2UME��0�Vc�飗
����Vyq��t϶���������Toa�x}1gy>nl$ij*qj:vz*jj�;5:=<�4���8=��6148�h������j�p���(����
�8�Q�\�w���]��U��9׃�f�J�uэsD'8h%9i�9c2ݰ��\B�'TY]2u��z�� 
?�R�SB��WDTE���@�
��Q*#a�9�\Il�L�_���W!�9-ZS�(k��H�f�P�+�v��y��>)�L���T���z���Y�*���B��A2�U��"����NtT��T5� ����zH��yP�! �טX��#����!��f�I"�y�xH
$.F�Dzm�e]2�>�	�5���xs���/�"�Tg*�5-���#h�pӂP��`��0h'x����Jbܛ����g��7��ϯ_ۙzpa�G�����������7�|��g_~���>��魧��>�u����7.>�}��7�x���M����w�]��W��/��~��ޣk�{�������G���>��>�ƕݫO_��s�ƹ[��\>����|��t�����ܼp���g���6��v��Ο�8��ޓ���ғ�j�����"|lL-i:�f�,K�!�؀�d���LL�NI���N+*�/��	K������B^n1��LP\Y%���jl�mj�kn���)��-������B@~AvLL����?u��ɓ'U�cͨ�����888p�܄�������@___sss����&''�������!^4ţ���P`/��`0�0�k4���K���lvDDDaaaIIIbb"�����A����DNU8��w����...���iii���YYYAAA���666L&�@ ���р��H$p�D"���\��bY���I��iPh��AC�� D4VK]���i�p$,J���4�qd�;1t-�~lc's���o��`�Ƙ���{��j�³#��a)��q��oz�0�c�b���
�f�;��٥Y�8醱��I~�8�i��E�?#�c.����4�ô0�.˗��f��M�1J�5L�3��7�0�
4�����rCE����ƀ�H��Hc^�4�L�(O`>?8��(�VL+
2�����Az����~Oz�A�9��Y~�i>�)^�I	�n��qa�A��ai�y��%c��s��U�M�2�zٺnٶaٮiɾyɱyťmשiۦj�5�MR������~8��a��g�\�n;�ټ��zƫ���o�_�yN�Y��-Ǫ5��u��h�u(_c�lJmK���V�kނ�p�6g���c��Uk�cnF3s���Z�Э�����u�	�XU�T_�z�:��y����SI]�m��o�������vgG;k7� ?��7n�{T;<�+������oz�ɇ�>�����]~�����������Daqt^NjQQ^E��&OX�������Z������adijʢ۸��{8�}\��}CC��ffT�����.��U3�R4F�Z���v��z
4�0s�X+�4R����?756x45���` �vXJ5l��%֤RK|��sS#�ȗ���5��
Ŋ'�2�*dO֟:�x쭶7����[�x�vh&7)�[z:7(�&�$�<5���-
0��0��<��4�$�LD�P�x�<ꀄ�A�<�0����K����Y2����7���w��}C|�C�G�\��]R�</�
���qEր�
��jpׁ�
L�@^���ƹ�[�98�uI���D�W��չ�x78�>f�9e��y�>��o����E;�;W�]v�fk��U%�nV3&�6x\~�¬�ʢ���[����֔��hPad���4/z?ASj�UP#j�!uܰ0"�3 �����4�Ӌэ�5kh5��m(L�&�W;��R# ��p}��l��F�*�[�`�f�na���93��=��5T�?YS1�X�S]�VY�R]�ZS�^W�YW%mj�yx�'޻y��;��,N���%s��"$M��O��15���H�xBLMg��qd�L@���$R�A��0��(R-7Hg��~����:g�R� �05LI�"���A�*� ij@�_hj@������o�0�\r�8=gy]D�*�6/��7���ή������~�ݷ�~��_?�u����B�pcnMF`V #Ņ�⤓��`c3]p�n� �|����4�'j�|j t4���$P %h���%eMU�!D��� �Ρ���4 iGA4��� ^!k��@��S�D�ZG/�k�<�$� ��y��y�����)A� ig$k&X��L����8u��r���5�ӭQ�f��K�W���˓��Iṕ�[;=wv�{P����sSu�W:��<� � u}od���R�م����A�R��`1`�+g�-u�+}�=i�5~�9v�1r�6�O�-65n���BǞ|��<;HK�)A� U��45��B�#$��u�櫌u�)	�+��)���7�`�� ��$�jwj�al��{��f��df�xi�`y.kn:uf*yz:ar*fr:rf.b~�����	 �č��������Ѡ���.Q�'N]�GE�WI�OA�Oz�g$����ח�c��Т�b=���(�.:Ilb��f��Z��F���q��<bj����RJ�t`E����":
��P����:
������-�	�C$�� PL�$���XW��@��h��d�״�{F�3���w�Hc���V��P=(ď"����� ||x��7�|  �<8@��$��Q��X�s�O� �@���S��c ���$i���y���y�Em�em�.�	�I��!3�B�iL��)d�f�eY&y���2�1��qC��m����+�c/�||���/���>{r�����~����~v�������������o���'�>����������������o���ǀ���������'���٧�?}t��wo����?~���?|��gw?����wn>}t��^�~y�����k�]�x�҅;�߹t�������]�pfgci~jdw�ڥ���Ɂ���� WG[3'kS����!ќF��2�ts�IJ�IM���J-(�).)*)��y��yE����B��_U-����o�nh�45ׁtKkCGgKsK}cS-(�����ࠣ��������$��ZVV�B���FDDĈ������耀 GGGSSS�(^4�5Љ 8�r�/<������N���V^^^VV�oooO�R�.p6---x�����<jjj����]�$l6���#..������ 555**����$�ɴ��066���%��D�B"�Ph-,�����03�h��� 5�Z 
����`�`��#��x,���<	��0�qw4帘z1���$_�Y��]z�Oky��D�\��P�`SQMa�0;�$=4?�//��s�|�#���=A.f�l�`W�(��4)�&;�%����O�S��"��D��0�/K@�3-�F/��4��0�CM�1L�5J��1�1�	�军�qM�#L"�
��y�fy�F�aԼp��H���G�����bZl(
����@#^�Aa ��� ѬO9��F�&"S�m���H�`Fz8����Ŕ�6����s��n�++6U+�5+6�˶��������ۮM;��k fټ^F�g�ٞg��w�������{ɫ��[�. $ܛ��Z�8�g=�v�k6*W�6ص��v�+֬K�m�V���hɊ��X�a�7o�>b�����$��-^6�N6�cc[c};];k#�%U�JV��|SS�me���>�G9UY�.	Gճd�X��[��3=9�p��8Wn�%���˕��p��H�-�o���'�}����~v�o����o���f�?қ��R��V�Җ��Z���ok/�hvuV�v���zEs������a�����h�;���������ކE75�#��P2�DE�ᄛ����R��J��F��X�0	)Vx@*��fML��2� X�H�!'�βO����[ᠩAbj�
�\��|��\��)�̉JY�zY��':�<q��M�-]ݻz���cc�$�5���q�X��7��N�*�h*�j(�4���]��6���Ă�!���'v��1��������&��$h?��#Pn��UP��.ʩ]Vи��k�%yu ȼ ����)9+#wAV��
��
a�/*c��:�B]5t>�I��j웦�[i�wӺ��.٧��=��;oṫcsZ�����i�m4uUKgJ3(�����	�铲���N�AS3*�M�hPa9�y��a5
�R�fX;����eH�8�ID�����@����ti�Q�f-T
ө��S���F��!e :��݁�n��u��ѭ��]!a���E�#����B8?w������ 65u5�M $`���nݽs��������F~�@�KM�oS��{��5 �T�x�'(k ��gH	�b���;�d��g�����,�`~!��A����7��AZS ���2s�_kj�+�(�&�Q�ȬJ��H�*��FZ6�s���~���o�9��o�y���?��������U�9AVin��l�4g\�3F���y�`�G�i~
����؟$�i@C��^
h< �F� o�������v1Ҏ�i �cj`�(��Q$�/9����:�5H��(������qg���k� �%��+MS�i���}<�^�]o��h��sS��0٢>�~�/��N�ݳ�7N7\�n<�\��Pqf���f뵍ֽ����~a�x]�B[��H��|�������3K�{�-�ӵ�'�6F�c�����������Δ�����L�ct$O�7�x7���؜����ƶ7�xcۓLlsc۶m?�����s�̛��s����]�󭥆���ë�w�lێ�����YY�
��� ��q	���ƛ�_����V����A
�w����
����%����{�X.2�u�sH�L��f��N8���f�ff� ���_Iۜn��vg��Y�k��:�٩D$�g(�W`��
��W���s��S	q}^jN�VŜ��=��i���r��sr�;J���t&�]��fM:#���
����WfH��#���؍�2M�ee*��Գ��L�}g��GuD�*��4�EYa���d��<3�M~�]����,KX��?\e�|�����!̝��HbwT��߯n��Ac��r)�̃�M8&�d��աaw F�ˮ�h�{Sj�c�Th�$K�dA���¼ L�G�Iϳ���& ��	��l>�����l5�{^��o������Swz�������v�����ק�{�B6���p& 6��zH:�e�-;�^�I6|o���}���H|��j��/K;I�/�C�>�p_zpt���zn���Z��z\)�s6�B�~�-��u��L��6C��m�q�J�w�]���p>��.�Y���~��T���p���|1\H�s�|n���`b��~ۿ]~�S����ĵ�����H�u���������LD��!�w��RU7#�)�(g+f���AR-�z��(��μ��P[CEME:K��
~kˊ�'��%��:7�<//���0��썄���,Xy �HYQ���IZV6(��������,���s�uKK�6w�'���E�О�cH#p��!h0���rhH1��%(�y2���2���UUUUT0		�-,����EE_�~F�XvU+���ƀ�ʐ*`ϿQt���B7I�{ijj�GO�`b������7���65�A�LY��2�� (c J����?�����^���ޝ�/��.F� ��Φ�X.ɫ(ˉge�]�dh�9$�q��vt�����s����ݰ�Ƶ�,3�\7�&ê T\s�s0��n��1��e8�Tm�Gػf���� il��V�ʾC����/���y֬[
�� ��S�s3����RQ6��`�.��Qʩ���,"�9�*�0R�I����]є=�4����k=�L�t,�&�<=ż�`�aو�"ip]� l#��kh�>PpFN2���5��%��P�.��wHo7JZB!��s��a��p��u�վ��xY�jS��R���X��]W��X�^]��d��h��P��V�c�Ӧ�2��z6Q�!��E�����5���A!���c�l���Xt삫��S��䴬�d��p�Q}�Rm��b܇4�x�L�ռ3e����^H9����48�7��i��pR��<L��䫬��7�B��1Ia1�t����e��q�����),ylyt�x@ԁM��
�&?��o��h�qVa�C��}`I����VtN��Êo�����q߲N�BC�ɖ�u������j��/^��;'�9�X]Y�9�׶�S�삔���	[�&}��@��`�Z�9��RMn�iZ7onA�B���M�J�w���T#p�@d( �7v��(z�y�9Uz��`��ٸ�Y�M���o����ȎEZ򙇉���w9�h�֗~1��T���CK�\<=��dV-a�p��Kϛ�r��S��)Bqډ�٤�i�(�dA�3B��W�To¼��6�F,�ӌ�i3ٸ���m����쳋�d�J�� �
	�4��l����"9"����]5��WA�u^i�����k[�w=�$Dr:�힋N�Z2k �K�1�����C��[��2$QU3�H@���d�dEB�B����R�j&Zr&:r��*�gj�=�j���Ul�����;I>��S!X��p�\�8 t���e��lY@�.��.��o���U^+�q<p��(��4Ƌ$��ـ��n$�!T�m.y%d1�`�)ob�l��KUS�>��a���r���ϥ����I���p�,�(\�7���`Byk7��BQ���:�s�n����K�Ų��آx��{gƐ�����W�o-%��I�(ă`N�ߞC��(�E��$�{eK}^�D\ױ�%�e��egBa!G7y9\]��	�~��X�HM���?��]�W�J�,�.����Y6�9������M�?�A6�"������E��@L���#���!5�Jv!��V_��o��ŗ�&Hz�띶�IY��7|���������e�D�Ą=fN�a��Q1�_����b�ؕ^��|�|�]|��4PC��]��]�i]�h�P��N�v��lDd�
ǂGVd\�����L��_12J�W�F�w�J0���j���ҕ��p��K��9����v/#�u��;����xn��l�5j�5
���cfe�3����yʔA�������ss-��T�O�6
�C����'�}���n�vr�v�L��ffŉ-�����Ď��nv`t���6�!QxN\p�9�����@�y�h�o���:�ߧ��N�yR\�XYg3+�w�j��l���ȗI�o�)�ü��,��{)1f�����I�b*�K\�{���c`�$�\�{�-��[iLI�7�B��9u�4�s(Ҡ��@i��LS��5����.e�Dp���+�EZ��]g�RX|D2��ך��Hũ�ա�����r״��ݯ�j��4`�h�bX�����Lǂ�Wq��{�(˴����R��+ᕾS5ؿKnk2P?��	�e�$�FRn��%��Hw������TN�S!jocq{����;r�l�v�i%��>��I��B���ze"��v)ޕ"���������P�q?d6�%��3�܎�Zd����x�_�������h u9�-T-��u�6��ډr�zz���8V�����L��������d��݁�:������{�coo#��8(e�L㕣2�cr����Qn����K�O�\�1M)�4���	ݼ8͒Z#t�\��L�L�MŤ\�<��C�V�Q����)/f(-���U��W��BQ�v�6�/[��,t��ɩ��ll�v�JJJ���\O���M���B0���@Tdd#{��ZZǇ��4�_a��&��$����,NDX<꠿������4�/#�O� ""�LO��������ׇ��i��K2������G*C�*ɶ�������d``����f�� 0u����I�my��PV�Ԥ�,9*�۳d�}�D:X��ݗ(Z�`���1�A?vB����������[¾��oo7����g�������2
.Ss�Ο�W�&F�7p7��۪�<����G3o�Wn�IF�'Ϸ��U��Ϩ؍���u�O�e^!j�;����:Zt7���f%q+��t�*�T�Z�ɗ�á����N�>/&�*#�1����b�T�<*f�U¶Y�A���
����4F٣��_�@-�r���(�k�4"P����߬� ��d�||rl��I3�}�d�e��@��_;��F+{�����I�JcC�n$�LYU̙n�:��Z��Z8.�%Zu�i��Y���2]3Ό�r��J='�UЍCxћ'���YG���5�N',¢jy���`�5��v�+Fw��H��5��_�:&�6<궋��7�e�r�V(A��G�Ih.p���ȃ�#�;�3C2��g&S,��Lͭ�
	�!�� Q�u��0&H�D���+Z�}	����b���iZמ/#TT���/Q��J�\��l�$�z)��C'�����o�ѝ/ρ==��$$>n�nz{l_w*�}��9�t�w�m8~���ģ^ ��M�\��j��;��[�[�M��-�<��Vv�W��+x��q	�η�Nwz��jg]r��gu��-��M�s��t�5#��+#�Cu���>d�#��,U�j�3�4��1�s������Y�CY4�����4�L����\�>?�/��_�������bpnw�Y�H�j)��z�Q�<&��C(%C�V42�*�W�����-�ϻ�b��c��)��:F�<��� ����sS�g9=����?8�~�B{�������ϻ`�b��Jj:)�a����;�V�TVT���I�a5��ezH{#�=g�O�V����$Z��7�4fV����.��gh�&�jG#5����En	Z���zkEMz�Կ���\C_[Fм��=������K9��z,��T�wU0�bX�"b�6*���7�f���_�摊Ìe;ᶀ 1>�H�s&�J|B6�y@��TO5�8 �m��:J��
�vi���/נ��XC�M���
풧v�(;*����乧��|���p�3ghr�ui��ni��)��_vB�����]���D� ��5��#h_=-m�����u�?#�OM�����i��3l!a2G�^_V�.��N.�p�};�)X���r?˛�����5��u�﫧����`��?a{`��\<�~о���Č;ZoZ��9>��	ő9��YQdR
�ڔ��� �o����� \��$%��U�"ӳuElz�u9����J�O-���<"���,�㧃��|y��ծ��/�a;�I1N���k��`�ɣ���
��4uG�5X��:���?�[D>8:�}�����
�9��&���iϱq$_!L��Ce��]'F��%h��@���?vDO%l�U��|��ݟ�U���5	�t	�+�0��\ͺR���)vљ��(�8�	(�M(����3�ķ8�{��(��R(��pwZ�D�@� �M������O�/а'�a��=�y���*����rS �{ 2N��U�,,8%%)���'-�s�Ż����c��ĴTgVW�6��2X �L����l�l:�P6Є�:ceg�(�\$⿪��N%��Ȋ��E��7���ee�n45�$���!��%TſV�yb����߁b�	��9���H��!�|E�P9�+Ļ~�?˿�kp批�P���cy O��a��A#�2���wIc�?s~�߹�1 ���Dc��!��!G�f�yA$'�a��2��Ax4U��a���M��wa��3�̉ų��f��#?r�*�c��bW�7����cq��3IV	Nyy88��\�O����6�5v��Nm	
p��|�o-dw�4����ގ��V�7A�k=0gop�v��r�&��+ܳ�,�˂�UD����������z'�Z�����	}�ZǓ�o�^�D|�N���˩���ͨ׍��B�>>uNV���L�F��ׯ��O__�?���?z��s��:�~W��7�jh����-�[y�pR.���|0]a�w��!�窕$1*#��c���=[��GE�ki	]I)=$)$������������>":);55=i������2~�t�cL���h_>�m���[�\WWWCCC���`08,,La~qiISCc�@NN.,,�}5=G����!W���P���Gc�i����T9\�tR=2r�nJ\$�T�^IFRe]]"�s�B��*}�NNN������������0((hii�����驯��gn��������<;�����Ɗ�mYRbQ\lIWj	.� ��@p�"Ia�W��"{�����X���jN���w-�>�}������m��5��:x><�+��+�&�Z��:�f�%⻶y�V>䔎�ZJnU��Ϩ���V?�����Ïϟ8�=��f�������j M�#�I1��7$b�F]�M�wL�\U�\q;�B�ޯo'�������r����pl�	���e��Q�$Pi$RU��ϓ�*��ǣDs�]��׫��X��,���n!= tbA?d"}�*�*J*-�EB�vzP�F�n�z�_�)���h�ܼF��<��cY5`�c��c�r`I�b!6��B�\�,#�.�u:�TX&�g����j݄3#8�٭֣3in�W!���wX�7�긖�%W.cOhޘ�������8Q�iEBI#����4�ɐH�d�ӏd���5 
�R�e]d�0�6�Zz��#�2+�˽�3K��c{���w��T�#IIR��5�b��8��r���֌j�̘�H}�ꉑ���'En�O�k=�]k��ޫ5��s:8�����:ng�W.H��"?T~���'IN��o��ż��j��Bq`�EK1����v�ua#UY�����um��u_哊�F�O'H�T�U[�h1M�l�<�P���K��2{�ۄ�1J�m�' �*�S+�V�S�Ӥp�Q9WIl�	\s��J]#ҌE��������yʛr���@g����Ս�hARq�pL�vN�?���k0��a�F��V�8��R�]��g^���tC���=���A�ߍ�^��%�W�.�9ۚ�UXT��B.̱�'*���j�g�O K�k���8*�ԥ���xe�<(�����d�����u���no�I������m��ނ�cţ����>O���̿k���s:+�|��u��vL~)�W�pT�������D~��!�-~�Yt-�Te��	�
~OO(��]!�*}�+XZ�K2���������K��Sc��'��I�++М翮@�$2����9/6Z���_6��	�@��<%7=<A��n2c���y1����4��~Bn>�c�Y�*��Z��c�S����<}�M�m������� Q�A&ޝK��j%��)@�#�'5=�)�b{H�~� rW�����q�B���
���r}�	�}�����Y��;�6�~UH���
���I� F����<�,�#G�@��'sػ�ӊ;�J@�A�E�Y|'��W�j|�'���Z_�7�X��P�_��tܖ[�n�'��B����/�/�}=�a�OK�Lr��;��;�~�Aȧ��I��q����'n� 蠲Yg�>9�~�f׺+��_�F��"*��uWJ��W^>,5O���LS$�L����쯦�&m����M ����Ii��d\B���~^�2s����,9�DjL��9b:'b�V�Xf�g���0Y� *[�)i�P!L��X6Z%�e<ɂ�7G�˨��2��b��<��wuA�?q�����g�gO��'MG�6%��4���Ru��d�kl�i�����$����ך	��u/L�΄��8VN���x6����!ɽ��n�%O�en���U�j�qw&��pyj��7�U�#�E$u����"3��;�h�J�����Rm��D��$��[��c������_U �*�b|,<"��s��,ޯ��҆�����t+��v��C�q�g���.Je�Yoڗ�r)j�,�~z�&�������f� 2E%eXo���DHF�dLW�ݯ1[3
�'F���W�k�x$�x$�g�$}��i�o��� =m>M���g�<;�����ӻڑƉ��V����Ή�GS'kOs�&��N��"��������vb�i��L��7����qP�s���s[�e���AAc}e=�<|A��ĺ"��|-����3z|�y7�Q�����@�����GJ��T�F�רGB{���������J^�FH��\��&5�������EGC[SQ_WUYQO_����� $?�l��ش�>
���x(+�-�����;�7a5�, �O�Ǉ)[_EIIGk����f��i�4-���!��Y+����G�����U���	�Z.���u^�����3��W�h��߿�[�O���aaa������C`������q]#��Q�edd���rFeg�+(|K���
���cyyimm�����Y�xƏ�Hg�����O��B)������%��������������z#Ja�+����m$�,���>>>�M���N|�E�y%ey�y�%Q��h�e��i��qŨ��X<1um�~�exָ�n�������?���I{Y��$�1���o�;�;�:k?n*�X��	��EN>s%����{�u��m�������E���X������=��>y�	Ew=C�Ȗ�
�U}�B�t 	���5�7dY1�����5�@(�5��rV�s,;�w��6���c���c�n��C��v$����^���d���&y�i�(+LlRh��w�+2�ӻg�;����H��G�y,9��(�TV��M�����젼�}ͯd�-�K�l��f��0�^U6�n$��O�w���)��`=�t-�}��`�C�o݀φ�O����.Xӫ�W�5�L�:�רh�כv��N֫��|�+��:�����54��3ฮ�G4�g7�����zY��YY���fh�3�c(��������O��CsAC��/��a�b�f��2��ʞ1�i�fIfgA�����O�)����fp�j������Gf�Ƚ��^��V���|���_B.P>���φ��&���b�����kk��z̋+��E��cQ���n���y��yj;-�j[�Z�r������c�!��F�s��)c�8�=�J��Pq�J>���	����4��d~�Q��}EV��ռ8�b�Y:5\HWC^�S����'UYv �ad���\��6RӜ[�,�=��Uq/,�a����$C��͡��F�[D�CA�VH���AhV�<�չ�go�X��Q���-5ҳ��t�̾�Z���{YV�� �����>��>!���?(4�J�ʪ�yWH��,��J(��秷2\m�EU�����^U�K~\CϞt�K���������Ӻ�	9I/����nw-���0�_"�H�ڥ<-y�b��EC�떆#�y�!gaa�ӄ��5=�4���������p�_�>��h4:�< i��¿�jݷ%h��!os)Τ�?��
�H2�c��g�T��㘻�8�ȗp��bt��'������%<�#���uj���^Ί�N��vmy�V���"*-N3m+a^�<ߋ|Z͛��˲�pѝ/�5��(82J�o��_�"�?f� ��{׺d4N��Oc�,)�-��X�-��CЄe|�T�u��R�˚����gY梵6�bq�/����'Dvf	}^wPI^/�^�}=_������_/�`�q��OE��)?����.�S���͍�c!���H���L!�����*!;�I`;��$�^���@�6���	�,���<�I)�Zp�!����+��n��
���`����P �s1��-_��j���/�si��/��85{�(yG:ᚳXѹ��}1�~e>\}��>��O8���
�l_pwj��?
�{݇j�+���%�0�8�7ak��;7�n�Ӛ�@	�I�K��kC%�w_""����y�����?I�)���sN�r/f�%)E$.�'�r�Lh���'�?eK)1"u8*:� <��#V�X�y{�W)�bW1�Tiydְ{ ����O���c�e,�0�2�r|����������	��
w���Z4!�lZ�Tz�W;�q\�*ٿWc�W�׮���.@��Z���]j�z�q���pY������UV?kN�
w9ZYh���Y	5�P6���C���3{~�RM4I������q1�ۓc��+Wc�R��\l@ �<��M����鄢Ǭ���-7!v�b	��h�v�'M$�G�'|0�q����!I�چc�}16��g��C�'�a��n[�蜝&t �Y������'�N0��=�֎Df"z�ھ��A�,��0�L���%��k��/��*�q+i��/㚯��],�,jֲ9�z{�:�ڹ8ٚ;��{x�8Y{��YY�x;8[Y�62�]��XA�=�h�q;=>_´r������u����@\`@�䂦c��e�ϖ5^�u�M�5qa�ff����Nv��#�u�nސ	v�12��ל�ߤ�{�0v��W[�GNj�w��3�#e�@F���3o"]�H�|o���{���1�z3��'�^�@�������#���i�Z�v���������!�O�`ccb~�����/�vss�����ֶ��66:
  �2�^�-v�����}�gH�/���� ""��o,.j�*c����a1�B:�����壣�UJh���A���=�����&�Arvvvm-;a\V�J)UV!�0~�EըH����^�O�o)2T�c(����_�!�ttt��Ԙ��z��"
KJJ���Sa88���^ �!m���I  PBKSVWQU:0�$`^af���uy���f?O��������4�c��Z
d'c#ӹ#�<'
��5st��=�i�6�|u�������3�h���������ݛ���O=_pl��N+�gcϞ�k�ɝ��69����8��/�D7 h����Wz#�_;�� '�D��y�C�e!ބ;��V��#֪f�X�)z�F�2O��x��u�L����f��Mgd�<ȁ��0Gb�D\+�W��̕�yT�]͌_S�P�?*J>.Mߖ��e����Ď�d�	��g��ߴ�(�Ø���s�U����8J�e�N��I����kr��=��f��6��4��t��'�7nN�]�"#=�rLY���~���n��5�rT��-�zKm;u��6����q�Z�{�L�T�z�'�J�4�0�#��ު��j�%m6�#�$�> �9������mlf�o�"@֚KWY�C��D���^��FESV2PU2RV0P���2��b�1D��RG?<- DPۑ��^�om�����l\��Om�E�)�΃
a��]�/�7��n\�ꍯ���^��=�
��Ә�Y=�8=U^�w���Q6��V�t��q�Qt�Բ ��>���KK[[ Y��3�ÞAp�V����Kh��aA"YȱdI�h#�?1�ƔhV���
�����,� UP,VP+V�)�r]K�=J�f�y.M^Qݔp<��>��W6O�P�����NZNH��}�wfM��oDư���Q<�q|�B'��w��;h=אk�h�(&c/�s�������<ύ�<�,�'4�@��&1ѓ�l 0�FLi��pl7R���J�kbx�a�k�c���P/��Q~������egr~kq���&�\�n��UZc���svp��C�"r�p���&�C�c\��(o���B��|Z��.|d,�v�y�����o��2np ���Pc�_�p� ���~>���D�dl�O^2k�~)Z	������$�u8�dv0����[p��V�������s�}N�sUE[gnM'���"/�X�2�miy����0�F�����y�4�y�sw4�Q��/2Oj��+����13���xq�u�Hb #�ʁ�ڦ�9�JDLm�]l�tM�#HL�0,�pFQ�}=�._�B�|�IH��P7^��W�^��j��v�s����fͱN�a�����~�M��v����t���|��+�0�����M��Ì��^I������X��gd#���yI��+C�|ӄf��A��g�@�Cp$n�G�`�V����k�w�@:/&5I*��$B(�y�	����A�.�GO�@oL��P�|�_���D��_߰k�Ӫ�Z�9�xV��R��P�y����	&ͣ.�jf_)��r/c�l�6��9�����eY�}A�k�	3\w����6V�����}t�^�нt��L�aW�K{�g�i2��Ċ����Ά^Ǐ�a}ZP�r'ݥ�%�5,-
�S�I��I��S	��q�[���MD�ٌ�����f�j�hL�,z������o,_
�{ˎTz[�+8����FTgf6��7dG�pOce�K;��M��uSm���	Q�0Ji����l%bSRU���g�~�p�9@�\�Tf؆-�a��&x�V��|3^OR �N"�m�z,6��?Ř/��C+!���	i\��%���C#~�ۄ��"9�d�gh����Έ���	ٿi��uC��_$8/(<<�֕G�v�����
VĵN�1H=��.<���8C��Yu��ԧ(P��N�4��w������?7t^[����t����y�9���l{^)΀R)�P)sg����zLwC��ɂ ��qu�v�q���2W���>�_�~�&�s��%������n-��x��i�u������b_��Zh���o�3k�;����<U.���R&���;�|���Day�,{��v+u/�3���k��/�/�>���k�/}/�^���'~8(p�M��>���L�V�������'��
B�19i�xiY���ܴ߿p������RRRʶ�@?# �i������R�HH.NOO��Y[���9�.V�S�Ӆ���ᩪ�jj.	�n�~���1�����VUU]^�3%#�www���� C������L��[Br���"���CJ��rw�jjj�>_�����蟻%""��?���Q4#I�I��/���e�ߐ5rZ!S�a,�0h*����.������+�V�������U?~/���S ��W��~�H�0�[[ym-��s��o}��XB(�ӕ\K]�C$��kG��_�R�6.��u�r#9e����:O�U��]]�hv1<���i0e�����Y.���}���]���d��?a�	�zB�������h�yXou�@li@td����;Y�����,,��
.2���WL�~�
1	��m����Q{��M"�C���t�@p������"*O1O��" G^T���{���K���E�bQ�b1a �8�X<�|?�-����Vd3��>�e�2�R%��l��҂����̽c16wбϰ��S�N�4gw�x��Rj���p��t[~�7�Rh� �-bѻ�T��b��x⽑Ʋ|P�ܽ��E�cg�!�X��~J�b�gB�SO��Y���%�b}��j�}��˴G���6^�6�ʫ�����W։M�uR��,�A�{)v�H�jT6#��(5��(+m+qziP3�ڟ�*���;�ȳ�C���[zB<$�����?�(pH�_���32�0�������c譔������+��q�9�NK����twy�2�@��ŷ������mD�y�#�b������Ng���6F���4���@tN��^�㵥ݹ�o�����3j+:x�c��2{�T����A�K���WI`��@�_�D�B�t����(|_�:���Q���W6P�� I�4� �sл����zI/���* �n6�^�to�>�]��@ЍPP�����벚�-췸���,	�(K`����q�e�\v��BE�$��9'"�:B�xL��2=��\�y �qlp��3�de����SF��9���/'_�꾨䷶�jS��o�(LX&�XYhxJh|�D_q ;��Y{��f��bR�{���>A�i�'
����:�΋n\^��O>�/ļG`���0����̜�D�]>D����8aA�_;$:H��-�_9J�><���'ჺw����*��i���]J$�%���,a�4��L%�i�c�B���c�'�Z�$��-ʹ��+
��-��Oqa+�%�y{M���vJBp��FxApZ��i��~��z��iw��M����r���o�㑥nvz�|��2�6�_����+�b�3��cA����y���ݚh�:Y�:�w�@x%�e��Ż����s�(j^Hj��*��*ͷ�5/t_>��� �B�0��$��
?����r�>�rI9llG���[ُGO=�@ Z4#ܙ�S�c晦�P��#}����T�cqr�5�Bv/�_#��Ľ16D�4�C�_׉����i"���q������j��2���'ҾhG���cY�/���X�l��n����P�e�܈��0A���빡�NI��N���㣶�T	�R�猄�:]�
�Se6�A�]�C��}�J-��3?������7��"�@������5��$��$�,-c�}����C��=�Kȗ4
��_�G^�Qi�0Sn������">m���Л�z���9��6�N?1������e��07�M���zamنK�6r�9ѡd�&�\6���2�j�F��&0�B������K��j%�`%�d&��	9�r�ӝ�զ��Zk�� ��jd�1ً��!vB\",f%��+��c�S'��~`�~\��.�iF�!�)y�x��Kʶhz��ij���2T��4������"6�6&5�q�~/+0H߅錋J�{�?���+1�Ofk����r�;�e��abwLvO6���1�g�=�c�'�\@ ��IE���Q�B��?0a3J���je�ba�l�QP�i,?9N�| ,f��3�s\QC��������� z>�gI~����K
	nm�\p����;ޯNE��j�k���Y�#	&�KZ�"b"�+l�'"����v�?!� $���Q��,>~�	�C��,d+����%��%�� b1�'�a�:d��}� 4�ǆ�	�WG��Q._W�HYE�P=vc����������>��3k��W!�X�� oam`�B-����^vn+E`ᝬ➩�X���_V�Z����6³�K�G(�+k�1�ɟ3�Y3;��uz���.w��v��(��K#���H����A[���ف>�{���0�RY��c+@���zI�ee
E�,4�u9Ć�R�{ss��/Ҩ��癚�>�W��g�G'�%.~�X˟��.>�^�
]Hh�H���>v�?�9������=��l�O�OL-�u! �.��
�Q���QP�1���2qP~���`�w=��¶6>�l�iIIɭ�-�&<�3�"����tj��O�}���A��O��>��?@a"�b�?<86o�ۏ����;0'-..����\Aqd_|�>BD������~��r��ϙ2W�񳢥�����T�bi�;p���)̈���|���Gg&�����A�
��;�W��/�ِϝ�Y�(2?1/)�Җ�B ���-!dM\Ta]��ȾMix��U,�	�1kh`Q�KPK jd�{8}�C%��8�*���~��o���`KT!�}T�~���p~V����zOo���vC�q9�����Q�)���6#�.���,>D}�����}��!�=���(y�����o�%�ȋ�?m��O3�E,^�-�`Rnl�Z����]�� �lf�����ެ�����U��ٸ�����a��T������U��,~+ M�e�u�q�Ye����\׺<���R�.�>�A��Ք�����t�K�H�K��1����K�yGL����&ǿ��=y�k)��$�?����8[%�}i�kI�w���Q�G��:���g���iG.l�2��2u�]����8	-OK8��4����u�8�78��{����Z.ɲ����\�)5�洂�'���ߖ��ˠJ�"G���z�����k�Y�j� ��Η�&^\�<Z�8�7��d�%�x�ȃ���^�Ġ@�P (Sjh�~(��}����������Xb*f^Ӫ�4����᭭��N����n^N+׆�~q��V���_8I�8��jjJ���F�������/����F�h�����������"�N:�F2�.X��R��Sp3�w/�0�� W�z��X)!AX�E6��4�fʆ�8
 V�±��eg�/5QDXI�'{����4X(��Κ C(��c8���A���EI[V��؛��jY���]X:����R��w5�+&�w�Q�t���z����.nw���.���	��-'�܄�J�F����i߭�����\�	�mȧ��Ʊ[9L��RH<�������� ��R.XR/4؈�SB@�;���V�Ɏ���b2|�ǴkyC K�Mzv`Kn��C�q��!5]p��Kû/��ݎ�ᢠ�W�����ធ��epe����u%k I�χ��Z�;�=���m�H�r��� ��Ov����O��'�!��o4𭲳��������$6��/G�/_^kI	w^	�,���.�3`r)oZ�@ �d�[�t�ܩJm�ʜ�MZ�) ��V,l�i���$2�+"OI%SHi��ܻ���z
Z3i����:��z�>�Y�����#��(�}Je ��q�f�Ӱ/�-�+-�u�Ig$��rL�Ų���2@�8�GP��N�/�ﳵ��@� �Ș�4,�4�o��pp�%�Ե�L$����'p�]vz���I��=0�[�BC����R�=��D����l�9�[O�,��$�+���r9�fu�Io���yrӾt(8� �}� �����A���m;J߃R?a���APJ���#���)���AGt��� �2��.����G����#�;���hCk�Tf���d�������v��%�B��ͳ=>���Z�ޠZ˫۶���N�o8�3-�ol��q����a�Gl���4�8JMqx}��M�� ��L�� ��ώ��]y5�XeY����M$&�s�<� �j�J0R�ɘ�K�}�D��N��]��*�q����������绲�1z��v�&�����X@��%�f�p��H�Fj�ej�GnyNzcy~WS�h�h���ņ���.�ܼ2���py�|a"��%�03���b��i������P�)��w�K5 �j�BoR�k*� 5�3�k-2H�LM�Qy�H��V; P!^�(�
e@}k0PTGH��(�����J�U�n�r��a�Y�"��-<̄�� ,�*^z��.��x~x	�S�*$��kx!�Z����R����,G�/u����
X�(�v���XiG�45�o=��15�V�~�+@�+×�h���V�ɋ��k�bZx)�91���	�)�n�>v��4G��!&̍��`̱��f�s��<,u �ֺ��f�/�ۆ�k��i�w2հ3Ri��=�8 ��~6�g�H'��~�-%�E���h�Q��H$z��"�m���ŗ�;�L�l�l*�ˎN`��ЈT��>��fNԠa��4�(eS�e@�1ҋ	��p�t�1����q��ss�qs���y��E�F���Dp�"㣣�D��D+111qqq���			���P����edd��Ɔ��xxx�X,"�x��	��@Y����y�7���?��O�h4�N���ں�����������{�����2�K`�/����3��vuuutt����P(8NSܹIYY^$4^�())�2


0�hbb�#}�
.o	\^\<��x�n���􌎍������NDD�a�R_WOK]CCEUU^������
@)��+��4�$��ř�1M�m�T7{��`/'s+�po���fAAO�`��������!�>�:v��̭3�w�-��_�}v���ԅ�q����K?~���w������~���W��|����w�?�t�ƙe�սŽ�ѹ������������?{��ȑ&h·�s��t˕Je�O$A��A�a�A���{�}y�ʨJ�U�j3==�3�s�s��.Q��@VI�������>�����*3���ˈ�#+�˽MS-�]%�I�%�,�'���e4ICT3I:6�"����B3��>ۑyr���T�Rw�ɩ�u��֩�P��#�ߘƬM�W[#�̡��ZsD�	y��Zi����H�����%S�� [䡩�:sz�>-=��<��_]�+(дm����G���EM�$-gd-��Z�(�����0��~J?u'��7%���Ǿ�/@��i��¨��u�����|\�|\�|TԴ%mڔ5nJ�VE����)v�8/����2�3TY�"K8[͈Up�b1W(es\��#�D�9�1tJ,3D�iu�xm/N�QS^99b�i���$-/�g��K��5����u�H�^5Y�_K;{$��fƉM��,���6=y�ws��oo��o/������/�=n�x�d}#mv������2���9z2��)@Α#������Օ����������锹������ጩ���s{���4��<$��Mb����H���H�l|&��BƩ)�PS��ƽ�Ԉ��"b��P.xij���N��8ĦE����(�m�v��,���y�	15���?q��¡C���$��=
�>�4����a�7�A��lc|���G	��������A�S!��a����w�C�p"_�c�������q�డ��%��u�Ӱ�O��σB>��<~A�>��>�Bx���������C��z����~���k�Pn�;�K�������T�}z�~�#Y�S������,�K��^Hܣи�#��&}�<��=���|[��m�����6�}[��ۤ«T��ϼ��余��7���X������v��i����Uo��M�|�85���#-���_9�<`�/pޗ<�C��!:4M�0�:@

��䈖5���������ռ�����������ٶ��Φ����։���>8N��15ϟ=������ן?������D��X�lo��@�b_�Bo�B�����Z�KL3�1���
�;��{���;5�05�y��vK&�>�]�&�O^<:������_ o?}�W������W��ܞ��̌/���ٹRj:ǯX��T����cH�!�NO}���I��E���(��j |h�	|�u~P��ԯc$/f4�9V�BG����P~zL�f\��S�z�c�M�|�!��S3U3[�P�_l-5�`L�t�t�M�ɓ�Y7��>��u�l������RY}JTCrt��Ӟª7���e���L�5��./�Z�̩�Ĥ��}~{����g��~��֓��N�\]o8:��6���i�k7-u%.w�;�m���QA󿠩A�l�Pq�v	�](��)��)��+f��bQ�y��p>k0��i�iNg�f�l�ℨ�4iQuVus��p��D�ѥ�k��>�6s���7����n��l�4��+{-��D�b��5��ư"]P�_�_�Ĕ+�  �
d�4|$`�14\H��x��Vh�^��87> Ww4A�( [-���?����+�3_�T�Y�#����{eX �6t+<7�	�sW^WϮ�C�%��g��p>7������w�	����$H�|�3����]�^�9�
,��=� ��=�@�7�ך.lLԚy5�ܪDN��[jd�b����~�YXn� �lq5i��,}����� ҵ�l#?/QTl�%�,�`-G�SF"�Ex�G����yx�O��Q3���
�XM���Q��������G��FF�:�@����Ƈd+�`Y�	/50J��<eh� �gx(�?�����ǽ��{)B�Ľl�>q\�O"7(E�0�hV	=IcG�$16�"a�1�P"7�"�
�q�JA�F��ʄ:�ȨT$��5�D��j4&�L�s���P$��f�%���9^������/8������KNNMHHT(⣣��{ｷ�zk�޽И��
,����������6������{y����p8�D�R���Adb�X8*�����w�ٳg8����x��M�����3JHH _���$&&�����lvTTTXX84(����K&��V�=���@y��
�Y�!�`�������aw�Cn���!���"xaH�~a$���P
�*C'�։�):A�����,2f]���:��4��,�6˘mZ�@�I�Z�4�\4X�;�R�1�r���_?��?����˧��g׎?�~�Ň����/������y~��]޺tt��|��L��|������ƕ��ա�������dM��o�3u����%�فZn��Gh8�"�1/~m���ZǱɪ�������3:R�덽%��,N]ZtM
�&)��Qk��u���Ԕ�%|��05�|=)GK�T���$5�"ki�-(+Ҧ��״[�$E=��uIݲ�~C�pTԈ�&#m9)o>)m;%�>��8�n9.�<c���s���3��=�u��S��C����u8�0D�s��}��q��v��z��rB�|\�r�]��)����ʦ�œ���ؼ!nNO��8Fog�-�|-�%e��B6_�f�sXj+��P�#���RLE��4bm�Z�W�ז��;Lc��9�zeN����^�o.6�7��[+�۫ɧ6m�+��E�⬢��8:�q����_/~���'�L=}:��a���m7��_�\x�t��[G�[Y[[9G�����޲�,e�.g�-ٗ���Sg&Sg�3�&��#����CS��*?�,Ӝ�dN�Z��$� E�&	K�S28x{,.+楩A^zzej
y�b�u15��+SS�%�r���e8�2M���t��q��Դynw;�~�<�������+x����O�h_�ÿ���yD�
����� �m��Q2�X�8w<8�t(�B8�R8�j�=�#f�cv�c6�S����r�Wb�5_s9���a>��=
|B���u�y �?�s_�3�So
�5.<vx~��A�/���-���(���~����������'���S�����S/zG���xүxD�|�x�-��	S������,����ƿ/�����3��N���oر������{���8�~�k��������Ԭ�yCS����fSAF�y�h��q�Y_Ҭ?e6 h8�O�R�)�����pQ�ٲ%�����Z��X̴��fNU�וO5��t4�t7O�4��4�t7v5����"/@M¹�\Lͳ���g�/�?�qb}lu�ym�f�/o�׾Л2�m[�-$CS�0`��15m��]��Լ!�:gS�!b�����qťG�:^z����Ԁ�7��t�;r9����Tf}�"�,8���������/���7�~�������gϮ޸�2;X]��.�
�85I�ޅRd�Z�ބ4��� ���S���g@/��3��3����#��f3�s��
����bb�=���Scj^ǿԘ��*dR'h[v�5 ���P�"���z�R�l�I6�(�iP̷jV�L��3�oV�?�~�T�٥��������uK6�.9��̨Ѕ�	�,�$�g����фH���T��"AOc������'Wf�_�����'���ｼ�pt�`}�cjVzl��֥���v�r�j���=p1?����1�����8��l�`څ����������b�PI�(�0Ǝ1��c&K�ł�\���w�
RY�&FQ�����>�<�6ֿ2ڿ5={������O��������镅�G��'��3꺫TZN�*�&L��ׇ��h�zj�_��T�_R���48H��g`��4͉���j2Q[�! � 9��I
�L�l����� Mh�@��-�K�����+�gM����	X-�sy �`s�6�C;2�y����
<�#Z��\����*���:����՟
<[����7���;�]���̮�b;�c�� ���ʎ��gr����,i�]֒&nJ7$��l��Dv�!���*I��$�J������7r��tet�<Үf[�uve{aBOIbk��1CQ��+�DhE��ByBt�2�@\a�צ0����#*���N��V�V�͑`	�E��"]pUbdmbT�9,��`�hc��rA��Y��)�yrr���-!�%�,1GA�U���Ņd˃�J�����S3��\Ml������bL��8f�<6 �	E����*!�'��$:�T'7*�4�D�.Ѡ7̨�q����ndddfe唔���L�ɬ���bihh����;���[o�������?��5{��l@�?��?��?��?��?���?���o��W�����_���'�'��������#(WA�����?����������
���~��:QS���k>�6��p8�������c����x��r�QQQAAA�۽�����w;jtZk��@F�,�^pDa<& ������u��� ���C�{`y�<|����:a�M%6�c�rfR|l�]W�c�ҋ�*^���_��W�՚g�.I��Tf�X�2����Iq���tM�E���d�3�%]�I�m%gf{o���޹�������~�ˏ/=�q�Ι�k�gήo�uo�tn�v�M�/��.�5,���6/�5�����Y��T\��a����@�j��%�ѭ�U�Ƨ��z+-���-���o87_r�j�'k��6X�j��ץEW'�k��km�u�t�t�T���R#��H(6��FB����#g���dE�N>����ߞlOO)����6M(���u���Uqæ���(@�tL�r��v"�����~�N��'�G>����0}�8s�Fo��/�!��}��ݗ���!��[N[NH[��+�٥3�E���ؼ!Vv_�����H�dD+��jW�b	y,��Ŋg3՜(-�*c��)�P��� ���T�Vm�Y�VS��׮m�1�����5�Ӛ�y��r��j��icɺ����j�\I=�e�X�,/�,/!�g�/���W�_~5������z��k�u��������M�����	��������X�X^�Z]�^[�YY�\��/Ng.��,��̎g�ں[���eyƂtcf�)Im5+��ijV�4<]��!�cq�,\.�xꥩAF���J�P��S�d:LM���%�s�}\��:ʢ�D��°�T�n�g�ո����{�u��>xp����C���ܶ��/�������&:����OC��т?��ݠPΓ�'qGq�cĀ��q*�D0�D�t�|�R$�r	�5���#��r��PH~��-~�c�e��}��~�$���xJyB�,8�S<峀��$Tր% �׸���h��'�_����W���I��`�������{� ��>����G��;�v���I��Ͼ�?�3̕��W�QV���e��o��Gq�ɯznH�#:̺���ʿ�gl��<�q65��U7od�n��Y��[�¬�V|H�e_�E?D�8Ʃ�}�i�����)?�T e2�2�O��������lSc<��r*'�TA�fnΒ=}��1��5ZV8R[:�Z7��<��:��2��8�^���0��<��19�=�߻��������7_~�������֍ɚ����ތ���.�|��������O���oE��ɮ������8[�.���15�åG�:�S3.����p�p�<No��PЙ�mʈ�L�j�WVf+O���?~���o��7�~�����z���#cS}���iM�����Y 	(���h)��8@���O55?IӠį��A٥���@�T �:AS@�k�������/5�f��NY��}�=����T�f�b�kx����F�|�t�I�i����m'_X.�u�	pn�bk<w�+y���U$��De�I�lS���v��a;�>`dx�9�h_3�Pb�,�|rc�ѥ�'Wf~q���#7���-T��*��Y�O[�K�H�LY�5�t��UK���:�L�h�1K7����\D��*�	l|~���^������R~	��7ZΟ�#/|���]6W%����
��%�&;��L/Jf��j���&WGW��G.���>�t����|���Z��~�ޙ#�7j:J���d�P���*�RQJ���DZ��R�Ɩ��4�����k�eZb���UZdT���sH���d��ZB�ma ����߅��F	m�^l�дs�~W~��i(#PM���Akx]y�Z�'
8O����6�.���P�98�
;W�#;�%�
~5�N�=�߯r ���������V�M�V��ws�S�Ȍt�0����b>`�P�_כ��Ή��V�gɚ���6n�)�$�Uj�-5�K�ܒDN�����J���R1�D!9��{|O�q��ڕ�)�G�+�1��Eʐ2mx�6Pi˕c�%R��Vo��r=Pa�jS��H-���q�R-nK�	���-	6�|P�Y�&��*��sX[*�=�՘Ue/Մ�B���ʰ-7."/�a�9�V9�$�넱Rf87���JXQJW#i�b��5z�ҨV'h4	:��dI4� ��$�9b��ج�i���9�Y�y`��`V��<��L&���Co�gϞ>� ʚ�{����{0v��۷�:VAʝ���g��8t���'�H��;���@��KX9���6���b�@���`G���x<��5��,�G��)��8�'>>^�V��b�������	�����L!7��e6#�c��qX�?����������^�<>8�g_��C�Cn7V �,��u��xvr3SîLU�X�s�R�թ��<�HU�`Y�T}�rG�R{�xMFg��6Y^aUۤ�Y��"3�-[ג��)L�LM��m���� ��So�M�mM���/խׯO4oN��N6/�5,7lNt,6����zkG�����U��p�$iF�#��4k\8X���{|%6�t{��Y��zn���B��@�\G�p��5�_��(���[��maufF���j��\�@.K��MM����'ek�v%>MA�q�%�����Ύ��ʚ����)C�82	T���aMҸ!j�7oD�۬�-F�FTݦ��z�f����C��Ǫ�`7t	��>��(�w��}��u��~��z��zB�zB�v\�vLP��-��-c��d�D�w�'5G��#���ɗ�9^,[ˌ��Ұ*f��(�"	��gd���O�W���z�M�R���U�m�J��3-���t��	�˖�U��J��R��r��J��Z��f��j��J���}e�<>i��6�J[DM-��NU��nl�05i���./%���ood��:����
�I]�OY��X���\��X�Z��^���\,�^*���L�j�5T'�rSi��ʒ(O�SU�4Yx� 8�G���b�9�8GX45E||�������JĸR�R@���x�^� �:�cQ���p�`�٫��*܁u��w�#
�>0|�������==����!�>���&��5=�3��'���AA(�D�q�w"�p��;�;�;N<O']�$]
'^	']�D"k���_J��($_J���������<&�3F����"��ia�PB�$�|��C~惇�@��N����"~�F�� � D���܋�Г|˃x�p����K�pW�ᮽ��g>W��_y�{(�ÃAG���7��L��Vw�cI�S�U��Z�a���s�0ic?SY=� �~��f��g�㥦A����f8���Pz|	�~��@�W��3�I�_�+�\^q��t+'w1#}1ӾP�3R�7TW:�Z7��2��6ч�������25/>y�>��_}�ɣ���[�ٞn\�͝�J���tZ�z,N��'���$S����١`~�;�����O`j
�}��ݽ��bQW>�1=��ِ�Y��5���	2��߽������~����K3m���C��dI�!�\�Ha�H�Φ�������YӀN�s/>7�G��G^���İK�:�r��s���N��� �. ?5�:���K��q�5�N�^���m����J�lg��=_�[�-�K�����&�\�f��zj&��f�����W*�M�vu�5��(>_fbz�iU�}*�>�Mt@CsO�I��p�+��:T�魕G��^�����WV�ON���)=:��9d�o��zLKMJ8H�t�p�����E�� г�x`��lj �k��|g���#�R�H�p�R�P���X+����l�|�D8R"�Tv�+l�%Il{���1{l�ub�g|e`�������W�헏~����}z��G���
���4-3�R��H��$�@/�\���વ�j-�J����u$��+��e���1!��D��3mVZgrD�9�� � �`ّ���ΠM�� �]z���u���&
��6j^�b �/Z	�FAw�e@aآ��[T�l��q�!�.��z���V
��J?��3D�B+���v|� �F�*���;�̇��[��
,��?nLX���x�K�JT�EځBM��'_ٖ)�I�&Ĕ[b�̬3���.I�-0D��ᩲ����4����G*��5����LlN�k�sń<	�,�R�B�TS�l��zB�
�u�H�9�`�6�BZ�i���Fk0ȩ���䚄@�i H�%��Z��Km�7ZC�.�Fx� ��
��V�J���x|�:�LE͗��E�	�@�+��Qz['��g3DQa��`n$M�5�F&Ad�"N�W*�j�N��j��ڀ�h�Y�ɩ)�$[��`6%XA&�����B#\�w���h��y���}�]hm�*T3����_��_��	��kR�{RPĀLP�����ÇA䀭����{P $@y�����������w���|@a�9p� ����U*������j���15f�,A��� ///��|}}9<�V�C�6�����^�H�������������z�;�h�����{��^�����Y����i�xf�6�@ϮI�w�&4۵�ym��'�:U�9Z�ԑ����+�<�l��
Afg���$(ְJ���n��S��m�Դg �����
���".���rͅ��괱�������ɮ����#��k������C3ݕ�5Y�y	Vi����S�c	Z>٢KQ3R5Q)J�EF�PG5����O�5���=6U�9T�ԓ1Vgh�T%E����,�j[X�%�>1�VVm
�2��He	Ē��D(4��lޮĥ+���`ED@Q�zir����^Z�^۝ӳ����o\�7�H�7�� Q�vL�FD�*�vC�yF9r]3~���:�|u���/p�.p:�s��rZO�Z�35��~�+8����AOj	I�U��źX����<)�ǉ�p"��p-��c!C/����{I�!qr�-U��i���imՆ��t�ܰ~a\�2���`�\JZ[L]]�X]��-�o�%�����fnn9����>�`�^ZM_XJ�����&�̘fgtS���1��t��B�����f�����e�ڜuu6ie:u}.cs`_����do�n-�N���u��6��*�9)�d�1Q�h��4����	15�@;���!��楩�bᵦF�/������Zx�ne�<��	g����C!�>�O���N�G��G��[��ۈ��7������||o��Bi_DF~M�Ӱ��!!W�A��ē$��@�� ± �vP���)���H'�
�!]�SnD}��������~�e���~��~#��J(��H��R��H�����*���_�}��ď���D��CO̧x��������%��_H��&D|�O��H��K�p�������:���>��w}?�O�� ��~�Ǉ�o�#�����}wh����;b�}��S��K��.������^���W>pC��ȚC^k��<�Y���Y��_�X�%���!+~K���w}�i08��R�q�2m2���ԟNJ��_|���je������|J�r�}��h��h��l��~�15��-�=M����/�~�������'8��/�~���˧�l�k��Κ�J��Nw��z,�A���-?5�f���{'���7�8i7 �h^�a�
�;��{��^�wjƅט��֗φ�t������nJë2�M���܇��~�����<��_?���_<�:>X�ۘ=ܜ�od'	H��4�o��{o?��)u��n?Sr`w�Y�@S�>
ça�(������Ў�n� �$ܨ�����cj��ɿԘT�����C��? �f�*���:�\�h�Q:׬ ,���ڵ��	�c�V�.oV�[�8>S�4�5ђԔ-N��Ցn�Ú����C�P7]��6�[寏�(�F.��*8:Y��G[O��||a�ӛ��u_X�=6Qxj���x��p��p��Q���jw���AM����A�$."�AՌs;�ܔ���ǘ��긑r�X�t�F�Ң�hӭ5�k���qs5��2�h�b�N�S,�N�)Mf�j��##U3�]���ӛC[W�.=:����ݝ�o>��GO��u����@�Zn�Ddi��U!E�ЊZ�!�LM(W!��FG T���Wn �(%j��Z�05�N���T:��Ic@Y���d�-������:v6Sh݅׵W(���vu.�v�]�����*��3s����@aب�v=[�\�ڕ����xΠ��ow�= ��f:��i'��
Z =�ХN�X��+q��.�b.�cj��c`�7/v��?Z&+��ʆJ��Ԁ�BUO~\�]Tie���VibL�)�81P�eW��A.6YH��ל*;=Rq~���p�d��?[ڐ�(�'W��fSD�)�-�k^o"Tj����F\]��LjM
9U:̄���%9�5%,�A
X6'ךH�Fp��ʵ�j��_�ҷT�]�����V��+�^U*��?x�@�4�A5���xr��T�
��G�k³�a~���Tq��Hqt��A�3�QJ!�	U�Z"����B����eJ�\�P��i��Z�R0�PЀ�A�h���	��Ls��hj�}�q���|�s��h^��7{N�9�_�?���`yooo�D�т��	X��O
:p��/X�ÁM0��kK�ŰXlTT�H$R�T�F�Ղ%<X�V�4�����H2������A^�
���)�<(�R�4,��������8��~�������>�w�x��6���(��`����3U���J�9$� (C���VDg�ٲ�$.)�GL��j�,,S�$+����ӽM1�i��|eD���n���h��^�IX��/ұsU19��(�_bU��
��������BC�}��fi�~e�qy�a��r����6��2�.O_�*O��Xaָ�T#���6q��ژ���|o�>u{���T��Ɋ�c%k�S�	�E����sp�5�69���`��7G�%�;�<45ŉĢb����%d��v!C�������4wf�v�/&�M��eY˺��%��-f�fd�Zt�����j�F��5��e8ӓ����8�y�dʧ��s���hL��������n�[:���HiOj37�ʂ��5O$	�R'���p�������b��L�*�(��3C<������8YTR�Vm�O(HIm�0wץ�f��3���q�ʴyeƶ8��0��0��8k_]��-�/�9��8����>�H�]L�[�26�2����N:��Y�֯�Y���G�̛���č�֜ecڶ5��5cۘ����WF,��i�����δ�&{S}Je�!3Em�荊���d[eQ��T>5�G���9<R3 /4��q��D����:>��O���B�������(�xa$$�?y�1�[W�g��g��{���Q�C��W�܏z{�����LzJ�<,�"$�Q�^X��А�A�g��(�cA�-
f��w4{2�p�A�����L'_��o0��Ƅ�cF�g���c��q�/��0��WB�o%���������'���'�#��iѿ�, ���q�w�c/�S"�	��%1�7���Q�K��K�K}���!^����s����>���~����S7�s��G��'\݇;{{ܓ8�־)w�� ��h�]���w�/��>�у~�{O<��{�jj6<_j��L`���!� �2B��Z⊷U�Ӗ�sYW
K��U\(�8��;c�N��K����U%#M���=͓����}-��M��m���׏(���/����/�|�����ή\82vt�e��>ӕ:�i��0�v���YJZ��Ԙ��dj�S��	�Ԡ�v��g����d�q\�`j�+�5�����|����s�r�=����R��Ma�ɼ�Ƭ�\��Ձ������7������/}����ʎj�`cVz|�2�#�OH�`��
%�(M��7�0�AM�����Ů8o���h�gW�C�] ��#R�{������L��cj*�35����Z�\�x�Q�Ф�o�[��/u�;�[C�g�.-��_(91U�6R0֜R��5��tO}��!��y%0�
�'���,�u6?��Q�xz��׏�>�>��������;�/��;1]pt,ks(�d$��h���9hS��O��s;��v�e+d��=]�����WH����[�۝��V�JC�r}�|m�x�x�J1ר,�ץŔ�Ėe˛jm�#󋝓s��3�K'&/~t�~��+N��wO���z��X[cjL��Tmx�>�DM-�Q���U��2%�<> j��T��5`Y�'���91�Pӓ�@��Q])�I��Ԁ�m���Ǜ�6
���ʹՂ�姚����a� �9�{�6���:����D�g#a'��.;2�WOP9�x�(���\~+����pV4X��G��E @f��|�
�
�e'p+�0�A� ����	�
3���_�u�b;?iov̏�+3zW��^n��w.�h��2�@���P	��S4���L1���rKlqBt��(2!�lMX�"HC�H��G��O֞,93\rq�l��ڝ��ՇJ�%rl�&�Qh26$����f3�=��j��t���f� �h�@@���ؚ��D�o@��Mh�ބTU��o4`��F,�^����4�J�\�/�c��H|M�!�\�%�Pr�\el�02��g�K��
G��*<_/)E�x�A&��eRI�L�P+��A�M��L}"H �#H''��%�����8p護����{�w��󳟁����������xK�0Xݳg/(��{�L�������?�s�;�����g�gHHX�@aB��ah�p����������P��!7P-� 2wl�����^��H��s��V��L��F�PL�G�H����{�Su��{
����d2�H�9��!D<���������?������{{���{�!����wW1(6AX����d�I��d!iB��dKC*��Rml*/0W�& &��^�*��!"҅$�)�Xc1�wS�O�2�9UT���6� �zV�:*O�(�1��~��W�,,����UJ��G�f��դOw���4,֎��uV&��ۺ�R�3�l�t��dUF���V�&ʮc����4��r��Xũ����uǧ+�F�g�m=�����R��FC&"�1���5CSTn"��H%	�R�4�T�@D����T�,!1�'KFSFb��оֺ�Ņꎁ��>[���qJ۴�l^Q�l�Z6%-[�#��#�5�ƣq��c7↮H�.�.)/;N�� ���Ҟs��S����vd��15�'��'d���UK̂����0K=��n(W懋,|�\&��9jSǏ�s#�a��!�l��KM`��dU,Q�+��7��
idR�Z�(3�&������g��&{4���A���ya�:;e��L��J��I_Y6NN�..?Qx�X��V��6 keþ������������������կ��L��y����9�|lɶ9gۚMڜ�����3���>�D�P_FkszCmvc���Ԕn��:�(Aɱ*�6qD�0Q�O��r�d;3 ����bx8��� 5ߙ�r1�#��{���4*���&���p�h(v���CtUp�+���ϫ�ۣ�����9�5o�c^^�������~�yX�� ����;��kԠ��i
�8��F�=p"�p�A�M�ʠ^�^�SnFQ?�0�1#o�i��L�v�'�������8�_�y%������W���R��2�f�6���P���g�c_�#� �����N#
��{��3B�߄E����C�
 E����!��<0���Cx������C�{{��y��y��ȃ�C��r�w�r�z�v�H������:����)��c��m7ߍ�^��O�����|6ܑ��O�M/�u��o�vՏYq���`�c�1K��?yڏ4�O����(�!��<�q]�����3Y�
�/���.,^MK5���ٌ����ɺ����������	�� �f|��,��=������>��*�o>�W_��ϟ<�s��٥3[��S5�]��v�D�e��6�g[Hv`[@bjV_��,����K���.�B�0���ͶK��҅61|�	
��& �4.��G� ���x���>輡�IGL�I�.%�ʂ>-�֢�L�Q��J����Y�8��N��@�d�JY�{	�o(<\;B;q���E��2 � ��=yH��Jb��0 	�
6��]��/5�E����決�c
�=���BQ{�1�]�U�]�&�Nm.Oښ��ŋ;�����/ܽzfuf�����:��<-]�0���4�XI*U+����TcD�6��&�#���Pk"՛����@gz��v�Pe�F����0W�1x�uy�E����ȁ,:�.0L Wa��g��N\�J!�K�����R-
��@��?�Ѣhx�C	/o���п�ʄ�;q��Q�j��p�u�� p/TЀ�Pм�BW�y�5��Z�l�p�������ի��#I��2�M�\��;?W�6T8֚є����MB��G�����#Y����h�^��ϓd=��˃�7��~uo�˟ݚze�Ω�˫5ǧ�7����7l���� V�Ջ��
d��z18aؔ�3_�N��sv~���}'.���8xP H;ڥ5�
�G�2R�-单��y�k�J2[-���-7�W����	�]���B�f�Hܒ�/M�7V�g���G'�'�6�|v�w�������յ[7֏�vf�bM2R��P�"Wik��Z�ZG�R�A��Z�w���P�{I�cY��7��PC@S�� ���	�T�fJ��
r@g� {�;��l�@y�]~��?�(��(h~$0�r0�5T;\�K$''�/�{�i É,�@N�`.}(� 	�ڛѝ֓ޗٟ��5�͋��	��k�k�k�t�Et�Gz�"
��_�ПїޗٛIGq>�]��Hv ���	�75Z��K� �`	�4�uP�/����Z�I���;�P���K�x�Kpw-R����]z���3�g2�͙������VBlݝ�Gy=]Gbjz��ݞ��#�G"@�@��B3˽��i}kh�iBe�<+3�4��J0������%[�rE�2hJ�����KC&Z��0Ѩ�)�乪Y� ��m65����Ӭ�*�����:����mꋙ��������?`%�zP	U��%݂�,�6W�4>��|~��Kr�$� �Z\.��$�;fxr*���-�^��-ۻ?6dy��}X,rA.h�����E#��QL�R���ԎNC���q�����|�Ӥt1��.����l���Kq9Aꭚ��1�Z���������(+#5
���t�s�#���.ȍ|E�~�cl�_�7o<�{n�:N%�~l�0 |��ގ�������(����!���l�������cO�;��ܒn�!9=�5Qp��� VMK��?�"�����ΖO#�a�P�`m�?�;A_vb�/!�	�ys�cc4˓�A ��`Zl"^mY�8I�G���+~�!�9&�Fo_�0��+^C����
L{C$�t'�.0Z�x�E�&|>n�E��\�_��Đ6��	h�U/�j`�{��nk��b�( C����aE�))%�~'iV�O�d]Z|���d�Ħ#=���������m�Ǩ!?��;#�4	b�M�+�LѰ�-Q�6O?�o#εʬ.I�0�b��՛�����4�kU2�N@+7s_;ܶtkѳR�-$��4�h��S�������&���vfz%_�j��dÜ)0{���Vрf��b��"���ϣƦ!�J.��^\�lQFnxh�Ŀ�l��т�|\��5K�
冶��oaZ{��M$5ܷ�d%tT<�[+��%O���
P�}9�w�t&��V��	Y�L(�*C��O^�|;_ݙ؝�H���HZK��aɽZ{O��K�5d�)��8,j�s�4�w�)��˩����v%��Q�4?�e툔T���e�K[�H�����w�������� }4��������]��X�p�h�sâ �.+�AQI��8���TO��жP�>�I%H�hJ�9=�럏M��M��+��5�fs��{��^Y�Y)3��n��it4���cQ��V<�C�_e�0fP�D��Zk��紼�d��k�n-�=a1E��3���+[;�%�E�n�꓁��\�` ��k+�N���oX]��Y�0x��o~E�_��y����n(s�������zaY�cOxį�h��1ܟȬn��.�sGoE�p��s%w(7����|z2��[��!��Jq� ,q8A� Y�6
\�4b�,ya�
�'6��W�̞6����&�1�]Dx7T4{ڰ��nO�۞���p)�m��i�F{����uW�n,����HQ`���������^�#���X���<�\�5��[F�ß��@��E��,x��O ��'����O�aT�&NN�e@����5�� ��׈wǳ�OD;d�-��]9�H�(?�2��'����s?e��L����^��8���Շ�՛����ͻ+_8��[�N��d<����	�����o�B0��sZ.Kv sr�/�,[�����8bh�gn�;����;!
��,�]��R��tU��e	������xR�hZ�����8YJI_Ɠ��w��M�+����]��hܾM���=�W�~O�����;�덚�����%Ш�q48��z �=V�ejc��c�I�xf�Fz����s��.����/����w����ݴ��� �kW�����\�!��&὿X荾�.i,̫8{\��݁��gw�o�%��H�5u^Ty�3��sd��ȡ�U;�TP���)~;]�^�&e|7M:Ϲ�C����C�/�~�+Ẏi�������36uJH��Z�_~O� �WD�-�S+�-�J ��)�֜���1�!z`Tgyw��Հ��12f��j��6��V����އBb�:T�X6�c#։Yw/��ȼ�4X��S��6��=D�H�X�*�>����G߽.�7%J��VM�건����AL��s�gS���+ިY�	��@��?������>�\����~���Y�Qa��.����x�����o�`޹�&l�LtD��x<�n�R �)�>��tG�^�
��j�����u�19�٘��Q���@#%Kͦ�d0������}�Mڹ�jf
�X������w��c��)8��(붿L�e "��忽��fYN�m�4Ԁ6�3D�G�������@����
k&6���Ӭ8��{O� �y�P�5q!���Vn�7�O���K4m�g���j�\F�������D�>��;��� Ts^ ����)�2 {���"��PRj=�׸�:N���-:��C7��g{Q��]�r�=0�Z a�!=n����(Y������j`��d��D�C{I�x�1F��6�G  {���f ~=�+������	Ti�Nn�� -����8|�:>%�5.��)Qv��`0�^bq^������x,�g�w�Y���"<�6�B��4��@�U�+~}����M��(���En�,U<�" ��C8�3��O|fťP>������UJa�{���Uy�u�a�e�,�a��>87V���ר�Ƚ?�������Wa~���Z��20Jq��\�8Au������P>=��F�E-�R<1����G�ǭO�e����V����[�㆏/�l`�%���G_�:�7)���C6Ɔ������-��o��W���+%T�奈�P��*�J���ͧop9��X��!Z&r�[a����N�Wa^إۍ.ύ 
�M��P��e�c$�Ǯ@@2T���n@�-ԥ��,?CG�$�41?�F|z~��r��y]��\�>o~踯�\��`ʝBFw���5�(�vw��K�/+s~�}��E��>��|�nk(�*H+�]qxd��$H�t5��
��H`|�0��xv�.G�@�g� #����vŨ���X���N�[�j��RoKkq��Z�L�m�<w��v5<s�������~�e�p�p���B����`����[��]%(l�
L�ֵ���)�׆p0k�k�B������2$� ����P�h�{B��Ƶ�3p�P�2�X�
�H�w�*���;���k�E~׊�Zp�y��֐.�0���
�X	�T�bF۔�_&�|U|U�^U�|�G}U�^����N�pݥ7<�|��$7<����<~���N��F��y#S����9�{�M1���A����(I!�����P�'�F�R�a/�������:�W1*��g%n�gN�$�X��)�*d�+eg)��k��ǋ�&~�Ř.�!����̸���̎��X����DۻSy�R�>�od�<T�7̻��ԙLw� du3��s��� ��t���£�*+K�=w�_e<4R�4rlf{Ș9�,��pS�b�p���2�����$��];���f#�0`��F��S�Zjh|
@��c��LU��v�ͫ�h��V�J�D\�Mؚ&q*�}m���p����-;�4\"e!��]��P~�$����ܦTdX�����]��w;9����pҟ>u:ݰʉ��O#���	
B`������k��/�$�G<���6���	��{��zx�J�{�Ԥ�~<�����K8~e��-�>9~][�����K�/�0��#`�<=�D�+��{�0/�^E�D��;)�߹BޛI����,UÈ2i~c X�-���L~'�.�%��w��(��{|)	0��A�{�2ET \�`��a7�
�:����
�1xc(�I�N@�E}ޒ�N֢;�`ێ^(b��"5�\���g�|���W�k���� �i?�@G��L���m*6��<��ݛ��|1��Ss�� Յ�����y��-���Ӕ��(��Λ~�Y_��ݛ/ցX�Rd��|����"��7G߄9A�)��R+�sY��
�����)�}2+�Ƃ��"�?� �P�t\A�g�Zt�Y��fn��9?/D�EQ�NY��0Z1�udNTi��&���2��1�E{Ăٴ���k���I^
�5R(-*>�M�lf7�t�}��`��BJbU�R1����}��dXN��E�)�>���fOI��G�G�2j'dve��$
���V:n���["݁E� �����A�zOO�v��b���wV)Tԗ��,1FI���1v����Gp!�� c�+Zσ����t.'��ي�"��H~3��%lgؗ 0|�����q-T��1�1L<��j�N
��7i��~BY�Ō;�f��¤��>�r�. W��Y�Ϲ�A�s�
9�:��
*�cٕ��ݸ	���|5�|9���~��lT�R�OA�/G^/�/�'/�7�9敛ӎ����%i�+�1��f��X�&O�=؅�6aW����xO���=q�a�)��BC���<�9���ryW3.a�(�(���fa�{~�@[���6:3+�׀'��}����i��*��+Z�Z�*�n����6��2}�Aa�����8I&"��{v��^����^s���X=��^��F�����Qt�`��Z)*8�Z���|wt��^�6�o_ �,��a~ډ�p��(�-b�db3�#�&25��[�)��@��T ��$���Ǘ�G8�K6M8��0�}6�H�I몸�`я�8��ʼ�ȼ�Ȍ�8�����%CC|@T�K1!uG�YId.k��-f�Ӿ�!8R��5:����E��!�h��R�������=��X����m�@48�B2����Q����%̢A;���[�вE�ۚ��{dQ����\R��]7$҅c�Ѳ�y��^F�O�۾�����bz�����M{��O�	�!���dP\�� ��1ec��^�ߟ�`G�0�����xə05n���JJK��HPh Y��,�O��^�It��o�pcVF,1���u��٪,�C����3dI��JW΄���j䨵��ă���k��O	�nD�]���x�h�܂�L��88?߿<��ڭ��d��;�����||p����7p��L�>��0�fԟxÇ�o�P�ŎbH�'r�Qa%wc��笚TK uתj�L�!�1!���z�'�3��`�NR�,9�8Zl���W��ۿ�"�(m�	�
�x���:��U��U�d���ÑшE����K�Μ��yB�I'�1��Os�r5_H#Ӊ�r�w�l��%��ƔsÂ��_��y�2��)⟐���!�9?��i�1�|#~�-7ާ�]��y8��t����R�\�Bc8D��ʆ�~Z��W�`������͏�^�����V��P��`@/Ag%�r�O�T�`0��n
n���蓏��Wl2�
Q&Ҙv8���:��1v���j��c�~Slz��[�k��J���4��
��O� H�dk��J�Ϋ�C)ێ9�-���r���$n�������w��nm������t,�O�H�.0�*�V(튺��[�^[�dF�m?l�	�B`��>N1�!�Rs#�'fK�>����_?������%eA'mnӌ�XL*&�U�5��I�ט���C↉r�9hE:퍵7���������l�����m�������t�Gz��4c��ؖ�3��Fǯ^��_�1��p����<�/�����sY��D8�TMX� ;�#�)�E['��	�%H���y�m�Z�%g����w V6�����ܠ"j�\à��'e���}����(�7�ȿ����{ ٫�ҳ��ŋ��}��͋=P���B�B�^�����;�q����~�H�6�u�a/��o��O}	��={I�g�ӖX���G�D�Db�DnID98�A�-}��$8Ϋ=d���0A��<�A�A?�-?V�}��J�+�����we/r�Θ�v� oij��˿S�h��Ga���^�B�ׁ1���
��"Wa]����ݳ��I^�D�n��Q�}�vKG�D��(~�9�W=���}������U�Fȼ��>G����,!�7_E9 ,_��²�P�-� ���q�aG�ѧ�I�;�"Τ
����/Xᜅ���B`W������=}�받^�"8z���s��TH��y��|���*6�(2|2`@R̯oѶ�]���<����:.���L��wsU@b9I�K�Q�˯�Է�"�ټ�޺��(�ɚc?Gbѕ1���/���k��g����1����y�#��_��/�r�IM������g9C'��15gS[Ģ���lr�rC�灘5�M��Ȅ�pn���Ze�A����l[���sss�5�3-Rrom~�_�5T��z�=ߔ�L��NN��mF��i�|>SI'������FQ��@S���:��-��g_+p�%���wR���ҥ�/�.��׳De�a�2�T�KIq�Jl�*� ebq��'�}˅7m=0�Z��sK������2fq��f�Dn6\����	�����qp��֥����?�ؒ�����c��Ȃ��[��[�գ��[��i�[�cݸ���%�J��x�)��������� ��E�ɷ���b:�U_��?��/�����"�0B�4������i�;�J���׆���o]W�=�_�+g~�4��q^&x�_����F;~$åI��u`^��K¾��a.Bqi����ю�n�Ш�������{�S��XY�F������r�p��ܨ��u�zwWgr�-N����3Q?c��D�|g�z���Q���ͽ�.,��';	��~lX8��^^��x��}x�b�%�ͨH�o��N�;�����7\g*�����\|"]	F&S��&�8����ZAFlˋ���_"9���s�~���#�=��D���s�P��}c��_>*�����"rڎ�+�1�E������ɉ�h;ǖ���q�f�1,�X,��יC�q�o����+~Q�Ѽ��0ҵ#���c ��t���1_QP��������ƭ��O/DK��$C�m;2Kyz^9��a6 *��s�tI/��E����~_�>�j���x4�jFEǖ������k��#�M<�,�ޑ�] �߃i����7�a �n�6C�;�
N��<ev�CFkT��&��P��NwC�@�/Ȭ8�J�um���6ȱ̂�Üp�ϕ�K�)������y�L\bM9Q']��]��=�1�ڋ�D���q��'���q���<��� �����j�ԢۑWt1$�;S��h
���ڛ����(�A��R�Ƣھ��d��E�3�2Ċ`�r�>F�^A,�B���l&�7�u}c��b`���@	5�iF.��4��I�+��4@q��y���D��Ӊ�
P�Z�}��}�x��~��x�{zQ�,��Έ���i%�}jk��x�����w]������lv����K.���^�0DL*���y���J�!�r�i_�`l[����h�+Z7�*hdi�<���I�xf�V���{�z\o����X��f-�b�������O��
D�aY붚6�g���#��甃�띰�}	���$���2e��t��/�Qa��&�Vm�6�q:-�#ى�O@�>������W���<h�T?�epo/��8F,�amr�Zr�����^��-&l#��cx*�y*s٪�8�(�O��n)�O.|��9�m>&l>.��/Ʌʸ��XǱ�������ġ'/V!�ż8p�����6?PL��݉���o������	������q���ȡۋ�:J�������e�9��Al���{�kɄ�B����!#<Bє&u9�Ok�e�۵��\<�_��+(i+��$�쩒��s��9A�p�o��o��o�&�B�$�:��%����`�a���XvX:ױ��ԽIU>����|���V�؍,3����u��9��8-�H��0Qv4�a�[Z����I�A����{-��m�K��C�F'ϖj�f�����8'{�mW����H/E�G��l��X�J����ex�a1\
ylE�sH������wn��_cW?��d2��ն=�Iy��@�.tl�쾅�~�>��f���#����2R%7�h!�c��Hs�Ɩ'������:t�"�Ö�e�������Y~�Y��:���6F��#���U�x�I������M�?g��}'�ld�N7祎�v��U���[4��4B����\�Э�^O����Ǣ�dv�
���dƏ�ε���j����&��ג��~12�����V��ui�+dV3e8T��9f_�e�;��?�B��c,7;��C1D:��fJ�o��+�X�� J��&�
Y� ,/c9A��Yu�5}�o�"����������P	E����=z0xq`.��1��o������T��*}Eg�\�I�����9�GQ=��c�=w��8��RS��	v�$mk��s��
��G+�ܫ<�]./KN2
:��j�r����{I��\��O��~3%J hKE8���^��F8~WR튀+L��m޴�m_����o6F�������"mY�-B������Ɖ�w������Y���:��y��2���ljE�����<�v���	�łQZ~TO�V�T�n���g2`ߵ��|?!�i�x�i���s�_��X�n��N���:Y��N�&�������y�m���h�Ҟc�Yox����aצ٤Q�y��˅*[�pO^e�>oo�V��o2�3�w� ���{$���"�V's�5`V��rm�lr+��e��э�E��2K��JxVb�#َ�J�:�6֯p�t���y7A��x��ݟ_jy���z��g�ZB~j���uQs��}�M�1�����$Q�W�H��I��d҆kg����^���������@�C���6�L�)���S`7��X0�ՋK��W4T�FZհX���X�Xt�H|Ƅ	���c��/-YP<=�5���{wW�WP��-h�y��	���ZPq�*#��i�%Å��Qm������ie�To�]�@j.J|ЧU����!hE���-�F���Lg���9c��3?����{kmAH)2c�4��g?��@S�ZHGI	��>$�S���WGjT#b��:�MH��ak�
�&��!��i����i>,��޽X::����\n�!m��i_���jC�tH��^ɘ׾�ce�Bje#�U�kM����nG󓀈S�B�J�X|d~HP�y�V�H��ΨgR��d�F�NLT>y��ת���<��hX�L��\��X�(f�Ʉ__�HҨ�ٓ Pe�1�#u%���������8�t8��7��#��Yr��ֲ���딘�Iӧ2 (���� H����z���,�0��WVJܬ�4���5��d�C��oi���)���a��u��R97����,��]EÓǑ��i���/�.��*����넁��k��奻����:�Y���`��sϤ����9p��A��({֩�!�b�J�(Ɗ81�	���#��R!w(n����� 㲯��QB�I��jrs}���%v��ճ�\V��S;�w���Q�*�c��Y<�C��8�ߋ�lRܤk������ESb�����I1���S_oM	��~{�����׉����g�r��[s��d��{_H�"j��H]˂<�����5��@���(u�s�O֕���ԏipW�[|FE��ނ�ҹ��l[�O�A#���O���Ǭ$�H�V&��*Ww���I���H���Չ��I$�ɫ�
&��)�ΌK0*��1�r<�S����ϺHJ+Z�J6�IfR�����Q[���t�� ����T�+��ϋ�k���X��ji����k��-B<u�@��z��0d�l��9�v����&k�E��d33>+���&ݦ>kͮ!S:[����;jS�:�=�h�M��͗8l3}�P���/?�z׭�(�2�hv�Xw�Lw�ԠIT~��W��6I�}�Fn��O�ԓJ,�A����c�`j���a�҈�r5C�h5�{�2c�9#' ߖտ���ʛB��*^dFW7��ׂ����)�����&���zc���1�3���Ν��އj���z�%W{�LM$��U�JUwK���#��}ǆ�Y^�t_�����L�D�Ê�ݦ��'�?����&{GK{v��;��R��,MV	ax����H�ҩ�Ji|^�%	:"��S��<��
�U���e�0�8�����r�o�$�شQ�:��[J�]���IE�-�Rm �6t��t����F�먡���5��%㏘@#�ݝ�N����)�` � �*)`����b����m{vNa�j���.�ܧ&j���7�R��.�M�3���c���+M,Mpq&��<���j�2���Z��hd�Ss����즨������������G��������A�&}�O}�����z��v��W0�hTD�ߔ
�)� h+}�Y��K���M��#��&-��u�k�͆�;��7���!B����ܞ�#)��R��fbM���0�&�	�*oNX?�
���L�5�݀��2z��RH=���q#�c�z���G��a�]�f���!�!xO�o}��'�������`b�W�?�ڀy҉	�`�}��q!�K���-����ËaP?;�ҖN��M8
�����+�M$AN�2�;�@쫗�f��C�-Ƭ���6��&���{�i���X��׺�ާ������I�B}���m�=ps͡ݵ���4��`�wK�Ө�������υ�������:�ǥ���n��b��x�2��R�M����/�,�'���Q�����V"^~��������g�Sb�Y|9�;��[G��}���v%*�T��F:ګ��-��ڮ�[�Z�J�����gr���K��-d���@f��j�7�}�:�"G$����f�I�Eat�4�_��;�ʨ���$�hH�hH�C�@4�5�=넼:c����nx{�)#+�Uh�9J;��/�E�Z_���p��Z �|5�	�zc��z��gαJ���E��B=��}w�[�RAj�xr�a��//�K��i�5�� lc<3�"�e�j�N\���Z� �HV��:HFL��?�&>����c�:4��gJ��&���濝�6�N��������di����Ș@�����Y�G�a�a�"�5+��kV	�f�D�����5����d�������ي��8���O>xWz4
��'~�p���<�'��r�2Xׄ/fX7"���m�~"�(�
ܧ���G��O7� έM���ń���B T���f�iu)���Umq������Orwxջ��@�8�X���l
�M��y�OF�xf�V��!�'i��+4�䪗�N[��Ws��aG���6�����6$�!y��'���7���)�E���eQo�L���R���`6s��o���'#�|5�n0�:�O��a�)J*a4�xx7�;4#�a8>1R<\�M��s7���G�����s�M޵�'�)�Wn�َ�(4�U��pv�!��x���a�����Y��q��
�|�2�j����c����V�@% QOJ�,ɞ�#I)�G���7�\�e9��ؐ�8���$&�L����4��Ս]���x)�6�y]�Qgk�*Cϔ�zC��:@�d�<�E�#�^A-��M%c*��G�2�
#�E�����O�j'�T�C?z�E��p{d�<"��gy"��U,9�J�1y�mo����o�<�x[eideW#M`-��|��N7B����c槒��=�zh��.�y��.d�~7��AI���v�'�.� ���ɵ8�v*�V*�6��v��V��.��6����X����쟍ّ���Y8�wp#���y��LR.��v��kV$�r���?5$��(鐮>��E
�<�gWg��]k��y�}>Se�i�v�v�Bkx�k{�X�H|U�0�8p�=Q-wǼ5M_'g���%���:���L��g�Tl,�fGWJ���:L<�;:l�F�VG�ܝ{xy*s�xƔ�p,d��#�
���}6Ljm�^�biS��f9x�,�I�cSf��9�­E�J�"�b�2E��#���"�!��V�o���#���������Y��A��x금o��D�^w�k/5Y�o�/��w�����J�Ύ�1���$͜K�o8.��8�@�;F�3k�?����jۋ42�����	P�Vpz�b��12�(j.��0�pd��$f��ZN`�;2�'b\�n'������\���#��pq� y��A8�n�������Ϡ���}S���] 7ᇛ�˰���ǩ�+�����m��ZO���w9O��v�{�{	�!4�{�p���i��'�5=�3FGҭB�^$
�tv,����8���ݴ����%)Ԁ� ������"*��?�ccD��ɵ���A����x�]Z�nt<��������������-�F�ǃ��bz�9�l��F(�꼸ԁlQQ�aj���w�Þ��r5q�<Ȟ�)�
���K��m�C�h@(o@./�4��u��ACo!�Y�p�&����/��������(TZ���TU)�/�@��}	$����H$�
#Vf�Jƪ$r����)�ߟ�Nθ�ꚥ�6���A�l3Mm�o�X[;RI�$�[��J�A�@�u�����0_�	����������	p]Yf2j�K��� ҳ;2�nY�wUH�p�L�?��z�N��z��P8��<�i�7��5g�,C��)��:�!�x�l�o}��c��s0= K���M.���������	 ݩ��DN׎~������'1���հ�`Hx��~m~�%8\9��`$Kj*wx��3[�hIǥ������/��ä��ħ/Bf�<��/������������8���);�R�_���;�s����AQ՟}�Yǝo���kyF6:�L$E���fv��{vۋP�(�hۋo�0� �`�-ݫ�8M�5>��5��6��09�����o&Kp�=�`�c<,K��:��R�vi���hp�2��ڴ�>d�.:؉��]�%&Fe燋k5ek��3�T�0*{"��������V�ni�e(,*�3ߐ`Y1�,U5`@�s<V8ߛDj.��J����鍙��C�v���D���&��:��9Ŕ��R(�b� ����<H�,k������,0����ݖ�ǃ� *�t��3�r2��,_mP�݂�������WrO����0����Bw��3���l��7�M����� �E�e�[���ބ� ��︂�����Xa��s�����#���4�$��H���ԡ	4�;��q;�!�M��&Q�X���t��}���P�d�;&";5�5�j�<�����O{:����d1��p��`�s�cm��UFA�а�~��w�@�/Ԕ`p�a���Yb��ˤzX^C�紕���I2|UZ�"Z�	��� �A�.����[S�c��4�	��Pf�{j���<*Y�QO����5��]��2�KgJ���rgI��8��?:i�O�� 4�f�O%��SBAB�U{��%wظ��8D����b��b1�5DrH�f��D~���ssQ�S"�O���G����v�I(ƃ7y�X1{.�T:���xH��8i4�A?M��P� x�[�)�-������M~!����[���V\n�d�3��Q��LY�܇�q�������ڽ����]_��������I�ŮF��#Qw�P�'�<(�uh{�lv�Q�l�]͒�:���<x&�MH��`��c��b�)F��2���2oU%LK})rZ?��&![��[\�����*��ȩ.����Ťd2Ƒm�wz�2���,5�o�M�7�8�]q-&�9�Ha��~ev�ˌ����rئ��������rh\�Hk}�� ���
�-�#�G�e�!1�O>����a�"�؈u�tр�\�� �1�0������T�����aHS��ZW�Ǳl�#�\��퀣�v-��?)���ח5��iWP�%��_v��}H_�ܼ��f)T���&j	�mU-#@�w����Aa������j�9�&F̡}3Hd�Q�z�E�Ta^��u�R��H[��++��3��˥.-�,�)�-n��0�Z30�(�;�T �k�m���H��Nц���2M����a'�-\�����
p��IMi,�w��\��K9E{�ҽ��y��8P	_Ip�l�WF���Vn�Zm���cf	���ɔFN��c�}v��z`����	Õ�R�aH��0�� S�% bd�!e��u;��Vu�{�P|�X��Ϭ�O���-��TO��@-��;<�#w�%&���������~��*�e����\��z���ޫ�˝�
��..}bƚ[�j���B?,����v���I�
*@1���⾑s[*�8y7�	5���8��J�̛�V�K�x^ZĸJL{�w�A�b�w��������|��L���]�<^�o\#���9��~�4�^"�Z:�~J�B%����[1���_������_��b�xN��y��qڋ�D�8p��Ӱa�r���&���-j��0���Y�G��kTY�T[Zn��ke�R>jV�[��И3r���]�c@[��] !�Ju騴n*2��$W-D)K��z ߝ�-P|�ԫt|\��Ld��wN�x��R�Ws(d�߲K��J���\u�ѱn-��O	H��?a�U��gV+�_N����\�z�U�i�.�O�^�����?$�0 �%�ǣ�s��Fn�J��15����M���R��#U�/��E���EWj=�KSG'3�I3
r>E�Y��Qq\kw;�C����wh�]d]ST�YD�M�,��S4�E�D���O'G4m�;�an������<����r�t�֣砋�_Jhɠ�R�X�g.P��~�c��Xc�Z��9 ]&���z�F����S6���J��!��^�Mb���Ҍ�}��?]=sc<#d�VM�q��v�2���9�-5�.ޭo'���q/��+����W���d*�"�BN���3��)��h�����wz�+���+����Q4ڲT�g3��X�j�3��Tq��e޲#��((���1� J�&��ϋ΋�Rͧ�\��|�����ls�۽�J@i�i{Txo���	ww�z�S�	��W��3���˃��o�����_W_�������L��+�R�L��`%g`EM�nb�YUu��oq�NIip%�!�TA����e�M�pVl ݄�����ɬ&E
h�1����,>���h��yg�
�7�#�W'���������)��ԑBR
����r���b�z��B3 p�p�6���ڡ�C�s	PB��*�_�J;Mr�8�m��������	ש,*����uݖN��<��2K�	w�.���p�O�l=������QQ/��6N۞��)?�">���7m4�g�x�����~!���bD%nr���?4�g"��'~;k���"mw���)5�m&�����hκF��V@=O@�N���C˽�mlp�OMA��a���2#)p���7���9٣�̚ܒ��HJBP��.�)�`�:�f�S"��PD�|ᨑ��z"������%�.ʂ�/)%�=L�����d�c��)A����ۛ�K�8::�DS@����/ջ��ȫ��]�V��E�����j���g���ۑR.@rdbaT@F.�;yV��I�k��=��16�8�8�:��5�w��!�����$��[�{}JGO���5H`��>#ʸ38޳(E��C��>���r~?�̀�Ŏ����@�s���n���ki:F=���s?C��ŉǉ�Y�P�j<(Ւ?�i�r�Dn�.f���ۺ�E��T��j���ݭ�����ܢ���P�s7��t����{U���{�'PM�z��؂0��O�)Jx-�ͽ�v7�`�Y ^9��`�Ao��?�AP������X7Cz@m�:��75D,�%�T���.���$\���\�[8��K3�a��K��Z��V�ߔ��Λ��1��W����F9
P_򚤿q؟J�LW���X[���'�&��9��;�y�N��NU��k�^�`����b�HT=2�>�׊g�
3*n-�6T��m�% yR��N�(��J9�X�M]J�Q����8��b���i͞�"J��Y�3�֨b3b}���~�[���@f��V#��Sg1�ڑ��C�f�x�REg��ݡF��+6e�̷�/:=�9�y�9��� r�����YJW��J0ֿ#�(A.V��r�+5Ax�Rl�,���;��g]@��6H��?����L9`F���aN��R���R�D*��,����c~���B�p��5�j�8��߫��@{�NSs���r ������0��|j�D!l�g�?��z�N=F���@�������oń��D��F�y���86
����������aA��ɀ�C�P�S>"`��0p*�~���������_hd@��Lhp��A�c�4�OHw<�/�s�v�纻�5O��^�k^ث>��~�+~ī�$�<������ŝ�%��C8�O8�O:�!�'� l��(�X�r ~�_"����!����s��x�s�Ą�V���{%wʊ��e]��>��}�0�Liީ�ʹ��z>^����J��<q�@�-WL�&����Ζ����ᶆך�g�|������㯞?y����N�;6==R�ے6ܙ>ѓ
ǩAG���,��V�"�5	�י��v�r�d��5���6�PPGz;��ɚ��ؙ�\��0,'+�1 ���;
�i��7ةx3�N�
�v�A�����N\v���a��u�8p��Of�P��4��s?93Z�t�ƙ�W�5P�8� �� ���7ρc����؁^w��D8P!�-���s�����<yQ��.?����ƙ��w�޻r��Kۋ�}=�mM�9�*��l���E��T��S��M�ԛ��1���dC���#���q�'��7�X���	*h~���(G�A1k$�pv�	:_6�+U�N\�A����h�o��޻Z g���Zg����� x��|ga~3��ɚ��Z�Tk��7��-4��N2S/D���֋�����n�f�i�߲5�|l�~j*��t.X���96��ړrl4��Bŵ��ˋ5�@�e���D��P�r�i�E3ݢ���-wڴ3��v�b�r�5~�9n�Q:� ���s��_6&��_	�)��+;�9��\Vx]L��;qi�PP5ィ}{�k�*�.gA��Ho�D8Y.��O��'*�����r��`鉍���'�M߹u��G�?�s��񱪬��\y�&�<��[,��0hj �V�6[p���j��X�-�&3ʚ���s�6��)��u�V�xCZ!4��U��H�Ԡ� � ,�ぢd�1��5Pٸ�A\�m�1��`:}4+f����hf�Dk&�=��B2������X�`>"�&K�3��l&`4'v2�;S( L�rF�X���|�H8[p���"�pnl�4�,�?^��#���|�tN�lk*#z,�1�J�e � ���p����d��~�[KP� @���]q�����/�{����r^;�Z��Έ�̠w9�lBnO�lK�@���vƙ�Ld)hj�
���p���Jzsy�9�V;�.�^j��(�+���	�g`*҄LU'^��r���r����#9����*UO>�5-�1)��Jk���$��s�D�5�ق����lC�� �/P�@EL�X��"v�f!�� ������6!�6�V���!CՔē3E�a���c�#�*6����"���iA��Pjt�M�1"yQ�R�����x|	|I�9p2�8�L����i�`
�����q������aoo7�C^`����b}q8?<ޟ@ ��d2.��$����` %0D	�� $b�Ò�kS�!:�����$b�H(c��##���a�P�@�;�qd?���� ��

	� 9�VX-��������~�ḽz�	�q�����������v��rs�t���q谻crH�����y7����������=C��'d	q�B�\�_��7O�+�ɑ�����2H������(
U�b�TG�X�%Z�)ӓ �2�����U� P �V�@�����33WV��5����+�)\)i�uT蛋U-������$N������J���@�iMs���B��H�l�m�N�_�^ h�b7�YM������Tzc*�!��	z�D�HT9�톀t��V�����
��+u�rmP�6�H��	OV��dt����b,)�)//ͯ�ͨJ��0�N����K��u�𕴭���*y�+��S��Ǌ�[Ү�q�W����n�w]Pw�ն��M�X��,�:�/��$q�0AkF�
���!5M�K�;� �Iz�
=�pw�mc�YY�D6��%Z$�Ijz����*��7�
��\�4W+�7HK�qU�*л誷��[�]-���ࠤ�_?;����-K�օ��R��r��\��t�Ԩn��0�k�H�챍��{k�M�񥩊\�:Ǩ����T:�L$�BU�P�(�$M��ŴIp�8�@D)Ex1�@ (��Q`L͛ǩ����O�|����s��bڒ8b�G[fQ�餩���@�A�G�p/ν����6��6��������q���#|���?�?�>�4��Ih����'��'Q�`�1�o�C�DP/E]c�]b���NPq'���#(7��w�Q$쏥��b6H_��]e�܌CčӘ5�DދFf�����qd��ꃰ��B?��>
"ާ?"��q��؀�0�����������r���COO�-�Mww�-7�{@n����u��뚻ທ�5o�+>��>�K�X4���+D�e,�"�x֏xڏpxK��C�Y�����0�m<�DH�)p�@\
ڠ�m�#7��-gU�;�T�IL8�j���u���A}��շJ
��/ȹP����dA֚�2�R.*5KrբL=#W�*T�F�Bn�fS�tS�D[Ӕ��Op����f���m�����p55�={���/�������9lvn���9c�#}�;u�7y��{�f��sġi� S��@_3�x�i���"hP�H��e�������;y��q�,���SM`��jƅ?�����O;.�nxg^cj��@��35̾"�@	����_"�/���H��O����,IeF\SQ�pk��sG?�{�����ϞY�����ik�˷�(�ZN�Y�&ː���8d2� x��d�߽h���V���S���?�������G�WG�|d�`gS.�����pmûޡ��\�[�,�� u�x�����Gcj�X���3lДAS�@:�$�k@�o�.6˗[�����z��Ȁ��p
b3�~|8��`�f���pƅ���s%��ό��9>���o]��O5+g��mڥ�B�j�A�ئ.��/6*�s��7�،�/����wg=0gW�����3�EР��f
���8�:S��A�~H�)�����my��y{�aq������͑�'f��>����GwN\?=�T�mʓg�V���̴kX��S��4/MM��h���dT��?h;��L͈cH`��*��b �.���hd^h蠬����������h$�������t�ds6������0{r���sY�����f��3���>�43����X&k4�5��D�Mw�X4_&�-M���wgA��O�B*5d�f�̩����XJ$`4�>�F��5�t��u�������/�ٓ���Wή����z�w�#o?A�������ԀM`��l��;��.�[l�X0T,(��zeېUgct���c��F뱁�ku�6���+�N�o���5��d�.i�M)������֔phj@��n�жT��ҿ@�L�5p �PS�\T�
�9	���hi�� 0���R��*�E�q������p�@�p�O�+�Bąè��*���q"B�a11t�Ŋ�����0Y\V, ��l�lNTD$�H��{��v���<<z��wK_?/ ����H@�lvj G�1�� ����0F���q9B>O��Q���H�#�
�z�߁	�
*5�z��pPӀ��VT�0n�	t�4H	���������q65β ��� C��y���`��<���Cˑӳ$��"r����4��\��7G�+�@A�45Ej\�_�% @�BSe�4���
�� �yq� ��>9r�N�ܝvj���b����S�GF��Ɗ{�F��z*me��|Ey�P�'_��:�\�x����Ss����`�L�e�Z�W*o��7e�6g� Mэ�QMiQ��Ծ��ph��� CCS5�����qa��AfU��³U����T5+�W�e�,����fVv$����G��Wm���eY�I���Y'����q��a�a��f���������璲묦ㄶqM���4�(l�8�\�T�E	b�U�"�����l15]�Oa^� ��iD��4�/�`p�V>�*�Z��ڨd�К"1��4�x�B��R4�VMe�����Y�k�V�Ԫ{ڴ���a��D�ȸz|*anѶ������������0��0�43f�7���N���u%�7Y;*��Y�&U�&!Sg��-�&6N���QH�($M�h	�@D)���q�h�7��
)P�Z�����̊h+�U~�Jl��<���:����y�x�������戇�%L�5��?榯��>�w�1	��Ԡg����է��#�GEܦӮE_��^��!�5�L͹���1�[�C����D��X{�øŊ�K�ǉ��5w@M�R�0h���ER�ݣ�!CYs�������5�������C��]�]���q�5�y�~Ňn�7ݽo��^�����5���^�}�e?�%�e�215�1ĳ�I��rO>@��ǯ�6H[��z4��F��P��a�uz�Zc��9&SǟI4\HK�hO���}���^]�VI�����g�rNdmۓS
�b��;S�K4-�l4�ξ��{��o25�>{����/�=����7�\81;;V�ך���8N���Y��~��i�
s`p�cj@b�i�'�	��bMV2Q�*�|��鰫��X҅�r�	���q�65?0����4��S�W�(��K{�%m���,62K�]X�_�oj)�w����<w���3��s3M��������L��$)-M�:S�K�c�Xh��ՙ��,y��Ad�<��>�����N��ىsp�y��q4/)f��\Lr�����;q)�g����;A%ŏa��7Uǚ����g�4�f9sM\��.�ɖZ�נ���X��B_3� �o�[�P���������4L:9�~j,��P�����ޤ�^�r�n�5n�Q
�k�[lS��ge��i�[hR,4���e�uҹZ�l2�rb;�	��A�}�V�����z`ή8C�����85��)��A��3=�5�ٖ#���:�t�c�g6No�\:��������<�s�����*K[~�]A�L��[�PS�f�v��6[P[R ��c�/�#K�op�������ݙ�$1K��L
�B�bff��g���)IJff������j��ow���+_F���̚���^[�����s/"�������1 ]��{�_>�<�gK�7���A5 �4�w55��l�V�؆��uK��$dv�uz`4O>�-�AK2���-TO���Ճ��A����OWf+�J'
4c��cY��l��,��L�X�l&W=�������ʍ+���
�|�a�P/Ԍ�)�rù�c������\��l�T�t"M<�&I�҄[����F m�N��%�૥�AѮ�-�\*;�Ul�r����9�5�vؽ�PЎ�n�g.Gԙ��ل���eK����΀F�Xg?i��+uc{�5�3�asQ���Mqk�Y�Jo���_9 �>���`���µ����ؑ���bMk��%KԜ)<��o�j(��L��5�]L�5@�3Gԅ��#������@�!�(� m[���$.�" ȓ�?�" �Ʋ�B�p�b���pf���k�p"$d##y�q�l�'��$�X$<�L�RIBYʢ�94�)�D��˕�x2�@.*D"�8��?P�ԩT �|&����}��]�w:;�pr�����e�H�]�}�|��� XO,����|�Q6x
�@��4 �D�� <���#`|� ��k��"8�	 ɹ!��!i0��b�cu*\��EXۀ" 6�R�h�� @ 4�3��60��y{z�Z���De�k`����������}�N�Ç|/#� ,�H���"#��L-
BLM�����Wh�)2�Z0��B�lAi�,_A��$@A%,VE��c(��h���5	��Df}2 2{c��(8Ԑ�9�)n�Q�W/u��+=;]uz���TՉ��##%��)�A�1��fN����2ښq�l�ó}7�����_�,;>^�ԓ1\�[m�,j)T5�* -y�-9��l��,YS��!Me�i�śe�kbY�jqL�l���S��+��Fråy1����ʜ���ܜ�}1�5ɕ��}�����V"��g�,~�Y����g)�ϓ���ߊ��~6��dL�����u2K�Rm6EDM�����^�e���I���gd�s��X�A��c �:��yn �ج B�����h�	|��@�	�D�"�dɪ����,Cx�%�42�41�&/��$��<��ި��1C=�c�a���������ɴ��̅Ŝ���CٳS��S���YS#Y�9�}�C�i]u	�E�e�a�a���4KJ�1.R��G1b�	A�T=3�����ʌ�2=�BO�B,3ʌ�R+e&��05{u�z�IKjUaL͒A�(XQq��>i���!K�������X�!_��0bj����O7�07|�ny����<"��i/DBhj�ʑ���K���"�M)�15�ؤS�9���s�_p/P� ���^�0���VzK%��/��]s 7��[�])��Lp_.| �?����D�B�}�5��$(k�����x�}���.�wK��� n�zn�x���D�����y�dn{z������捹⃹싹䋵�\��_�/�H����D�y"��v�4�q��q�L?La�����Ǹ��<ު�wX*:�/;�R���0.�E^�H���y�0�jaε��;�+��U߫��SYz˺Nͩ��CI��c!�1�~�
M̈́9t$<r,5y��x��~��y��m��}��c��c����	�t�������mS�ɓG_���jj�_:97?��ߒ;ڑ�]L�jo�j�T45�=�?�Ԡ�֠����R�v@Sc���A5����1�u �z���7���X��7��l3��;G�0(�J�-�dj�����T{+MݯLM}��&C[���̌�/|���=���k�/�<574�Y[S��h����A�=�$����������N�i�Z�o �y���Eod�x	ܻ���05�N���y��0|�@Y�W�f�k�򗊩���A%�[Q���WBMckj �-ƅf45p&�d-�x�f�|�-4/�����#�6�aG�c��į�&�N<������i��7�������`��4��Ax�i�V6v����a����=�M�6��A;n��r���/S,рd_�)�3�-��]M���*��d���g߸���/�~��G7VFd������x^c"�`�%�ߚ�kK�Y��iN�S�X�)̶TV{:�#�����o�mckj`��f�W�l65��4��]��45��l��5h���0^l�P	�(T�W�f�����l�D�|*�0��+P�igʂ�L�ՖC����,�+��EA�ڹL�|�r1K���=� XH�OṲ�!S����X��P��P��T4����QM�fr�s9��,�\�|&]:�.A#kƲ����
Ĉ�n��b����}�`jj`�v�����O��
Л�aX�@��@�� �о���N���l8T��<S��� �t��{��������PE�d�y�)r�-�hg�Zw������#�Ǻ2O��,>�W �G{��b��,=e��9�-j��f�[3E x�;2:s����Γ�䃫�ǰ�lP#��� �A�<d�j+�fCӤ��$���|4%������(N���g�j9�"���-¹q�ܘwև������x���|
AB'J�T)�-��|>�4�b�R"���R�B$��	�������q��{v����CG�N8���������������������zb�)oO?/���Ī��@�,���x,�B�3hl��0�'f2�$��&ĘX�5��P��S��[E�kx
�<�8(��@Иpr8!֏����v�`kjp;�y9���遢����)6��M�b=�Ā-1��0Efߢ`?Dӄ�@fK�#������(�ilȃXߘ�mˑt�wkd):J��k��Z�@)��h��ٽ����q���|��P�tG�Boᩅ�;�z��\?�rq���L��H�LkbO���4��(�%�j��|e[��5Wޜ-�a5P֠�TB�e\�f�u(D�ık�Yu	��m����Ț�QN��(!�$=.-5+$.+�����|�TXìv�lh�����!���W#��N=ɘ|�4x;��JX���c1M��nUt�$ Z���̉F}�^�ePdDyFA���of�YyzR����
6�%��5z/$����r��9:B��������+��Մ=5*�-����$�CRU�麰�И����������]���1#�1���cG{��`��l��\��t��D��D��L��t��x��H�d�`sFkUxQbTnTtz0���jB�qFQt 3Q�J����[MSa�CGc�4��1aJ��r3��L�T��:5�LT�~+��@T��QSӯ����+�!�pU�]�1f�I~��7L��'���|���~���n���>�p�kX<�����M�c�#���D�T�l���VsO¿#�ݒ����3\�i.�,�vQ̺,� ��y7�B��592ꊈu�ϸ"`^�n�8��\T�ܓpHSs_�De�C.�>�|�N�O%> ���ػx�}��35��AM"k<�Y�aj W��.{�]��������b��q����v�L?A��fq���k,�Q&�q4�њD�"���kʓ��uC�Qc������J���)+�QVp���~]����wk*�T��,-�P�{$-i**t�48��3/C�������艜�Ś�嶆����΅�.�l_�tO;P3��:fe�uj>�hc��Ûg.����h����.�f�?�P����j�إ�(���Լ!�z;@�v����1!K�Q��N��YL��cj�ԌoS3X4P��2t��۬��4d��fh��ei�5%Oo\���g�\yz�΃kח�'[��3�B�T�A�� Q�Φ�9�әe/kz�
Hp�Rx/�`��=p��[;c˖��g�Ԍ�x�#���+�5v�p�f��`L��*)ކ�:-�h�`@�2{@�_h3��V�15V_3Z�ߧ��Q���5����tFj�Xm_i�Xn_<:�<�`�ho��T�~��0Ӡ���!�9 �����lSc�D_�7��<�fKl����_*���Ye�dC���z�U]y�΂�}Ɋ���g�[.�;sh�֥�O�^��酧7�>��<ќ�Zd�
�Ճ!Y���~G� 2���.^���tf��Y��yP�b�-�����6�ŀxts��mj�����d��-�p4Ū�dr`��\y�l�f243��"d2S>��Z�X):Zb<Vl\/2�V�UKI��\�!��υ�N�i�ӵ�i�c)���G��+I�#��|��"�~$7p5K���Z�T,d!�e�ә��L�����y1���V�5�jƎ�Tޖ��Q���15�}��f(�[m4֛'�γ�4X�T��'%A����@g���@��TU���bSġ���IGړ��IKM�[SN����?ޛ=w j���_�V(;�-�f��s%��Y/�<�LiG��Aҕ�FMO���@E�+W�l`'k`wȣ�����D.�*8�,<�"iJH�L���	*�8�F^��*��(�B?G��#�Ǖ��A�xQ�|h_�&`�$����SpR6S�e�x9�����|�H�A *%�B"����:������=�k��������n7H�w�z�qx9xx;z�:{���`\�(O/������\�����yb`dp>x�L"P�,>�ɣ��D��W�)ܪ	�7�5�.���Ʋ2֖p�[��c]��"4F/���Ԁ//����2��A�A�~r۹����*�q�ѳ��A�|�0�Z�'��q&L�ů$S�)
�@P��8JSMTF�P`��X*�V�4�p uI���tP2͙��B��RMoi@oyPO����V�F�"�����T\?�tf�����/�������w�_���q���s���.-՞��<2T0ז:X�Y�o+
h�S̑7�*����� �i�Q���6eH ��4�.dS���P����$.x37%	j���b��ܼ`v���n�f�Krb�qsTtjaE�x�б��Yc�|hש��{�+-g̝��羅����>x5��h\�J��qCF��P[C�N�f�2����&Q��_`��s
C8�j����
޺�:��s��%�c��FR����ç��	j��_l !�g���-,s�%I	�ɏL���i/��F����i��oK��m:��ݑ15�7=�68��V�0W���we�zq�bf�l�'��>��X�d�HNJ�$��bM�(-#>���N�32��,##��@5M��Z�� �6��F|�	�-3����r���4#T��lj���(�m*R��>c���U5wIΜR���qv��7@��b����~���.�>�'1~W��[D�="��x�{��?!���i�y�"�#��TM�}�ஔK».�\2��g�4㜘yN@?/d\���ȸ����٠�%�2�q��!k^E���Iـ�b�U�<�3���VYs�b55D�]�����ْ�~ސ�^�}<׼=nxy��p�� 2�<<nzz���\�����ho��^��<} �=�O�`Napgp��$�9
��~��<Ag��p׹�5��L(Z�J�+����e�xE+_7�
7�3��/$���ϸ_^x���NE񭊢;{�5�ذ���W�O�&�G�����}*ՐJ3hZ0�̙�G-�#���EyK�-v6.��ۙ8�	��Ԍv��t�lS���~���O߹w���������΢����bj��ؚ��O��w55 o�i�ԧ7�Ԡ4h�jjТ]�����Լ���Cn;��S3R��ڂmLͶ15C{�Uƞ
d�Sg���Dה������Ȉ�-}q��>~~�ҥgwｸ����\SyyR�!N�L2ʓt¤ ��M���O�i�V���`kj����@~�ho���� 4c�J������Ѡ�o�.�}����_*�7�J���N;Ӏ�T�XQ��P3��+N7ۤ�s�@q|�b���V�(��lC `�Q����lY8`Zh�,�o4O����Nlh�TS�dC�D�n�6p<�: �Ѽ�4��� ����ҏ��Vl>���f�^�XL\eк�0`�T;X�_�]d�N�쏿��u�H���{�W�xz��g��_^~tqv�`VK�!+ט$j��5'�Z���t dZS��I�˵�����t�s`��A2"����`�` ���g�8�i3�+n������lh�ʹ��\��u��<��b�J��Hw4?h-/�D��T�� G&+�l��r��bF��Չ��ɱ`�!#g9�9*��a'�I%a�?�&��h��
?D[��M�?��MU�%JfS�s����l�l:S6�%�Ȓ"gI�`�J�5�)��z����I���
���@�6X�-A,�s���bj��d3��}��7���#��S >�F�@�;���ؚx�~c�b�`����������V���%nM9Ԓ|�=m�3�pk�|c��>CU@g�K��9G�ȓv�˺���%�rY��lyO��7Wޝ*_���Byo���\�*4� k`�m=,��n��9�ʵ�J�$s���
�`��9Uz0EҜ"kMS4%��F���d#��Q����=TO'��+�ǃ����aX���0|�/��ǧ�y4
�N0h"C�F�CAw yp�A��<<������3{�v������c��s�������*k0?O�]� 2P��z��	~D�L��E"�?����3N�n;>����?x����)����k�#h�l��������jݫ�ۺN��u�'w7o��6hRh	 ��$P���VNH����+��0�3�5p�'��{\w|�}���q����<�$?���(�Q�t�r#��K�1�!��)�!X5Mi��T�P���(����D&�.��i��i�H�7�r��x͙��\�F���*���P�]n�l�9<�sf���у�/~�`�W~�p���ϯM<>?tvvߙ���c%��C5��e��� ���kZrU���Դ����(�(�id"S�`
hΖ�"8Z�&�J��& Q6�&a,ko�<�Y�ȵ�r������`E�Yo2�G��T��ͤ6�G\��>�1�(j覥�bD�դ�ۙ#wr�o��Hh;�x`.��[W��4$��u�A�o��A^0//���-00
4+��I��X�!1�|#&ǈ�3����"��L)0����!- �����i	��%�D6��A�1R��K.K�m)��N���U?М=?7����ߕ96�=2��ݕ���||������#u�sUS�%�M��AQ�qA�q��pU���OIU3r��#�H�5��4$z�@�4P�T����j#Pe�U�q�L�����o�j�ԙ6 yPYm CSs0�Ү&0��N͊��(c��f���a�i�Q2f�5��<����y��N"�!SR���T$��HzJ�<e��sXw�l(kI����=	s[ʿ.�\��g���"�sb��e)熿��JtK!�!���hj��7���b�	{Wb�4b2J�z(b=��(0���x�B�05,jd���e�h�z��{��vw���mw����7<<�{x^��\�����s��笇�w���ǽ|��0'q�3d�*��q��Zg���k<�1�pM"^�ˎ+�OhT��� Ū^u4Dw*�r:6p)-�VA����;���
o���[�~߽��7J��d�MJ\
�v)���~%bj���CȬ9|�2��PU��^7��8��:��e�l_�Lo�d�TLM��<�ռEL͗����ӗ/޺}y�̱��ڱ�ⅱ��bj$H>ԟdkjްK�;�(�������شr�m޶�&G��物��Ѡ�oɛ5�?lj�y�';A��15��U�� �s�]i�,7���r������"��=�}�W�}��ʕϞ<���/��JKc�Z�e�^���40�35[�(ܚ��ʶ�ǅ��W�����":�ن�%���+U��U3v�~�6�`���_��`L��fPI�6L�i5s����nT! �vk��v�A:ۤ�i����4�f�m�K�.��7����K̋M���Q�8'N�&u�����~�Tm `�&0���ۤN�玾��K�6��l�m3x-�� ?r4;A�b�5�bkgl��������N��f�H�W�Wj�J��$�<�{�p���{�W?r雗�n���ybd�!�@�.'f��lhj:҄]b �@S7x���-������� |�@�2�/�-�_; �Y� `~G�ƛ���%;��-�f@;Y��L�X�D�
0Y��.�̔j��L�ȧ�s��|�d�l2Er4Uu,^y8Z�*�7qft�)uFE9��������V��_�]��:���ޝ��������M���M��S��ߔ��7��M���w��������t�{��1cr���<Ș7�&�٣1�x�d�p*U'@�e�G3�i��U*�A���my'`��T^W
 2H}Ə�7��~mƮ
\�4��w�3����ol��n�Rd+Y����i ���tȻ�%��)�5#��*�H�~r�e�.b�>r�1z�!j�:��(��T�Y"o/���[�Dm��9��t�w�b#�'[ޕ���S���ogj@j>�-!h%�������X�>�7�~jJ��IZ��-i��i�PL���1U�>FCv�:�=v�=���ɾ4�7���ӈBAH��>���g��
�kU6MȤd<��������ø��������n������w��?pt����}�z�q�����8yAM����4x_�"
 2�נG�J,	.7Ro�����λv:��� �{� e͎��C���]N  P����qd@Ԁzx6���R��I��� EP�������j����V��"n���&�v�o�ar��%��� ~A �8�Z��0�h�,[�-ÖD�E���!~e��(��XJm"�>�Ր�����8*��(���T 4 ����$&�9S 9���d	�@0��/�t�;�4]%���ᚰ��Ƀ�˽��rz�&Z����V
���+=4\�ܛ=ݚ<T�Ua<X�i�W�����O�Җ�FLM��5[ږ�l��HX�iPSӒ�  �����N@�%�k�9��pn�kc�{�X��VE��4J��O5	�����!a�1���)�i�3	�#����>�Yy�>�4{�������w����]J�8��4�ߤ�RFX�!�FSj�6[�o��&~������#���,2�m�"�`p�����o����C���"��L,2��'#��HʹВ,�H#1X�7�FEk��C�����)��[J{k2ƻ2�ҧ3����G3FRz��{:�'oߚ�y���ك����sZk��2-)a����U�E�&r2ع��� V���k$�Tj����UzJ���׀�J�` �Wj�US*���*�^3M�~=�QO��f0�9k.	���e%�Ǧ3D�e�ǩ�Q����Ӥ�3bjp�k�צ�1��,RC"?�Q�0鷸LT�<�rO¿/ޕo��We�K�91�~J�D֜�SOs)��57���
�몘}M�p]Ⱦ!� �Yw$w%�{R6\�摘�DľǢ<`Rа��䍰�~�[r������;ಧ�%׫�7]]n� ��uW�kn�W��׼|�z�\��>��y��봛�)W��nk^>�����p'I�S4�)&��s��9��p�JDG�u���Vu<P���1iW̚á����g�#ϦD]LO���v�4�vY���B�����Ms.+�Bjʑ���S"n��z��C*͘:`B4��1�[BF���Oݍs=MS��:5���L��O���t[S���g�~��7��|���k����O���NToSsd ��վ���Ů�Έ�ajPG5ܢ�{?��L͟-��j�I+�A�S������ �E7F>����J3R�o��o65C{�����rCO���*��2���ܐg.I�d�7��=�u��_|�����?���~�����%�1:e\�<3X��&0���7��]�۬?�]����ͦ��"ȣ��-���6���/SM��!����G��|#�j�;�����f�N;ۨ~J�D�@G �up�n�j5��������Z�����&�|c ���������:�B�a��e�y�&p���q4����������>`�& 2�_}�����:�� Ep��ن��5[��r��k@�%Mc]T�7_՝���J���'�Z�x���B��ˇ?r闟ܺ~b�ʑ���I2rt80$k�堦�;S@M	����RY�����T�5	���d��h6�v@��*���h�������@�I`/T�@}���y�-�K 
�р�W��P�L�g�5����b�R�v%_���^�V.��gCa�AqH���v�\��u��U��?��?+��p�/�K���ry��}Ǡێ~���v��a��i��i�{O��������:`{����Z�?<��A;vw?�m��5����hS!��H�\�p>A<�(�NO�J�ӥc�ґ񠍑��L)«��l�,�t>`ê p�S� �*[S��v�n���:�9པ�PD*���Lg*w3�	n	|����A�N�15�AS��cS#n��f�[2y��lQG.�nz�}E�#0R�(��j�����j�@I@g��� q:$]���BEo�? �5և
 ��|���v����A�P� �^�������頲�=<#�I���Z�D��|�����-Cё�lN���
2u�%����C��Itۅw�E�v�㼸��I��B�C�c�|���!r�$V#d�adjj8�����k�����vvܱ����λ]v;9�t ������+���������������������F�؆� ��k���;Fa��� �xa\�=��r������R���];�!��� ���j@
j�\����<�UPm׮��0�Kp��m�!8	�<��w�Kpw�����	l���g}�U���O_���Z�����q�v���oՐ�yՆ����<8b,$�tuHd�;��#�q���Q���j_ ���2P��Mxc̋:��{���>G����*4HZ:��7�xu�J�1�T^ƌ.�3?� 	���P��/��.�Ʋ��
�C��4R6�r�c��0�~b��=�Y��8�o�	k��'��%R�,<s��hJ+ug�l��av��T�$+T7�}��/ӗ��[��=������y��H�h���T2^0�`�J�ΪoNL���;����u^q�&w�?�ގ�^�����Rt�;��㝖g���������/����1�٢o��a�����NǠd�Ǻ1_�\�Va.�τ�}�(sx��������Y�u9�J�ӜZ���@ŻF٫͖��։t�Nw��;疍��~��O��Jr%��нGx��j��ĊB����>�K[�0���`��R�Oھ]*��O�#�Dc;��3�>:��Q��a���~A{���'�ֹ���O�,�锹��ߋ�8�l_n1zXW����y԰�4�q�}W;j@��N�L%�g�E���\@)2:>���(�{k�f��ȸ�q'V���NӠ/E执��ͭ��u/FJ+lH��+������� ��ͥ;��cJ|u�5�"#�ѵ��*]�������Eo� �fʭg��u��:�����Rd8�)��S�P�Rj7���>�<k��S��N�H�PF�e����a�󤲮u������8�39�����ş4��r��sX���(&�yk��Tv��\Z�2��[�q�1b��B��xJV=��Hk_�#�X��r��:{��o;ϒl}Cn3rsk�>r� r���*HĔܓxL�~�`4Z[4Z�������6D^�6}8�<�C���~���;,�J@�Aa�w�p{Iu
�ڴQ�����?��n���n{Ič�n�����3�L'm���-=�'!�;��yPr��`�;u�o��y57s�z�g/�%�P:�yZ�猇i����Ϭ�����U�!{J���wz�0�Vlp�#�qX�ľ��&�w���?�|���;������h���]jf	=w��\3]��Xؖx�29�uu6=2E[{�ma�Z&<	���4������JK�����/������@��M4�����>�q_� MVe�g$�}�u����8��\�!��.�%+�4�bk��JP|6E�jDtEB��v�e��1P%�+��lc����=`	�#��I��c�,W�?�,W�G��&���ݭ�V.*Z��(���r)�IE���t.Џ��T�����"G�˿E��u�VhGG�� ��e��N�l��}K�M��ͨ����?+:{�NNwä��������
��:����%v�("��t ��;>�xl��6]N��\����oh=e@8����zSZdy�(���5����4���ӚU��Ɉ���$r�I�J�Ĉ��Z�I�V]V�7Fr���%�W�C��F��((�L��_�?���3�P����S�~n�)�,���W��"�KH�m@pг 8
Y���?��w��?Eil�E�,L�KĶ&���mы6 ���SI'�O�'�%x�`<���:�1�1�9��R��I���+�GG������XC*�d���#�9r��X�k����%�JD����<�z�(#[X��pw-i�${]��u���q���w������%�O��4_�%SK�TY��J���2��
��2�jŽ�9������[R&�N�)x�q��¦�K���`��n+�`����oƵ�BG�$���C�T���:�Z�n"$�iH�CT�G�,vB�FlB�+�lZW8�r�Q3����JS�����~�)��q��rn���J�i�c>+������Y�6n��P��j�n�Y�<�ܶ�v�ش�Xr�Y���S�����#��2�C�=ڤ5�����1��M�g�����َ�93�7�G���A͙+��H��<<��l��J��#�\�6�K��2���WVY�LV2\���o3�|�@g~�Z�Kon/���@�IGk:�g-���e4�<��(/r���<^����S��Zj����NV��=*/���Fy�R�Db�x��A���c�-�>��ʐ/oO�)�w�7����P��G����OН3'�)$x���۲���O&�K+��ZH�5�������&����XL_PEm�ٴу�^���Ŵ��,`�PL�L?͆H��(������X��؇ٔ���D�g8�DX�i��� ����զQ�r��S�Ժ ��*�e�S(�$������'��}~0[_u?w�����<m��S�9.��9-~)Y�p.!~�~�t%2������ ¶�͝�tu�@>������,�n�����H�f��=:ޟa���e?`srq�i���[ƛk>qZ�Ł'����t]E�՘;a����iHF&A*�CQ�)o������ɴiy1+v�����T��.(��_��C �`�K�е�;��4Fd���RWd2�n�܎��1��%Ht�ֲ߇�2�|L�b��5g!���P8 bY� H����kP����!�',:w�?|��Ocn@����< S��}��E�W���Ǽ�jЊ�	6��Q��jי/h�{�0����V)�4��S�֫���I뎰�Ii����EÝ�e�MD��Yv�h��$]���~E�N9�A�Wi�*�ݓ��D�8�:���H)E������5��I��|n?�y��}=�P%�����z�
YtFR�ug-־������h/HM��ӛ	������	�~g��RM�O��G�k#k���$ņZ�$��(O[A�H �І�0�Q�7�]�nF�c�-z�@�6��^<�w_t��hd=ş��X�ƕ=$�kK��V�ΒM��Xm,��e��6��N����@�S\��?��x����������ߑAZ.��=���$����^�.��h8�ڊ0]QN?"�n�X�1k����������V��c���NI���/�Mp�$�a�?�̲�~�I���}�ra�1��0�7�[N�2Cp��y�icН�U�pR����DC\Ho��.�rn��Ԩ��4��PC,f���2��\%|7��t\�P`��ܲY���ah��Į�L$3~-5(x.A��=�����AȎ)vDrl�_���z���y��27�ε�>�
�;�ȴ����J<s��L��=���s�QlVe\�ݪ��,?�ӭY��so��N��,p$���SV�S��M6�d�����TP���̏\�P4��r�fy8��o;��=�M�yL�Ueƶye:ދl�7�uSP�Ӻ�s�%�NZ���Ey�!TX��Kv��|�G6E��q~�H��(���b����>f�����`�pj��(տ��]h{�uK���,�~!;"bt��.D[�!���3��Q��O���mXf�Z����TüZâ�[��]�?����ٷX��]o��e�r����߅���KFϏ������E=�0i��{Q�P�+>��[:��K|�8/�\�`������x�� b�@��n0�����=9jp�o|��F�P�s�٣��x^؝'�Iy@�g׽(�IXv���ޙ�����!O���\?D�[5�5��0�| �4����z<������X��a�HZz�yf[�_��(���$�����a��tV�A��o5�oaу�ILb݌G׀ ��̎m��
����Q$#a ����*1�ݸ����ń���Կ��U�'C	R�,�� �T�3\	|��Q�>���\ � �xY6^V����HKVV-b�W}���B-1_6b��^�<�+�@�n:r
���J���i���e\O�%t1���^�oW�j ��\���G��f��q���l@�v�bYUL��(t�E�s�#މ'���y�r����nz�=�D�\�{�hR�	��X�鲖���;xTe�ت���m@�ш|O�x`I&F�R��@�1�]�M5�
��D�D @	K�?(�uYe$���v�}��$���w��� �vܧ�#+��O-�D���r�e0%b<�%#�|@�H>,���͈�������/|�75�2���*��y~�����[d�!vWX�&��k���?��~X�����z�ע���HMz哓�k�q���%������,{)��JBJ��Z�Qt'"$m}��^B�"M,q�Pm�2����^�C�	U�ñ���#:x{Q�3�t#��6�Ɯ�tʩ�EJ�<{�zu/���F	�-��ڹ�:lO^x�4�|B���_?Bf3�si�W�1��M&F��%�ˀ<�K`�ژ�0$л�+��_�8�1��yI��M�0m2	P��� l�ں.ޭ�p4�)Q��N�6��#�L|T������d��\�t�C-�bI@=��8�e�ͦ���}>��vDa��f��du��(dB	}�9� \"܄�%����j�<6d4�}Ӿ~�t����ₓ���c�+z�=����i���ϝ7�I�^��Nv��O����#+.�����\��wP=\�y
�t�e�����@���l
މ5�[�=��v�z�쒋���T�8�D؋�ϒl֍.�W�a�Q�Rd�eS��� A�R�����ڎYTes� Hg~E�	�*|.7��V�;y.,�ф�6>���x�(����̚9�؍N��� �/2�OY��r�͢�3��+A�a��ƻ��
�Jʩ��1Ȉ�
�,�5U���?���4$r/����%���fL"��ŵqP `*q�J�24xG�\���џ����B��?�L2i�x����73N��mn.�dRx�>�`��%{���U�B�zzn�ߥ��͍��;Q�B��R���hA�s��g�\z֖�����jѿG�9�w�I_�����F�z~3�����֨~��K ��䷐��hG?�&���M����`�B/ ��`���#�I �����A(e3=@V�yU�b��t��.{\y�*Mບ��o��	�#�|~�z�)��{����%�{�ˡ�q��uk�R��r��)6�ow��IAmA	�\%SP+"��^yf�Âw��]�C�	�O	� �|E'���:y�`�t���D)���[�)��BO�RK	!:�)�0�qe�.zG������t��?�.1;�#����N�<1+Nq3�l�������
y�}�I;Hp�/&ϴ�^Dk�Zw�\�A�N�⌦֐8n�r�5��#���י8�����ۿq��<Q|'U�N�r\!��Ţ�\�c���7��G�b{p�φW�|�Xxq� �K�,��v��O[���U'�(�7tD���b�@t���/ަU-O��wB�N#�ꟙ���Ϭ;����Լ�)�o�v���r�7'9��\{�q�p���+4P���v�&�3�������UJ�2�� ̡>�ynY ��FQFR{�_�X!�#9�,�h�6xڛ�V�@: �����҄mR�{�/���L�y��v�	�_��'�'�o~P��hn6��ĀVgmǒ�
J��'|Z�/.{�}�u�|�I���Gn⨦48�m�j��k�ͧa�CS�x�g	��Ҟ�t�_���QsK� ���'������p\��He��o{:� ��
k���*�$I��5V'�Ҫ���?n�O�����1���ߩBX�UUM��{���D�~7���;�d�V�b�����u���J�CN�&:���^�����<��M��TL����H��9r1k���S�n��R'�q:���'#�����`e$R��Y;�e�{]W+4�v|�?H���uHڦ����r*�y��2���A���`�W������RoS���8�� 𣡊[��B��=�C������8M�} ���Y�O�,D�H$T��!��>J�$dQo8;��!�Kf� ��2�n�#�(�~=}������	`��xj���ָK��҅�����/S5�a1���*�����S��f���q���z�56v�AN����@���y����R
�t�ӏ1��$���㓼��ZL��}�!�{�9�[�P��M,��h��4D̿��!���[b(���I�4U���U�;��7IN��n(��ch���Zń��9R����}�**Б�1��Ζ8E��b����`p�lݰ�U%ߓYӛu�_0�jA��[9��{�#t�c����V!lyלlԉ��.��!�!���5��A鮋���YH�9v�������^/�)Z��];5�I�b�h���_��P�S��xo�>�NK�-J�w��X	E
'��(����VP�:%fYL"YlJU�b�v��S~��/�|nY���
iq#Hu���r>H%�Y�)��j;7�uOZz��QΡP>_4ǵ�Z.�`�"���Ѵ��K ,�E�Xð��#��������#m�i�8�.�ҹH��L_�O�(�AdK����~K�>q0ݕ&B�bn��N�I�]���a�=��lmcĈaTVۏ�����"B:}(�_��	�q���a�m��\{�&����GE�$%��P�>�e�D��r�m�®)ԉ��M����?���S1:0Zs�3�#�ǉb��d���>Q��:�KItO��6��Kf�)�:_� ��kp�����0va�����Ʊ�&�n�8�
0���&��}��/"dy��{��n&�d�6�����,�y[�;�"�2s�ay��O���o���>�5��x�GJ�~%}��r�Pͱވ�F��24�Bzi�V'qֽ�!vx��f6Zޑ��d
���GI˥�Z7^�Y�.-�(7ȣ�qd�"��G�8h����Q�Զ�ڳ��p��S��x���'�������f�@iE 6P7>H��HBo6{ǟ�H+�?�o�T<����,�O�h=�ʪh0Q�\F�����Rsy �N�/��T`�r��|�=�x��qp��_�"ίOi��� ��R��V�A����M����T-�lB<ȁ�������6� .9lnzqi�I����j *j�d*%�V�J�cV��9
(f���jl���e��*02OzV��ߣ�ׇ��/ST����^�����D�w0�&l�:��ơ2�(*�����W%F�!������+n\�k�b+Ć
�DPp8[`?[�GU�V�|Àĝ3�GM�{jcQ��N�����\��dO��a����8�C��LYޱ#ͣ��s��5�(�H82n�yG]�i����Ǽ���Qϙ�I�s+\8F��N��dq�ߒA���(��;�_a�!���8hg�8��u��C��(�|B�:{�Q�����F��;�ѷ��T���<��&�sk�x�u(�m��䄏����ߺ�z�韌��3o]�2��E���{V1'CZOv��I���#��eի��(J��℅�]�W�`a�$���S��ճ2��H��aN���}yY��$���8H�å��tw)��F�hfN۩� ��]�{���L�"�=����Q嚊���:{LE�{�k�#��J�s��d1���C�(�����ب��3�{��t�۔9�B?^;��ΘLŕ=���u�;���m�8����iV�p5��V_0�߿Ҹ���OWX��{���"���E���B�+�|['2�����Lmj3�9�>\v�Yx�ܴ�6�0{0��oS�����E��� 9�Ձ��\��y̌�^Q�es{�����v��0�;�C;9W=��4����-�ad�`k-(;Z�(�87�p��5�1���oLR�+â{ɢS��QXT|h�e��R����/�F����9�z��x��_�G���`@�7�0ļ�C(��$= ���DZЯjO�'�<���K00��W�1}����?􋖐C�ֻ��<�f|,F*�E���+)A�W �����<�s����W߾���s%����K �Uo��@�F�1%�x����ZVʛ��&�~ݍ�5wR]�#2��:oR�E�n�)�$]�����A���`0�������bڏ���q��kN׻K��/�vI�X�>��W�t8�]���Mh�q�d�����n��1Z�`$�O��#�}�
b^bK�g˕�j���㫣�����^`|'aN��-&a��He�N�hF�SB/��ֵ�?�%�:'<i�}�������u�,ߞ/��xR��9cQ+-yג��l���y�Eͱ�_'8�e�ɒ|�)�洽��,�F1ہ���q~)S-��&�����b����m��xS����5�Cڔ#[�ny�u���ƕW���&�^v
��"#����0�c��ro6�~�,�shhJy$(P.��M�bЍ����J5���L\�;���R�f UK�)����lƭ��OA���鎡�3�#���$�%�'oO�O�ݞ)�c����<ނ�>d��-�;�)�M�'ψ����
'�
��Mff5�p�w���z�C��+�E~n�i�r���^x0�0��ͨ˔c,hV�342�ޭI��՜f��s�yb�Q�
�qu�[���W � )>=>�2D�
P������k{t$�fG���r�*ŏ�x���..��Bf�d3�ήܗZ��a�e�%Dm<<�[����<>&�ĉ��$�Q���T�N��K�����pT;-�D�p����j�U䀦,�L�w�W[X���MC_��� vk�Aw>�d݊ݶYY�����_�� ��>T�^i�mp�m�p��g���j�V����SF>���[��)l����t�t��Rv�7�0�F��}���s_���>�):�+1�_�Z�w���Ѕ�q������Yw�/��]8���G?+l�]�nb��N��P�M���G`��	B��� 2��r���U��>c���m�)����%��˩���K# �OU��`�@�Е�����F{Y�\�lHڰ����j�����4��8W(��ù�
�*���4\e�b����]�s]���g�M��9`]�^{��v�!+D�w؃{G��?%������)@�S	�))K�WH��j��-�������F[���V�!5vK�Y)�X�V�䐨��l�k����9A-��߂F"�+"Ob#6H9���ª�����}�ٺ��{�VR�P�FA��w�A<�%�ŀ-&�omQa��첂�?��r�y�*+�	c�h��K�r�u�*�o�~�;�)U���&��<Њ�����T����w�c7���p�\|V!g�*W�q�^�ŉS��'���Ҡk��$I�P����3G��Z�n9gG"�Y���Y���m������3$��K�ɜ�Z@�3�Q�#�L��/�8��8 �q��˓6q����Lk/'��	!�G��r�&rS*���G9����r]� 1J����`�=�=b{F}��٠3�������J��d����,�}gv�o����O�Y���[g�s^S?f�ʰ_�q�K 9x紺�n��z[�9�	�m4�k�Q_���ǜ��E�+�Iދ���gt��0��L+�L��/3+.�B�XO�4�$91�?�=��B����Ջ+�T��WگP���s���	���`���o����h8��*��M4�M��M���M�U��=N�pt��\lM�X��L�,���czX��YM`Y�cYWcX�a[I@��rn"�$=�*���6��H�ܥe�7�����l��W<f��+����Y�?C+n�-U?F4��n�m��6�\���)�X�a��V�:ǔ��0��۳��w	���Z��4�ᓟq��\��$��	+*���Z�x1H�2��M�������5+}�Y� q>)��ò�I�.���,�'���>�ɛ�Ž:�����hQV����������v�B�$@3	$�::���/�f��̣7�,�T�-~e�1�^� � �Z`4���,�6T��N-bNѱ�6e_��R9^��Av���k�e��	�USn�E�\�=��:�Ѻ�D��j��A�������zN��!5tjn^�j%�Ȉ�
#��?\3���8�OdW��y��S���;�H��%Qw?�/]NYBO��5����C8=E�>.ې��<YD8�N�Wu�S�tfVd���dOb	��x���w2�=�j�2wNa�d�v��	�dn�M*�YV@�Ip�ۓ=d�[�~/�e�g��ݧ\��H��4�G(	�T�x�__��R��|q��޽*�?u�FO�jY~��p�Xޚ�c��Te���BW�k�ȗ��7"�\���Z�M�ꙺ�D��nO�ɥ�--��c8���	�Wj �5R���+N�<^,�$�YT(��i
;3�Mz���Hm,.fl�*{D���]����~��a��&bI�A|`��55@�G��'��D^��[(��H&+�W���-V�8�X�c�}���,R��M.���y��L�كjBR�E{6�����H�	q�ИV�{�~��e����~�H�vf�>�Wj��xY�K)����8>�s�zl��5�5��Vg�k�r��$��b�#j.�+E�����*��7|ka&B���;��%�@�=$V�Q-<0��'u�4�W�4��Ni.X)��E����Y��b�:���~ݣ�����^�Z����]�gs�yh�թ��es��/��ϐ�#��=��S���q	NV�~���u��!4�n�	�#0ޯׯ��U�?7��w�;��?6�G*�[mu��Y6װ$"{���s��k϶Z�Ee�C���F;��\��W�.(FD���� ���$?�44�l�oOTE܂9s���L�0&EkO�y��]�9��;>�J�e��jM
�a�0i�l���GTU��~\Nf�����x�]!�&m���(��2%�c=�s1-�E������3{��q���hYy���$�M6SzK��'M�-KKC�qv!�7�*jOk�����|&-�P�Av+��QSS�K 5s���G��MV&;	�d�#ide�dTc�T�D\�EH"^�ÅD�f��0r4)�ު��a�m.���h���j������O����a�����ceyS,f߼vQ�|Co�D�0?djr��zQ���4��Z�Y��l�}E�\{T�$H����9)a����m��T5�8��ɴ���r�%*k;���1<��f���k���y�s��������w��k��G��I�#u�}�Ŀ�	��Q�(1-
�����K�Q=��6��4g���kIR����!҂�4��(�y�D~Y#�p��3<���ՕY?�GIM���Gƻd������o;8+x 6 ���r�?�v]I]h��o�����O��l&R�)b��?��lR`z��Hߵ�^uH_��^�Fܶ^6G:uE߶�߶�\���E];��m��Y�g1*f-=𨌃���s<UG����R���-��`�A���O���n;lk���G�z��:Ӳ���i5�YA�VF������dL�5!ř��TIn;�b7���Kv0�ҫ�g?D�s-���ߐ���/C��f��������pV%kV媰O���J����i���u����|����a������n�_.+��&����G
wun��kχo�T�ɪXV���	LV�#�W��zD�ݓt������ot[��2P�L��'u	d����ܗ�^G�a�Vⷄ�ϑ��?a������3�L�����m]�n�g�Z�O�d��`��X�}�5��z�٪K�*����i����#*��&bpM)�2ڍ��fGh�!�3n.�!3��b�A!�d*{�*.��0�#)�����ܐ2gWF�����?��^��W��# ��<:�36�v���o���a�	մ[�T<x��_9侸�[�����g 9� �k� ل!uH���n�wK8uF*�GJ�p��+č!�V/�8 <&US�%���-���?��1��q��_G�������v{�Eu��>��S|���7/OC�NF���f��E�.ҭ�S�;����&�霙<Opd���^2���a����U�,���V��g}Г��`�~|m#s����Z���=�~�s�>o�3� ri6ԩUk������]���R|'��P��W���Z�e�R�5� �!T��!{�J�dE�Ѹ�%�g�tS�?ι���s�%��Y��9�Ë5ϑ��f|�=?Mw��#���ҥ���O⠖p�Ct�QM�m�/q���|K5Dt�)��q��ؼ?ڠ{���U^5�a6��v�H��TD��˼v~!!qPU0��K�G�s�2x�.u�_�H�m���A�f�5��v �k��sY%�BUϾ�Cv�>OJ���ᰇ��y�A���wx+� (9@d��E�08�HE��t_z-����I�j@�j���J�p��X��L=Ⱦ�K�:A��A�� �t�V�ͼ�ǔ��{n�+�
R�>|0��\�2�
�A��5�9�'��K��:p�h�մɩ����
<����[��t�c��2c�WC'��Qq`��u������O29�s��������r@�ߊ���W��B�w@�.0a�o�<�Q�O�P��a��F���J��\���>�8����X� �P�k0��Gz��e2gc�ݯ�4�,��|��_#��v���n�n7<�<�F�ɼ8��]%N[�:��A:��y:�qZ�:h%�iD�.���pÞ��_pb��%���h���dD�aH��K���V��������i��QڷD����j^�>����*o1$s��0�ͬƦ�\XV���5��P�4��<��Lo�]{6W�v�!� �{����p��A�UY�h`t��5V
�[m:W���	H_$t#�$I�+P��I�a�s�e��S�,%�QJ�0�lC��K8�uԃ��)X�!I��sc��O�ߩBG�v�[�zf3�KpW�f�����g�T�"zR/���h��kCp�XQ�R��F�f8?,�G�"m��C�O���b�$L����BEy�ȈK#�U�+��:}c�u��ŝ> *�4��������GUM��𥉉�Y
��!�k��w^N�_���69�{�r�+�n��V|�<-;r�,$3�L�g)�T�==P�S�D��ﺒ�g�gֆS3葔���jG�E>��H%\�;A�r ���>�4�u���;�CY1҅ؒ|�RI�3گHa$ILo*��� ڱp���w���+�$�3�-���I�+W�k��C��U�ԝ!��	G���ߩW#_��Z.r��K�1�{�����sm��f.����$����暌HX+7�n� =�d�'
��f(QH�o���L��(����""��*��k�Vt���.��`a\���<�6��9~�#g�%�_ԶK�r��m��m�̝�����U�x�F���S}U3���{����ǁr	j���]%�k�Qg,�ط��O���}������_�����N�n
Hյ���6�"�2��lgp��n���b*��3����B9@?�ѿ��9���ģև�U��w���-���&J
�,8R���O����NEW��?sX6ZD�æLĞ����/��q�d��8�2~�'�ndq������R��^�6B�?�1��XRuq�-��~d�/�ꛕkn���`�@*v�_�a�HpcS_ճ���}S��CB{�n vF�铗[)!����wr��3!�y� ����mт;��d"�콢}�䗲q(��z�
$&R�@D�C�W�l�ҡ�\d,Y�Uh1����Q!��en忦,ئv�nbT��ܲZr�8�a��ʲ@��\�2_)�ls�ni�یڦn��$���M��S����o=ש��AYAb!І[��f`JT��IR�a���)����G��Z%ta�6�c���E���8ؿ�}g�\j�2���r,Q��w'u|�T�']%_�h'����Q�l%�4!\M;�W���<9g��������kϦ��P
I����#�
]�$dn}K�?`8�����~7���Aa�P�������d k�?��\���J�6'[����fimο���Լ�U���n�����v�u�}y�ޝ�f�=:(uh�`Q�9��"�;!���*�c@X��l6���a�EV$�L'
b#�=�2�M�\,��1��G,�-�֓5�k��Q��^�H��G��QoW�LP�C�w������[��}ڬ�P��"�{-�	���^�P��G
�k���к}P��4S;3�����a˦���+a�0��F�Q־; ��E��pq�
y��	��̾G��,/ԋ�.U�N�q�9ы.��l�Z_&�w`��̀�J�'�&o&+������ځ���j]s���J�չ�x_�
b
��� ��5�a���R�ٻ����t��7*Q+��ʫ1�$Z��������gy�����SW� v?C"��'�4|u.Jv����N�Us.�_8��*b?6���ZiR<�ot�V�[��vj�Ư�K@}��Y�׬��X��(��QPH�CD;�����\H�W��|�I걓Z$�]UN詹��5*!��� \�}t��4��$E���5:�d����on 
�&�N��v75)0�s7uV<��.6�O^�6�W�K�g��M���?,T��URA%�󞡖�/��BO�1d�?=
������<6זt?�n��;z	kt��V�4�/�b6;v$�]�L33�Nn2�����m��5&�>��5*�\�X�J#ι�ճ���L��67�>�T����=Qϝ������}˜�1-��c4�c�wX�{����<P军���˕�H
�i�%��=�?��d�� @A����`.B ����Ɲ�����U�����4惕���߄�41fA5�^U�~k�~��]w�D1�����'U�������yK��[�#��C��"'-n)XΌ�X���M���E���a�|C��c1����=�)iI���v��$-k�4� \�y�훳�s�3�/�����4 �_r���4ѤQH��#�(���u�H"~$�^��d��Vu>�m�p|}���86D!�qu��zk����ֲ�ɪ���P�2[��l���^*����,R�,�-��vj�I[C:gu�A�m4�l�e�(��l�a��~�*�o$3�����g����;G�c �-DK%9X|<���"�[�*����9�0Տ�H����I����� �U8�®�A��O�Kr�_������y2�&,͌xk����}&�:�zx�:��� ��HI��	\?��C7��GF��(]��)t���d3H/,I��ҝ%�{��6�s����g�-�E*��>4��ۿ(��㚛�D���n�����Ւy�UA<d����Qf�4ǂ��T���á�F�k~@~'���0�si��o�����x�!:.�a
sF=F�=qMu����x��|x�t��W ���W�(��y�W|J�����K��o��8BsQ�̡p�D=�F��,��=�y�*����(�'�C�eF6s�	_f4���xC<QʂZ���zvv�`���p��njϊ�C
��"+EE��g���?��W��[�	����w�{�=��#�ѯW�#Rt� /,+�.���P�}Ԋ�g��������mc�Lֲ|ɳPF�o	hT�����G>i���V�posu���_#� KWq��6*�jr�X~|�<)I������o�������Nd�O4T[S��m˄t�R@2���<8�in~��g\�;�n�qE`����`��$g��xp�͋2�y�To�X ��t�?�B�iޖ���+��>����"/w
�30%��f�.�����ZS`*ٍ�I�^����u%΁��V�C���zkc>�w��R��i{x������.�7�+-��\���|[�	pTg�X�n�@3f�y�r���.[Uh!�N(x�V�1���R�{�{�]�"��w>,'�9�w��rH�q����|���έ·��]P��#��
2kU��4��\
0X��=���.[֚��4��A�#����تP��_7���`�m�<VH-5c*!g�?[i�"*��@�d�=Ij��kJ��(�y֬��h�.�7p��fw-9hUg7O�?7Hd�G6BiR)�|���!�GL�^,��	����15�0��E����Q���"�No��&\OV<+�K��AB�AA�^�b����ky�����չ�L*R���������f�j�9�0zB|��pN��\�9���ȑG&�(l�CP�Y�2�Q�O�����iy-�TU\����������ط��0��	���޳(1�]��t��p� }5}���B�7 
��#�D�v.4���C$�������3�n��u�������PNO��܋��#'1�\k5?Q�e�ș%j�v�閆28c���B�����b3�����gx����V��\�O���o����5�Z*A���s�������m;���v56�6��qN�$�۶�ض�������73k�̺��/d���S�L>�����#3����В1��~� �����/ߺ�~g�b?�<�EYc��ڢc�A����-^C4��B|bS1)Ja���	�� �����UnUU7 �C�
}!5�Y�"`�菅?��4�]2�7���	V�����L 8�1�ht���H(�aa|��^��t�b�h�N�4����7�s=	�~B�����x��P�.R����q|&��r,"�,�?��1	�qR���ECz�����Ju������L�x����9��9������ j�-�Fˢ���Z��-�flw�NFU)���쬱:�#7t��ʶ��CHݩA+�$���˧�^�A�p�T��T����ncSơ-HIEHҔ��y�I�c��m
.5����
�U=>����)����˫)ٛ*{�(�{y�7�QR�+6�(`�T"�u��1}�!daA�K�r�#U$K�7� ����?H+�j�z�,-��йWd�P����\đ\)`�N^^N3�#��S���E����}���}�F��2ߗ�I(���ۺ��f�qaf��+);�U`��Ozu<B`KV7g�ۿ���q��l���:[ThtT��	�.Rg�$�"�	�,$��4�ɺ`i>$��^�.s:�[v�����l�s��$ۦl.H>-\P�U�8��O����!O�!���W��j��&��յS�s%K�y���kiT)�Xu�#��mXp�D4�	=ݺ9��}�i�*<B`����� ���y��ƞ��u��TF�u%���g�Q_�]W��G��W�uJ�<v �dj"u�J�ݔy���f����!�jŪ�)�_<�Am�E<�A+�Z�!�UZ�A���)�u�<�,���$'E�e !�[?�wAJ�	����Χ0��k�������$�H,�7.�5�`w�8� ZE��Z�(>���?3�����~�Br�� 'B1mo��G�0jc�ԅy2�q1{��&�I�L6}{ڋ��j�x�L��L�S�YeVL]��;g|���*��CCgU���
�@��[�J����@�e�����������m�݋�ʁb�`����b�{9�ds�������r-�J�2���_�̲�.���ΪP+�g���X�Y�������;��j��V�9���,v:'zS �C��\:[�?�T0��؅��@���C��[N�,��L�F4������3-J V*�d���h�Oǎ���Z�a���:��tg#Y5s}���񇛆ճ�:h�v�d�~���:��;M(��,BQp^�"�S�������Bw��Uv���.����s�oN"߭L��`H���/g0��`����A��<Ԉ|���n�� �8��>�=�M�;�H���=Z/�<�
?ʂ���ŦX���������������� 7���j�7^G��\���������^�W�nQ#G�
�1�#�A9�@ϸ�\&D؊�[���ufMh�1�	�X���
�eڲ����1�l�z��?X��~3z�����!UXrCt��V�	O�ց}�3�$��L��:?�.4�V,GODW�\S����w�����v�?��}~��}�g�S	޻�+�	o*�ͥ\C�x�W���&�����8�������Y�|O3����(�%Xogsc�i�{�נ�.����Sjr���X5Y:�����8UI4��6�i�7��h�J9�����'F;�pZ{#e%G nfEoO���(ی��C������;Tl������n�8�A���=hR�S`�JZ��R��`��b�s�>��:��8�����ɓD�p���#Q}�!���Cr��{{����_�^T?���>q�s�T&d5���~_wwd� ���J�X�-y���� ��Q�ͩ��7|��Ũ
V�i�$X�Ʉ<E��-�͘;}Q�Ȧ�9��h.�S���X�ƙ��1YU��m0B����(7��M[����`?O4A|:Q%;
����U��VO \O6��$�@�;B8�X���.[.E�<U�sdk(=q�*h���@�e ���h
�֘e�"�T~]�2P"�p]1�
^�|���_�t	ԃ�C���P|���)�@r3��Ќ�T8� ob6#�#y�C���8�T�X_�E���9���7�Q:���6�gXr��Ó2���3���ZIIyI��Z7�0DQfn]Nwq��>0�������m&&����$�A��I����I��F�#���AM�����:�c���7�ʊ�6�����1�c>����x����]PPDE���JI�����Ҵ��O� S������y�X;�����0���w���"^d�e��@�8e	���KTӧ)��lҜKW6��ja(Mf��;���U*��8`�RkL�%�Y�bv�7�-2�����ޤ7g�F�uwYVXM�h8A]&���53�a9�l�U���u���0i�)���c_Uc�mfde�c��T�������m&;��>>+�e<�e�_�pg��/�?���j��upB��?x�T�f��)`C��B��4p���9A��q2GՔ��(�01�YWԥ+ރ�1u���S��C>8gL`�HT��X�>�9y��"O��{=h�;�M�X�������sv��]a�}�eYR�G萆���t!5����A���q����d����;"�4@����{��H(�rF��E^�Aܿ��e
�4�z�Y�?�$���m�(��$���ĳ$��NVG�_��z�"���v��c�\��a�s�8��}a�Q�K���A�C��M�Ɵ>#�
K$=�BƓ�����`�Ho�"����*5�~���49��I��#aO@�*��[qG�JV�Vs���xON��G͡�Ә=d�Sr��J_Nɓa�)�LMF9��ѓ�����9�gRb�x������2"��sՊc0����吂pǎ*�q���@��p�� ��7iʷP���w<�֟�q�-?���ݓ�2,W�|l��v"�>Y(^]j�}$a<�6,���IDz�b���;J��ÿ-j�K;���QD�ܔ��"&r������Oqx?,����f.�U�Bb�J�bX�@)�Sy��y�T	VT�`3˕��j����]�H\CK�NZ+h`�eꞓY���v-��M������W�v��v���ڊL�㟚0���*�:L@��.Fk*V�7�x�`B��g�u�Ӹ�W�??+͂���XQ���x�������`��9�\[R.���co���Ko��5_e�Z�P�S���,T���� _s/��L�zxw^]�g���4����R5pБպJ��*�6�9�zVӰ:~�CG��Q'|&�=���Gg���_����_�v��E����2��q ۳�ik���\EƬ���*��wASܘ���ΒQ
6K��i�q�z%�;;��*����Xt~$��;�[|�@t&�F�w.�"�'Po{ț3��\�4ҷ��j�Ka��^t�aͬN��xz&������{���B��)6����TO�[���}j����+��s�J�~�B˳:P��cH܀������x�d�,�}"��s{�5�i���0/�z���H��ջֵ���Zc�] �Fʈ��m�:���U>Y���y~9A�-��WH��m���s��3�e�&�C� ���J}R�#H"���u7�4��^�Y��i%Ox���֋ɤ=���'��:]F��/�I �#"ܬ��5e�g��	�Ǩ���Zugm�`��H�`)�<���N$�֔U���d3��,h�c�O+��<��y������\�&�I �������:g6��\�.�-4�Ɍό�c{<�;��;@��V�u������[��}��~~�j�L;�Ev_�!#��İm
�����gI���r�Ǣ=�����)�n�-!���q�=�Z�/�%_���Հ�
V�[>%|����a���9����6q5�۩�mA�~�U�k-j$D�Q�j���|�AT����N�]�,:bJT�����;��^O�rЧX���Ur>���4@.b5��4��b�i�L3�Y�̏��J�¨��ä����j Ƈ�S�w���Q@ܸ����;�#$������E�y� �e�Q�eTȩ�T7Ө�	�ʾP�Ey�@���C��;���ZbS%Q�Ŕ��vR�E+E �숦9��}P��=�!�P���h��Q�f� �Mr)�gX$qhx�-���c��(�'�a�cBiK@U�FB��:����:�BU5��`��@���p�[�n�p~X�J	E/z��c�&�fO;u��O����fIDt＊D�ݬ��
�Gٲr��tK�g�,�/�����������s.��;)K(iO�X�s�|N架������G��أM��T��*�4��|���s��2#�JE�I.��iε��o�bWӨ/0۴��W����Y�U\J�H[���42���_�u��Bj�t��o�p��%���J�8�����Kj͢��0�@EtB�58]�X�|�6A�ͨ!���,�-�ܜ]Hr�����<�Q��-Hi>��E�ܦ�����*n��|R`�6��Ɖf�2G1ې�O_C��xQ���/���_�KX�ћ쌚����U�ꇀ����W���g��O�W��߬��%��R�k�ڣ,�'&�����[�g���U�$� r��_����S����YbZ���a�`���<ռ���K����K���2�t���E��F��࿀�~
R���Mʍ���j�P�,������x����{�Ղ)�C��$�D��->�.����&p���\�M}��9���~�^q��
��B���`�ʶ{D�ޢ��K���_�C�0����^g�m����O,q��j�lVɬ)=�����Xg�,�j��a"�#�s���`X���^���m=�s+���c?nŅ���Z��T�A�g���X��}��| niJ�zH�d����i�u��2�D�����g�58W�a�l�#9�#8
�u��?]滭	ׂ���<؁l�Y���-v����
;0�Bu���_2��)�]϶d�Ǘ�P}�jt�d`�YR[���n��]P>6�']�n�y��]<o�-SK���+��a��#t��5N�����ų\:���'�i�D�	�{����|CX�R� {+������ Vb෥������[��R&h��
]���m���<�j��g�h$�;7���W�D~�
�	`�U�,��2�S
�N����wŔ����i����<�a�@��� 7�8n>ָj��6i?)̀/f��3����u�ɰ��rzK�Z�|���Z@�|x��ؾ	xҞb1�;���R�V'����0�xE�[�ۗW-�\@���� (�T�I-Ì�-p֠ p?��������|Z�L�*8�`$l$���s=�i�fCo*�T��;j���?A���׆}���xq���ߓ��%]�(:(���Fs���q>�,\T��:�pX�^-�m�2�:�]T�VO")'D
	sM�d���B����h҉B�x��5��u<�<9m�Ge<"0] '�+�J�:�v~Zj	!��P
V�Q�|/�w��o�530�e��;\Iu�c��)�7ZT�p|�Q��b9S�z�m="b�-ǑNw{�A�ďiȈ/`�8"<�{B�@����(������@���+Tɀ 9����`@(2��x�M��zz�=��+��bٛ��ξ���0�`�P�����Zb
g���ZaQu���W ����i.��w�6z�|�'P
��RC��'���YG@=D��R�5&7����1RO�Ե�jr�HCj�a�I��)�36�ekY��,�A.�PG�f����#T�
B���J��HN��m�B��BX^á�2�Laqe�­��F4JL�A��2��mIC��?��9�Vw7?N.J�1)�.�Q6@��:l�#����#�'��QHY���{2���%=r�x�,\�R�� �
wMn�l$�`'o��:0z��ʒ�θ&�^k>��F�t�ƈ_O�QM*�����!�[�_��	�i �]}yp��"�)��f$�DQ����&�)�6�Z̵J��NO�KaZ���G�Y����O�ӻ��j���@y˞Ĉ��OG�[r.���o:�0�t͊�r�c^��1��!�6��d�VC!�N@�BD[��%ba�K�@�� Q���q:=�Y��ߪ�3q%����A���E'��1Xh��7cC]��y��h��y��C�y]�'��:K��'����a
v'���}X���ک�e"�-<�-<�"q	��5�5��p��Uw!���2򉞻PK���Y\�N�Rq��>��}r.�d��M\7}���j���2�E?�_�����]�Uw��ٗ�+����"吟��O������.\ƀ_��jE��Tϊt>,؂�W�Q^h�~権]G�I�����A�#V9�l�F�����X��� ����3fY;�<�������X`N�Ff�q����l!�]�2<P@y��w���_�^%�E�~�U��R��d�=�,���"�V%��w���S��#�Q������N�4��JهU�3h�����s��C����L����R��~�2w����Z=~y�M�b�-"�%�9H�nD��#�����z�S��l��O=�����um�a2%�� �����l	{��≆!0�3�0���`:*��h!55-�,�m=8n��fv*~�j�|�����)�U�v�����cc���>�o�V*�7׬�N���m��U���wDi��
P�
#�:��Y�j���M0�s��3�v���7ޭ���m N��F��� v�:��U,o{^�ZF��/�V�+2�TS
��u�/�bO��cV�l���G��{��X�z��j1���	�CpS0�֒��5).E$~%�AZ0h��$�o�)~Q2�TU.�g���А̞�#��E��{e!V�B1��}(���zQ�,��^�Ԟ� ���+�Pw02=����!�-����VX���Xdd+�̢m}�[��ːD�'Fp3㝫.k���!��������#�)(N�l��}z�������3�31i,p�&�P֟��twQ*,�|��GB��p���������4񏟿�>�y>����ch���㥁�$s"�Z��"��j-8�+*��-ome{УVf�_i��
�����[��w�I����.M��ty��d��x'Sx�%,�!�_���A���d��j���acD;D͌v��,>Ш����1��xO?��_�q=��\7gL|�&�6�ps��׿�y7�X����u �q!�z
���B�l�/��� 8�H7����`g�̕Y�WyİΠ�C~��}����ke��H���
_�>cz��݇�����+����~*R�A�xO��ʠ�4K'LJc�VI3j�EU������G�Z&v@y΍���,�[!��
T]�W���[��c�(�x�4Q���=Vl	S�ˏ��]��Х�A��Q�^[yː��h�v�֙�������4@�A����?�R"�nH��$�"��7E~~�����,u]	楹~Ր��/��RC��@X��Ա�_oj�a�h'?�U������1�h�]^����`��XVd`�$
��cn��5� �f@�

,�3#Y��ש�mg��7Č#fF3��CR��F��VK��c��jFu�U�㦪�=
��q#~�����YƊj��e�"fo�?
�����Ղ��S7�#�����!�ݛP]��@5C�QV��؎�,5�l1�l�D�pӺ�fe��韎Uay&�G�Aq@���	l�|�nZ�JZdj��í�Cǖ������uȔ��!���J6�Z��m09�}�]�i�3;Վ�V�L`�r{��%�j��* ������[#��m�h�����E��\�>�pr�Hmf��JB����7jm������!�C̿ʬ�>��:-]\��s:hl�2�U=A���������؀�������g��Y��vd���V��e�瀶
� pC?[#��F�'#3|@�!+���X�D�!�%�E$���,��D��\�`2a6ENq��-�C�ŏ�1�ej��j�R9���,�����Vh� ��{qrR��<9�Z�S�+�OQ�|6v��\�bT,)t����V���>��+>���D>���]&~��lɡ{�v�՞ae�Y�/Q��_�T'�q�a=�������1��ɂ�#x	�bjK��W79b���;�=��5��=��U���i�
�3��Ӝ����(A`�7���'��!��A��a��Cݕ�NX����yK�{�ޛ�ϝ6�@*�7�ڎ2��.���"�gV��0���<�.N�@;�n��W��KJ���W�ʏG�A��	#Z���ؽ$VL	a�,�&���^�k�@H'�'s='����N+ts�IcQ`>�B½�J\4��"��ԠZ����eJ�^ ���z�[���#�hzZ��DsK�ýqܽG++��,������]d���X�f�a��Ǭ�_b3��|ݛ������3���Xy����ڰA!��](�(��s���> �iŅ__���h�n��.3A�m�뙄�-���jw#/�%B�Q��jS\��E���@�f��"�z��������b�N�x݃ű���Y:�&�T�=	�[�A8�]��~{1�Zjn"�%t�W�3�Y���p�zk>3JV^�z��g2�Ƒ���Y[�!�f�����H��D���r����l\�%��b��9���2B�]r�^�:�T���y5���Q�7�Oao�0^8�fH��K��~���p4�;r�=�`�i%U�V�~������f����Uby��3_l��M?Ȗ0�q��6b��r�h-����<k6��l��=�Z:���g��ӊ�]��}����8��.Vx�~	�ְ���xY�m�.N锂i��Z��R�O����@}�&
*aÚ7A�[Gp['��u���X���ƴoR��J�BX���O��(N8H3�Ĩr)5X~�W")^ ;��u���Z�8�Q{��1�+߫��S�{�cKs��n����<<@��'}h�z����-�Ggк.Άn���s�D�#�z^+=��(�M2�����P�ڪ�[B���|q=xY�]���o�s(R��$Y�-0<t���Q|h9=��Y͡k��h(']]e1=~�	��楲OA�+g�R��b���kὖ�q�U�N1��&�*�BbM?$������A U�M[�ѐy�N��D�"�������$�zz:ؒ�S��yQ���~�7���0�e}ym�~"�2�`�ݪ}�wZ%��n�����b�������$1HRU%�r��"�5�_�0�S'hU�Ц���]3iQ��C8VE��B���4D�0��O��߲���̣�ӕ���uǉTM��b+0�f?cr6-�A`�#*-Cb}��p�8���'n��F�C���ʙ���i��5�YP`(m	e�:�%�9��z��y(�־��b�"�b����ɍ����zJ��kO��]D���e����U^�:a�:R'�_��_�%�h��5N5����B	Bҙ�#�'�����(�lh��n������S'�ۋ�o�o��UN6d����;��K����d�
�j�Phjj�"���(�Y��XZs0��c�
��O�.�楿1koH{�w��擭�Ohk[��Eyqk�\VA�h���!*eI�ʖr��RǗ�ח�y�}����!$Ɏ\X_T;��tD�㮄]�ʷ��
Bw	��V�I�s�P��5��,�e"�]�a`�W�g�l֏��-r��Q�����c�Q��e�n���Z�	M�<�X����KV��ɗ�Hrg'����Kcۇ�Y;��"B�L�NCї� ����00�>3"��jB��r�_6��f�L+R�W
�6	�H:,R��${����5F�'��N5W!�M;ݓ[�E�*Ӝ�l^��"�^��]�⵪�`���,�2�-�=��ʓb�r�#���<�?����|�'L�>Ť��Ǌ _��~��]�)��Rކ�5�k6�.��ZF.b��3���R��$��+�]�Cv�$e3+'�_\]}�gj��$�qE��urx^��9��!�|?ab.-I|ӂۤ�6���Ƽ�ʩ�l���U��4��_�����!?�g ?�����Pf>F_�Y�g�_�>�T�=Ղ��N��_��y�e�����RF{�`��*�p�;���Wt'�3X�KP��V	ø(�$�YJ2)�59�#�����f6It-�\�N�4�D��b���QL���S�h������&����^�ׂ�§��"�����'��;�յ��X�]��Q�g��$�a&9d��9��{�X��y��rx͈涪7g��6Pzw[8o7��m�7����7�N�+����,}U�YP�^L�&ps#��GgT<�:�ε7��/7}nӬ�^m3hA��9~;u��Y��Y��`l�i[p�]iD����Ꙡ�Y%}�42�-r��AiphCm����\��(�r��%Xb�E��'��^C#�B/sǋ��B�]�0��0�uD���!��K���%c�-W�#� z7k�{�vuLԻ�;�������r����8
7�Pr��
�(/�/�f���feb_^�rb{�J��R|�1M�5}����O�fL�d���X��Fa�nA�B&0�(r��+�Eg�L�!|���}�ҕ���ib�#��!E*M<��<4�s��qǯ@0�ð:<t�Ξ����|j�)U�F�|�y���g��oW&D��}��/X)8�J�s �j�Wљ����a&1I�Զ&�E%,�X^~<QG�o/ �J7�v8���͹ԍY�6Dz&�0sK)�n*:�1v�f���5�Y�޵�9�-��2�x���3or�>�f�&P���<{�b:>��X�������ف����9+)*�Z��	Z�����J�E��	��>�7�>�LnU&.g��WJ>�7�E9�ۄR>�=O<_-�f�W��+��fx9Wͳn�N)H���pU�i*OF�����^G�X����sZ���6LwZ�.E�p���k��V�)Em�H�+T�תZS�#t%(t��_JJJ�5�� Q�Ӵ�er޻h`y��+���n&��D ��|w��5p��Le�t�?(��n��4��4ho>�R�D��g�g9*�cj����%	f+F���YNF�)#��2ĪQ�����g�X���
,hBt������x���b��}���L�xcX�:4����
bzr�Q��J��55��(4�H�]�yi�F`��,��R�����Şu���C)^t;}d�P�U���xϪ��9Go؃�c�+`�����Q��1x޳�q��Ӭ+B`]a���A����#��r��-U�'�O#��B[j�eD�.�O-ۅ!�r�q���#��#��3M�u���L�_ӭ�r�`�%S�*a�à�a�2Q�)�j�A�%q�' �@P�6�ֶ��V5A�E6���_\� �8��@&���0����2�nP�9_���kd4B]�5����0a�'>���SSÞ�(�N�>'��:�ͺ�Jit���]��3+�����nX!:٥1�څ�x�Gp��8Xp��W���1e/r솒��q'+'�^��T��!+�v�e����r1!��#�1K��Sx���w�'uU�I�Fy����o���{������������Q�����r<�^�������e�S�&�W�N|�^�rF���L�#���N�J-�S�c��o��fM��O���G�P`jjT!*����@w ��aY��	�亦1���yd�s_����䶛�ʻ����O��C���{V�_Q�-}j��V��D�otzު=E2��_���[]~�W��A��j�	<>y.O9�EM����eN����B����͢?�2LmE�;g���ưP�|�rS[F��s���:5�.��(=>d�A�*>��7M�����ȃ�a�L[S�{�ux���9^#���C�'�!A�0s������|�-��>��������3�r@�����u�����O�y��|j��wB��<�p�G���u����βyM@-�rЧ��ؙv�t�w�����e+��iu�e��oa�v`ˁ��as�cr���t ��7s�s����Ȓ�����U��[%X�71�.����Z���P�&5�����r�7�]�����P8��:X帴�q�E% 0����<�����<[/c?�.�:���6p�R��q�I�m(I(�m���w���S����ט�}�ߟ/�%��P��q}N{��!l�tWV�N���-�m�l�.���lͯ���t��Tm�pc�q3w�o�f��_/Q
+bC����k�Я!�o^�X3,2�g3��O�er�~�׆9{ ����eV���6��bN��*��a#���L��L³7 ��/�%��Aw�[.])�J'C\��M1�o�^A�}Z�=��� R5�P��>+�ˮ����T�Y�
�y�/ �^�!�ׇ�S)T�!�v�5�O���T�
(#4������(0D*�D�^�r�վ�]���x�N{*��i�`��R�(�W�u�L�}<�t�w��z����S��H��4�,��T��q/�@����%�Feq6a%���#b�i;H���Ϟ'ǆ3�F(�,�}(F\��q�r�p����hZ"b�w9�'�8gn��w>SgMP�E�=�������=�M������4�>L\�g�=
���dY�s}l_�K ����3"&{*�������u�~h��	������tY�>�5Oq����$�(tLBU����Y[6J�;準@��V����#���G��N��钀��	;�
A�!�|�3_X�^Yv����{�����v���waXwaZ7%mגP�� ���@U�A�|1-.� H�2t��W�;���=t�I$32�v��F(m2Pr��:��gc���"�⧷�~c~zIM��)r���tzI�fDDrD��Og�
�v��*7ݹL��{C��]T�Bju�l� �r7N��L�,��we�2��졏;�鿺)j5���	I!�rm�������94�Ǣ3��_����;�`t&�C �U��H�8xq�=�˺<�M<�g.�Ί�Tcd��s�>j%4E�?�G�k�t�a�|�~FR�&A�1��E�ހQ0��5��֐��	�	�0,�IĿ�/��9���P}U+�V�s��p\I2�K���0V#����T)__-l��ek��Ĳ2Ū��V
?�#|�����cU�P�\�6��[�('
Tp�#j� �s��ʹ,�0��{z��r�ܟ���FlI�8o �d�F��H�M��@4�$�HrB�����%����;�W�/�cS^�iD<���ܪ��L�S��}��v�a����q���\q�p��ٱ7��^�ҝw��sy���Y	�����h�	ڙ���ߓF���V�����^G62�H�[4�b��S^ꌦ�*^��lV���8�1T�&
�܎�W%/�z�tR���˼�ȼ���yϯ��e��`�aZ��3ZQI,��nOI�%�Mͻ��#BY7����Q�w��E��>�Y&2�&�{���-
űS�/9����n������g�?(~��i�ݨ��f%��gY��c���݁��\n�|��~�����i{���\��Û�2vs�]��8=d���/<d�_b�Ӟ�Ȱ�q�>CP�jwgw����1�/w3�{���mМ�_��yW�-����m���\>k{Y�)B�/q�\���B#3�����ܼ]N ��n�1`'���s�/Ӌz��$��M!VU�S+Wy�x䭶���Cm{t�{L�g4-�K7|����g���ցB�>I���CD�,K�$S/+�ޣ�����ڡg�P�-��h��K��-��ވ�:�K7�dH,��{I�J��W鹎S2�c۞��>$L��}�	jv��|�;i^��~�'�����:��j��������ޝΝ�7���~� �;�yf��?f�{nj#�7ի3q�P�߻2A�MT�� �3�gS_J��V���}c���<ɾܛ_v�	ÚN�Ev�s���ǂ�ImAp��Lv`�j@/�ʴ�٢�h����#�y}�i���z�]��Z�w��1rvj?�,k�@�y�3w$&�3��6.'��1�6�ѹ�0��.f�.�7R��<hhq�+�n`���ͦ�opi@��'e7��Y����2y���[.���q�蟽��qcj��0�S���gX�?��ל�t��I�M�sI���OS�$�I�^_�QC���g���~Q�sMM9j]�LD}N�@�zA�s
+\��{[���M@"C������I0�RL��6̈́��|��,ؚPT���v5Au.I�V?���CT'��������7��OՂ�ש�����9�-��}WW�!�_�{�+dW'�w6��>�9�7pp���OaЌ&����p"�����|��EGc���6E�"�J�ф��v�\�τ���%�O�>�6";�n�]St\ξ:Q&8����1s�����<k�}3�>Ƙ޴t�c���u�s]Xtz˝0���|\Ѐb�p�,"q�i�B~-rF�'�����{7�2u���E�H5���`K�-Ü�Pl�{qN"쿇SY��%c�25���Mo~�H���|װ�N�H�)_����x��J��4~u���q�����t5�.ؼ!Ȉ�[uS�0(0׬i�c���pވm�'�<��t"VW���m��ˏFU���5�SZ�~�\�m��{T���4��a�,6cqP��LRkF�X���Q�}s`>���@T����C��0����;ؒǁ4uH�ᘓ#�47Q��Z�Bi~�����)T���پݐ;٨������M�Upj�G`؟�ٳMn�^�<E|(Hso_����u� �A�FPtJܼ����8iC�;iצv1-R�o�:��K�j{R7�9��9�#l�w���C�������2(E�
�2.��� l�+l�c>��=ɚ���\d� ��W" -$�+d��fBQo�< q%�e��>�������UL��C���0?���R
��$��A��1Ή3#�u	�k_4:7S}� ����t�
zw��#/�e�8Lr�,��T��V!*�/�k��Ю���W�
z%��V��B&�o *ܯ�1cT8島��(�N�~���-����Y�#���%\ِ�}BI�EM�O�-c����QV���+�S�36�a��h]�
˃9�F�5KV���Si{),l��c�O�x� �qm6z��3�ph�d|:��l@Φ�v�������i�,�F���<�)��{�V�q�5�	NB8ۙdI���,��v�9��8�L��nڊ0�E���h(#��u�l��E}���R�E��#@�4l�x:>%�|o��_=��@��y��Y�ǛRtO7�-y�(���[#F�BE�zEr���5���̬�aSs��Zz���d��d�@�6J��:�H�$+B�݃���U�i�^2�<$)7�Y���Vߜ�Ad��+GzM>�=6�{�L���V���n����d��W|�L{"��m�E_�-���?�ח���`����!�����^�x��Z�'��^�++���R����~�QgP��8�cn�D�u1V��$�۲�oL-�:�	s�tX�D-�Z��X�y��Qi���8�~w��Ш�|q�|��t+d�����f�_�d�͹W��f��9���ӳ��V���VpOk���C��C+��Og�\l��(�6y�6�)��)���ۦ�߽5��i���N��Y��|�։-K�� �~���!��9��1��%��������,Gi.���F��X�/�B�_�3���QbZ�&���+���C�8i���<�Tr����X~�̶�ɵ.#��"��5� ��,=h�g�8�w��8��t�r~�M�><��0�u0:��|���`�H���fT�J-+�Mꀨ���0��E��CٽC�}4 �!"	�ړPB����4�`��a�^�����`��
Z�0L����!����N�V?d�B�ȇZ6�/H�e+i���BP.�q	���B�`���,��+;QPň��c.'���F��\$�u���,�w�u��Fƭ�����zΥ��b;��w�CrF��"B���Aw9�غׯ��M�]I4!�ܨ�d��d,�7�S���Do��=h���$�r3�蔡���4v�b�clG�g�M��M0�
6Ms�`�V�,T�۪�X	�j�=|�K�4W<u���L iNv��nxʿ�r��Ό��G�[��u����@�B(PZ�-����^��Cqn�kq��-���^�8������d�����d���ϵ�:[�[1���13��*т�߯<e�|ľ�v+DI*��*����ȞELht�0��u�[�>N��}�����vta��l-?lB�3�/0�Ƥ9	r �UW֫%N˺����f:x�B�
mə=d*i}�}�Xz����LL��P=�_Be�b�&~Tp����/?_=H��!�CE/u^��k�(� f�^�=]���꣛�<�`�C��pP��M�����o�_���8e!�A��Q��U�".�9B�A[�k������P���x���W˩\��L�Y��J�!��/1o[�b��"�%��6�q%1,"c�-�}-U�M��c��,a̅
bg�=L�bC�C��r������+�[��ϣ�z��cV��l�`3g�I6�?���s��A�am�@�W6{c��o�RrL��/Vy̏��ܜ��uH�O��a�
������k?V�A�ҁT7���W�wc�o��rs��gLA�F�Oa�&w�'R~�n.�f����w��P�-F P�-[!����3��G�UR���_��/���4�=�n(����Q5�m��OVΪ��`C2#�_V����̀T���22P�7y�*���.aoMb\�w�_A��4���U��69p�H�0�9����V6#R9������,(��E	S��0�ļ�<����7��luud	
�T��ŀ�☥�����1�\�n���l
_�M�8i�Ơ���C�;��\�dLJ�_�0���j>���D��3	R)���I�F�����n���l�`��>~a�uBr�V}�|z>�+��m��a� H�f���l��?���=8�v1��|��:�B����ؔw����3� �� L����lqagl��z��ڜ����p��A�(r��}�hC�=�CGN����E�ry�hp~ZԤ�\;�P�n��G���@�؈ʲb>ι?`b���Z�������5��
B/˄]��@.�n(�y���������؋�� =̽{��]��O!OP u#��T�����O�����xh�۬���]ƬY��Vŋ���F���^���a�ʀ����|~}��^�z���D\j�䗬Q?8��dUȐ�9Oc��fSplQY�5.>���N����9@�7�O����6	wlj���ސ%��%E��j�|���s��9OG�c����G�X�3�jԱ��M۬k9�xvkֶwS���h#�(��$�|=�ts��]��C��G�/,Z�]o>��J�<��6ؒ�8Oۡ�$�F�+����#���Zʮ�C���ɋ��H�Pg�?t��A�ץ�������%�YI׽�����xn�3v-B�c�u�f�r����^��:T-�ꢂd�a�9��W�H��J� I\\��P�/���9ҍ��G�-��GG�n�Ws���᳛z>N��i<xX�Xw\�����y����lv�19R^#�l��x튤�������04�A*7�ZC#I����Ko��T�#9 �;�MSԾ�uN���.�X�����/k�z���Y��j'1e�������F���[��E;�W$vzj�4��>2$My���UPa? [��h����iL5	s̙�2?��p����Q+�R���1��}�5��(�7=󺱥79\%ڡ��C��rm+�3Vn�IK~�<ǬgN�}3���M�=���*��҈hÌЊY�D�:��� N4A?���qf���B��ꄽӄ�ox�-�����������h
���>V�G"E%�'%�����-G�-�ZmɄ�4�z���\���������(l��������P��D���Ur�&�<ޘ����{?b�R�����<E�x(��P�P�
�L�D�����R~Pϋ�,�(��ۜLڞ�<�c��h�zUH�1�^3p��nf��g[r�y�#I�$B7 M�).����_=����<���5�u�2�Z��Y?J��.����_jZA�>ǲ����a����u�M	����Ɣ,3�L{��`Lپ�Y ��W"����YA�!�Q�a�Mwu�8Y��',:MQ��
��r�0Ko�r��?U�4�k��~�g�P(�Zу9wT�Ą-��1�n�!Gw���^J���cޕ��ԋܕO�Ga)�d����f��j����[&�`�oVj#�w���S3(�XvBY9�F*tu������2�e�f�AxN���� �t7NrW=��{ݐN��.5��ѿB!�"���Z�R̰򗼪I��պ.F!���B� �A����Sӝ����f�X���i�~S��ӊ��?D�Ġ�r�]��C���e ݣy  P�)Z�>���"�'q�����ޙ"tU��a*���(�]��x�4(ϵ�+�ㅱ~3c��;�����p
���D{��xQ��y>}c1'�qG�sn}Qm��Wpk�#�ս��y-�x֤��
��lT��{�����J���s;�	�����Mk�k��P�ƥ�~*'�*���О�[���Ia����|���X��P�Ÿ��`�Ʌ�s���t���a��;�y�HY%��Uþ�wFf
)�+(�P��Rj�s_�F�$$�8�ך��+"��)�YS�����������H!$�r	�f��t��˽�X��!ժ¿I�"�|��L�Q+Jt�/)S��
`F�J��z~��M����v�M�IF
�d��<�e!��C��)vNS/GxPG
k;B����8o���.��-a��j��8#HHI��0xH���kLa�""�Ոq"�u���M�N�]�������k�]wO��z����Q٘i�����c�U�vw|X���.i���/�5�;�s� ��"�"3�Xg"�͂	�&���3�CJ5�,�l�&5#�0A�ZJ{��hW?�e�;l>�������A�H�BNz�U g�O;�9yCN���b�ֵ��I��|��:Ь֮���%�-P��^z6\n��l{/�<S� ��ȅ�;o��.��m�t��/E���8�轺����ٹ��K;\г��At�p��~t�>g�O���\��~�Q7�5������Ϟes6�k�ǧ�!\R)�G~�S�{��'�g���Y�i�8=���qI�F���/}��R)�t���R�}I�b��w��r_5�������A��0n�Z�'d̐�}��BW��dG�6,d�������}�,�ѷ ���C�ᤝ���V! H}�-�	f�F��h(L���O�����tJ����j��ӽ�@���:V� z<hL8�E�]����C��r��>+���aс�ldV���DA����s�����A�8�^5�^+�F톝�䡍�h�R��e�c�2�J݅x��?fy����l���tCõ#1Ӄ�ә��n1�NE��2wR�g�<%̞0L��u-s��Kz.n 'uEE��Ó����!��0[O��n���e�ϊ��ȬYׄF:dj5av5uy�׾Q2[Jc�: t��t/���;�&k��VP�s2�pY���M�$�=nL܉����?f�����Ɵ
%@�L�AS� ~,�;����1S:�7�$>Kq����?�����Ě�j(�����&�ǳ];��LN΃�n�� �²���\/��������I&��:���?��!>O��O�As��.L�C� ����[��[�OFRH	���7=��_.�(r �Y�PYbޥ�� �����݅�#�P�H�� ��nT�9�[^m����:;��,��kap�^2��/���t;#�I#�ǐ�?Қ%ҽa�G`�]��r��z��I�@�Ǫw�y��y��O��W���O|���ǣ7�G��zXC�����������k�Ǐ��mƓ��Ģ�/k��Y<]d �&q�������3�{bU�"�Xo�e�\�V=bWw����ϱ�[��gf�o�~έSc�e9�Xk�Z3l�^={��O��g�m�a��oU���Hn����70%�ȑ��P���x��qFV�'E���癞~|���_%�@�!��r��40fc�?�ۗc/���3&�S�R#�+ت��c1k+l�
���"�}W\îUő�T��uP�I����r�b�����;�f$2�D������o1���@�P�N +�o��m��v2���{(\�3Rג���m�_~�d��2ur+"�ԝ�/d����T�a�.�K_����Q�(�[yW �!�W�ǈFK!�'a���pG����>��:$dj�Z��0�		�R*Q���tkY!:�h�TzZ��X�<�/��[��P5�祡�_�i���xA���<8,�28~�H�ގ�Fx�`?J����q��tG �ek��YK��7I�_/X�P {hD9C;�0�-����j4�O���&�?����p>�ft�E�L&��Q<YR�e9�p�^�wm�i�h�ݔ���p]�߽�11�y�KW�r-��>����k�w���!8X-�md�L���m�eU���^���N���h:���*u�H�S�x���h��蔾�N��x�P5�4
^�:n�ܽ���P���Ǜ����H��U}�Zli��׿��?��:I�8���k7y��ݝ��l�w��]�������~�d{T/���GF%�9���F"��Y��r�T���&cņ́����E�1��E�91��m�f��WĝN]����}
l�-�$n^4����e�=ݐɑ�/$� Y{[�}��=j��r�{����?G�������EM�X�Y����ǵ�O��_d>��D���v=�GmNo`��� i?�B�V��Cf����1}��>��j[�M,+�k��U5��ؓ-���<��"P0���x����9�� ���3� �m5��VeǇ�l�-�}�L���f��"�ϔC�C�g8e52FK�L���$9�\��Al/TEbMߪ�ȝ���8�u���;z���@�P�}�:��b�wI��������.�:��-�O�}�9T�������O��֞�g�46��`o�c(�u�T�}Al��]^,/��@�S�o���t@p��9e�3�Ec��n�J�!���by��#�F�ğ��fP�9G�,4Y\�!�{��ғ�z[�Z8)��s�d;�����0$c��������̏'�+z'Hx+�oR��t�;e4���들*DWd��x�ޓ�"��K~]���3Qx/^��Yk7h���^�y���$!�s�C�YO}es �sĲ/ϣ"��c�3�X�v�1?�*n�x����kg�i`~z0���&A
��4���N�b����T\�c��Έ�n���h�!�E�FTyf���8�b��__V�_@� �>9a/j�i�S8p�t$)�cڿ��Cs�KC,�S"r���r���x��,��i�ˏ&�W7��~�{[��[	��7�U0�7R��������� yI'�[?�oO��y�N~j`XH	�`��̿#�U�������B�*D	.��$m.%�>��q����<��2���FQn��l�i��Ӗ3c��#�~ό�^�l��� �l�����*���.��6�(�Ɔ8+O��Ū�םS�_nK������O	�%��KJ&jHh{~U���b����o�C�����$������qQ�]B���}7��͙��%�7v`�����1�6o��T�U(ϴ?Q&�;-۸���л�	ߞa�%��J;{=���-z0�i�H�:Q ���ǵ��+�	�(C�جѿ�$�2�Ӂ����W%%ӂ�ƨC�\�t}�~�Tj���Bw�j��uɖrW��Jд�4�h�h$�=fs����߷��r�Bn%�հ+�.$D�Y�w�Vq>�#E�[#9�I)�MS��Ȉ�SО��瀛Lڡ����`��j2Oz�w�/�]����r
��KZ��}���uo��N��:	:� �� �ҧ��A��&PN%�EZ_`G�_���y�8g�Q��6q"e�u��o�ȧEg+��W&2�$X$� j,�J�n�N�O��.�6���k�G��X|�������<no��ڎ��n�����v��#�"���)�۷hqB3ܪ�[Բ+���Oh�o��R�i÷��G����>�t�Z1�TQ�ů�-k���^�L^�2����eA�,�|������7|�y��dp�wp_q��F�Oa�����σO������,8}G���m��h�l��Kֈ�?o��Q�B���� ������y{c�ϩK�#���1�xMS
���|��+�����pNYw���	�sby�Ү�d�������p?��J�u�vRw�m�g�ɏ5uW��P�W�6:&��Q�0��-Q��E�"!o˯;�r�J��nzd�C��xi�"'��<,<�{Dn�(������%��
�o+�K����V�I��kfDen��vU��z�K^|�����p��5L��%�@Tr"��YL�Jxii�Ǔv�TL��$�t�4����8���2�p��B�_'�ȩ/9��6P��Fؙ�"?�.{�T�KG� ʦ�u2-��c-JFHҘx��qv�+�eU�xT-�ҧ�|N�Ś��9�dNۨ�a�M�{�� ��^?$i�>p���-L��*b�5�����_l��$���/�S����f1��N��Q�ym�i$B�A��~��-Um�}�ǫm�)^�H����,�9�F.�".,����Z���ݤ�":�4��ٶ�ɿ�鴁�sh�>�)USͫM��L xM�w$��P��v~�����L2�7� R�W,��E���������ԕ�����掚T�B�<���1E�^����\�̔�{��И�D�<��M.����[N���N$���y��K�Q_��𜊣�{M�bʎ&$�N�rK���	Z������G�4E�'PC��|D��*��J�}�>x9I���Op!X�M�xI����/�N��zPl�*{�ҡt7T�&��6�φ�C�NVˇ�c���W�/P,�����Wk%O�0o�=��wޤ5���/>������n���+���~d�`��.D�2��ZG:��(0ʮ�I��|yҨCK8�˖��9O��� ����c��v9�O8�8ڴ
ڴ�ڦ[�Ki_hg�h�L�S+U_��ά��h,/�m�p���V��j�P�4M��'lM��z������;H@p��1�8J&X�{�+��Vm��+(����;|�p�Z��]#�<����! ڨ���H�_,{��L�wcg��=b�� �c���cC�f��P٪B������ʠ�d�g�T1F�~<���6gM���b�L1K�8�o=�of�#_kt��
�ܛ�K�+V�&�Og�ß�F ��=F�?SN�o�œ�H}΃�GUd�$���#I_���j)#v�o��Dl ��w3�.��"�۝�������
�oQ��	��ղc�2D@�S7{\��S�)�2{�<�TK�LM�E:��3,"���ޖ�1�����T�ԃ��2�@�}k�(����Dx�H�U3ͭ5�}�ʛ�C�;ŋ9"����j�
����(��
d�2���q�@+c��>�d ��Z𮤀����fdN��:��|�Vǒ�څ~e����������+�U�OG^p��\l0�m���#�|V7���Q�P��&g��ke�ie�\�Ƙ�/�#�a�M1ȧ�jNU����>'1V0K�$�d�Oy���W�,<S� ��ĳ~ӗ��e�B:0��B߾0�lz\����������S~�5H����{v�+�#]�JS��5;!E
L�Ƃ���
���]W*w�f�ɟ<�t���e70"� J�TʼctF;]�(K�Gڧ]�Ƈa�]�TQH����q<��^�:;3�<w��5)�j2r�2�����g��״۾����9�t��t|��������"���Gq���/��n�DN�⾾�Tu�=zDo ��b��
�`L4��a��H`�=�nP���{�M���Y�.��X���%De��R�7C�����}�ӱ��b��ڱS�jD�Z3y��h� ��X�l*�����Q+�,�Nh���֙Y���VM��_`Y��b��m�Ex�L�W�-H�V��u)S��(uʙ�u�T�rY��lm�БΤ�� ��,o��wH�����b�\q��@$�G��_�N!%r�`��N��o�v=M{�?���]X�����4Eu���4'[���7;%>�����G�ne��n�qd
�C��zhK����S�(S;������ I��I�xS����Y�^���|b�$�&዗/���'p3�� �6Z�aOu����?n(�SLu�t��<��*X������i�
��[tyI�8z�d���N$6�R��e�$��CY�����.�����=B>��)zPzy�.�6��P�0'��bD�\H]�C���!����q�8��1k��̚�z�#�]/������([�x��'�[�|�T�B�a��(<���d�/L;_��Q�]�7�櫷�����%�i�� ���������?Ѥ���B�A�ӂl(R���IG�R���s�D���7|��~��6=��d|/2�>z+�����mKw������N7-�"0���[�1�h?��z8�1!l����Zv�gF�W_^�Ld��iq�xÞ����}���	G��a�L������M�E�h��X�^���$�]��F!��bO�Nc��^���ͅ6M��L��Z���y��X�|�9[�_��$	R�=��b�(u�A`ی46g�)RQ�%�Q����"m?W�+H����&bFɌ,�����ߦ^��Ɯ���� s���|�݈��!lH����q�o蠑�6�s���l4Q?�J:���[0e�7�`��q��1�`���Q�ձ�����lR��Q�p�%��B�|7��D�ы�TJŶHK�@�b�A�oe0�E��w�e6�3.{����@Kp���e誏 ��4�|�rZP�S��\ҽ��D��B0J����乇`nV�<� �?�DX�}�����@f���/ّ�,��y�`�@V�xIB��d�
��^|��\����I�Jq񙵉����[%�ܰwj�e2�H�v��;^{�����{�
.����(f���nC�~d(�)�.EY�
C��^;��ɩ�m�AM~�/��s/��hI��]�K���5�WU�(6��V5b��'�R7C�ҟ/�W�Ï��g�|��b����<���Ɏ�6�ŭa��f���+�������*1S ��*ƫ/���@v��������l�D!���ҁa*�T����/��FF��{���t�n�D��z����4w���_~��"����yh˕���/l��>C����O|�ʆKNqu�fH��C�����)Y9�

?u�S��RI|W#nm�����`u~��j�Oq.�WD��e���H��P������PK�o�P���4'����GM��ۋH�n��9������2z���15׺:��g��g��D�>YK�k�n��"~�/�(�q�.�H�=��:#�X�d�s��t�1'2'��<�N��"�q�y�)v�l������V�é�P���~s1H��o�V�@�ѵBw/ن��zJ-�#�)�U�7"B�Ue<�P�h�NK�S��,��t�o؊����GT�L�>s�ؿ���d����j�gڎ���O���K9pХ���Чd��fQy=JUъ�(�3Q���̞#뚅9f�
dʑ�ν�%����u�Tz�3/����x�&
�6��t{�R�1�6?�N��AJ��i�iM+�@9��I,�`(� ~ǧ˺˕��ن#v��Ͱ�U����@p}yp*F�@O��O԰bԋIË��Xx�bl�0*����g�dXi~�� ���a[��P�ڢb����s��<�.��!&��|���Y$���A�+��9�R�a�m~��ͱ~����U;�������IR���m-�l�P������:��� ��-K�w (]�CsM`�[*"������5��:��喵�X��m�x݋�%@z�pcx�]�_`�����0�0�h�OB�&��'�����^�[6�K��-��]K ԍ�XF�]ot����1SI�Zz��u�Gǻ`�W�J>��e��Y�D�g�B��П.0�SL?,@_��72�^����-1o��-��k�����q�yN�@����x�$��f&t6uw)gm)�h����	b�k+h�q!��9c�^�-��;fS����e,xQ�b�)�o'��Z,ަ�h����ǅ�_eT��z|�r�ZM��͢x�NA{�")�yqn�}��M�)�O*5Da��}`I�L�0�~J�VrI*�qa�\�^r�po���U�*�d�!rz�zR���n)Z���o9�����}��}���Jjj' ����x�]�Xzz���&��򲚼:WYE��Uŀ�I�i�B(�Ќ;�̳Q3�Zy�?�s6���}i��\�(��҈��9ۧD�h��9(�����tɾ=}}xT�-�$��E��ƚn�V��v)�or� �� �9vSN�C�>Qc�}�����E2��ȡ��G���mm(~��	����>�K����6<� �����S&�7»kK3Hw)�H�M9��P�k��D�1���Z3�4��iӼp~o@�򇣵�HC��� ������ᶛ� \v��E�28,��]�{
>�h.�G�_��aa n��* Sc�i�"�ju�J|����&����Y���z���%S�{M�c�|�I�o���������u�Lv/��7W������L����Ƶ3����n��nAw���Z�^�1��E��
zt<�Ii}ƩL)�F)l�;6��2hz'~k�VǹS�u��e���@zF�7�Q$�a�갨tƌ��&<)]�ҁ��O~5�E|>�7^�Q�b���^�B�+H�:"��"M�j�8��I=G�l�di�Ob"� }���]�J<us�K/��[Z.�N�gqb]�����O���u&�ђ+΢�J��J�f�Ж� C�[����zr��*31���##Ӈ���~3�+o���0q./�]�)�˴�K|s�ǮɇO4i�/[�������5��Һ���x\�����'\��;��\mnaM�����6HU��>�- ��_��3��L���N7z8����I���q����wݧCk�8��k��D�(��8Vj�|e%x���-/Z+f�i��f���x{���PO.K��D�Kvj[Ŷ��]��4]rX�v��t��,.�E�(�֬*b�c��LT���gG�㛖D�G�y䶆�p/��͂�`x�Wqh��K8�8H�en�24E�j//kOM���	���>+ٺϝ����Hߪ�6�>�dw䶘����ژHu�,g(d�GQȸ{{hr��"
��~���إc���.�S�2�ͩ�����D��̼7��d�]��������5Ǽ�M�%�=��HE��� z����p�`�z��n�*k8�n����ӡp�*w�I�~$���FKq�YJ-V�y��$�ap��K̋����%�d�̯�4Dȿ'��*�2��X�g!`��������e<��ɾЌ4�D��&B��a�S�&"Í`����[z��f�"FG�_lK�=Eq��o2�D�RJ]ͩ���V��!�����H�D�]��aiZ6���l�a�ǭ���[�9%�������M��Jx���ad�eO	~��q��*���l'bs�<����ZX�}�*��B���ԉC�ȇ�-9U@!����@ȍ�ޮɩC���sT��ܟ%��=����ϼan���U+�l�>�ׅH}�ǘ�S06������t���hwֻ��>�6��_-�������\g6�x���w4!e�!-ً�uOBM�:�Dcɠ���{�8��#<�#��!�Ȥ*,u�p������)�u1S[�_[K��O��0�7t�8��_i,\<+��,�}t�ˈ�8!���E��DH�TsƂI�rP^#�c��Q0�ː��4%���e�������wg����Ӵ�Qy|�;6��r����B�m�L���W�碹D>���bp/?��q�HrNN!�4A~��m��ߌ��������G����wsK&{6�1AO�]4��g�E;|8��7��3�����;^��&X8��j��Z��ZL���*`ri9��)���%YjD#���'�u"���GQk���CS����� A��-o>�u���t=H*c��,y��i�͵Vj�:���n~�ee�G4FԱ���~���QR��=8�jk���ߤ��ˈƿ�
:vi�,
��#Q:��K+�KgC*n�`�$
`#�@8I3�x�BI���)h}�}��c5��)!�F8���8�L��	�D>c1?D���	�j��!�OJ\�Y?�>N�D�^�=����l�k��RzB $�2��Xm�'{����Y3:��L��Wg�)J�)Z�U�m���O����vB#>|�>R�s�̿܅�A�C8o�t[?_�@��ԇ��b�Y��{+.�'��Ǵί����,T���P�4����7lY��	�0���A��+�M��J���>
��xQU�%)U��8xS�2]�J9f�ģ|��qJ�������/#��
�I�Ű��Òq��6;�ܣ��)�Fg��?/��]T@���
P��U�r-=�n��ֿaKFi��ַ[�w�1�=Q]\�]|vD9��;�����L�����T���o��{LfB�R%+�h7���-t션ǝ�$I�+����N�Gb�?��0�F���I�p��vt}0��ƨH�Gb�\���7��by��써�rJI���/�LLk�L-�M��L+�L����3?{�(
�1k�6��6|<~���O������͝��^�ܞ����˝�A�2�md�ݓ� F!��'e��t��Zш,`�ԜP#��E>Y'�����	W�;=Q���S��J���E�׮��1s���y"Vr�?$����}��;b��~�? ��K2C|��P��5��g��xH��-�l}!w�"+�T�&� ��O��7kn�+������P���z*_���(`,����P꒝�/̆!����لn���j²L%�[d�^��Z�I:���5��M�<5���I��G�0����@��U]��0gڐ �w���Z�-�����P�%+�� �J��y�E��}?�ެ"�Ʊ�;5��,9-������Cj(vT�M��Fτ�f���}2�"�n��v$�wՈ?ZG�f����]K�3���`���O�� �.ɷ3фq�h�;��{��}����p��@ٓ)Eb�܇�+����gag<�
��Z��J5�2���;���"��;fD_����Op�}H��t�F׫�n�y��y�����&�X!��ǥa��2:�="�D����k�s;��y�fD�(�ب�"��7��htU�誧�(%�M�M�>M��x���byw�\��?4����b|����3g{�uۘ��jv�AUVí�hT�#h������ކ����b�ʛ�Z(k������t�xy%솛��#M�?���|�M�}����=%�ƅh=�>��`��"����F^�w���P\��P�o=X����Za�*:�����g���:
��o� V����V�M9��<����e�K_ȳ�d`��}��G�"/���*�Nv~�؅*�F]
'�����!LF4w3d�=�u_M��%�1������J����o��^~�QgH�`�E]'�9�Y�Gv
����S�<�}��I��	:u��-8ؾ����a�Q�-<>ja��ic��:�U?�����x�g���TH1ڴ`�^(���p��|X4�N.�(��}�ʽsԸ&k!NtjD�QD�A��RrVTf����8XDb@ߎtE���� �Ɇ;�O!_���������J�%��I;�;��ݑ�'#Q�R�w���ɥO.�[.�z+��n���oH�rZ�X�E�[y�mZS&QJ��E6'Փ�g��Ck!�A��%���t���F�=�I&�5x5��KĖ�`�}"W�� O�vX�b������ĞJN��W�'g>ҫ�*�W'%8���k����G��:c�Yf�����_�j;�P
دh�"���y"�L�9�q�B)����"ojuv���%dT����0R�BaiFo3��j��n��e�b�7kO�o�Ge`����3�z5ַ*Ң�Ix�L�
�?#�=�����tәb��\n�����}4M�y}��dKb��s�S���gg��Nˏk��ѹ�=k�%� �WK���3�9Ie�,J��%1�+��̓	����>�#��JUQM�����!D��N�+�l�0��+�� ��a�n�V�7�/�]$�Eǯ�لV�c��[(B��,X��u�6^F�X�v/�FO�Yv�$/P%~�gL<���-6�-~ҙX������^�dH<��5�b�*`�\g����9���f��7�.��o��ԛ�����@�ʛl�ô���e[�q�׃>"K5��|��ol��?����8�Z(N�:ڊ��U��.����L��O3�&��:����Gy�V_?Z�%�^�=�������XD��bGc�u�g,�
�_5��$@Or�=���R�<�#�`5-���+yhw��[�_~~�F���q�vl�H���Ku��Tw�B>[��GP�VyŪo���!���*��T>S	i�Ё�Ee.km�>Û��Ĥ���e(�[���-\�,�,���to&�{	�s��}��2h��R�&xo��味&X�3�dc���Hal�/�ә�i�U��v�N����2�uo����DRkƫ/nY��ȴ���{�"z�~�|2��񯗏r���3qϚ7�q���Gk�#o�y^9��ؐ�+}mx2�A,uK}$x�Ǵ��O.>\��� WҬS�,�?����F�5=&��B�I[h�r#�K�6�����G��{��^���l3����K.�c��<�'�1��F\��{��!r&�SR�>-�P�჊�@��7���_�oy����r��1/�6��=ԂE�=���*��pzv��_̪���	ߺ������T����~��e�a���X�"���T;�P0eRp�@��k��;{91*�[���c!^���+1�D�h�>���^���6��O�e�{95�gE7^�\�+/f3�U�#%$$\Q��QG6��+����CjM�e}��B��x�M�i�ؤ�8(@0&��� �b*2(F�������;X��t����s7�cq��B�>�%Cz��}%�F��u2"a2��y�
6-�c8^7U Q�kWt�L[ajW���wh�<y�5a����(<b?=U���xI!����2���*ť��M��Ç˦!;[f����gB��#���JS[�[e�s#cX�t~��Q�T�bF�6i��<�!�S��T1�`�c���3���;��rQ#�I����	�^�������r�uw����%
rŉ��)�`��+��A�E>%�Cs	V�_����-�*����)E7S�o��̈�����s��ic�c��G<���� p*�n\�n�Z��E�C�t��`�@y�$o�$��idK���
zIq\+���d6��A�{p�99�	���3c�"+��7�3,c�K�~��~���v�c��m�+�Q�n�2sU�&Ru?3c�SS}87�ߵr���9�?`��f���A�[.wB��6���d7'�8nA/���xp(<	��E2�D����|%D�X���|�����ً,�8m��#����vTmיYjMNj�ixp����f���%���kkeR���
cI'���C��W���k4NQ�iG����(8��pO�o��,��vy�`v֒u��g����ӌ�o�%_�����j������Mӑ�C��ֽ,!��A���xZ����CW�=n���:[�����s��{n]���CE�rS!!�x�\�L��Z�7,jH
�c�x$���糎0ޫz��c���~��x]EpAH�����b{������#?/\��4%��C�
_[�`/E�Q�v�J�J��g��ƛ���&=��:�J��^�>�)x�����n>~�:�=}*D��S�ѡj�?ʾ��,~h�A3�m_f�����r�qƻ�����)c�W�k�B79 ��M�t)�H�ºZ�"��,��.����y�{^-ޖ�G�A�q�K���:j��Q��yܯ�����>_�_��M�=�t�f���<�-L�`�.��I�YL�DD�e��T���
S��7!�c[n����}����M�����V��y,t��~�֠�I�WI���-n�}�=jg�t�`�haR ;�GU�OU�aE<��鼖�
z�ˬ(��v@�:+h����D�;>a<9m>>e�6�0����Z3_��L��W�_��A�QBJP���T��Cj��%DB$��k`�����K�C:.���{����9������lΤN@ !U�[l���ҵK�U�_x��>��q���@𝬷氡�Ni)��(1C��t��e;���7V"=Yu65�Z\��0�'0�)�TE�@����
L�Y�"[�M�$�0�b�{b>xF8tMb�R��w`��V���g���`���g��s�Z���z��Qr�j�e�1H��E�vy0i��KDɯ����e,���r��1eM�zT|n����5TC2z�O�b�<�!�NUvB�!N"�B)��=����}xug#��$B`�ԮU0��7��Zx��JM?"c<Ḧ́�پ
׾*<`]wL�4wg���ue�Mx���0���ٹ��x߀�H���΀L�'�r{�V�s�˵DODBDBm�{����R�qp3��>��>#GTܗNy��]d��
̪��K�)x2܊�30_5�`�uN���DƬ�1�0�&��^�)�8B}n7b��}��Nܼ-]�U]�^ߨ�5��� e�H���Hf���m���C�qLYm"e{���x��.E8�)7)X������?S&��&KP�6%�V��Qm�S��nuT~%��m�/��+m�������(à�[nt��ZQ6y�� y�6�r���5�%�|h.҆���kg�Hp��[�T��V�о#Km�h�\pt��_<v����Z��h� �3�.��0����X"�L(��w�;R��ċ� �&lK]�r�_ź��@��V�A )%X�"t`���e�;�2e�T׹f���9��7n�0U���:N ���0cL�|���2fN��R�90�6
��}b0��	O�blz!��7�?3�d��l���b�q����v�u
j��&\�tED�`S���L�0��3�65�)��OL��	�nL��Y�zZ��Yl~��y�����z�U�v�Jdf��^�l�Ce2`/��j�?ݾ|v�F�J̏�q����[�љ>�]������}:����L�-.)	�7�|#N��m5%VE��#�An �"}�K,hG�z)R����O8���	�x�p���%�`?����]4�������ݟ�f�not��,`m΁�tb̴�e�g($>� �h���	��\>���Zc�!s;�<�a�O�%%�3�h�$ѭ�6����}��`��y�B��qw��n��48�S��������}[���� � � ~A�}q�k�Ry�|���:�0�5��9Ų(Pd<����U����X�W����ϵC�'�P�~�kl&g'���^��M���<�������$ )Q��0[QP�e2��8L9��'�;RQ����p��rQ�e;ô�P $sj��p� �J���l�i����@ww�Uũ�i�Q9�C�Iݗ�� ��ʩ�J��3� %G�������� ����/�1q`� ��kC�)+�iQE?�f8C��={=��兑�PH#�YM��i��(�5�`�Yj/eH�h��ʌ�����+�H��s��4���۽Eft�0P���Tp/Lx]��IM��¬&��/�"xNW��J�)�!�2�7�+��k2tV������@�.�'��t�e-K�&BD��A�i���.%�%Hɼ�����?�|EJQbU�*i��,�ݺ)�f�*@�@��Y5�Ac�r̥�,�#�7(�˙J��%��}��蚜LMk�9^>��=��#}���U��q,�oG̨�s����h 'j���;��V��}zߘ�+����?��!C"I�h`� 
~�̎z�(��>����5Gh�(��'���Ǆ�l�!�E�������FϮU�[��Z����OcHR��ܘ�o����'ͻ��:�M�
�AM�|C=��jL���z�;a�'��>�&ā̶��jLO�yT�p
��(�x���������9�F��4�*�ůN�|+m�髃�q��t0��QDT�a^�E{o��[�,�6����&=��f��wܱ~.�-��ߌ�l+(��7D�Wk�L���h�F&�J$�xXW{��vL��I'����o� r�wTx`Jb$7u���Oo9a�,�yM�]o<ہ����>������*st
	�'�M"����*hvH�ٳxk�n�EX��I=�ٷ�ذ*[~�RM�e�fO깥f;��?�#�+!3{R�	]��ka�?�5���Q�j�����AIu��|K��ȯ,�5�SBaM�2z�ƍ�kw�협o�ɩ���u�o�.�)�l�ޏ�Nʏ����[���0���jw����\hۤ�84�8�V��E�l�`!�s�9���%Se	���ڢ�D�%����ʜ#� <z����V��bk��Ne|9��S$Vg�%CNܕSDNq�j-F�1�l.��]��2��(���~%Ø�O���9J?��Iy-��kV8�D�&�"�#U:�`��>,oV[v�Yw����̊2�i��
߬�������L����	�q�fY|��Ps�:US� ���^��q����	������7ѦcW{e3lUt-P&���8\�ߨ�#K�?[��Ik�<=�c#���*'矋Lf�S9BK?���DU�#Z��/�)����Y�N�)M�+a]���N��^���]T�yws�T�[mB��w�unXS&� ʪ����� ����dv�����V3&h�.�-���:���A�W�B�1�8v��TTL)�Ԕ��ڗ,��7�s4QZ7�Є�ˬ��{�`�m%�[�I:�*u{��-�Y�}آz1x�>�]��ހ��ع&�i$���*����E%�IR��3��\�O+X?��:3Q�N�i��87��$S4̀��vՔbt�;@��F��C�ڟ�N<#Zn\�����k�.,�(n�(�@J̮�unkݜ)��IA��g��ڡ]����ٟ�����������د�T��ِ=��A�&ٷ��K�,r/�w(N�ekz�����ɍ�w�a����8�κŢ����0��ynD��G��i�·{�Q�/�i�i��7��F�_]�d�^AA��a��N$�&"Z���g��Q�?H�'����-��p���t�r50��Tr��e+�p3l��8%I��:�d�J�@u�륥A2� �� �Eʒ�����E��%��3�čL�
��
�/�k��M�4�yl�~�7�����:�!��6���L����K>�/K8�"&�4J�JG}GĩGq�>�vvI1��\�w����}�( dgBA���V9\����)ܝ�9�ikf�C�u���	���.���t�������Ϡd�l؜f�[����戸��OMA3�aq,]��t�X�#���0s�6W�6f�C�9�B�f��1k�L4�r���Y��U��o��w3<t��������<���%��W��K���]S�&����`q)>g�Y�"A�f0�C<��=Ђ��I�����2�v />�W��[���G����"�)�P5��g+Dm��+M�y^$��|Z.�kQ�nS��Z�ZgŕR�7JA��M2�sO��g��:�&P#��򖐵i];�c�{S|�f��.������°��T����ޣ��f��"�<ڵ~?t��6|ǳ(��?K暏�:��hOK���/�س`޶@�Y�oYe���ʼ7��2Ի��+v������	�Q���<����� ��ۣ�r��
-�}�$8r1=�Gkڟ.u3��@yJ*����=u8V����I���t&�a��ӟ��������+[{�8O�q�ͷ�t���9-����3�WU��c�$�83�sF"�CF^����%������]X�`�#�_a#�3_�'K�`�btF��L�y��'r:�݉Z\P�hzW�ST#�T2������N�˧�hr��ܷ~�uj��0:�O����8�o�~�n8���G���Y�_ �l�B�+X�#U����\,�Ϙ���JZ���f��0,�&������qc���@V�N�Q��������']�G��;_��T�z���C�LB&�s�a�M�jl����	2�����3{k�^\� ���R���5F?cA�9�mK(�J,Pp�R�o�66*� ����݅��!��?wl1���Ȳ8#���ѯ؂<.�+3�W1*u>��l,\�3�x��y���?A9=E91���H�2uTr�4�4���j_j&�a^����+�'^ "^�	���p��@z��\{�/����o���og���>#3��l��/s��K�~���)RYe��r��B1-�
j�&��^Xe�h�_���#Bb�!�XK�vd�Yb��)�E���H����aJ�J%c��Ӡx��1���*%�����f�)MI�OjȆ�)�PDQ�W ���?�Q2�j6(��~�ҏ���u��%CI����SGɳ�1��2�ť���L��˧I�I��%B�!�}F� 餰 w�7!��UKZkh�8��D������I�v�g�;}M0��#�A�E����|��E�ⱻi�~
��Z�ڝ��" �[n�J��e��z�y�y���uF�����u�_���x�
�}�Y.�Zf��
��Y�@2�`�rp<�Q�D���"{�+�����_��W}�I1c�3Ѵ!��>w��BgS�s0<I:i�w@�n�2u�i/�=,�Y�L�9���p��b��hm�L�d�ٙuom☡�Rt�9K���MU���)���j�n��ݢ;��;��%�ϕ~йw(3��tط���W獉�z����_�:�<�Q����Nn��+��9(�C\�ԧq�Y�:���|W�u[��f�\�P��{{�.(�T�뎅J�Q�O���y�+w��#��n�f��
�M6f���f��^�Tcp�٬�o/p�0Q�u�	��D�?�H@��(2�)H���o19E��g�s�ئQ�:�i�AU4��y5�ڨz�y��r-1�2��|m]�M�ᡇ�)v�"챯-�B���ِ��*G����K����j]���-}QY�pR��GP&�#�=��\���pe�Ⱦ�8��:K�z2��C��ʿ�a��a����e�vM����4�����9-y�/ޮ�x��6�e-}��}u\��׾�JCY3UT~�g��b��?����h>P���Mw'٣8� �0�s��L|����i�PCH#���r�=�+(�O`\��e�t�BFʱ��	����c�=`a8�	~*5�ugW6�^;$��8@C�F�د!��X�ָ�������G��(�[�����,ȍD����znzm.��$۸�W�jزO���6kz;Wߎ��y�����[y_B�Z>w����vǬ�S�Z��ֽ�6����s�6�2���i˚�Y+f}��N�[.�r:d`�>�|�sٓ�P|yu:7-��x�On��y��H}��8�p�h���C�@c�}8��<�zj�Z9d&���y˨�b8Up�!�墰lE�;�|�˟[��3���FJ��U�u��YI�&ۇn�`<���z��z�"�V
X<�
8ty� K��%H9Q<������A�F�z��E[���g*�ZI����W�N�����	ڙ\`v��H�Ȱ��Wo�N��<x؂|�}�i@�7/�}A�"ķO��XHf9'��8U�O^�xޡ��(I�蠴p�~!9a���T'���ވ��������U��H��?�����E�D��_�]f�b�����ՅN9�8��ƌz֭� ��(�5�K9�[]o�LQ�k�p�vT
�j�������:�H�L�#�J>��.���)C�OQD�痪y�č�A1���č�O�j�aaG"D;�$��
��z[pgcz̳�V;۳�37�xfc�
V���b��y�j_��ƽ��z�~݁K���Q�tUʟ��}����EE�,<5;EɯX�B�� �yR �/f��/_~��cxTv�Zj��MO!�.Uҝ�ݝzW`����������b��������{O{�j��»>�=U�B�u��F�g�F��.���yg���>UI�|� �~�V�XoE�ʛH�}I腅�)�Q���|�فAӍa�D-|�;�9��A��Cg�c2hr�l�UHJ#���:ԯ���x�^y�l�ぃI�0�@viMuk�0[~�Z�	��#�S��(���o2�����t���,����.�v�6�%U3f2�g5��"G3*�c��o����4d~���䶤f�7"�hI|�G��nl) X;�P�'���S[��0;%Wa�%�G&0�}&j������gn;����r����4�&��E����ó��	o�Mϩ󋽔����U�Ŀ��������;%86J�ޱ�NU�U~���N����F������!Px�0a��Ѳ���pP(D�Y�<;z։�փ�|�=�I��P�&�Q��ᇀ"0�����!l���[ȳ7:a;1v8*�_ɯ���י�J[�P������6	��+�H���d�������0&c"}�� L��Ŵ���s0ߨ�Ĥ��pNM�O>A���g;̥�B���Ɣ[o�w}�w9�sn����V�7n5wu�u�%�P�!59��:�jT�P���[�LTu0����&R��c��?cr�0�~���B!��S�y2Kl�xl�3癛#�_*ɹ�
F��Y��L��tK��T����7��pV��u*�x�I/oSf���D��-��c�����z��R��Q���<A �P1�����/(�E�q�s��֒1��Z�E&�A�,+Ǌ���&���ЖpC?���&cc�l7�t��6��8����YëٺԆ�7��#��.����ޱ����y��~����kFZ���\��R�  C7�P�=˂-��g�Y[E�o8�Y�n�(�{���r�th�դlPW��R��$X�>���]��.�ɓV�u`��d�Mؒ ���">��UB@5��ЧyS�^��*�}�]��U7�,(g�Hz�,��������<��l�E��Ⱦ�ux��;�ڮ�0�W�(��6y�,�7xh�8�mZ��7{�d�*��8�mG�����$@l4z�vR4Y���rL,���)3����U�8����^4���F�7q��{?Qq-�|���3��S�&���fI<+?\�Q�4�BFq��܍c������D�^���܈Jg�ANf�J�P�)�T&�k�̷r��G�h��Dw�`�%��M ����e��M+���{!a-2��u����%sz=ΠtT "�k�.JDʤ�<���Js�]Ƚ��$eHa�Ĕ��Ľ_�A��y �c��J��j�/E��XV1[fͶ��ٽ�%ԡDK0��$�Oߖ�
(FG�����x�����)�8�_���>�1���1/���=��K ��e`2��0�v;�o����l�Ӡ�
!ϙiKP�Y_�Y�q����UYj���YM2n?_w�>�_�^���Z֐��^�C�@h�雼x�����I\�2��1 O�˞�Wl��v��_f'�1ɑ]^6���z]#t�GWX-Y*^'�m��-3��L����~g�ˢ���#�_��v��P$���F�/���畝@抠�H��x����EyIk��Z��*3�4�)�Ŷw���d�c�Q��|��g$�.�|O�&s��S��wdx����2���7�PWoQ|��ә5�� ������@U�FA ��F���J.P�����Ř�����jn~�o��j�]EP�Q�����W�3cp]�<O?�M�u��P�;UL�L����1b�?q�6�k$���NI�7@��JU����[�j���ն���T�k/�����a��u�.�9x.�/Stm��7}=���1�������g{�����k�=��uA�e�����?.����`g_�.u���Y_-��rOt��5��K
POO�LN�
"��Fi&�Q��k����A�ƴ����a�H�N�d���:i��»�0(m;4����~;�^�]3�$�_�7=7n�!�2��C3����2���[���)�D�zMI�C@/�PfM��W�-]�����'FT�RT�%q���n�Q+6{��#]	X���ޭ���g1��`�h#��Z�#�ȇ���SU�@=℀���	��~������f��󢧔�;��۳"�&��,�E�㙡����վ��TXeY�̚�E���C� �gYۿ��A����{�����@����������A(k�����2�nE#&23��;Lmdr�Q�aѼ5c�k�_|�cNH����;��Q30�����a˘�0���8�gB?iS41��.��R�H� 7�`�r�B��Em�t��:ɇ����(�Pr'�8��^C��Jk�NĲg��Ja�m���$�p���CJ���KJ�g�t��&���~����V%]��v��vԟg���P['��"����#��RV���	鱊�۷�_1�Է����w��朑��M=��Y������j�xk�/(���������| {V�������mg�+�>-��~,3ѵ�^�n�����!�
{�:J�1��E�rM?���ďq�ו�:g�x]��cݦ]b�]δf��ʁ�
f����V4,��w2����)�"�^*gS������o��ɣ.ν�0��޵�.z��CO���n��S��.���k���W��"��s�<����`��<�m�5�EKƋ���6��6�i�ze�E�Vuf�T��L�q�4,��T�M&���a���Ѹ�?1��[�9�ڬ!:6K�1,(��dZ�D3q�sq�7��/}�6�������?�l����B�%U���&����Y>1 ��2�5幤e=�����p���zѶM�uC仯��dH�|�o�m�.�_�&�2/B���C��TŐEŐT|�t������ZaC`��XӒ˰��n;�.�����-â��fr�;��0��@�I�#u��=��A7s-3�n8fwA=&�sփM����iRڕ�T�̓N�$+j��D�i�'L@���?��*���)����U�N;��f����jzV���ȕ�����E�Ɵ�+�8�%��Y9"M�X�(6A�ؚ��o4�,QF6QS���1��J�X�`ϋ!�d�s{�d����VHEUDIYH�[�*�
�t���;U�äc:�#��G�}�� ��o��c�=�������S^��Z��7�%�VRÈ���3܁�ʌ��zJ��۩?6���Rj>K5�eY����%MÉ�"I��~�4�]�bR�N��)�4c� eL�a<�/���pU2�-H}EJ��=#�5@�ں��lQEŇ�E?4�pt9/@gl�P T�pF�0���[DX�F�B�
U_{����������7T|�!�~���\�̽�|����ᶾ�������tܫR"�N�)������ܺ�����Q��^K�����]4����`:#Y28W�� s�zg���-�H���������V���ι�k�_�j��:c���$�J�v-r����~GogFy��_�kj������M��z@Y65���_�^\��N-�����*1O�/�?\E�%�e��s���f1��y��å߮�L,��*��
ۊ(T`�h:�a��������_�!~�X3a
��	�
:�;�ݦWB�s�h}�=�[�뺣#}�8��E����������)Z���A���b��2�Ͻ�p�
hWQU�%f�$���_��} 3�!��9��MJ� g�߱���X J�ʍO}z�!�or���B����*�l}���F���i{}�2�{E,�e�6��+C%W_�`��ז�y����=R���*��L�dʞ��ǧ����q��8I��]㉿�%./~7|����i�-�uֲ7�9��#�&��tn�蚴��lZ`��ѓ��{���(��}��b�����D\�V��e�U�A�x��B��:M���^�+aq��?6����p'O	& ���cS�/f���6��g�U����@����d�E�S�'��$�R��pֵ�-5��և��_,&��^U�2��2����PS�S����Nψ�7�~��T���CL1���ۚ����r�����y(j5YM�G��T�f�Q����w�щ65�#��;�r1Y�U��r�\mIʟu'��Ş�����7m�p�!-U��_����! y�$�k���9���΍���&��&)Ɗ
:E{�@3����	t"���7���-�c!��	�"������#�w*�7dH��ac�w������ࡲO(����^�,���?�?6nm #���)���xշ�ނ������6D��v��(�|u7�[�DJ:z	�w���>��mD�GC�8�@	g��w��+hC��r���5_�d<P�@C��q-��J��L�{x����ZF��_t��J��T����� �XWh)��l���O��7�����c&�ޗ����6�[��*u��r'�`>ݿ8��nǼ^��N�B꣌��p���)t�؛�8�ȩQ�{i��z[�<�O�����X�/�C<쫎W�f��/�Kؑ�Z��Fk�Y�-�ޛ3eI/�D�Ng'�3�O��ɟ~^�C���YUeh9�9R2]����0�;�˛`!qȧ��ۅ��R>�t�	���"���U|`�W�˱�mڗ�M����4�櫣W���Q-�T������i�޺m?g�G|�p�(�ctS�:r?��1G)��17�"ϧ�2 7�^����7.�3��b��[x�[�I���z�5�3W,;g4g�]ٲl�=�����rʦ�HYݣd�����R�n~�W�q�s/�/�O��%?K�H�����N�%��IH��!2wɼ�����ӣ�Ȭ;@z��~(yLW�4*#~�S�;h`kN�hM�w���
p�n(>.���%�5;�&1��7dS{�@�%C.����M�����xA��i�����l,,z%����W[�O{�BCN��Χ�'>n�|/YZ˧�FՉ X��,{^_�$�����&�X�'�S�?f]�f�mPKh>8�{?��s8Ez�&c��8d�@�Z:V�Ef�x�	�E2��B�[K����ת�܍�R<"�^7=����Pe��qZh�^|�~� �����l�{Fx0f`]V�0��Q���AcJ�)vA�a~�J�����4�>�t�J-8��;�~��P��с�:�����Ld��+�b��j�h.~��s⯑����;��;n�U���UlU��#��R�c���W3kU?b�l�o/W��Խn�Ӛ�6��9[��g'#��"-��]g=g2������~ϳ�c2N�Ӧ��0U��P���`��T���W����^0X E_���O:�����w�q�*y��b!�b�@�q�y�?���.�#W�=��A@�ݡ��Y�o���H�rZ�Og%�'#U����bb�I�v����q�l�+z����i#FG�(�+��z�%3"�'����l��<9	δ`�j�vO�W�%�Q(��UP�y��BS�(p���i�h��Jϣ#�g�=�#f9���R�j��9hc72�^X2���9W�{+�Z]��huu5D�������jr��}����3��5V�<��]��f��%^!��&�z�Wz�"���om���6}@fުf�otLO7����g���9�܈""ITK��=�~dx�vT�?C�>��7D"��g̦A����o�����<�m�?����Ǒ�}��[���-�@#�0z�@�@�}�`��`�ڹà����,+m/]MEu4��U�B����}
�e>lb�T������>���*��iie�Z�?b[*B.kN��_�ٿ鿄��f�u�U� ��
ζ��`S_p�\�y5hȲF��͒��/�p3R��D�C�m�.ۨ��\=*k���&������e�U�`�Y��>eš��� ��>|ȆcRQp]�jƌ�-CK�K�-��b�43���R����d���co|�R)���*��4e`��Wy ���^D�J�k�fx��]�@�]޸� �{�G�R�0���.��������@����9��vC?\��T&;�p�gV_BH���R����0�V�dް
΋�����2����>�5�)�� z+L"hm���P�X��͟ x,Έ���D@Z٬_n��rY}B�TeW�`��<�鴙����Y��ZN_{"<P������\��`�/X�)���+NsI#��O��S���K�R���pD�4�Ar�&�h�h��LeK��S:�])2fX�i��'�#�����*�4�r�	�-��
t�pKG j��l9C�,���g3`��|]5t�7�����&�n2��ʗ�%-���di+��+}?��>������+E �A5;"&Bn��7]�cP�)�v(r#�埐�)��X�7�����d�z:��sCo;o���3M1K��H�G��<r��G��r��-��bAEaQn���+�8�Ew���>X��	-��pl���a�vR�N� �P��U�V�:ڄ;G�{1�Jn��n�kv�
mLىt�L<�~��UfgGN8p�ŶMU�
*�h+������z��	ʸE���W��N�ϱ��ЮP�7T�߂���,8l���tI�՗ �a�[�zeE�@nt���^9>�@��쿤�7 A�EtZ�A}:����P<#�Q��ӓTL�YW^@G�F��S��d��h@��7�ʨy޸-K=(�Y=����]٣�Z�<�y(�B%v��S� a�%�\��y�q�R��W�JZgh�P z�>�ߘ��9ǫ�RR�%��5_0����x#d��	,��(�{�-�5�&zy�p��v���{�^!X�i�O��Ǻ_�_(L�$:{n�JI�r��*m�%�za�NL�Ɗ�ç��le�q��_��6��̡ѭP�������y;!��ݫQq��ͺI���46�k��Ӌ0,�{�C�~���PT���zD��Z����w$^�w�!�+D���t?Y~ē˅�|͎��y�'
�{��GbB�jG��2� ����'zcʻ��i�BtU�+�M��D��[�X�C�����6X���:�����*��:�t':�� ��
���⼊��7�SA��K����^����4aǻ�մ��l5k��U�z�t�5�N��kɫ9a/K�5̕���.��ͣ;�^|��19��e��f�}���>���Ԉ����x˫�6tց>��L���~�^���{M���Ɖ��4|y�1���=�>c��B
��P�#���_�	o_0�|g�9�m��.Λ��.��߅l�Q��N���>�4�	�y:�_�8�Ol#�r��S�����j��#�r�4?ú�8̒�>X�������7��h��e�:���)��'���Ő��3x�u39����7桩�k2�Ä��"G�[pxM]�����0��ٸ�4��n���.y�����=�5pH� �p��#��JFc6��'a ?
Q���#Xe��$��@{�	=�HC92�����dX�WM�t�1��f��g�b��~ۯ�-�P(�8q��|�P��䧙�F��4�I?�1C (��T���d����r�J#%�5|�)��'ɰ��~ f]C��GXY�q}ˀ_��1���oPn��"6������c*8�b�V���8�H�m5�N�GP��8�)9��T"�6?�jZ/۩��8o�����=ew09��2Z�D.&�^9��T+
�NpU-�6������P��؎��Esi���c��^�[��J�y7��0��do}�/�m8�%w��7o����ud�i�!A�����~�� ��o����K���f�C��;~��4�<į&��\Ԉ�J�w]���W`ɿLZ��N�Og�$���_+�qn�(F�}z[;7t���Re�C�C5#r���h��}Ӷ��N�W.��f��8�ܾ�-����+Te
�fr���4���t���cH��Z>˧b�<�+��#�
�[YƂ����՗xs&�i���Xs��-����h���x����~o|�Ӻ�-A�"��F0�>.E^I��Lo�R������U,���Q��R�O��ך{t<�jhڡ]����њ�UbU0������2
3��S�B����3E7�:)Fŏ@�Q6��Y��#�{1��������1
�_��zVt�/�T�D����:���1�mQ�/�K��>O�i��'�kE�g�A�p7����̹���dc
)PE���V1Fc䗶!�{R).����ʽ{on��.����B��o�xcB����*��#��/UEf$&�����~�+�H2r9���2�xFr�OJۨ��j%��\�O�x�w\���?\�jlR���Of��t��5�2Zע]�p�L��0T��Ln��E.�K����P�1�	$A�Ʌ~�����*�4J�ʍ�n�3qZ]�Ә}.��D��|�u���7����g����Q�ǳ!��w�}����YCl_YD�/Y��c�z�Ӿ�C�Y��2��v2"c���]o�b��KƓdwA���BkG�{��>S�I컥k�}WdV^� )�� әF�hL]�+�����@1��7�=	0���z�b�v93,��~_Zq1�c�J��O
;J�����3;�3��+v�o\s,���^8h��^Q��>�Nx��1h��ew;���������_��q�|dd)�x� w��dzKi�KJC][���4q��o=�����Q6d�(B�|����E{Q70�����w�V^@�J���,���C�1y�?�Y�A[x.�O��}'���Y%|���(YOl)Z�W��/5cy�)K�4��"�6�d��6b��+l;\ʍ�N�Ni�,
RJg��+Fc$����<�o�א��?Gѥ+{��@P�LR�����P%$Npo�=XlvޜLJ�B[�9��_�s��^�ji�:5�V��S�f��H���?���Z.~��������"�S�������E[���ѮY��$�WqU��}z�_��"IH����]�Ɠ�s��*A��O�O���إ8)x�����4v)94:JɥM�V׈���d0G��k�)����鋒�ƨbą�u���D���q������q�k���;�mc�\{W�N�qj�	�5{��j^�Im_w �\|����ARI�w�C��]'a���j�yH	�T!��`5 ?�6�*N�V}G�����gr'|ʏ�}��V�v^|}�y<k���}@�5>ֻɜD)k�m��åz��,��y��.>�����T!����"1�6�>���\XO$Q������?�^�Ga�#�T�k�0jr��*�HJ;J�Δ����R�������(�g����]�$|��$_�<������pRk6�@AS̸7���]"W}'����HYݑ���=���29k��B��� Z=n�%��Q+���V��X�O&��u�@�$�gۀP�(�?�G_��_�a���T���?-��sL5$!�ʪ�j�h�� x7��5���c�_y�\bQ�ͬ��vNy����>Ԝ|N��J�C@cO����3`KbF)s�H��@&Y#1���C>8���J@r6&�����|��F~K4����AD�{e9�-Ejx��L6
��?�������(��mR����Y����y��)��?Q�ȃ	�O
p���!.����@)�Ե�	)-�v���Jk�����;(�/�![���Pb�֌�_
 ��7Wu��6�tI�N��W�o������j�'W
��ه�Z�=�j���4��%�<}�Vmo/�於.�K]���n�p/	�x���;Eï7�aj��!�>�J��v���"����m)j̹H�}z���qt-��[��[��u)�{%ݍgTT�a%���7��5aX>�ǖA��w�-�+1-͵�vyYl�v��� yC�����Oh�i��lX�_M �0���~��f��� g*A<��"-��f�4dX� %Dt��vũ��'P�5���,�V@a_nD�T�lUN�ӟ��"�4v��w�]l�*vC�v�R+��~wMU>N���-�>᣻��v����.�ϴE[��[������:p[�kB>�f=}����f���aw>���;g��[-}�y�:��[��q��fu������m~�����r��Fw0�'��{�
�6&�Ï����C!�uS��9�h��������ob�V��^kC�[t� �Hb�ٻ�
�!Z�T[y,��?�$�w<O�&4��:0�{C38i��*�l,I ~�G��b����(�a�"�l��j����"��;�M�Dn���fWM�ZE�X��I�.�X�4|B�d��n�ޡR�u�o?�s\xt���ޖe��*ڵ#{��s���h
��s�W#���Y6�G��~�tw]��}y��E��T`�o�˘z�x�U�p-�ޘ ���JVU�2̧�Es'�<��>lyN�>���CORa$.��'�G ���"���A��*L�a���Y����]�S�Բe&�`�nOnf�7��(���h�d�ܜ|�^�K*�C{z]X�	f��)������@�����U$��O$��A٣1o���d���2,��a�4,! ��ҵt����t���]�Jw��tww��)�H7�����q�k>L����9g�3�Y����XVPUFw$6*�{b�?D�!��B�)��o��~�E̲�rjgU�	�s��𩄉�K]-�n�G�9[.{v�3�
巙�C��jFM�sM�Z��kMl�7�aG%�f�I�՟��C�{BFĥF���d�4��hi,_�� �i�N�8�.n(�v^���@��{W5�re\��{�w���튷�VM����\7����Sm'���P;SY$SY.[�C;}���AN��'�1�?c��4�M�w�m/g�6�0�B~��/�e���u����^ERն�C3q�^Lt��0!&Y�s%խ���C��4��B���C^J�H~l����@����0?���Ʀ�z$�zh���aD�� 9E� ��9�%�u'��=�o6�j�Z�;e�M ck�[���d-�V�AC޳�h��8�*� ��׉WNJs��,�����9���ib���Ɠ�=����G0TJu.%9q��[FC|F'-F��g�<�t�������s��7G��&`ȸ1I�V��E�	�V�.7f��,��w;a:w܊s3=�!���N��9@�g��q�
('@I�m@^���oc��K ��y���MR�&/��l��C����7���J]�  �k�،w����^V���3����>�Z�#R|�N��F�~OmR{�4�D�2�cd�1R�{���8C����,���ɬ�p��tE��C?Kz{��J<7ع����e�"�U��[��jڱ�.v�A������V�:)#���}VRK�c
Kڕ�� 5\�Èu7Tm$�Qm����u�l�KMNE]���na�[[_JIӈ��K���~K��4��##z\��R}pr����k������^;N��3�V뉇���P�1t�E�K{3�L�Yǂ˶��n�\i�<1G���v9��<�v䧥.{�Sx�4��T؅�W%1?e>�(SLWh�h�P��_��.29;�OnOM�R��w<��g���A�uQ���N��Y�>��L����k��������D_hLJJ���S���1zG~�G)G+�����4B��kf�3�MU���/fK�n�Y�3��o���G���oR���4'��h\j�I����1r"fÉ���K
n{J��W��Y;���6WO����,�,�h��&^L\&8��ytUG"�����%����0����i����=b?��<��59�08�\�3��gbٔuҞg�ȫc]Lv<U45:�&�z /�ѥ�!�t _&M�������َ�[�~D֝t��i���mz[�&�4�T��2�h�Vc�Yctt�E���q�~�(FpT`d���z�PQa^��3v���u����aޙ�3U۶�*_�8@�<N�4�_oH(�noh):^wIb�_�O�������a�����SP�T�E��<�en�-ث��͗[�]q�JY��(=x$�����j��AS��A��e���X�=�,^�,D��P6<ٷ�E�<�����ŨwzTߍ��)0lIni��l0��J]o� ��)���E����Y�Y1��n)����c�h4���w�"5��Zd.�>n��A��
��'����L��x�Gu!?�$��GaA����tb�x�eX���ʮ���񻑶����Ө�c,c�V�*���%�h� ˩g����m<�[�_��}�R~�/]�o�l�pL;2,]h%��W��6��o��� k��hNf����XF��
,���e3C*����*?��ϭ,����#�WU�c1��'MƲ�b/E�hbBg����%�~@�m��ɓ��j<���Oȱ��k}��ol�=V��A1o��O>��+BM��A�h�o�!S.�yP\}[H�ؾi���%[�%͔5��ޣhF;M�ͅ �a#�++xK��a��%WL�U���L�F}��NQ��L�S��5rɦr��\�O�"�Ox���-pz�XQ�Щ>ߦ�S|�*Ja�Q$�n54��k�v���چH��=��]��f/��q�$� ��nQY�o`YY
//��w��mlK-�~�)�Z�y/M���>(���/C��L�eyN�y������d���	�m�vl��s��`�4ā<A�_���^X6Pl.�14��+�I�J�������FQ� �ݕv�§��%+�C�<�ko�-��+��͆�JeǊp
ʥf�1F�\�:���=2�,Cb�����LEQw��`:rS�~��E(�N'>��1�K��_���T�͇��T�V����}{�5Ŗ����{Ȓb�k5TUY\���-fT���n���2����(�P������;_�}���p;3�h{��!�=��~^�.���_Cw�	+����+�+�0#HR��Y�4H��XAD���K�-�k����f���Q�*��쨆�r�$�la�{AEMqi-��|�Z��{���s?/�dxY��8!�;X|����on�(��ܤ��!�����d@@!tY�g�~C�8s���I�?Ҏ�xA ��(�P����L�NXg5
��ћ�ާ���hv>O~�����8h� -����q��L�9<�?b�!��\k��= �����W��B`@��N�����x�R���߽��.��\b�8;������q�I���D�������/���/�ug�����z�z-]��l	Y���Xױ��`]��?�j�a0l>R���ܥ��U�/����'�aP�#��H�
�ұ�_b`�ږ�8R�kJ�Q��.
��={��D񲩆����jf����ռ2���G���E�N"F"�8�)�5��Z�R�JZ��S(T��~��J��v�O9������[�F��˞Г^8nZ��񐑰SP��P����q���S��.�Y)���ju�)DYL��S�c�e�b�MF���o៌i�pW�z��hhR����xu�����n��a~Ţ���W��o]�����$�K�����s��9V���XD)'�k�͑�ڞ
wl.2��#v�"2�,7������B���h�^�{�����i�'�M�R�tDK�n,?@p֫����IN}��pg�\��/h�j>�fC���y$�^eLg@T��FH3��Y����b�Ef,ۻ�ؿF\p�Io�[@�6�RoD����6eȟb� H	�� �B�V�ﱼ���B�/��ק*�zv���V&����
L��ģ���'s�w�7���N�޽4��+��km1a'�`���K�d�iRk�2�����{�9{s}Xs�Q�" E)����P1'�'-�_Xx�Z⻧������%����߃�~� X��� �C��" )i3=�]@�}��F���&�1���{���@"��>c��]������	�J4�b��:���mU������ZB�F�� �1�ɶz�?$eUt�R/%�ԘE�[�4��Ʈ�`����G�"�\g2���_�!BUOâ#�xx%C���0�c��ql�Z:��7^�q3k�W�A&�u�L���O#@9� �
�-���<�܅�R���ҫ*a�޹ӥ"磚?F��9��8C۷�����Ug�sM��?��+m�i<�EZ��+-�2����,�J	ײ��S���d�:�ќ!��c}��^ŗF�0�_z���@QD����P�Ž��A�Y�����o�6�QD�Ի���w��#4��r	��g'��)���g~\&f�1��n<XA�����O�n��K֛��)�����`�����O0	��~:��L�����E��a���/�����g�Iې{[�֤e�iË�����h�E�E݄�h�b��h>PV��e���z�c����筰�Ѹt�u����yY�V"U,Ĺ����j���;������2w�	�[e�rT7b��i@�@v���b�?cN��$+��d$���l����^T'�y:��xBnޗ¾5�{z��Yy�z/wcc�6/�Im^{�~��ye����wV���M�kDi�n�\�ޟ�CX��5c��R �䜓�����W�'�.���{���q��{X*k3��I�������G�NS�L���E.6qܕ����S��Fn~�y���g.9e���Z�J�>�WO��6p-�������@Y����iH����eESf;#=h�N/�"�{ƇzԕsE����c��vA�G�?�n/�V����M�@��Ljk�`�>��4�ų��o������rr�؃�'��|F��(��ƴ/���Y��c��R�a�G�J��rӐ�u=">�<꩐�)9�Q�YT�x��������o'���۸m�~B���=�[>�X�	���$��F���td�3�12��[���X��	ws ��!��V�/�U#����l��}FEt�?q�P�/�w�p��&����݋=��J�+�'�QӪ���F�;.��{��&!�����};6/��z�(���ڠ�c�io�n��\q�3;�l�]�_���m+���y�"a�&���J�˖�E��;=����y�T9R�r^h��;�iܚ�bx1�K�v��`J�nB)S��X!���} 0Y��^�
@��#���6O���G��|0;r٦������Qӎs{�/b.�P�a.�6~6�'�d�O�=u�7��c��Kr���sww�3S���J�����ʮ=����)X���]�w������Wat��z�$t-F6[��v$=l��f���"�<�q���^�d��X~�JD����o�1+B���8�LeĒ�w��u�y��ߝ���z�,NB�ۆѕ<$��X��z�r�K3�s.�]���k�,=sRNT��n���5����7nh&��<�:-���y���W��ɬ����O3�,�I� =;K�3�����!?�����#�~+�a9
���##�{��c���ڥ���]r�s�<��>R�!^#�M �d���]��F�J͸L=l�ܪ���<�=�ThkiSPLr�;%�j��=��u��v��p6�vf�es��v����a�3}�F�D�9fX�)<�O��D~�F��C� �|���a
�6E,�$��d~~kU1��y�����ep�6u^�^�4"vӨ���O~X�IT���	(��P@���w8.X
ueci�W�@c*����3��7�2�7��.�6�ݕ�Zw��wc����n���ﯔk%�Ñ��ܭާ�ȥKSMʻ�b��q���[��ga�M;�C3�cL{NN��"V�1J��O��'<��1ٔ�������yc��V�[;��9��9��2�#B�L���1�5���z���Ϲ�RU�{��FE���(JQ�e͆	����D!-QMH��H�_�(X-�����H9P-%M��� �����\E9���T���T#;Ɂ( �I�����[�m�W����0�������>���M�N�n�g ��,���a�Ŕ[c���ag5��;���^����l ���\�u�����%J���p'*@h�����&D���GX��H���`e��x�~M��\ 
����(�fZ:��J��;����w�xB�wr�e
�;�pg	�����Y����8u!���u�6WO�A~��N���Z�RƁN�_���2�\f|�Ƽ���u�M�;͜��b�.P�����T�g�Um��H\��N	Ǫ�#�8����Q1��j�������[�Y]yz�z�w��~7#�{v��m��y~*��m�㾼u�<R��$
��EU����|�y�FN�f.�F._����ҲRb	�z�\�x�"��X/�p{r{ֻ**�*�vi���w8�$�dv%�W�=�G�Ց�)k2}I�-W�×|�&�XsjXS!��`��O���f?O�T���WH�Sh�Q؞7�Se��u��6'cһ��o/�MMVč�"�����+2l�y��m�U�c5�)!y�����ә�#F��{�/�2���L��uհ?���wB��a��:^�`e�M&@��Pq�Gh�*�w=s@g?�QYEl̎J��_�Ϥ��yq�`u̹g�i�$H��~�k��u��J+��L�L :���II�U����;���	���|0|l?�m�WQ��>��e�M� C.2<ڃ{u�v�Q7i���#B\�U��V ��2�{E�c�Gu�o,�P���7^��
���B�LC�!�{�E�=*��┆���9�.jئk�69��	�	v�RS�{4T���ԉ�*�ڨ\s�xh�;+r�-��Z,1��"JɍIS�?.��]�&�0�h�[N�fM� \� ��N�zz1��,"�8���^���w��(r�vRDPS�a�F��,D��u�Pψe'P�B�3G�p�j��$Eބ��3�]�����9qj)*,�Ɓ ��ڼ�H��)"1gNEp&��[�A��ԅ�Tл L\1W����c�MX�?N�<I�Šd�u�}܈����o��%��C�Q�ג��մ�T�5��_ÒV�C�sy� �/��1�H��U&��c����o����H�3H�0UD�yR_vTBq: ���|(�	*�AFb�|~[3E��C��6�*�t��4掓H
�]�J����T(~��U0ԾC�R���?��v�m-~;~�*k�`@,����99�����ek>l�c��Uѣmy��Vpœ֐l𴠖��-' rS�>+%M�y\�g?Kj_V��Q�i)t3�[��,o.j5�X�6��'<��_*c^��<U�0�-�{k��|�������uK��@��n����񄌕�{-�{M�;Mc����k��Z����}V�}�2]�Rk�������80�e�F*�2�.�TT��f�WӍ�.��	�I�i��hkJ��{<�I�k�2�fe:�p6Y�ź��0�䑄-TXN���ˁ��Bu�rl�%fD%/����S��M��q>�.��d��H�v�_񍽓�0��&wfm*���#�]�&=Gc���ѥ�ݵ�Wx�n��/��믫�.OM�
j8�e��2��/�v�r�p����ds�� y@�zh{�?�D�	��8��4�e-4E�@�DZ�m,��B��`Cd=�u~��G ��5l���Q�$蛘��pEQ��$o�5�3�o,ek�e���]��[�wPֽ�y2Y�zle�io�E���YQ,�u\iyh��*��1?I��朓��p���t�y˗E:]�XKg�}�%-���]�z��}K��UB��������q^�̼)��M���{yk�m�
�3�x*�u
� �䭡#�� $� ��/��Fn5��N��I��u�z0~�SO�rV[u��2���_3}�U[���Q���M�e�̹�Y۝�����x�q*�0���P2��F�Y��2�i�9�	I]ӦW�b�v0�/��%���^�����#,�Ap�k�����h��n��Q���;�\�|�L�j�.���r����`]1�GK΁��sf����'+�&��nқ�AMe�wL���wr�n��M���_H���Z :;'��� ������s�,��nN��Бl��51�n��zb��v(�:|u��m��t�	��-ffQ��Ab�.͓n��)�q�ě�n��
b�9Z�<�<�P�R��3Ҿ�N|V�4܅>���B8�j%L��a�xA��*�hi���W-��TU\�%���M#4/$�p�k�NCl��d`V�+���|��b�Bv5�8f��6|��6������G9�7��ă�'X�;!=���7���������������<ؾ�&�s��� ����]��R˫�:
 ,����a����5�焖[�]Fly�z���%G��0+Wk����2���߸��������� �đ!���H�q�n�0<;G@��?��qN7�L��Բ�RFDF��v,�l �,Ϟ�>%j\^(���t��o脰��g�~(�e]tw��0��3�K���xvv����+�������B0�rs�d=�_��u*�\_�q|��해�[��z]��էm�ac�E��8�J�ĝ:
�r��V�\��?6��m�K;^j%ڃ���g�aձ�a��\^�^�Y�\f��(Wo=3}	,z���)5��vX-�9�`��W�=@Q\������ �yVfN��h�A�Ե�Vo�?���i��5�e�r�,�^+Pþ4?�V���Vp2ɦ�@w__!�Z1Ä��ƌֱ����޹�4�	�ĭ����~�-&��O��{w�F#w��Rn_H����R�bJRt��[m�W���n����,ؕ;��_8vƺfu�7hli���^:�h�nX���!���ۉ�|�h��%�:`��m�W��e6�i�/��x��1�tp�r��t��_�:�4��� ����E�p�8u�-��/��<3W1*����Rj�fi�-��25���t�`�õ8#tlz��8��N���h��N�%�?g�<�'���`�`�Y(�}���50Z��~9�ꂆ0Z�~?N#���������A�ʁ#۶]��c���]��`rZ� ��<��M�Q!�Z3W-� b%�WNe�=�D� �<�/�b"��-9��u5�˺�oMb��ӧ�N���Q� m��2�9��>�n%��-��Ý`Mq*uݻܯ����Iʈ�(�!��$5���;��rY�+����j��wZ/WS����w�ͺ��۹�$������$��&զ�����fab��xJȸ����հ=DBz|x�ZE�FlG9��/��g��V)XN(��۽ӑ���?�q�;��=�i��˲}��O�}#����ݵ����Xk�*J�q9��Q|W����bK��ޅ��/Q����I>� ��1����k�}����q������� *���i6c�q����l��%=�&�<>�|���m��m��j'u��4���2Ϊ4�%�38�Ɨ���%�ۿ�0/h��yTq�������̈������+k�Y�E�׮ N.E�n0�Ԅ��3(�L��_�fF�-�ˊ8��w���R�1�9Q���Է�v^�k?�w��訊���U����,�moӋ���l;1�-�]s�D@�L~�	Z(G���g]����'A;8J~7��>���]����� ?�?��_Rve�����.��B�J����D��MP	5&?����*�ͅ���[�I�i̽;�K�k��~�7`�� �mQci�4'��_0��?�5��d��$:��/�T�����d��U{���m<�H4,�aQ�܌&U]���V�_�����zz��h�\�[v�]�&� ;��f��7{�ۅ�<�/������ �-�i�=��f��mL��Uo@���a��	2�3P\�P	��v�B�m��9�����_�f�R��HL��/у��_p�[����e��K�T�V��E�'kTRT�p�@���}�ؚ�<��~�%�C�h�7&&�Jf�)��� ���Ts��������sW-��&5��ċʅ�	�戱�(�s�adqY�Vc1������������T:�V[���6�,����c)�~#ձua�or��zdt��:b�P��R#���Bs=O���~v�mX�S �K�Zdh�4FVL�@�t��ᔩx)`��e-U�b�?��|����f/�|"y�����R��8FoWy�_������t~G�.�P���Rd��Ǟ�Em��/�>���7��i0�ؔX�so	�H7�\U�v�y���5��o��YXX�$�m�]�X^����@`�Ą����e�v²i�'ҦM�S&~���t3���iDp�Go��LG���&��2j�ju���7:v�Z6N�v6y���.���~}�<��j�K�F\�>���a�G�T�SS��#�����f5�p<��	�]�d=��훷a���5]&:�ܫuı�K������\��E\�����b�4g0��2�c�ce���`'nyx ������9p����"�T�^.�%Ti8Sx���~�?An�H�-J���P��k���Ŀ�{��;�ɇO�#��t%X���F��cܺ�n�Ŭ�s�d�G�MsWy��g ���س��Tc��O���
�/��� U��!@�t�L�˯N����s����M���_cS�x�?�����O[]\_�.���M�H>����᫠�߶Jw�ײn֒��O�:����4�ˣx����Wg�r r�dFKi��F�]>m}�|t�� ��r�]�i����O�}_Z�ܘ��匢���K���o��#瑎��Û�,�.�߮�vӁ8�e�?o�\ť󲶆�D�~�Gղ~u�T���Ë���x!!1�~�{Z������������~_f�F����{ږR�F�<����\"�#��K�h�H�7�E��.zX��9 �2��{6V���}E���2�(ḭry3f�5�|���LnY�����γ��D&eˢ�3�^@�L��M�.��L]n]�Ο�y��>A�=j�x�x�eqq��(~^��[��;2�c��醇k_������L-g!�N�U��n0+)��IpAJ��D�+'=�|_���de�D�G���뾵��+�)�+���t-8=J��[N�T�
�o�}w[�JCxy�L[:�p�8�a�ܶ�Oα|c,E,�qx�����P�/��ٵ]>��t���s�bp~�d��%�]�壎����n�	I��ml�����v-����̗�B)��ِ^YL`\cƻ(>�ϑbJ~������-��5P�l-|���Rwg,�^�Wa謑��o��������T��I�Ih����!��y�@ރ��^��0������$J4!,�S�8\s9�f@i/���F�"��9�%	����!�2N�N���0LXEme;��\$`�o��3��(�t���u�ì��;[S5sё� f0�zD����\/w����^��z��MZ{�^wn��]{�
]����E�}Wj���cĪe�қ�����v����bfV�F����_{\H�ÉSn
P�9N�P�����7���&����=�Њ�����]�y��=��Z�N�Zz�s��`*4���Qz���s����e*����C[�t]���P�]��^�ޏ��hH�Mo��c㉅�V��P��D�g�ؒ�MJ*�U>�9�nマ�o��;���8��A?����vTbf��-LTY �=H��W���p~k��T��x�xG#/<Y�;�,�����_;K���Ӝcy}~r�L�.��	p�D�9���Ƨ�t��8�N����G6&4�?0�|H'�H$G��5��,�O�NO����կxGx#���ܽP�S:��"�TH���Uc</Y�-;wqV��2qu���X��߁����t]\���}^�+]�u���٢��⸜�m�@�/�p�F�~,�QRw&ͥK����ww�b"�r����߇L��kQ~�J^�Ӽ�_p9�s"�$3�i'��a���1ƿ�"��"�IH��	>&/f�aH�4T�b|R�NR Nu��/���Ƿ���a3.�6l�o�[�i*gK?f����z?�kH��ڏkɍǅgk>�kO=�q����rO�������E�CoC�����B����XBS^*.�(.^�lmiT��� %//]��[�7D+��t����f��Bq���\�ͥ����K�]O�/��.a��Fـ+T�l�l���3�)��Y���T�����m�T-�s)��/M5t+�#�  ��D�Jy*��^�r�̚���]"'�h��`�����*l�mJdo6f�vj��}r!4k��O\��Okk�P����^�=��5��"GA@���Thgi��1ÿ1D�d4��ǌ�W�V�^����<��'��A&E�Y���Mr��h����+k��Ht�TH�V����|zsM�7i� ���jh�	�-���w���b��AA�NJ؂��v�̳oHt�p�bW�!5��K�8��A�=���W&�'<��q.uz�f�N��Y�tx׮~�N��*�n��A0܎��ɾ��`iڙ��� ���g����瓘������uJ6���?�����zK����N+���v�-/��/V�,t�j?�]>���˹p�����i:���3>N^s<������*?h���j�X�$��_�So�=��n�=�Znm�mc��͕�2cgM����KLP�?ߜ<U���N%G��ܝu�1?��/ե�?8������djv�Z�?@N���[.;��`=��&훆��#{Zs���gV�( څ���@��}D���D���N�*}�]��p�$��m��g�!O�����;���9q����n�ym��1u�(��׵�\��\~D�RZ�K�d|`.�� p�Xi>$ڹ����ȡ��_��t4V��;q��<�
!b����N����X���T$�m%	���iQ��=;J~�����#��G������˸���ёU7�w����~)������;) �q4f0a�ʆ��#W�30�X�uU�i�9.�R��,�O!To8g>]���`}��d��cd]��Pά�=��2��,L���v�����r4�q���/:���&�Z�<+|���A<Q.P�г���٥ !��:��-�K;]��r�#��1f�e�X�����������v1��xqx�"�l)2�x����F��]�U��K�-���e��9f���^�2&�A��v�r�w�L��2���Gܿ�_\nSl�u���	~2�5q"l}��}�}y����N
��*�Ƌ�EA�+\��}YF��I����+%��x1���Ҥr���5j��Z�NB��;ڸ�ޛ�tYb�4�j�k�R����b��������E/�yڕ"M�>c��5]B�ѫQ�2�ś��D�3;��
Q���wDh
2�:ݦk�
CF��۩�`j��!�D���DL��<���9�+���R{pd��A����	D<��L��.��T���v�$Y7����9��,:�!~��ǆt]��lAHYk�.�W���k\��oQ�"�7�G�:d�r+��wG�rN@7[�<�u��H��V��v�I8~r�i67p�t�hr��u5����йM=g��M���9M~ߑ���7�ۃ�w�Z��,½%CS�柨��f�k����.�X|�+|.�~��q�:^��ݶv��z���_̢�T
�����i�@�(��R��r�v�dM�:���$SQH�JY��b�t8L����%�n������}�R9�*��Q��p�JzA2J!r�7�٧���u�Y�"2�D��D���LJ�Կ�BFpEJ�E�@'H�ҋ>;�`�h���w2I��+����cx���j�{���ߣ��-[�3EU�Y�R���e������\e��U5��t0�O��65�<�ox�g}�ۮg�05Z	���O��<7���,y3B\$��[b��F�}*���`)#�Fs���ˌv7W�=��^�j�<��~d�;p�z{��3#���虙�<C�P8��3�W�;������1ޓ���S�ab���(��P��t�����b�����8�|�)���Ny��'��+��c��'��� ��T�7w׈.?�����j�����^Fm�Z��,)Z_�*:�6n6��������K��IU�+��Ed㗣j��qH���	v4��v��3Z���L *�KO!��9+r����;LŇ^o�����v(�][�W�|<���ɦ���r�,��9OA)�o 3�/�-�W�)eV����͒`<U�l�-<��^[��l��.�]�yX��+�.�Kx��oʳ�Zߩc�?~ �Ndͱ@9��u�R��a��7Y�D��3_S2j����hta���߼9����s:���w?����4�l�������kl�Fͷ�#�i3e%T�=;5fzȈ��,ęν����]�Y�x�K4�p�Y@J����z@��w7Tʅ����w�B��}Cf� c�o-����Q���1�ᙹҜ�s:=ڭ�koG#�P�@�2��S�
�%�f^|�A�~���7;���@����d�C[)�| �M�0Y��~K�AS��ҁi��D��z��?ט��of���f�\��6����5�q �������2�4 c��x�4\n)E����D�=}�L��(`,dhP��Ҽ{��@�o�6ƶ�Z_}�j�К�~�צOE�o����zt+u���'%,̭1)��y��(�4xȟ}qկXC_��Қ0�k�)�$Q�
��t��^�|i�[��:>岶z����h���o�� �4ܿǉt6�<%��$��d����ω�&o�zGI��3�9��m45�XT'�0s��H�e��8�Dq61�Y�;�ҁwG�h�`���5A{�D<IB�#�^�b�"Ȗn�T���g��ᒑ��[sF�l��.�=K����v��X�N~<�;���?��
7�;�8�jM@�q�AxIhٳ����i�t�f��}S�@L	�$�����K+gЗ�՗�W��[?vwF�c��)к�&���k�{<�?��5$J�q�^�'4��4�p�}Ԑtv�1psOU��ʹ��5Bɱ��8�\kDG�=|k��@>������ "��ԥr;�������t�~�
{5��d�����i����-�ח�4��Y[����5��O���xqk����^��DZ��G��wH:���O7~ͦ�E��|2e0��š�'D����Ã[:����'��h���P��<�Ƒ���l߭g����M��/v����Jo
��L��Sc%�\��l������d�)�e�Q5��{�!fٻ�)W��?X���xJxu0��ȷ�-�Ƈ�G�z�G8	Bsv�~��-��SZ�Z�؄�&X���(��gp�
�h85��!MZ�|�Iq&]�7rA��=�55a��l$'��bt�]S��c/�0���+�!�����h�%G+W�����ChS���>B�L��e��b��ߖ����=��uc�	���;�)�ש ��bJe��ҧڃ^ڪNG�	Wv��5o�N�����8nK=�ڧhzk��# Ly؍c�󋑢M��8P>��;f2�'#,�b�%D9�:	���)t�dk��ʽ��ߎ�b��jk�*s�E3�8��:B�@;>���	]�9h*"%��~B0q��������������l�a]�7�������N#<z%����]!�!��h�ym��l�Sp�Ŕ���P��Ae�*���O��i�.p:�J��<����x%��ܯ�ȶ*~5y4H�4kdm?pH���<���#�/��UY�j�25ǣ�cJ�����L&Y}��HA���ŷ���c�b&�u�3���Mu�y��K)*ogο"_�"�7�1L(�\���XhH�j�/���(>�����U��:Y�[��
���[I��J��c�0�*'>x�CQha~��	5q��D�>d-Ї�G�<�.���7m������ $s�
�T�"�C-1l�ڮ����͠�u��s��^��{R0�{(���NLG�4���g����g9�[!^�)o/j#_��G�p³���%���.��K*���Z��y��p��i��6�~�V���ny�i�v���͵��顙��h�=��e�h+�be6��^��>O���g6�ƍ�*sH��B�U��(�>�h:�w?C%���wT�@4��&6�:�������Fv�/����BE_��mB��4�?zu���櫙�˘��z1��G�wݔ'�����B&��Ъz�B6k���љd��R>��.IF�*\s�Zrk	�zZGo��!FbJ�f��r�q����R�&["Q�;�S#z�ݒ��;Z9yG֞ɷ��#�K	�v�4�0+�S3�������L^2�
(OC��C��T~����5Hg������L�������^_����0+T��5�(���Ije�?���G�zKG>�J�l�/.�x������S)墘�Hl��M~�-P �=i0�v�P�[A1s�>9��GP/Ay&�h��Ώ4��OE_���'��С�Y/;|j�^�8�����Y�p4���l���[)tX�X�n��{Dl�jc��
�}�A�_؀s���J��N��u�4���k���K_�f�qUa���g�XL*�޴J!^�Mp(YS���2������Ӹ����Ʉ��sE��tŪF�w-�0�	x^�QQ�Kh����N���d�r���rMZ:���-&o��ގ�L���!�p�9p�\gg���tK4C~S9�0��{�>UV�،�!�`8:8�G�l~�4�G�� �h+��*r9s8��z��x�����35Z����cܓ�h�1�W�r�{p]�z�C��NW�`����v�HU>����X��Y�,�l�z
Z��+́�Х��Jӡ�Q�hU�@�9S�i~j��&��ћ
�)��$���&�}���W�g�W��{�񟁕�G�Y�EՅ��n���T�S�!�nR���E��A���������{��霏{>��u���vhj;3�	��c�p8�d.������|�"�Vw��f�7$js�&�pTU}��Vǡ�)�e_���9r��	6.����AH1�#��?����o�L|�۟�qp�t��R:4�ŉ�*��Y'��Q�}�֟z�����AF�jhR��X	��,ʡ?��zX>�}�Q����6P��e��?�j��|����X�}�]3�����x�c�.�o���M���0Q�fZÂ�4B_�x]���]�lY�\��:�@��6D�hs5�����o:#���D�K�;�1�6��Y*�� �ۺ�����:ga�`^u?DW��:9.�`���ι�6�+�V�	��P&/Ck8���s���l���3,��@�~�Nx��V�9e�x��Հ֠�К��"76ȴ��@�Q���-Z�ț�QoIx�p84>����X�M�ж��X�	�����X��(�zR|A�=S�A�C����ߦ��ϻ⡖�Q�?��Jϣ	j�2F ��[�8��v,.�D�[�b.�mлl�Y<�5}�������g2�H�r��+��LӋ'�K�b�����o�P�;Oߥo�I�6iԂ�O\	?hp�/��T����V{Y.&�a�YQ���B����謉�K}&|�;�;S�@���3��5�?�B�S�fba����,i�ī ���M��o,Ü�0tE3�$'Y���{��]�#l���h�pH|��-���Le/N��3ż����ܢj�U�n:���R���D���p����5�P$��B�����y���7��:�Ee�q��
*G�#��x�����Ր��{��	�`�{�j^5{�9C�k�/6o�"G �-D	F�,h��\쾳�Bo-����ݚI�D0�g��'�,�ju���|�W[�lK�w���
�l�p��Vc"�n���kj���瑞V�(,�f'�<�<M*[��a��f����n�U�.��G��Ƒ����Q�(ծ��RJ(�҃j���&[;�+�@�� i���F^c�(�q'R���B�	���^�,��/W���������B�¼���$v�TR�+�c�����{��+�4��|���*O����Iq�6˜�AAcqL�nN̽T˖<֝)�V���B�����?��#��o���^�hTT�v`���f!�[�ј��a; �8�$4�Y �b���~�|=\Yul�sz7�q�Ԣ���D&H�j�Gx�Ih��H��h�p�װd�H8.�Aga��4�s���U-�y_$MѴ�`�����s0�C� r�)?���#�X�Ok�cWΆN,p�g�8�{����jUܺ�S�ZF�
7�ID��1��؟Q��J�l������(��ۍ�p��]Q��1��"��Q}}|$���)+�j#�o^g8�ǝ��Ur)� Z�����&�R���ܧ�c�w]��/oDk�߷T�(��(H}=Nc	腐�A���50s�����%˖feox�7P�6+���|�"s�O���rR�/.%s�B�7�N�H@��M�Hr�m�>�C�c`u6�HNK����l�ɞLô�@M���׹�BۯZ^�z��~���uC���5Mk!�B��U�A���y��A�Ū�2�,5�$i�Xg�La�q����z��z�Nǭݠ4�Eȹ����)��9w��N�w]�|����6�,�9�������Z������ǝ�֗���M������������Q������Y�\N��3�(3�[l���zD��.!�OV+k[5�8�ꣻ������o"�ߔl���cm��u-3�5�����g����w�k�UHՓ	-�d�}��$S�s��܀�]���]�Q��V��U�cȶIȾ	��8�Dw:�F&�*~u���.�����דQ��A��aG{g[ ^�?�\�|�\�T���ik��Q��c-I���EJp���]�����%:�ui�QB�Rd�$�B.��̨B]<YAކ=j��x�͎ߖ��0��p�����͔.U!�N�_{-q�p�����E��Ű�����������kw-��Z!�,�^=�^�LAx��\*m��~^�{�� or!$�|���I=����/���o���<?��-����W�C���[d������� �^��*�$��(�qZV�&O���|��~?�x�C���1�r���cy)Z<��@Tw�f_�/� 3f�|fisK:�Qفў�1�$C��x=h�p�!yl�Ψ���z�T䱐�Jpu���B��� �7a�߈wݍ��r�$�_��y��\����Y�z�7���\fV�K�>23��U�K^���6�o,`ѵ�& �jTP^�����λ���X}��i��n<ы����YJ���������
�b��I�	�tg
�E�pV=�Tq��a�7K�����Y��2;�s�oW��w^��� a�(�I�m\%� LD��A�Q�)`ӆ	Q���O��z�b��D�F ե"Qn��I6�ů�Y��ܖ�^�����Ut�'׳�[�%yK�[�A�$����T���sAŪ�NH�O�"��G���������-,��h枳l��t��D���W_~~E�䞌���r/�����w1E3�$��{J��ˤ}�����X1�Q��lꕰ�T��T_��&�����H�dl5y6��<����N��P�=�ɯ�{t.�Z䠅�.ܜ"��z8&Kĺ�Eǰ_V�Ez�݉�o�R�0E�SL��@�S�<񧞄���w �|�Z�9�N��9�6=�"`�b�'����##%�������L�KٟӇ�N��/ې�����Q������n��ғ�9:�91 �|:�@$�F�&�[��9����0QV1!`�]
 #�29c��{N�׃��ڍZ<�=B�-z�-Nw���b-��TR�pep}�h��zUoj��b�;�IҰ�"�����4�n��̻U�������]�5	���3mZdwG!� 틝֘,�����V0l�!zԑW��
��Zw�:�'y��b *��:_'��]�tZ�%K���T�*Wi���.?�m��C���@�u�����o���n��5('TYg����@9�����-�z��M@�]E�òCeli$&�&�6���!	z�,�y*��&3c�H�\�)�@�M74)N��w���,�=ؑ&�5��L������G\�$��[S�u���0��ŧ��3�����;Ʈ��6"?Ց��HV��x�W`k38�u[�\�to�0އb�&���`�s�-f�����،��e�E���K蕥{k1��| �]���2 5w��y��$��ئ��muж��Ȁ�xr�n�Zg�Q�#I��+���8�F�5_��,^��з�\�������p(N;/��u3�`
��,N8"��{����[��n��'�3q=�<X<"�ޣ���8�����~{['���G��,&�2�o�m�>puP�dK�g�|�3�֢*F�������*(7/�L{t!��	�^�([���y4�!������A�z؎�4���O�Cy"����<�8S �z7��3�J;�XӼ�ۄ�)W��!��E!m֊a�{B&�v�Q����~��͉�S�����������֣iD���߆W��*R\�Z>�.+z��p�E�WYYS)�B�6�ퟙZ�#�/<���I�TM�?/ķ��R��C���g��@��%�I*(�NP�5��J�oHޚ��F�����6�D�=��x���?+���Q�fng�}l~R��V\Þl��c��/�Um?�[9�ce��e�e��L��A�0}�a���JgjЇ�ĩn�E��?p�߳Jg�iE%S����>�����|�#�n�u�������>w�$%������jZ�,7�صN��ś�Y5��ާ����
��e3T�'-g�����-W�%�W���^[�S[�Wf��������4['��������H�y�u�֖v�%i-}js�� 
,�-��2��VY?��oJ+C[p[h:����MI�2���E��w`�X*_��cP���0�����I  7	�_��ɶ��wL��0�h�� ����'�?�K�|mz
?��}�a$:��Z*�L*9�ZD͕ڗ�����jF*�\��~���m��ݎ�ާ�P��M1������~?j^�����s��o�vAw�J[uocmW7O/ɯ>�\�d�Q���#�ȿ����)Wx4�ov��]
�(��ՙ�ơ���EN�\BK��f�o͢�/��)��wv�(�;�OB�\~�2�{OΕ�$��{BS��14��?��˙���Z�����T]����������W�ŜG�>�M��N�b����E��m�v�$��Jb>��9<]:/�]�m�p�5��@ށ]R�C@��JJ��|
���wTMt'�&+��;��"�3z����Gʖa�\��5|�7!�7GHV��44i��Zȫl��Ǎ��mO*���n����e�#�7	���p�6�(ZV��̤�k�/����j��LDוv1��a&���R����h�N����G#��̀�5l�Q.i�������'T�f@!�
�o�Գ-�՞�^��ݔ�V�s�7�ǂ��Ƞ�htP	��5o��\����X0.�-��7:���� (< ���D>xi$�Q>N�7��VvX��l�T�v��kT3�3��ĸ<o�����Dҝ���{��
nX�Ӈ������K�\#����~��7�z!Ɔ�Zg�k�%&%����/$��T�z`�� Ą��߲yB�f�N�p��c��)a�`H;�ф�
�Hm���KO�����T�J{�L~�L�L��5�(���tygbq���4vNKI���: q
��۠�N��n^P�7���~�ʫ� (�^oAycE��(S4:KP(�)�g��Q�g$�T���6u��-�����ƶ��p~�+&�:���`��6�c�[["��у�����@J��K$o\1�N���k;� �:�V��(�O�P2>N:�#�l�YE�� ����{�9h)ԣ�U6Ey��aAU�Qi��V�v���/�gq+�w���'-�|l�6�,��b_K�>T���uV�t����y�n6�M�����X�#8P�	�MvѵJ�s���7ShҊ_މH �7���óY�Z� ��O�6Á@�L��([�i�]����M�(��1ϹS�[�����#�l������b�}�3{)���j3o�8P�o����)f�c)�gj�mޯMvO�~��@>��mi׏���VL�#s(��2����U���T.�ؙ��G�6֦Q�/�֢
�%C��<�o��PTk�OA�#��Z�Ʋ�	V��k ��N���#���@�J���k*"o*"�����to����[ux��,4@�C7d����!�l�?R7=�I�]�M�-mnA�d�A�6���ojP�Z�&��1_Vo�8�a�vf�{G3��u}����9M;iy��v�;�뻙I���������H���l t6���%��tA�{/�;;���Q��p}(�G�R�mnˆۿ>U��V�pp�ղ掤��R�-����,��� ����sthtm�2����������R�Q��K]�Z�4���(P��b� � ��~�0�˘�A3�"��:��t���<ߟFoj�0٪�X�1�±H���A��4wk;���yU�d��E���^��6c����u����kf����\����Hq3*r��/��ߍ��uOϵR^w� ���w�gqq9��)|A d�=�ʛ%	qc��u�1��s.�"�ĪR5<jS(�M�(�P7�7Ʉ/Gn�@-s6�ւ���o>��	݊��>�-��gaꕥ�� !{{��N�=�t]`��4�uFR�A��T�oJ�� ��tZB�~��H�-YkQ� ���Q3�F���a�}�|�fw�l�&��J[�9q��+̔�וv�T��O r^B�{p�aRG/�c 5�� �כ���?��z��ێ����P��]l�Zui8_�&������d��gC�4Ȏ�4R�E��d�o��ǥL��I1���2�@��J�M':��7h6$���{�x�~9o=i�Z���Q��^�^?�>]=yϺ��`��8ꌄ�D��FV�^��Wed�W�ˊ���RA�b�h�܋G�� D�Xd�f��h�z+js���h�Ѹ-�S ֬5�o��F���>E\X�oG�z��&?�e�B�����1�K�*�9���-Ѵ0x�4 "4���� ����9��ͯගt2�u�|x%�5\��gl ����#�9��vM|g�Y�0X���]pE���yc�ح�.\��,�;bY�w�X(
� SS�*>��H��o;�������v5Jٿ~����F������8���YX���=�xw�2���E8 m��9�:ٵ��������|��8���C��ɮ3}��O��ɛDsW�߷�����'(O��q-�[Ge��b\h�;"�f>l�`�"�@�J�L��~���R��F�ګ�.����Ɩ�o��6c�şVόTb�{z�C����g�_���"���g�T����^e��N+H�m���;�rᄈB<<��&~`R!��7m���M	kB"��xJ�?�P��H�ʢNk@�6G�"ʾ����r��,�@n9�C��ۺV�c�*��Pm��9j�|T�����.�h�W�џ�&��냔_��~k+zZ��R���d�SE�Yq��͚�U���'{��ZP�S� &��K�b}@����\6�y��K�J'�#�ORh�2E)F��g(���f�N�aA�pM�r�(^�0��C�5q�#ZhV���/��0a�<���%������Mf���YB#*�k�8��H�σ~�u��XO(C團0�u�;p��,>�ݴU[�P^�C_>�ç˱x5��x��f�}���ɝJ�����'O�Sg��B^�Z5�1���TSS��Q� ov8c�$E����i���AEq}��h�*�<��	�cB��v\�db%5Xe�@-�ߞ�̮��K����=�`��J��� ���!�a�������79]���y��y��^CN���}��}��}�p29Hll=��U���JrEHM\Ru�G*�Ķ6���r���8ߗ�o7'8����PW��%�W�w����̒ä���@���S'~gl�	������2��
̦��u\��w6	���O��O��כq��oޑ���p��a~��H�r��y$D��F��Ǽj�RXk�q����~������S��퐊�c�&UK����Ҥ+�0-���+����α����.� D���"k�AI�Of��9/�_̢x	V�0*���[ޗo="0�GgE�.�8YN���P��;�<Դ�Դ2�m����nZ���J��������  L��ou�Es��Q�)e_1��jh�Y��Ӽ�R2���l���Q���uG"��[��W�qY�J�F&���"�b���պ�d�=��~�xk.ܧ&�?u{ö}�]FaB_��\V�3�.䰘��p�DS��\�ܿ<�3ʜXX�GD鞟黝iU��X��%�#Yp�^9������ժ�m�U������D����DZ����J���5P$L��Y��d��?>�M��ź���ل/fD���(�se�ܸ�@6$����䣥�f�!����(ج%��/�_8F����Y��=:���l��Ĝ���M�ו�WčtՊ�P�r�?v��ܹ7���O�+���hX�Ŗ�Nq��� m�\ن+W�D�쏃ǆ��j�S,�}u.6I�{ɓ��	�1{���e&�i���1�yWY����|��t��k�kDn�j�,X��Y~;w܉aݿB�:��5��r���k���^g�6Yqp��9��e������߉1䳃� ?	��4'��kr�N��V�&9�A���ݘM=�/��%���RW|}n,O��G
*�No�U��/�J�}Z&V��������9��W}J���Α�e��o����8;�9҅ɍ���'{a���>�(a#�`͇�OHoq[	��!�U�Ѻ{I��ȸ\ɝ�48Ą�}^��x%{�� �~�_
a��g
!P�u�7�̺�u���]ˏ��V�?r���(_�B�u�z⣆8I���~���ܫ��n[��Vh�qL[:sHJ��C_��i,���|�F�㹦�C
|?p���F!ʓ�d�������,r��Ip��l��":m�Q]��0���R��7o��d�hc�;q�:s�h���{6y�UIw�;�K��	�9t�
;�g{*7'C803d+'�����	m���x�H\b����&�������g)+�8ofUBT_�Jgl�铫蔎�1���HQ�ѯ�Iԓ�����}C�F�������,'�aϷQ�L	[{� x!߂ɿ��-᪟%�g)cM�<�J_��,E�$�%�56]�G��`ݙB,��܏,Ѵ� U�����Z���N4���m��)�]�Y�0������*2�����j9��;��e�T"��E��A���sn4>�4��ZN��KuKXuk��H�Ѕ�][�+&<<mCN��O(��
t�7<�!ei�:�m��x���x��<��F�y:-�~Z�W��ʾ�W� O���I�`���y�U��Rl�~���&}�����H�G����t%E�p�@���H��o=�[bۈe�Y��{;~��X�b�=�J7�������wf�]ޜ��I��0��	��{�m~�ٹrO�ؾgh%v��	�5{���t�l������������-�80[`#�&��:��I��5�Y`�k�1�U�q��I)����K��L>��]F����s��d�1����)�ݦ+ɵ/�&��������h�c�*@�" �1c�Yy�Tb��7���J��,G2zO��%��ABc�zU7�w��!#�2��@����1-��7)��*�s�7��8N�8�J����IG��杩U�eՇ�צỢ/+c���ֻJ���ކ�<쓂�>����Û��f��w)����Ή (<��{��wqA 9�X�B����*�R�AE��U�b2i�f�)�'�X�R �a=l}`�=��
/4bz5:�hU2�I�Q;lS�n��T ްe��}k��4n0F�-�/{�U��_֗G��J��h�l���"I�d��&��T9z�=9�̖�e.O"ZmR2p���.�Qȥ���ɰ7��X	>�f:N���p�1���ݠ(�Q�?�u*B��E�CdZȩ�]_�1�	y�ut�TWo�����',������[qcDg�kB�ƥ�S���u%�-��׬/�K\���匼�FX�PWu>��z��~���R�"g+�M�!�	��Z��C��}��Z�l�aG�G�Xg���ߌ3O���eg0�y�Y�Kyd����D���W�(�a�١���`�My[-����tz/�J�Z�5�$<ʤi��)j��4��^�KZ�, {o�H��L�߲QՏJr�v����>�,��D@9��Q����F��$�l�_�^Q�v�j���z/����B<߾���A���=U�9����le75&�A�#3n�e"��{�T{S�����L���Z�j~�������>c�g�O^� ��_�,!E�o���R= zzS��58���H�?��2\>9%�� V0ഃq"��H��J�о���,@\ч�B�E�� ��n�H���E��6��Xp���Ԅk����b�s�b�1G��D�!�ǐ��-2�5�laIq��\7��|e�}UHޯ�n�?�x�	�
"|�װg��I�b�G���;}8i�3kl3o��7����ګ������s��o��b���_w޷Ԫ~��8�bY��0I[����EdǍNc�;�%ڗ9��½[��1~lb1����jn��c͔����(C�o�R
d�$f�[6��&��cU#pD��j�-j_u<�i��$	�����q�$N���ǯ������A*��������U��g�vߤ��~T٘�W���;j>O�ny7�;,�zz�����|2XL���	3t��<�U�}����4�ܚ�U�d��iA�|���D�]�#cTW�X	�7������ϡ�����S��OOD��F�Q$��A��E\�RՆ�S
��S�u=���i�w&OC��'>���������a{fl^W֣gVn��N��n���%�����[��$������RH{k�)WR�o'�݊�VL���g�j|R���w�b��8=�Y���l�bz����������ڙLt��V�H���o�}����%l�e����I���s���?��s��DsNQҼ�e�[�m+�u�ve���ѐQ�'"P�.&u^
��X���)�-�x��n�%�j����j�����)ĩܫ%2;M����/̼�iO�"�Ko$���Fm_+B�-�0*6�e��`��%[M[	z��w��x4|�����8#^�XjA��+g���_��@���IA��Zm�����M�0��!��U,S�,D�Z�d���!��Z]V��m-�jq_�����D��4C�`E	rP*���w��?9�j��c�F�Td)���&�-�6Z���� c�2kMH�62�A�>�����f��FF�`�����	$E�6c�r��f�T�%�����Q-�a���㏏C�D��	�(ݴ"��i�w�p�)Yi�C�Mß�]�?(
<|X5
6ň&��J��-Zm�Xx5�_�ˮ�
(XӃ�g��5h�.�ү���7�뭢@�e��eP�T��"����	]�2�󹧝��3L�O���O�ξ���R�l7�De�=[��?8����Po&au&<��yg}\���߼;x�'�`Dt�ͺ�tH�m� s!]��%��:�A�Yy2��y���G����<l0d���~x<�8�F[!:��]��Xw]jO]�yr��$?��_������I���Q\<��� #�P���Xr(<Vd�~�d�E{��:,��[^l> \�ȯ�k�ѫ�J^B�h��!U!�NȻM�S��4^e���ji��âu��o�P�ǪcU<����0kkiN�oL]�h���<7j�"��NVL����ta#Y滟j�=����<8��L�E�6��H��zjT�F�u��X�b����Mr�{c%wi��i��'�7�W�����5��$�����BO�����~OO	P�I �.0���U�9�>aE�gŚ~�|��[�U%�EIQ�[��[T\���[z/�t�~�_�q��L���+��%�*��f�.��}m�Y,L�=���X�{ϻ]��>'#o�=ϗJ.��L��v�@�Ik�A�Z�Զa��(�T~��5R�,�W¨�&A�&��!���R6 aZ��$�j(y}�*?� G����Y��_��c9C�ךL	;�|�g�S�PɹI�ēξO
���w.`Lcc�8���qQ��J�|�e!� ���ǵ��14�5���n�Jm~�V�����,A,8QN�)����K�[ ȟ	y�	s�g�Z+��j����4��B��ۏ��"�R%�+�9)A�T'ظ��O�b��<p��3��;KA׫/!�
�V��^ȠIO����[)[ů�=�/�E ƊŶ��dq{��o��|�O�5���SK;����(c�݊�.��N�^�BFڈ������U0��vڃsd"������(a{�� �c���k��
��ZS:Y#���H��1Ż��ɽ�h�1��0�KFH?���8�����+�;|�:��u����Y~�P"53����lb<(�0O�BK���aW��ޗpv�[9�����k<��vM��gi�M�7���ONf����}s������<K�V�oq5b�5�g�2��3��o�s_:��<J-��j&2�N̸/���~���2CUr}Ipk:�Z��^�M�2R�hp�q�xd[��.r��`#"��k�M_zj8EK��+k����$�&l���Y�>7j1:f/�׀����� 67��3��Y�m)b_�o�[�oLcC�$��q�kx���$��~�(0��7q�yk�	��ؑa��
�L��b˯�ψ%]��߂.��F�HM#3��������#�F��Kx�`.�x�1�J��y�Nx*S���RFH�"f�����k���ABO��7k�/;(���;��X�ؚ��m��6�L�o��y���P軙|�*��|څ�W��z@�T�������7��W��|�;���0�bs	����w"�.�*ئ��&�y��&��Fr�g����D�\�_�/BZ�a�|�$���O_��a�.���Y��_���X�p^�d�Q%��e-k�����k�QbA�LU�)E֣^�C�~���4��� �*9�9E��Z�mX:�ao~�I�b[A*x<O�&ᴦ�sB'�������lS!��H�]�	Ţ/l E����eܗpK���44�V�T=x�l���U�'��t>��q����No�N��.r�_GD�ɣ����_�ie��	�e%���.V�U�*a�R�����ܮt��c�N��3�叺�o��uX[yT���.׬��a���9z�$G".ݮ���;P��g�{+'t�IC�\V�	BԒ�`@�XAa��y�s��2����WW�s�Ҙ1V�+�o%Ǿ����V}ΠnW^����3��{T��f*�x��^�{"�8i}�f�n��l����[�,s���@lA7��U�9�Z�F���_�mL*N� ӏ�#�aZ���O��Y�i�!��T=��qX6I5��9S���o�I�!��s�R�܆����m�+�e��;5��$��0z��O1U�/�`$����f�<X�6���V��sB|.q���o@���b1^!s�?Ŗ�	��R�B����S^ ����W�_�L�	|ߢ���W?婶m3D�#�%~��X�/�`	��|&*d���>�3��=N{B,k�K��N�k�kȼ�|O)�`��z�K#ڗ�tC���J���� 忸����֖��iR�i�2�gʙ�%��8�5���gR�������������DJ2YNڊ$����t���Y�ف}��4�z���P���W��+-Sɏ@���������֪����ۮ��7�s�&�YO~`��e�t/@7^o����I����,0��2����1�5��ऌ�n^�q�|8h/� :u^���������q�����_���z�8a{�6�K0|�1�jZ�ޕ�k}����@�F�Q6����7庇p�s}�)��KR�{_��|G���RL�jU^�݃�Ԃ����R� _�����iv�°�&9�r.\L�v�9h���	$��@`���
ۂ�YM�E�ا����ږ�!�����8�ڻ�8>q?��V~>C�ǂ�9qk�e��S��OM��lCv�;�~���k�3V�R���Uf5��ln��~7�(��~�Oɺ�-��F9�#%��-�ˤ�i��"֫���U��1��J3�W!L����-�k.;�ÕڞZ��F6%/�!Z<(�p��\�fB�`>S{�Ef�V�ipQ�N����O�;��^y���,�P�^J���:I�Х"� �II�;'�3b����
��D�>X�H�:?�,Jf��ɷ���\�Lۢ�%f9(O�U�/wn�$b�`��g(M�w�y3��*���bN�,�Dx��>�ex�h_l,�i�� ����ȃ�F�Np��y�A4$�o�J��@x�0[́�x��9In3P0�D�V6�gk&����9IxZ��B���v��Ef�"Z���-���F�T�oK," w�\�N˕����,�5���n��~Vq���.
�ۓ���4����x�D�Uo��br)��y�T6@)N�)⚾4�S��W$�6��M8�N81�5���Y�z���'u6��.��GQN
A��Fl�2-�Щ�Bh~�4r��j�I�m��Ѿ��i�S��5r��Jy���HM��r�|�!T�V�U����J�����l���"mbac����|:�j����@�X�}�ﳿ`A/��x�(J0�s�\�����,�g׈�V� �oyӏ�I�hd\ 3�+��_����s�:GBG?�d $9"�8&W��ޢ�=T.���k������b�w����b�b����5;ɥ�ӕ�	��t,�soJ�8�Ƒ|]��|��&mұ���)>��BGS'w�L5�_z꼹���0OC�NcH`;Im�O���l��Q�t��B[W,�ٱ����|ƄÒ�����+�����~�t����2هfٗ_��TN��Y1g~AQ�4&?�!�!Q���ײVH�a2��YX8��G(}��̯n��Z�� @�ߖZꏠyZ ��~ruX�f["{�d��=ܶ�-{_um忻23T4���6p~���\)��]4x��β
!����6k`B�����a�&pҰ>��ۛ$&���d�ĥ*�LI=�r�?�'�ʟ����+,VE��-����_�S���l�*�r2S��C�$�f1&Q�u䨍����}i�p����]p[��rm�;肨[���V΃
o
;�4�|8���-�e_�@;X,��'�K6����[G���I&ڽ;���,��	�jj�hg��@t���hl��)��pj�����x9�}74��;�� ���cSr�Rz^%��8�wUs+d&k\"�r�;5"�|<���d���e��y������[��`k��r�'�0�5���p-� �
9�#Y�Q�E���j�����C����FfݖL7���`)y��
�,�����F̩�X��YÙ��8A^�tk9�l:�����n��ʺ�\��b6�KC�4��,{}�\�p7����0;�m:��Q�����4���ޫ�,��/!a������G� Ш9�䀋��7]�Tzd5�xq�q���U�H������j�I�Y�vJ
����o���yI�5�cg�|.�Sҋ�'ZJ���L/=�B]Ǔ]
�?5����@��ZD*?�
>ݹQ}���	��/���jM��v���6O�o�&^�-�B��&�BV��)�~��:�|����k)�J�i	E�.r
ӫ6�<Kҷ��AB4F��Y��5�Y|*�CI)��4�-�8H����6�dD�������vSfg:(�\����ӏ|�� Fv��~rc�� b�$PbO���mCkV	:�h�L�(&q�"�1����p���� �;��<x�`
�S6���d�5K-��<_�/)b����m�\�ά.e�lҶ{ɽ�n�+W��k�S�f)�%?`��d�a��%��r8�sc)�@�� 
� �;�(��AQ�ٕK:���EKxJ@떥T��d�飡v���n��motU����!O೙l:7��me$%&���z%q_Ί4=�������B��U�A ΂*�q�	�>H�p�Rz'!t`�zy^�9 �B�:ݖ��gtC'�Z$��g��Ÿ������`����<׵��s�%�0Q[���.�CIb�v�ֱ	�@�/6���M3[���	��~,�9�~�����In�;�C,)#�������2i:�����~�92�
��1�y�ε�{ap�l1ZO����j��aK	ߨ'̈́/Âa�A^��l?�kxɁ�	J�1ZfA��Rq� �Q�	]h�T��S�Ӑ���.��K'��#P��Єn��[y��DE���Mo�|�_�&gB������V��1��3h����HN(v���U�e�&}���垼0
(����
K���X��nl�.�?��Z,�)���0/�)�rMFUE������8��kXw����7z����z�cSS&,�,�z{`Q����A�kE���w�/�\�CزQ^O)��Sy����B�k���D¦��,����4� }���݀��b��-�����#����ab"\�<nH=����L�M�0����Y��-b��%8�M�y��6�]�zB
�ǒ�i����O�������,{6����~;V��r��������(�G�1��u�4���pLM#�q�0�L�u���唭i��3�M� I4��4�`S�����r��܏����ѫ�m�w�-S���_ܷ��=C$��Aga��]r��ܼ����O*��6-��Jѥ����/&#���k�{6VL.�v]1��I}G�1���e�J��h�C�i4�����i��i��m&��V���}@���-�mѭ}���Y�X/���i�Ok�'�UwY�W3+/*�s���ã��筑PyR���<�5���PxH�EP	'������s\���R#������0��������Y��|�S8�oZ����gj�z�<Z�[���W�b���}��~�f�9FF�`�����xJ�u�A
D�I`��`�1	�v�Õ{���n"�^�F��Z�H��i�g;7�n�_�e[�S�&t�#]�7����ھ���V��!(U�����j���5^����-.���opw	P�P�ݡE�[ ���Jpw���}����33;�I�z�u���Y(��o��kG���7�U�hY��8�8�r���X�>��^6'�Loh	ފ������z�Y�Qݰx��$uk�x�b��D H ��
5k�	jM` �	\�79�` ����O�ϴBb1�]��5��)I�� �a��Y�E��\�q�6s���;;�շ�*q~$U��`v�T�)�fV3 o���s|o��Qo��`�֨�%�0�\*�*�Mr�Y+c����h����,�4?�E�`9�N�V(ilkݷ�8�t��:s���o*��ٲ��3�J+0�R��$�6 ���o���e�(l`ΣO߿5bS�B�@��a8(�Rg�ހ@�3���G�'0g�p���)�~�ͥ��ɽo�C��:)D�� s���jH��������z�����P���Q�w��w�ق�{2oT�g0�נ����,s�EPu�����ZX��^�g�Y9�t��ݺ�����8[��*?߰E�{F4�K`؛�v7�b�)�&(~�t+`�E�%W�=�x�`��/xS�t�e����8�~䱜bգ���ˉK��j]���UP�U ���)g6Eg�Ϻ�Y٣��F7�w��#�4�/J~XAၒ	��O�l�����Λ��OcO�5��ڹ�'*���Av�	�U����57i�e^�F$� @B!��V�Bp���ɵ�(b�V�mU��f(�n�y,"@S�D�ןV�{5�B�+�����_n��x��|�;Ux��y��p��y�$W!��K���tC���;w�:�3����$�!��VG��_y`D���0�3�7xT��μ�*
`8= ~�m��E���r��KA'�]œP��L�F��`M(�/57�� ���W��90�JDb�^����� ��R��5Vj�ӑq��wr2�_�	}:�{�x�/�TD��8��7�hK�e�0,�~��-o:"���#�֒(b���Z�7Ȫ4��J&�~�T�ofzU��%t�]���a}k�=~�:P����K�Gn�^D�����w^ӵ[Mn�XXZy������Q���&�)�X	1�H�%�:�]��b"?�Lez�+E��:9�^�G}h�o�އ����Z�2{��͠��K�x�����������˵U�����_��u#.�C2��:���
a��*�L!s����;?��ѷ�OFk3ύ~�Os9nǯ��lةm!2�U��{����t�x���͎��bGqOL@B�l�jG��T��!�XN�˄鴤��r��jF㣘E�ko~"(׉��m>�t�;,/�x�R�*KT��C9R�^]�Z�m�Ш��ҙ�_�U������� ����ȯ��;:�;��2A���U�������.6G����H��9(�������4�G�Q����`�/�~p�ck�0*<z�L�o�D����K�ӏ�-W���3�d���v�W)�s�F�xs����TV�{�ԚJ-;J���k�
ӦT+��U�IV��5�L�D�@hג&	�̕�����7F���$8c� eT���k�t�MU���˨9<-3�(��ͱ�<�	�˦Ը����:�q]�5�L������0��a�Z������d���"xK�5���%,��/�4ۆ�_t�·�~�,�"KY`.�$)8"%��y��G���oVN8�8�#b8�)5@H��]M�m��;tJ�v��^��*#�����槀�n���n����)��)���NǾ������m&�ygwN�J#\���E���o	o��P�A[d3NoQ�9e��jy��Yg�J��:\���z�r�:��׺{�E4����AX��������m��g-)O��cf���1�`׵�¬��p�l�,@"WAq�ߟ
�0\R,�K��\"w۬R�E��g�i�i�`�56��=��⒖�.�'�0���&BH;����?�Ȧ.�T�CP��.V����3����C��aA��(9��q�ų������+@Y	*NT���/��q�o��Á���JB���뻽^Jۆn�=k�2;W.	,M.�?�(D�tM�޽�8���D�W%*Ɣ���5�����VBOd�yX�nv�{����Li�-����R���ޫzi�#���צ&y��XoR:�f�!��<��7S��шّ;�N:-;�/9G0��GJ��g	ω	e�W:zXʭ��ݔ`��v>n��ݏ�=o���M�2�ȑ�S���e��1�:�ɹA9�@��br����
��
��
�_�q����N���S�g�H�����
�\���\���+X��D�?�O�RN!ju��e�{��^�Ŀ�u������Bv+b�Q�Z��o���׉�P�|��TdQ���E�R�ᷟ�1]�q�s^�v�n7Y��0a��5̍B��|P�H��E���f���̓�-���˵
��C����zT��߹۵��'1Fq���zd���;Cw?��r<!���־��8L��J����d?{�>�l�?����ݽ
뗮,,X�|�YSM��Z?��kUH��[R�V��D~�����	���İ�9b���`�΋sQ�,M��.�iwb��jF��-ɀ��ې~}K�nj�%�M�^�i��ַ0�%Ʌq�lO�*�bz����4%,��N��b��x<#��]|$�4B�3���ޛ��EY�$��]�o5Au#[cH������c� 1�� �o���3!�܌���3��$ȧe�Y�!N��T��e�b������{x[�������P�7������ҝ K�ó^�x����|MF��X�)��^�-
�
����4
<��=�=�:���""��8�?e�$��$�$J]Cv��l����K'��m�m:��*��=�Դ�h�����8kx�3����F�S��{̹]̽��n;+)�X�@9BO�hSk�� ����ؤ�&ןG�k{� ��N�0�#�E9���UѫMz�X�<�l���Zᖈ�K���?dz�ra-��C���G�bdPY��T:�[	�!�y��u��}x=�|˯8��Q�?;�\;��)p�.dMf�<=��6E�xL4!%�^3j�#t��_�qJ����z�vK�)Y0S[�����΋��C�T�It��%|�U�������t�X�S=h�>o6F�;6���1�hx`��qGx�&�(i�BFA7��|�����!�A��ﾻ����wya��AxME�C �p�x��7����6t)_v1�?/<���4E�����[����t����'��ri�`��`�|�ľ	�:��Ln��z�Z�W�|ݐ���Ԕ���h�%U�H�j��9[���3M�
��ְA�
t|G���t�34Sޔ <��Ʈ�s�XQ֒߬wj\��*w�e�S��
l9��v�j��>�	V߱��g/	'�q�A���76�����ˁ����deʾ����*��z���:Dl�[�=��:~�j�S�:	�53��<֟MX���BPv�-��=Ng{�9t�?g���}{��p�A㟢(�Zf��~�n���� q��3�	�
����|%gd;�P�<��~;��Q�)s,��Ţ�� H���=]Z��^t
Qt��76������nS��{\Ȭ1Ȱ����}���6����Ͳ4\��??������
�"vm�)�Q�d��h��cR��t�YRKR7��RŽ �rF��U�U��e�N"���J
���e����u��u�8e��\��ӯ�9�\��$]oa�a�m��@��2|wb�ɕ�$�y������)��L����V����4��f߮_�k<
��`��}�x��k�aQ�e7�?���f��� ��[��×R�� �4��f�q��ʴ?i�}�������dUЄ�sO�l0x/��+[�}U�2j[u�W�u-_����ę��1�G�շ�Ai��H)���ϳ�%\��o*�tB>�u>��A�ed�)M�*|�D�&5��̉���(�����%ƌ��C�=��җ���A��ma�k6���}_v��]�{10z��|XQH}w=*�7#~��bV�e��5,B/O�Alx�Fq�"�j��3N�8k�9c�呄�`B Bj�l��D?���
*gM5��HW���N��N+7UO����3s:�b���,�Wm^Ü{RE��)��sɊ���Y���&���FѴ㈞��X=ƶ��ǘ�D��ץ~�2��H�
�1��|Bo�G���n��=����)���PO�2CL��P������޷�jn+8���6*#Z�:��,�A��h9�dp��Qk�1����c���I������~R�����-�,�?�	�N�g��v��#�hI�0��+�.Y�I�o8���"v��k�w�4�� �(��7�t�s"D���&u�8%>��n��k`v�ܿW�$R�ʵ���h�VM1Y��e�qݭ���t;v��:��(}���WtS)��1�<xM@��o�@�EL�����m���� X����}�ݞ%��9��C�q��nr�uэ��w@��>����uQ¼��	m��1h��1�����[�8��d��`�����L���V$e+T�W"v�o,��}D<����W"f"�����2u����v]w	��c}�\g#F�\��cY%lGFZ��wt��!�&B�jī 0�,�ΛSh�2_�JT�	���*�Q.z$�JL����H��#�U�A��	��TEp2!N�O��:��K}�^�-��(�M�C�+f�B���Q-%9�zw�UevcW�pD��s;��잉� ���N��N��-dW*�����xܚ�KP��ㅭ;塚@+�B0�\�%��0mS7S��/��z��?�wV�Uq��Lؙ�:XM�]L�\�؟wV���U��ΓRc��(4�����#s�P��7��[�i�Z���E�����z���T�/�1U�ؗ�.=xu24�F���X�� h��I�TK����'
��D���L%�h�h΍���f�[��Y6���آ�ھ�$D�nU����,g�򜉮>v����)�M]||�3���ێ�a����˨�J�qS�\H(��&X�{�{�ӯQ{q��-��7��)��={�r�Y��VѪ��\y�aåg�s����\��׮®�D��°~�Zգ5�$�"._�Z��u����:�*�&�ڥ,7�:�Lם@d|�m��:��u�&����;�J�L>@���?u.�)��Y�sm��[�3��`93{� ��IB�'5*p�uĈ1(�1F�l"�Fi�%�ɢ�E\&�Х9\���@�ݶN;zA�|���RB���u
�����(GBt�> �?�=�MGt���8������O &�vL~�P�8f,N0p�k6{� ��Pgց���G�z���Z���a�a���8��|5���|#Oϙ��>uw�������Ax��b��.�7^��Z�m����� ?�q!��Iz�������ᛝ�V����e��f𥕆G�&�� ���ߔ<�?�%~�p�����r�7�1������|��fn��4x+�z��l��r��L(|����ɿm���F6 է,g�ԛ��J���@��݀����?�	$�	�/�-k}��"ߓe����˻j�A�HǇ�'x3��v�V
�`��O���U=^�«�y%��	�]�f��,vˤZ�T�-��ބ��S�A�����`��Yy�1iҳ�Hw��R\�z(E�:�$]`�s+w�9ɢ��EHyuě]'+,��v]�ϟ���Z�-_���,��~y�F��CW�{Ŝ��������0y69���ϯ$��Q�H��t�E_$��f�s�yL�����
L�}�a����	�ö�������Pb\��[�5HF��c����[�.�3h�-�x�������W+T	䊡q!��] ��f�w�{5r�g_Íx1��bo����?�������)P���?L�m��enh��-pxpX���zRh�]gx�<-t��ūe��W��7�~aӀ�E�|B�}4�M��x����os.����ASMr�%X̼�9��P�����-�{u�Ȣ��3�*��Z�`Ki�=���OHw�� ��ޑB%�W�;ԖH?< �<���?�D[<�h�J |��-vPHuP�=\�g#!s/oQY�_v��qXŚA�+/a��������r �R��>,n�W�`fz�A6ٺ�f��t��}��B�'�G���
���dC�4����+<��֡(E��w�0���C����"�:H�@#���0(��(���j��{��W�B���፯�{����~�@�_z'�8 �n�"�Tp���L�=���%O�1 *���eD�����s�XYSl4m��{W9�V>5�k�4M8��N�&���}տ?GAw�e���w���:����.{��T�;�E�j$����}V�('�[���ƈ�F`��O�萧����?	�\֪S	��g�J>q<w'~����k�u��ٍ�W�Ms���t-�mhf793�1Q#��.[[0l�P��E
���Y�jjG)�b�-4���R�%���O��01��<z����㊚�(�R� ��Fˉ��]��ˊG4v[��r��ޱ�s$=6�&3�̒��&����cUV@�Sj{Q��.�QF?Os��Jg�R�:���o��.Ug��O�Kr�Å��2މB,?v�!�U���S0����I��`��Q�����9jb�b�;;f�Deޞw���oP����'ΠK� Uh�%ë�vK��3޽��~�jz.�)T/���4��"�}-������6�M�Iת�`Nf�w�>J�|g��c �%=��~y�K���#hz%�B2M�-���e�z�֚��T��!P��^Jq"���s�$̊_��k�V־#�Q��\�M���#>+n䍓Ǡ~��ʗ�bA�R�b����}=�x]������H)F�6�9P���џ�U޲R�S/��5eX����=�{��ԙNڜ�<��dy_$x�hI񴠥�Π;�0@�Y��ˢ+Z5�[�*�B��{���/S����§��������q���N��g?'O�!�U��#�N������ґ)Y��R��}ed�GO����8l�JI���iy�x�_xڰEڹ�s�q/)%�0�^���Y�>D�����#�$=�����&�9XLw�������sS�]�����n��i��a{/��P���%j���}�wy*�ԏQ"E2 �]��k�
 *���h��q���o&^�C�͍^�����l���Q���Bɋ����Æ��Ǎ�6N�n��6cu0/���2qBA\��״�g��W�l.j�8(6֭/���)�7�1�0�
�T�`��?	1�F4�~� �_F��/3�@l4.�`�b�ԕV���B81�S��p��d� q�g!���և��w?�`i"��
�U���=�1��rjԺ&�J�Y�YM��z?��Y���:"]��|�_��/�PP��B i/N�,m}�U�y~�S�r#��S���l�wt0���<04rc��V4��G{�`��̕�Ԇ�y�'���eR[�g� .�!(��uxǢ����<u �z�o1�{��2x���������bJc=T<�����U����W#�-L�FK�VC
:��3%�:�eh�b���$<��dO�e4O�M*y��v������QxzFW���xF���㻟��ڃ�8t��,��ol��_L�=�T��Ff`w��B��^��l��U��U ��������z,����b�����댫GήY��bL��8�[��S��@���(!����x�`{&m:��ڥ�e?n��`��p��@��F��!�(�=O�6�Ǧ�!�G��X��T��6�%����X���ӇyaG\�����{z��\�[�����D��V�Sr���C0t���$��PܥN�s1��eH���Qc��+�V9�\Y*����*9x���m�c������8��#�����4jS!F�*���T/�(��;��V=�Zy� �w��oΛo}�V֑��\�/��~�S3�S+�3�9#_��׋IuU��5�C(�$횜+]o��ด�C��|�����a˪��2i��ɩ�	1ڻ�;hs�Rsȱ�n�ꆵ�9��p�,����m��b����lӆ�M9S�ʤm'����U8?�kk-ߥ����{ˣ�����ԇ��{��72�����P�)܁.�0\ul�T���3c�78�3C�C;	�w�C?|o!�j}�
`�CK�r��.?�=I�@� Oʏm� ������\{���S�����u���!`^���P~���C5i'S����t�e(;:q���Xi�{=ol>�3Թ v4|U,Jj�������-�߈F�/��{'>�'��� �V�ΰ�?n�߮z�x㣯�|��J�گ�])�I���#����\�w���c�����
�'&�I� ��m�hgbx��Ks�/�G���	)���qC�u�k5������Q�*��*���B��LI�r�]���)n]Rv~	P�'?e$�n��`����ɨ�/�$z� �B~by$�W ��x�P�`kC����.Y-T��F){�Ҟ��CIv�ё������o�1�N^�5���F`���-�q��q����PD�P@s���X��A�'X���M�5X?;��Ö2����w�T��J^�^DEC����9w�� ������+�9X��
�v4S�;�:66t~P�t�fe�P�}������;�w�j?O�sa���P���/J��e��S�,�8RL��fWE(�c:��(f�TQ<��\1#��@�/)�W����6�,3�M�Dw��}�y��}��>A�M>Y1�#�6�w�l��	1������a7��Ee��z�ʋ�*m��$���u�E��E'�w�o�<'�<��ݦ���f��ڐZ�j%Z�G�����Q<פ���q�R+��rXn��+��O�	�Y\L˰�(R�ś��F��"��V��R*u"dNIw���Vn]�	W�C&�Y-Hэ�ÉG轂V
<�(�E(���f�u�����GcK��;$(������Q��9*�B_޾��|�b��Æ���E^���=���>�Eb �~n�\K��u�F�������L?�;1�N�8�N��sn�������܀!"�X�\$����������Ts���O͊����nP����1���337.(����,b5��ʨeX��$tXWD�H��-�TM���}�$Bp�5���5���bL_TM��촪n�������J���"��wMm/ ���(���Dlv
5�ŇHL�b�(贯o;t<�S�6�)��,����M^�FYCQIQ&�}����o�T�*PS*��5�j�j��W!69\�<��u<�XW#�V�"�m^���S�?0�����W��·o�mUy��k߄7I�7G�7C��@q6��O�~G����NX�E�`��3$��&Yޡs��F6w���.x��{?Z�T��� ^�.�WD���c�Y���/�i� �����	�ь��vցj��I�u��<?��x-�v-�{�MG~��u���maň�aQ.��i���d/���
l�����Hc�*7���iC�m]�YSAa��6��(I4�	�ɣ˱�Jz1�9FI�-����ܸ��~����¨��Ò�Q%���u`��߷��#vQ+������s�ʗ%��_"��*�O�}?l�xT�+<)jߦM��?%��Y�����"���>�;�[�\�������v;�h]��CP,�8�1߻ꪇ}p���2�8,gkwy.�ݢfߎ6(3�M�ް�VՄŸ4T�/�E��nc�FC8y�s�Q:���-��F\G���b�V��C���7u���8��Ci`�d�b�	h��Ki�K:P��2�-�1;��W	*N�Z�9e�P![��mժ`�Qd���z�Yy�31��<)^���(5`�VNb�Cq\L^�� �Q�g[�|-x���!�M����~�JEz>��]���v!������%
Aq�Z�UO�~��B�� Q/�)���<t�Sl�cJʨ�;7�c~�p	�
�b�F�.�U�>�K���f��ـ���-�h��J�ѫ��>��:;�>s�~lh���ZM/��Ju6�*z�&z�* }��p�0�����Ym�InsjRm�VB̩����3�@���`����5̝�F��"g��y.߆7Vfm�q��� &��i�N��uP��Ң�D�Km/g)I;�k�3�KVL�H�0���w�)����N�d��w;՟w�.���CB���y�� ���%�O�;6���Z����j� "�|�Nܼ�	��<�A���چ�rAe]�X=��A���|�y���ojN�У�ڋ���O\��II�l�7����W�&t���
�4����������B �WKH���f<�G���P��6Ui_"8=�� �hE���	^8�1�-��LQɽ���7c M��]�*�79).
���D#�˫�N�[ܿ�2���ݜ��p�KԻ�ϧ֪��MN��a��>\j M2�Z�BRv���a؂�9���9�A��TlN5����a
� k^�ޛ(b���с��\��Ap|���2�/���٬��()�ދL�-��hrf~��/CՈ�uns
��)�2��]ޫ@���"��Cģ��,ϰ�kd���Gq �߬����E9(��AT���e1�����qǥ����:�5CnaR�s�#��� ����Ǝq���ô5�t����z�B�egSk���mG�݅���s��ᩎ��S����D3�V�.��V��P�يަ�"n;2�Hw��7 ��b���!����g�q�-�Om�'��r$ݸ{��J�����qܴ��9[{�����A�>�%^ i_�5��mC�«�B���g`宱��HNDN�b�$(�^�m_�a�4��<��	����f5)���_��avJ���8t��i���P�ņ�<:��JR��e��U�:��z�6c���g�5����&Dwmd��V��E;����V�:V^�U�r~�r9G������jt7�7�4G�kyeP���6�{�3�(N"9��3�ʵ�\z�Uc�Ni�L{������t�ph��
/G����Z8o�ʥ�k!˱���=s��� >�G8\��C[3�|q��T�̍4���.B���\�:\�6\I^�ަ��V��EM�����Ir�"�F�0]�������7��a^kTc��A��Io[��;v�ۀ'��Ӿ84����ګ�E2?vQT�s�E�2H����9��gzD���:���4�eM9�QQa�%��BB�M���9���t�4�c��
h�՘�ԉ|Q�������l�QK~�;q$Ò� f[.B`AfP G7��?��J�GQY:�3�R8�㙘�N*>��0v��f���z'wv+�V����@]�ƙ�(�g���_N�^�X�o�o'�x�KZ��ƶa�8
�(H�9	&�Ax]�P�8 ��ꝺ~c����j�v��3�"�~���m�绻��~�au�A,N3�n�}(	s�Q�����GQp��Rb/��	�W#�_Cgۖ�U��������մ� �L�nDf�Z�NP�������"��,\�1��t�	���n�7�R�m�GI+�V�G�Y��	��2���D���2��Bkpv&��Ҳ��o�t�6��m�&�<H��|#��F�nO��#C�N~b�z2F�8��?�f.X��N��R��0J&�
z�d�!k�%��	R�vz"jAwM�~_G)��fX�ERMǚ�?��s�X�����,��ڼ�ǵ�|#��m�����,d8�q����_A�a���W���4?�zv��KD��s#}��f���܆�ř�-��]�F�`�������$W����`Ć̅̍����I֋2H��4���KI�	te"�ܟ1(���WoErfv���}�Zj��.�0(�OYmz��G� �;��������c�Z3e,��в���W?Cnr�!��i�?Җ�>�T���R@�#p~��Y�5�I���t���Fl�P������m8|bkf5m�d����-J�ޏ�{�Uj "�8�[uB����F`��x��^��K��K��m���k����)���"n���tw�v�8ta���d^�D��$�D�7�a6�F�-��v�"�I�X)|:�}�p'�����j_$������&z��s�҆Ƶw{�~	�����h߲�"=�{�{A�w��+��f8K�u�T� �d,[;=�acq7�xR?��|TD��n��Sq�*:��j���9,tgb�0��w���aV�F&�TF3˞�D�L+��2���HP�d!&���⩤���T��2���u����������x��n������ ������V���]2�cϝ_m�xMAo���<�j(Ŕ�� ��1�K+����I�H�MW
b�D��~��0�O�����\���i�+�;��f3�ީ���{�RRq�-�����G=�b�x`��}�ӷ�s_P�(�̃�b-���������ЭT�:�;�S�*�|�EZ�3���á�������2�p(
���B�Wj7����&_�.h�3	�h���i15C�ȷ������և{��FH��?[2}e���qA���Z�������K����	U��G=+i�7�ggl�cW8.'�e�d�o)��\���[�c�[� �����j���We,�
��&H�~ضB�R�p�N������8
˩���@Wa��x̳_@�H�pg�Rw.b�o��W���\7tT�?"o6v�i�l(�d*o���}[�p�-�2�7޲�LF��ڨ�*�I:IE�½(��@Lv���p$���Ɵ�׵��,:�bZ-E�f�C��4�>^}R�ĲS;�WEe�dT�Է@;E�W�(�6����zLӾ��<펈��3bfк�ҊK,;���j����Dp���c�d�i=)N$@��6�{&�\JE���n�v��l��5�Y5���+��^L*֟ +J�#��P�u��}佉&Ĵ�ڐ�Wly_�u>�hu��Xe��ꥒ�g1Q/C����l�uhv"i,$���T�;*3H�!(��A�&?�ċ���U?�����nH��oV�H܆�~@
�h�MmϿ#T yւ��W��+��}�Ug^��1(W��Pѫ>#Wu?���v�o�A=�ߝ4�Ma�ϩ�z�	��M[iZ?<A�#CsYP��L�r����&w˰���hGlX'�X!�F���:��L��2�L4!��������+)�XL$?!	����YP�-�#�Əa�@�_�H���E(���X�ԍ��ͭvb�Yl�I�1�6	/T�OaX/�#*�Z��/UBq,�#j6ґ|�Tw�]wB�-��?��d�W
Xj���Aat����Z�LN�Jn%D�糳��W�^���
��F�+�6Ae��$���M��576�}��A-�ds��{��'=l�����BI|>w�a�|g=N3�++���s%Q�^���y|#������ �_�u�[�=0\�꟞z�������\�U���̭�\��{>��b��|�6�տ���5�R���ά�5n�q�i�)��_��hbHX� Ŕ��Q�z�JX�6W1pŊX~ݿQpAFA<���[���c�l�	�X	��wY� ��H띁Q��[-S���;ij���1�W�iTqNq[��ơ��P�
�a%Z���j,�M��SV��E�M�G�%�6�!.�$)�lf�A�	U
Z���R�!f#����Şف����{Q�L�Yn�S���!i�sS%
�v����E�m�L9K�QЫ�k�T~VlS�5���q��3(�����Eؙ�~�лi^�����4U�<�D/EB�"��[b�T��M��H���U����Gخ��V���0qfZ��W���)��
���A��{�Sr&vA��f��f��b�+��qe�Q[�+R�𬝀ZYmۋ�&���v���6���So`C�}�"��¤�m$f���|q�3M=��|rU�w.*�$��V��t��b��7��(��C�Zv*S�ޒC����M��?��~d����:��2t���Z�D���g1�J㝍^�$qL�'�G�u���!;
��ρ+�R{?��X#4%�����P�����os<�������e*8�1�Œ�T��%ԯSH��r��!$܀v�)�BNkPC���$�"�ГI���	���x�L�01�d����MF���"kv�w`��K쾗�*�/66a����N�9�$# ���͏܀���۟@��\��N��4܏jUK+�I�*��W�Q��}2Q'=�.�����!ƅ�mV-�|�]0�{xm��2Ưr����+$�x7���o78����N+��_�݉�=����/!�"�H�~�ڻ*rrY�u�%��(���d��6��7����ᠯ���A����}J��L&QJ������K�\�;��ip�ʬ����)����������͇����m�$.~��e������>�y�6u7�Fh:��T����%�1#����;t.����B.V�W7Hn�rU�2j豣�e1�p�u�Պ|�oԣ<��Dգ�ܬ��%��	�щ�o��G;�1�ot#��O�����q-@֧O���_-�cN̲��,샚��(�҄s�k�:<۬$�ъ��c�X����B�5z��L@Uڧ��+N��Ǯ�����Y?��{��{���k�绣�ǻN���3
�7�;5�sӫa�Fb�V���rKW�3c�� ��YX�uz�`p���� 5{H&K����3
K�gu�p�UU3rA���_ì�Hh*	S�nV5?�5
s���& �B�N�_�#��Ý��.��O�`��@����,6W��b�Al�R�Q�s!��V����s6�3hUᬈ��(t���j��ںE��5Wh�53c(z��|Q42�������M&�9�j��jk�ݑl��&A���=��U��cCT�������C֝΅fT��QFF�b_C�67��?;�<.ٵ�!��f,�a��a,|�l?vy+1Q!1Q[�Fh����;�{#Am�r~������J�J��3�	=�W�<��ڕY�ͭ��9�&5gm��*h�p�� �a�Rq�t��&�:��~ʾZʶF��^�{X�F&������/�Y�B��\�[ii�f�Ɂl:�$�f ��N#�L`O�o��������/g.�GP�ٳ���9�Wr�D'���,95T����ay狈��L�,	t@L��B�ļKZ1MFr�Xm73�#NA8�(o�k�U<"	�kP�d�;V���?57d"�A�zJW�t�z�
FI��b �Qcݷ�#�Sbt	�Z��є	��.��/|?�?���Dz���京Y�W?# Ą/�#�#�4��VE���_+,1�Kί����?�y?-Tv�����`Y��H�rk�x�^��\�7�f$��F��XȤ���gf���&�'��.�&^�TR��
fH�@�[k�x�����PnU</�S~ ^�����>��2|ӟ�Ū�P���XWH��@���F�V���_>��Ų�*�4$�?�����o`�gd7��oo'���F�<��os�lZ�ƺ- ��ϋ4����~F(�P��k�����H�Y��J|�˗бڱ6�L8X�O���E1�r5z�m UY�!Б��O���l��}�M7�ɀ�K��5�������Y��O��m��^	/�DBɂ\���w�ѫ�0&��Ta�Dyt�M�-m2Slk�� =��TpôH��sͥo�����}6�Q΃SHH��v&ξ�`5�j@,y�<���swqB���d�vV�}���^��Ǫ�1}���,�����'��QP�	ଲ2���	aM�*��*O�*۽b���s Ҏ&�`�x�0<�#!�;z�W�w=u���򊱝����R��3l��}2����L����Ou���9�:��<��s���c�V����U�C��US�q���,X)�����]i�J�V��g(�$� `k�?��7�n�w�&I��70�l��;#��Q�=yr�s���V-�ZM/e%�>���
�H�^I���!�[���	h�7�m��km��F���eP���5���F4~�R� J�|h��,	��>�h��U{��W��#T.L����$���T��R�=��K���V�*M�؏H�g,0���)����Iwc��İ�XI4dލ�T��N�'
7��jJ���O�ӟ{B��G�j�/����W��?���R��ҫ�e��l�[��֛�4�dX���d�)���+���T�@����ܶ)J�B�@��@���76�׶�o���N�&�	��ƺ������3���YR0��)�G����B�+Un*�̔Y�k�YA_T��t<��}*[흴y��@��ۙ�1%X�m�z����j���vqw)�w	����R�x���N�h��P�����\Z�ݵ'���{Μ�|��C�{־���ޏ�h�M��o��;�ʔ�9[
N���kY�p߷���X��I����ĝL��Y�-}��ЃM�ѻ�}����� ���^�u����6E�d!������"c��yt%f����P�����~��}�Z��B�l�h2ŌU4��Y=��B���e�䰐�b-M�Bu抱^"�����b�_��T:E�Z=u����}^��]��� GT:fԬ����寧�+k>'�<u�ղ�8ԓᕹ��e8�((�c���R�Ѳ�"��!7�^�ǲ��_x�}Nq~n����*?P��[�7(� ��w����*8�:�`��%h&���!��:�ʘGH�7�&�j�N�&n�vD�t�<YY�U����yF��B�k^~�����\�e��ɰ����ތRgu�@8?�YN�٨-���.��S~>�;Ug�É���8X
�`��}y��0��y�{���͑����k����趧i�����UX�������$�����->��{�3ʆ�)F���͊ݠ+��@�	%(y�S����հ�V���8�P:�b<Gk	'��lb5|bV��Pp|�7�9rr��ȹi�ᬋO���pFY�����ʵ���we WMPa�]N��W��������i�����Ca)��FCK�](�K�Va�#i;�x�p��|�r�z	Խ��;��I�֟��6˟1-h����ޖ�"dEJ0J���!B���R����)���!���n~?��ß�+�e�Qo*����{�a(�=�����c��c�]AY�Dn��Wv�T���;գAvvx�fl�1r�4��;�p�������!_}$4?٥@ 0Ջ��D�N�;E��#��[�����ۧl��l��;)0;sW�PM� \�wk"��oxm餍� �e�l�r��x��ma�ú<;�"z'�e�u�i~���+r��~��8 ;��_%�e�� Ԯ~���©ܛ�m��@3rQ6Z�Q*���ɗ~�ʈ���؅�����u�YL�"Q�d8)NB����߳b�L�����V���urLj�qwS��*�+y�:��e� ��+z�C{Y������ �N36"�3����9�,�
p��C�������|�*�AzD�#��յ�a���j���-���>5�Gl���`�Y��|��}u�}��}��x������y���L�	^3�?Nw.���՝���~��}�{�`�Q���~e��@�%�O�r��@L�Ή����Y^�	h�Q�>����I��b�=�GSM_)�bD� �Da;k>C1O��c>��{T4G"��0�>o*��RSK�X��n4�Tl��1�!N����B�M/at�@'#�E86M�by�Ȟ�H���fC��i��f�Կ�䢜6Ì�)6n�-t����S%�	�aP�^�{��d�L
����V��QF/
~�P[r&X���*-�!�x�DĦ|��R�J�٠�D��S	W�tme���\2�4�&�F���J�C��) ��p0�v@��M&�]'�;mcno�`/���8�}�~[g��c����藡�ζ%O��TaNBpƟ�w-�B$6A��[�M������y�B�T�e�]�;rI��^���/���:�Ȫ ;v#40
W�1+�@9�*!����aҊ�ѥ`�l[tK�Y�4���*�E�pu�PҔ�<�����OS�ze�)� ��,X�`��פ�ۖ7��G�LxÄ�DҰ��a�ц�gS�L���V3J���8���P�D�?LoB�r�O_>߸Rͧ���%��j�!�d����ݑ�����&zkQ�52�j$�K�̛)�S�V��}�ec���Ľ-Yj���2Rp���iN�=���]�a��7�0�QL����ts؏�
�[�1�L�x��)��u�m�ю^o3�V�V^���7�F�p� uZ���1 m 	��f��lm�}.���)r9CWT�hf|��L�����.��V -�]}�N�Ȟ�ϔ@�K��Y�*w@��0A�������e)ke����������e9ge��SS��bM*��o�B�=���?#�#M
J.�ISI�\�"�*� -��!C��/���c�<	r,w|�l;�;8�[Z6���4��/p�KO���"TӇ��ʭ��O�����y�S\�X63���� @p�7���)��2@sA���SZ�&ziqB��Y�P�;���a� D��T���ݝ��p��;-�o|+}��:%
�^c@.Q���eu�Q(�x�N4�^*�^s�v|(�c(��
њ��|n�nD�y�"FH�+H�w��N�M����X��x(b�$Z'�
B$�5`��*J�K���W3�9v䴾u�V����I\�N�B!m$$G�c��WM^k�"5
��DMBA*S��x�͞�h"�ٲ(1�!ٔ��k�W��XU�Y�3u �O���f?>���W=!��z�J�u��*/^#/^�&d��L�.�n��g 3��^tmf��������$r�r1���x��c6хl��l�~\ҭ(��7Ȕ����xM�BS{��q��&�_�
��"��9P�_㌿8ڿ������ե�7!g�JϿ��!��?1`9[��V"��{rr�q��h�Du��e�M���
���:4�j��χ>"}e���>bW�#Naz��ӽ[C��ù^�'j�[Ư��QKܝFr�D
U��|��ǢႮ0������[Aĥ:JhZ-e_�-&i��=��D�_^��k��ⴓ����&NX˗7H>rD����n�"��_o*l��!���D+�O��D�4�-l����<�eƵ4���P��>P���\����dW����.��׸���X,6��e�����ټ��ȍ�c�ZW��wTt�k����DL�9?�w�׾9�z���T,�	xX��K��M˼.�&{�v�b5�|����o�Q������E|�z���+�ȶ�5LL�Nd��w�&J��B�>/�� �YJ���/�<0��
�C��s&,�s>��D+w1��yB����v�P��3ĚO�wx�Z\#�!t�A�q��J��vr�L�#! �h�rn��̓���%������W��2�l�����r�PM�7���{��#I5�E*��ol}���?he��&�־~tϩZ��3��sv��Qhhlj�`+�`�v�I�\ra]�-�6�3|-�8S����e�nf�Y���z�mQ�i_bj�%�ؠ�u $��2E��;gZ�5�1�D�H��a,��_��:v@/̳����8����J�<�<I3�Ňl!��T(̿�*#:��,*N�[�t��/+���=)_lʩ�@�t>�t����Ө%��V��5�ӧ��a�:�+�z$�2֭�C&c~=1�?�5F�:B��^i������!��ϪQy�R`Z�M�����w�8ǆ�v��{���"^I�3я��a�2�:D���m���d��/�ᷓ.��v~Iܭf���HP-E�����n�[�L����x�}=��?l��09��e ��`�'p�щS0�Gcpb�
o�h���ӄ���&A$�j}f(F=(>r����:~���]n�	Fw���|�1�s��H����YK�NKE�\��F-I+�f� �E��n�'I���d���V+�9��o�P.٣�>��H�E�q�*�?P��D@�/T���F�f���s�&�ɼ{	KN�[M\����j�k����A�"���MF�f�[������?CצB���n���2�!o�k��W��w��wE�c�ZҩC��4<��_��3�L I��L�ZfY}f~5�{ZD�����S}mda�rc�apLօb�����j�C��-�mq�"��u��{F�	J�
�P �؆�H�ђ���zD�Z���{�	h��VL��M���#_� Z���}z�3G'-�aW�XE�B�E�Q��sx��E�l�(b�J8�M0�~u���s�:��]%�T��9Ӟxs��]�b;�<��@LДQ 5dq`�&9��)��s�M�`�v��#��7W�ҏ�9���{���>��lA
I~���XNR2=2��{;c�@u�O�ސ4����s�Za�`�VFUv���i��ˈ��w�[!]:���]vM���H��f���N��wl/��1߽�Q����m��D��w7F�xz�_�j�<���!��/Q"c��D���dڔ�FL�O.i��Lj�;/�C+�k9�vC\%[������>Ml�v%C1�%��<WD$��L��nk�e��M�cz��-gjE�],q�V{_R3�J>(��`^�J=��d�����L�IT�N���u=����(�W"�~g,:��Y�I����[+��;q�0��[�Dt�����#���+��O��yի8~�����}R���T@R�?�+[]��۪�7$z��B:״RˏtLK%䮮�3g|�"ŝ0$�`>{���wm�P�4Hы�M������7KK���;�<�F�e1Z��U���8��e����Z3��)K>�_���{UO#��˒�j}��C'���آ���;��;����fٍZ|@�~��Ǐ-�1���v���"E1Prэw���8kO��+�l��,��T�
������iV��Z��k��U�,6��R$��q��b"�oy��jgz69��6_�ROt��5�׈�����qyQ�Ñ��*ײ���"\B����¿�k/|L�\Wh�23�Th7��>���7Z���.�>�9Z�L4^�̸�0:)$��V�7ػW�☸�?��p7��p��̙#p��Kr_���yF�ok�����VBF([�	0����3�h{X"��h����!t�v\�dR�dP��Cc����[`������5��c�9� ���'�@��V�1��'\1���Gl������vb�6bso��W?�?�շ�_=D��:˙�7��ʰ�r�ٜ�>�N\_N߼���@R�Er���O��OIԈ����Ԉ'Ri7Jϙ�m�<M�����J�N>�Q��ގ>L�wOe��.T[�(,�+RK�9g
o2-{	EՃP�F�j���
�+`�ƀkҷTI��ZPk{?��^�?�/0)d���.��x����ٓ�'iY�}��h���4�)Aն[�)�36�^��G����6��@�Xa:s�/�T(=iQ���+PzG��JON4}��
m0T<���4$�4L�������x�)�0��� B1;]$�eT��[��3zZ[�.��U&����{G����>x��Ţ���#��5E��v��MoxQe4K+Z_�3S�DeBB8d��C�~��J�J��зb�J����n�����
 pWyE��0Q��2;���t���F�_i��"�s�Z�K��txr��\y�(Sef2�9�2u�l&�x��
F;1|�u�Z��앑3�%�,��&E�
.���OTJx�,*��nEV�}6�w5���!�]K���|+��o�$g�{�qs2zn0_C�KQ�����=,�%)?-���^�ߕ��Q8�;j�ucʫ�u淗/
�޾���E^N�ZN��R��ཬG��b��]��O�"0�Q>���%5~�S��ͻ���Ӌ���'rG�e�~��WrVM��I�l��>� 6� _���v�~�̗:bV��D��v0������~�+�J�&�n��(��:惰�P��2�*oB9�n+`f8�� ,��oC�7F�o<��uv�[��4���1��7wM9�1Y!�bK�q0-.<�	k����wݵ�!ss�YK�v���r}�y�]=���.�$-�������&fD�g�3��Ӥ�E<�)����j+N[CĞ9��s[����0�߉��d@��ME�@m9"!=#vT�	��E�$�3NA�k���9�0�����R"Q�k�e�)<P.9�9�/�"ť��Eϗ�h�j_K�ωѣ�|��2���/47+/I��|��G�<_�Q?��*���Yl2��':l@��y%�܅?�2��2��|�*�����)�[�i/25i^�������}�F�!6L%�uK���P�^�T��V2��ٯm�W&�B׻���q��R}�y��F��\�!W�W�W��\o�P�F�����������+8*��a����&�l��^�YU�xUy�^|(��fP�P1,e���2�K��{�߂��L/�������E��;DY�"�y"cX@aV8>�3|��=� 4�uS+��� u]�dz�o��$@��uyӀCu��Y�J'�}��*G�8㓢Y��^>$�V��F�0�I�z����P�ˁ��@a���Y����k`.o�.�
��qWїz]L�Sư�pW!pP{θ�]�Κ�>��O>�,�L3M�3��j|~�Gp�{��*D�E���w�j�7��b2v�H����J:@绮 �����E��g�aS>���X��V��Op�2!9���;kr�PV��r�/�����m����:ӏ�Q]�F�a{�v?_����n�q(�i[�ڄ��_�ehp��귽k�.���%���������=tY���L34�uDp5�/���PZc��V��sҠ��6��K�& ���.�g󼩂�/�^#�+� y�-=��w��"��L�J�gS��f�v0/�����fi�>�]���"��{����Ƙ:aqVy@�a+q��](�[(8,Gd9�e3����Eȱ`ڬtںh��8u�B󏂤����_��@��Qtrݮq?��F0��#���^���Bm����͓���H�*�>�?F8��|�	K�n-�^����>����-� ���.�%���獫� ��1�r*���':�4�|��\c�|��0�*�'MB����)Ի������Q�����*6��G��O_⑑��MD��d}T��K({��j�;��O�+N�w�|�	v����nZ�G�Y~U%�2N�͖u����%��az�*�U,�E&5���+��i ��u~1�Ҋ��Mo0�H�|�tY߾o���k�ofn3���Yn�r���cm�~����@B���:��O���]����p\bf$���܏X��?hAa�]Jf��)l��)�C��%�����=�)�b!b*�,���ǡy�OT�����	BՁ�����nX�2E�P�hnWYW&.��]�j��x^�j��ý��AA����Ӧ��*��w5]}����^����S�JA�45�h\���_����
"6m� k}h0�Ѝ������곂�36U�⪗���ER~�5�$�-o�x~��8�����pFN��/UN��	#>��,��,�1t!KZ�x\�/���ե@��R.?�������q�ު���%��K� �OP_n���!�*J�NaDav�L|������r��� "7�5�5����dgx�Hު)�����z舠-ؓ�T�#첑H���,��۾6ㆦ���8�S�[iH;%�ʮr��4nSdĲ��Ơ�*Lf�wW���s�v\q%k P�.a#��#�E�Od����: 䊫��L�]8p6��d�����/o�����]Wx$��+������6��zqU̖��.<��[�z	�[ӱ�(�r�o�}�Q5r��~)_y
�㦁?��Y��\bnfZD<}�)�����P��2����B����Qx�kk��Mb�����F)�V"���:W�7j-��b���F��l%�&�Ab��8V%q.���boq�O�1��I� 8����R�[�K~��L��k1h��kGN��AX��@�����B-�Ұ�g��z���)������on�:{��9��op!�p�aK�gS�%+��<�Z�+wl~͞���K6e�p�b go O�>H`yڞC�X���)�=֌=�X���Q���S^ ���S�Z��I�M(��� "��}���H��Y��$\�,��C��fxq5���b1�`F�|d�p��vB�oI�J�$��-j�"�?�_���R(���?�T[s�c��M�gK��ӏp� ����t+���=g�\����D]Ыs�ܧ^���{5B?nx+k��jbv���b�&��c0��?቗�T�0�i����xK��;�}=���`�~bov�2�n`�Wj�lk�4�`"X�Zu����P,�X� ҫ�K�M��@n�W�i�y�RI�ݾsk�h�� $Ɉtr����d��M8�b1Kci��g�J�?:��`O���۬����bӅC��h�U�бV���H͍h�����S�ǽ�{����N�r�1�a*���F幏�����K4���M�"}(R�Qc�5u����݇7MOS!!6�~�k�gi�V�K׻\&�~�F��J��ғ|?�2=�����h`� ܌�=%��QBfc�����k6�n�e�$76�ֽ`[�ߞ�@��
c�q\p�A�h�Y.7S�H%;w0�8�D���-�ւ���W�:��H��Ѓ`�ȏ���8�1Bx��
�M���v&�f8�`���6�%>�m1ai�لҩ��0 mB��Xl�μɓI�sY��Yu��s˹��2����,���5���Z����Ӂ��ݗ"��~�x��*�E��H�����l���]��:k�OHV��wp=�SД��g�@e��|�Arg8u�𜍍GF\�w��ɝ{���"I�o�y;nn+��/-��g���Z-e��qhlC ��z-�#:>���N��yՁt��ZHi���m"���úB�8�&j�l���r����66얽(R6�MP�F�r��YU����D����x��7k\K-�K��	x6a{�N�>2b� `_��Ee�XlJ��7��1k��]ƥ�7?�����Zs�
�k��J���$�x/�����M���8�=�S��l�T�q�;^��Jл������99�g�B�,������JUBR*)T�� &�9Y�ߋtz*i���e��A� ���Wz���.3�ν�� �������p"��;]�J=���y�L)�V�`���"�.?��g֟+5I�@2G�Q
�Ct��ssȩ�Q4c�ɝ�0�J�o����?5K'�QONG�1.��=19NE�ǖ�c��ӛxO�T�E��殺�v���
s��seT����3�E�/�v�Gv��TN7ct���l���a-,B>ʺ�@�AZ���dQUa��l_?f)7Dd�A��3�	VJq2k����X�6��f?>���>��:%�r�L��w3��,��	qI�o�-��h����,^O�BE�E�ޕ�����ۭ�����؏``�/̐�����J�����E7$A�����Ô��
�FD
σ"�Q�M�~��hE��x����Vȸ�~R#�R&�*Th%�}<�F�1~Y�`���(��kI?�˦s��3 kHV���]�Z;�Ѵ��T�ήe���� �:�%��&�<_� C���'Ik�_J��^��e�u�nf*+�nQT=y֎�F�	��{ic׎���'Ӟ�����A�w�d��^���D�p�RԠ�G�������ܕ\�n��ۺ���όN����`���Q��(l�^ Wk4�F��:��H�δ����ͤ���f����ڏ���o���n0m�DS�\}��塡��R,Vc���P��}�oC��ڥ�ۍ��q��)֥QI�X��i� $2�Z�l�w�2��L����3��!u�6MA5�r�F���k��Y�%���}1Qe�#�"K˳��j&:��7���̄➧b�Now��v����h_�ƀ��9@SOہwk�	Ok�Pk���֖@u]�D~����5�����6��o����<?����-�Z"@o!?��L�i��Y�X(�A�P$�H8��WP$�&EH ��a�-��FZ��q�� ��K�Q��O�kF�@	}E�G��'�� ������+j��~#��:զ���\@���E�ݨkod�0�U:�"%��[�{��sn�E8څ0}��a��������eG���)[���
���n������>��k�'�Q��&�${����oy�Lo)P�Y�Mh���+�3Q2F{M�&o���D���%�g���Tr�òP��͹���m�a�I�^��>^67�67���˖��IC�mh�m27R��R%�X3�ͯ�_N���?>���=���,��ꅧ���3�C.Lcݗ���IVO_���M�?��ҥ�<VOb���GPQW��{J*&����i�v��hqM^ϟq~�b���C���Ia}�5^�}�a�!��VL��w���`F���e�QA�(�5w���'��=4���c;!)]�jA����3�٫�����κ�yG�S5D8U��
	��*6�U<ߐ�q-3 ���%�Tք�#��6/Y�=Tn$��(����;�����8n]`��w
��͌�/Kg�B���M��҅�ڝ�$�Q��b��[�H�[$� �&�G~�K�uM�N~Kv�~]���,� ��@^p�b�z=Дk�C�	�|+��1==�Q�%뼲�q=��+Ђ)�9#�E/�h.+k�L\����_#!Xh	�N�0kyF�Ғ=�A1���r�d��K��P���n[0_�u�֎��矽 ґm%j���tvѤJ�B�-��@C3�� ��Slr|�"o����hhk�������i�[�����XjK��;���s�+Z���~�ʦQ����/Vh�F��O�!���d(}%]H��L�L�ٍđ��Q�e���]��a�3{Ӂ��@� �Fl�������~�}9/4��	 ��+������
9�I�Ct�K}�|�}.fN��Y�m����~���|�M�b=�΀T�vfw}Jr��*e��)��ǘk��#C3����fƴ�	p�������^���q�B�h
4��~����M�,�w����㳔c� �5C!�|w�1t��*bx�e�����pQjx�i3&2{̽B�,<_Na��f .�S{_����?��J�DU�7�w���,��lI�GV��
�4�V��^R�;}������R@�u�m��Cl�޵'k��!˔�ō����մ"��q�]�_�̉�2l�/����D�noS��UU��s����4�6v]��ڞ���vE���&
��'v�(���"�����e��kS��A�D\�5���a�/�?Z� �t�x��'�$���H��4}M^�B�֝,:3�'zI:�I�e�!��"��=��T�^����4�i\xO��!|uZ�-�&��6j[q��cF���1[���:�K���� ������~)�ٸ�1��/�ڭ��tR����~���þ��ҟ�ӰA�Ҹ1�����&��Q�<c���2�)��ﴱ�T_y�F��T��n��ϹDҶ�b*9*`�h
���N^�a��b����$Uv��ӻV�L�ɶ���U_Z���_�S�V
ĥ�e����������Zd����S������q�Ҿ�!��Rt�%��W	�;C�([�܀֡n�vz�Jt	|vN�Ļ1�����	sa$��S�E����4a�������-q%�(R�y��s2�s g���'x'x3q�����=��>,�ia�������ʤS���˼,@@9y)F$!>=5���P`��l�������q{_iQKq���Q�ztW�<M�!7X����X������=�G:}��\p������22�VwQ?�Ȫ~X�����C��6p�7�Ey���/��0	����5�w��B�B6N��qE��#����`��0��2�K�$��8�e9V-���bk���!v�'6;`�6j���E�N�I��C�Tla�`�ױ�f0������E�1� h/9K[0I��a`F���ppo��?*��4��`Ļ�I���LwJ�50�c�5N$�A�?!$�F]�N��k����y���E@���m՗.���@��E��ݕ����Iw�y؇H\J}\ >�<h*qk!{o2eOM_�*���3���D��G�:ԡ�I"��n}�І�'�� ��O��4���^y��,�Y�K�)��6��҈W�H��dE���$[+���B�8���X`�� eg��Q���2f��դ�5<�$�c�m��aS��Ri�9J��63�ZA�F���QP`���AkP��B���o�W��t)�a����Σ��$!W�>gz��8L��'��?���!x��4��O@�S�b�'���赢�䚙�.I>�~Et
�"N�a��>��^�[�&�~[I����/11iv�5�6�K����ٛ6���H�:5W�<5:;ї��XN�"�5%�R�-�ŭݼ%���lX,I8hdS�Y+H+G�QÅ�����#����~<�x�p����rE��Y�E�>��H�Ę�������c��_QD�(�}W�v��}��`<�H�S�L� Q|�����u��3��<W�μ���z��U���{�ah��wU:~�龻���-�K��}��s!�aϩ}���8	�E��&*�-X�w���˾MQ����t��i�8��dtz�u4q+ϧ�r�g|�jN�A��^��� u�8%�Y�m��g�^HA�j�3��j�e޷96������ӫ�+̷���1��=���c����s�z��d�\�L����j����k,��g�~�'�#��'��ȉ��ʧˀߥ��u���_�}�N���D�K��P���+8[�`��-u��UP��bDN~��U�ʓ��*�a�7��Ǐ��ø�� [�K�qYR�=H7f= �#-(����-��5��k*��2�,���_�͠OY�����Б�L�/l�dL�&�t�o�K����{��R/*���Y�m�z�B�
=�ga�N_a��5c&�/�a9�e�V�>� �DgE�[�5'�m;�a���^l�����5mh?�O��Z|Ҽh֮4L�f
Uʳy=ۺ��]��u�����wz�����g��#j~���[�:�[��,(�#�L=�����J���y5�iҎ��� � LJ���J}�*�J���C��B�*���
Z�,N.�Vk��dD?V���B��|���6�=�M���\t��4i���u\t+�%��Zл�`�Y��ٙ��Ɍ��,�|A��#�r��x$�f_�f��f�;_�H�������L?�G/<��q���S�x\�\���t1 v.�qF��+ȡ,/����"7WP��_����D%�р�����f�x��P"~h��N//�\K�w�� ٠]�7�mf�ˡA�ɽ���!���y����p\�W�)0�8��4�\��7mC�U/�ջ���Zᣔ���o�E��#�Q�@Y腠6����B��]:���ϰtۘ��6v��l��_CD�T+ITә�9$���YD�i/��ћd�~H�|�<@��οV�v}_*�~|k�{{��1Q7soу�R����jk�#x|��~/��L}�V�g��o��`�IJ���奧t��ܳX���xc��A�� ~���'���K��Mt&݋v�_jB�:�>�H��~��A2�����vO)7~��
Aՙ��v��}��8����nEh=���{	� ���}�G��Y�����ך�yxY��3v�ؽ���e۱�)G5{3�I�i�֪��,N�
P0N��j��m �qf��F���uK:��{�|���ٞ45۟i��@��V`�#�x���?1�i����S������H6g�eݼ�#�`�]����Sc$���X\�$����C���-(��ǳ>�Ƞ檢�ګ����K"�U������ܑoT��P?d��h�oO�A����]�N��}7�ï6ʁ��Jo�6r���qs��AB'0�7���'/%ҍl--s	Tְx ��o�ߛO1�W� �9��?:���'�����3v���|m7�'�1<ۭv��}[�1"����X��=v{ʋ)R���9�;L���D��<]ͺ� <&����I
1-�}tu<��'��C$�x���k��{cQ�ia��NJj K��z��er��s]���V*��#���Ax���k��joL
���z�~��@m�K�Iv;_۔.,�#2��!�����L�"��HNo�>p�����d��/���P���!�=�ѱ�l	C��:Y���
�u���Kx�0��B)&}�3��R���u�<�@��ld�v��R_P8�ֲ5��F�y�����s׸يl��)!p����F96ǖJ�Vn+(�����G�;]'�$2 �9��q����C��}�����H?�زwy��R��������X� �_�ݦ�
|t/��.��3�z��:?�TaO9eP�L�h�A4��P�i�?�@�p仄�P��8nȨA�q�N�]#ʴ"�u-6E�p����ӻ�����=Pw�B��u�6�B�ܽb1�{�����;}��C��!�cV0�v��^)D�1��<\��ƾ���?�Ʊ QH��ğ�Yd

 �Ɂ�`f��-��w�wg-�3��i��ԣ�u'յ�ھkx�~��(ާ��Dd��p�=6~*�(C�,�p@���%�^��^�o��,�V9����\2�M��%K�=���M<�%ʘ8��@��0�j���s�F'��{|�������)���s~����=
�pf���������1
�܀�;}���m��}�5R�m�W����%��&�^Jގ��"�ê��5�x��e��~6��?�D��<->�>$������C��]%$�`!��y!g�-p(�Ѽ��<��#x|�V PUX��m��
wq�hC�D��^���Y��&�}v�M!=�L����໅$����WPk}���S�o���Ss��L[�<tĠe���=.����
�IVrv�3K���l�*���UQ��ov"�^�Gl�D�Jh>���D|Q�\���m��0�]T��b(�D冽#��@�Iro�Ѝ����9������R�?�R�:s�~�IF���[ć�#'r(�L=t>�q�V����HNx& �
�)��(�4�&�`O�гy�O5����n�Y'�}`4���;���~�/�oA����V�'��^Y¾e�_P��?F���O^���-��7ES˼�T����Ji�Ü2��a펰GX�!���$���0z�A������y��zj�AmP]$4�Fl�-\�?3S�Y����1�k��ʟ�Q��W')ej���(?�F����|v���=�<�	�EhQj ���x�$؁���H��/ l
��K\�X� ��W*6c��p�G>�C<��1{�$AfY}A����7��7�� k��Tc4���{�v�R���V�1����#���#��S��ӢR��y�Z����Ң(�p����'9�+���Qu�v�K�3�P��g:G���!-�۹��s��`ְ{��?�{�e~B��\����@����ko}!��d�w�
^K��H���8@� L�V�R���_R�(�zE�Q���n�7��f8c�(/U$o�oFz'P`����z��/���:�ay�a��<#ϒ�a�p��U*�̾e�4�ժ�5��LVl�h�]���{�(?չvu|�U��̮TuW��~M1��1o�3MH|ƐCG�I��(���M�<�]}޾�ъL�`啙O���8XL"g�g�fG���R�RjŘplG�ة�q%�s%r �8�·��1�ɲ�)+��;��S��u����@�錎T]�����p(ꜭ��<iM�|	5�uH|���)��O��x3YdJ�ۑ"6"?Ѕ���n�Z�ak��,�
�2���e�zaz���w>���u�K���\׊����
!�|漢��׼��!\eӐU��\nt��\r�\c�y� �Q\+l���:�-4�	)��]Ȏ)���NxXV�d��F?��`pNЎA8����w���g�ʉŭ7l�3��"�������F޹u8^�=��~{w���*�4��?�t+K��V���f4��^=)a���ȿ7Jؓ����J��/�~\HV���`��@1 �r�L�`�/�(�y��AЭ������?iR����:�v]}��?_ �
���lq�t�X��lޖ��l��4�C�Hq8l�ZO�α����K_�pR`�W�/�<�������5���=;�J�V�ΫO{�R����±��j~���\��R�a�/�\y��9xkf�{�����t�᱆&g亭�{%���4�V�n�4��A��A��x
V�<P9�Q�6۪��D2Y����Zs���a��%�jz� �{=���"�9�A���P��ԛ�������M�d<�M�]�E��fQ�*�Ω~�Wj�<��4����$M�}[/�v/�0��鶴�����+���0��$��j2�T�rsk�x�a��2^�1Jd���Wu��B�& �u�H� j�<S;z��3;b��B� �Hf�X����xZ"^�빣��˦��!u�ڙC��*�C',�ց�7Oc��S���:�#�8���b��s��S����a~�u�ӯ��4�??��]�Z�ͥ6��Y�O���;<:"$;��vm&������:��7h��"�@��X)R��@q��m��{pw�R��"����݊{p��wx��9�yϙ�?�$3Lr��>�{���aq��*���N��N�XYӮZ~�Ʌ�Ӛ��JA��#�56�;qu&<�����Z0�J��n&̽��T�xۖ���Z�����K�����8Xa�_�,L�9���CM5���a�`4��B���U�&΅k�e�B�0�I�<�4���F���O��v8 nMJ�.M0|�t���DnB�Q�E/�@=H"�E�A�W���f�D���+�sK9 G�i���mu��"�wt�j�6O�T������U�X%q����F:��e�@�B�B5ŞTV �a"���+[X�c�y�,L N�.^J#���5H��~bT��V���58�I�w�g^�-L��9.Qa���ý��<y�C�BL���Tz�_��=�|	>�7�Eg^ΥSl�h|������xD�^m����`�D��^���Y�uZ�8�LJ���j�"T�f�5��jpsf�	B(OJ�-�D=�A�V/9/���g���P�����ɢ�1}l�b���"����wa��C�7���&K�@`��Ier9�,����4M~�Ӏ�yL!c�G'��W�5�R��̅5���K���k&;����\�2��7a4ԂV�}� ���e�ħ9I2�/�5A��p�e~p��r��q��Ǎ����ᎀ�z�-��c�Z�����2ؿ��ʸ�ߪI��o��7w���k���%��߱���u�n<w�������U��7��-"}3݅g�5�%���	��iy�����5d�8� ���8��vKk�&��2	��O"�}=����7�,��f8�>`�t��\ ܧ84��5>��Ɣ�P&W�C'�C�M@�1�o���HH=J�0�rQ6{l�"�h��dӉ��������/�QŞv�ǈ�

$6��=V��K��+�7��M��ؑ�G��*7��Ym��[q-sV�٘��ޠ.��_�P=�Kw²��#>%�N*�7q.S~ٗWh�p�ޣ���ʌ�o���OO�X9x�n$%!�N��Fa"� E���)����|^�8�j�!�d;���`b⤃����e<��]{�5i����?tr>�ނ�[Cp�����P����22�G[��ς2k�]���3n}����b+!���%��7�lJ�� ^��IX�,��,X#l$������lCfvT���>��h�fK���K*uRJ�EH�7R�����b�T,���B��v����Έ)PDÑ�N��c3��Er�jr��3~$R��c*�y�y��'R"����lg�J�p���U��r��&k�`�˰�eߋc�Na�K�h��\�l���l��X⌺W[9Ð�6�[v,���OiF�.����N3:M�|A�qh����W8�uW��D��c�!��"�m�1x(e52��N���.���z�Ec�ǘ��࡯<����6 �+���C�N�N:��o����%�H��H� >;���y��F�23y9�Q#�D$��=��/��Ws��گ��6�/��MaX� Fȩ��h6��8�w�������X
����:������ȫ�A��Ā"�j�)|l �@꒿��S�s~���@�Ʈx��[�+'�jHl�����7<L��/�h$*c!E(ʱ���7�4:(�9"���DkX�NQ�����O	����ϸ��@�s���2�5��?��������V�
�����v�����I�`_�!��s�`棟34a���"k�5��U�3�:{���+*��{-���ϋ)5y��8��F��;	�5��,�I.���][� �В�_�[��;j�黍���>�yEC�É5�UeN���!n�^�w!�~��W�k.*a_8'�z�y���UEF��O�����Cn p��I�g�Ш��-�?N�~�k&����~�|
ߚ�[��nC�$�h�w{�Q�i{�;�ᨂ�g^�;�,{��=_P�8�^��϶:Tz�Y\w��t�]�۟��l��!B���b�uIF5���+{������2<�;�%>4����N8Ȭ-�74}�?��p�?̮j(�D˘l��� K�2��R�	b��UG�Sq��2i;�6>83=��Te[7�Z�浖ڶ���wA�S�U ��ۇ(o��XRѡG��w�^�NΆ�����Cx����m8����B]T&�w�L�v����Ս�����3�9�#�Ԇ�/8��N�)y P��Qe�&�l����~Y��sV�H��-j �`�� � ����g`V-�E�v�#zl�.A���Oj���ϱg�
<c��j�z���/Ԫп�J�dW�#@G��p����/���IˋCN��Nh5��yP��P1����0�p科�����W< F9��f��FM���Tu��t��GSh �7��?�R:�ԏQ�Ʉ �6,��vy:�qb�wY��=�T��Z�7��;T�]���&���A��.��FɌ���Ϟ�O�"�j#�	�_$):�4�x�|����������B��])�IZ�Q�Nvu_`y�� ��L�]���I&�q��B;����K�[;�:cۜ���R!럫���)�&9̞��H�x��՜��@O�2k���6K�Mư���*��*d�����ѫN ��o�@% vY�1D配x�*)X �X���	s�g\60ք׃�,̔x��0!\�B�n�S��q�@m�N���QDT8�&~|������dyZonr{�/�JYd��¶������((�g�R�j)�i��R�����t��Ə�+g^��zч�"���E��39q�и���Ab�.��f���q��y�^Qg=�+�Ϛ�D�X���Ż4~S{Ӳ6��RvXH	z�!�2��:"r��/�'����6ԐV���ym���i�P����σ;����"3�R�ϥj���M�x4������%�-�oDK	$7C��+4-�"���Mw�z�����4�1d[���n%M+������j��\�Yɸ~fr�02P<�r�G@%��8�Q�"�x���M��1���60�
����}&����ܘR��`�pԪ��r�Ѝ��׸fĵ��uӎwþ�`S�l����mǽ���S�ɺ��� �O����[�����Y$�]�͇L���d5c{��Ҍ}����{�������ԉp��ة�qJ���
iT'J5.2��0�� �d���-)�L1nk��q�?��D���VG�H
ބ�ya�@/���>9���R$窾���n?C�w�����t�kIK��8߁��)�����{�Jуˊ/q9�!�#{�={D]��#�����LQ�L�N�j֧��a=��yZS2(����N"��9\<;ͺ R�~yx �:��ģ���͘o�Q�>��� �r��'���l'���>�@)��bv����:���{A�����z�9���������հ�;����D�{�VC�rDD�ܩ��sмSǜs�3} <�|W���c�U@��ȵ����.����V
������˵��3��l�[@�<�y�ꎍ5v*���	2����=4�����A9WŲ�3�w=�؛-J'+s�M$悸L��*p
���H�A�������ذ7�s%B�q�;�q����+��L{��Ǿ��ͫ�sC�lξ��Zh`�w*�I�?�dr
>v����� �(#�Хqb�(�^��!���_Fh$����b��Rv)HzZ�!�,��iA��mBjOi]����/����q�&3S�Dc�#�%��a�/NJCb����ڬ'��ob�<�tm��|����h}\,���+b�q/c1e�\��x�|P����
/f����=��@ԳQAt2#�ź��i�\P�WVa퐥��$Oo�Q���4�7�K2UZy�u당�nF'���[�>,?1��c�����֊�Ѿ9͜�r҂p����@Cb�)iѠ�:ʮ�r�� ��g������rB��D/�l�dw`!N��Q�����洩�g�����* ������ ���9���Wdw�a�%�X��
�.���)�>��i����٢�L���QW���r��W��o�ɏhDz�6U�j�}��0l�6��/W�F$��>��Ҽi@!�h8fi��8�e�T�	@�P8��+�/�Yk���c@%/�������y%o)�p�\��/;�&��2ˑ����s��?�7���ӷԊS;���C~loE��f�:�UW��V�;�G;���v~6`��%�z:�9SOU4B�W�&�D
���Z)N_I���lZ�;�$nH�yfg|�-0ڎ�1`P�}4�o�Nd��m��.�l�%�S�`�Z�v�a:ڲ,�Kd$�7#�[��m�c�:�K'��W���I�N&�]^|w0c���U��w4���{�b��9qa�����X-�,K�LUG��N�!��2��譕�TY�
Y�ح����V/����t��ð�:튖�����'�~JA��ˣ�
�w���`=_F�-,zk�Ŷ��96��跦%���[�R�ca�iTNP2�O�aZ[/NO�X�vOdr���W𙽄��yj/�T5��Z�m��o����\�++�Ж��kPK��[b�rTg���c�.���O�8t�W�=-�CZ�҃o���DY�g{���\r��ě"YZ�d|c���6���Y�ʎ�	{�� %N���M�e��֢A����?�y�(t7Ak�a���Y�QW�s�@���s�S���6�k����2�1�W)4���v�����9��dK��!��GL(f���(�}K��Om���Ϻ���OL��'$���W=����u��WXt�I�1��V�b�E  	H�!py����div����k�,���T{9����2g(�c��I	����X������9_�>����g���x%��g��GG5�d�? M�e��Nh�q;�[�\t�)2�+�pM�yܞ/L��X������˧O@&���
-h�֊�'��'3� {vR C�$��{RK<����cp��GE�"�7N����vtX�"�K����0����U��o8�H�IR��ϔf�vm�|���k��O�a>�q�뾪�d�� ��X���x�)z�I�F��^�{\;�G�U��Ws��[Ǆ�5�� <0S�'BU��>�N���F�I�g%��6�����O��2& ��άWp�������]`dǽ�<6IW_`�(*�4��0h,!dB�����:�r2c�LpRß�ܲ�w�� �Tt!4/���ͪH�r��ls�[�m��T{��*�i��Fk���=OJ��h���	�h���l!�!֗��7;	a=���DǛ ��J�D�Q���_�?�|,-�ۊ��)J���9&�>��Hپ�1��-�fy��q�."������n��`�N7��u˳��.Nx.n��~�i@�����o���q����D�j���,p/+�`�X�$��zr��Bݯw�h���:��t��yD��:�;{��9nѿ6�%�Α`f;FK��C��e3�F�3�-_ʱ3/�E�
o�)��j��Id���k
���0��I���{Vox��_�yi+Ǻ�����ؿ��r���l�J��Q�ǩ<ɵ�o����.�[R�����F��zqX"�A�G��B������T�wC�Z����6L��$����)!@����*�l ���`rgp�'R��y�T4{�~n�>%[���Øc{��Tr�3e���3�~�[w�����@�y�v��}|�S�e��z�Q|�X'}X��V�N��y8&v����4�����	͉M���Y��5m�+u�W��,��,�
�Hq�*q�t,��$L��Q���q�N]��ȳԏ*�Rl�#2:������k��z-K�d���2}��,GQ�t����j
�Ǡ�4S��ZT�y9�58ϱh����� f�A��6n�Ck�s%͎�=�+��zOah�%D/�ѷ\b��\��X�_��&� �J�8�f�P��%S���F#Z�s}�<��&J3$C�S�����b~����_|�R�������J0�LB��L�(V��-/x[
E�M��'+�M[� ����(%�:�p�.;��Y4ԁ& ����:O�XlL:��y����d�&`X��"9�J�a������b��ͧJ��jsk��'��w��l#�,��u�k�vM!2��i�����n�Y������c*���ڷWn[�:%{өԺ����*KR9�k�n��a�ޟ��E���YX����` 8�E��<��3hX������CB�o�v��
� I'�Y�
�{'�x����G��-Y�-|��y�Rbp�k'�i��� H[��S2���ڳh�x�OJFS<<2b��d�;2}�vI�{q�-�̳�Ԍ����<��`Kk�5�F�~l��D��L�o�(�N�r|H���A���kd|�gn 7��a� &�}�n&ٱkdtW���>�Y\�<g&���{�j�z�Gc۲���ۨ��#�%򺏊��)�N������jgh� �'$�7u�9Cg�	���j�6�j�K&SV���d9Q�G�'����<mz��#fh���w3$sua5(�|e��ڞX�q�-5��b�����u��-?OQ�)��Szн�q�w_�1-I�-�O6��)��OH�%F���v��bP��i�l���T�2�J� ��2�#%��k�e:��%Z5@�.�j��M"��)���2?x�L_���]�����I�R��2-�Yh��7���?W2ڢg�]o'<ݲUh�˱|��f�E~�;�����&6� �`J_KŜ��(Tz{6�v*���0�n�)>[�(F�K���u�JJ�̓!5VP���ڶ\�*�0�2.X4����u�l6�T"�>_�����ϰ��/��?�	���:��TS�߀�6Rb'�U����]+�c�	��s�̝���d(�o|���i��P��J u�C��j���շE�~��2�5��N�@�q O9��􀉾HK6�|Q<�M.� ���9��p����*�"���'��t�K=�t*�5A���N�;�gr#�F\}�_�>��v��ǯ�f�Ek�	6 i�L��s�F�� @�_��Q��<�e�f%��-��8�<��=��O5p�n�9.�߄���=H�ڦ��Զm�dxfl�gL�5�a�Kq��A� �������D0�T䅥�*)P4Kv�(�0�B����ח��&Q�}�������8MBw���[&m�N��F�b�u�~'�v8��ڀ��gIΒ��!�]�zHv1j�>��Qs*p��޷�n�
��y%9P@����į���9��$�������^��� B��Ag"�[a�=
��^�k��"��|,�0vK0S	< Q�x���~�Ȱ��|��'jb��^/0V�%\'��I�wI{�O��v\k�V%5�se|b��D������wx&֭0IX�:��(f���E��l�����P`C���%�	)hc���>˜XxU%���m�jd�(]�	m�:L�}�r�xq;��V�ފ�~)�ק����S7ҝ�2�	~�Fk�ϟ��M�[�>~�?+m����>1V�&F�	���bL�j�e�%��W
�Q4S���y�f �U&�k}gh��@�I£�K�Y�v;T@�=H�=H���j���X�b 8x�`���W&nL����]�.�D�y�n�Lէ��{<����Q.j�W�T7��q��NO��]^����ث��y2h:���ϗA+lϖ����PR���4l|	U���]R�ǂ3p�^�̺���L���ǫ�d�����t�$Qf�v_P���������.�"P�-��(���b,�V�m,�O�ō���d`W�:�u�G:N*�����bh���)l�Kw�����U��_�)t����w1��$�:��կ���� ��:���-��& -�}�������h�e%���+��VV�ا�w��v{/-G��.�{O�C'���d���
�f�ŠW���ۥ�̝�56˛��g;��
�6
��Ɠ���y�=���0ђ	�{ՙ�/,���H�Y�B������E�#U"4��c�t^�P�LW����x��W�)QչX�It�Y�dk筃
�x��x��Ausǋ�~Gh��+�{#$��Hqx,�u��:����;�ǈ��͠H�6��J�R�1͆�I�L	e�^eo�-���qߘĭ��>4dtCx��K�Ҧ��Oe�j�R��������5+{�^֓h0�su3�)����o�,�A�_�zPԱ���k�S޽K�]�a�UMW���sO7����%����8�N��]S@��<�C�?c(��Ճ�
��q-��g�<�V:싶�ͨ(1���`+[5o�8���(�ZꩥwY�T��د��?;�d�JZ?��iC:�"׫�����cS��M�m�ެ�Z�����u?�/���$�P/*�hk8� U���7S�o8��	���·�L}j��4`%U��&U�G�����@+�F>7�����$��);�kVPj��-fT��G�6|�mkm�]&a���1<R-]oF�ȕm^�0�kL��6BPH-: uZW)SRЎ��p"�V���Ϫx�s�b$QJ�w�L�(/�~b"��0v��Y����0.	qs�0��k�4�~�,_��H�U���n�� �b��RZ�����+װ�>�sƎq}�d��V��jm@��i�R��Z�z�Y�:T�w5 #GN���o�(�Ƭ��W��Zv�,^
����&�ĭ;(<��[p!8��(�,�
���G���W
|��{g]��d0�SZi	Wvh���s���?�N�W-_������TX�ܽ��2�ܝ�,l�T?���T�%.��p���u3=w_��$�|�s��s��ǆ�7O��_O֌��lͽ�~c+Sȷ�_�=Ͽ��b�p����\[2l�P^�?D(%�@�L7����Ϯ�PW1�@�˵y��nB���g*l��p1�9 �u|�7C�|7m	}@q���f-���ƾ�ܧ����	Yy�gr_PR�)= �A�$b�`F��\����ٿ��D���n����[���N��	(%�C?�?M��q$������Ǿ��PH�����,�L��`p���׻E�dq��",>�~���TU[��=��B)���ra��<� Il�=�F;3��1�m�}��Ԍ���"��/^(8|�FeY"~�K����ҍ�OB�,J�q+�r�
��	W�{b&x�r�Nt~��N|X��;�FREIO5<�)����7���μ�n��fV�zv�� ��=R�����2bU��������35�3�����E+�<,�gm���et* �mp����7X@͋��ٴ����Ӏ2��>�w]���h<�D[�5�1⭱�n��ZZiҼ}��Eu���F��G�F</2���
��W����bb�\$��`��;�;��u�����պ��h�A�i���\�@�U�	��l��/���?�Zm��̕�S&�S���a�z�V�ͷ>���ݩ봗.~���q�XyN`';�P�,�d{�Nb����_�q��r�����1��(k�3+�B���/���^�Nf��ŕ�t�3���DP�q�@�?���qB�tV���ү���	ʬP6�J�m780 ���$MrHi��%x PxQ�4c��^�T?e�F��*��3D��s����KT(P��&�"�$5T���PX�úS?���"�A�.~��]�],�v��È4B*N;�9�R[5�}���s��~�
�JB�D�eZL�\8z���iW|���fv8��sg٭$mn�Y����ȴf�h��/�鍮6�\
��m
.R�u�k���E� 1ub$ޣj�E�F�ff|z�����9xF���K��֡����qq��ۚCჲ�:�ޠ ;�{��"E�MB�d�D��j��V��/h��E��]������J9i����R���p�K��u��R�曀�l���y�:߅WG�LWGSi�#|7�A��W��ׇps�䥲%��`��r���=��a���~#oDߎ}x�"mߺ�b��ʵ�V���+��g�*�˧Q��0�}�	�����U���KЖd0mM�����5|��A(]Ɔl��m-f��å>�ߖ�\���	.۸b����F==��>n�x�Y����B�vKRx�?���go�����G�����l yXl���6m]�[o�����^�u1��_����YRh�HR��UH/*�X���`c�|�S����;�ܜ��6Si�R+X%�qGN�E�kR�Ds���$!���C̨�@6��v���?��*,���*�`V�V+#�v^'m�]��ŭw��NF��尩F�S+�Q&?Xj�s�>�%�}��4��a=���KZ�NTM<Ƭ��L�p������ jA[=�#��\���jF�9���R~�r�5�����I$��|,��i ���U���}�J�{8,���e�����q~7%K��YS���e���GK�X��j	g=���UTA����e7��K�>
�㦋��_������|�ow�8��T��6Ͽ��ݯ���?�<�I�V��R����!�}�=V9�\�17������]��v~p<��ʝ�*�@��%w6��K�]���[��7�����l�@���l�`l�������V��[�;oeR��{�m�������Q��m���b�����7m+��O�8�L����&Xٞ%��~�1.�YѸ�RS6Lc6V0[��"��Q�b��E��"$[d�lW��`O�� 8��^�
�a�͜`���+UL"�h��g��)�?O����SKk�#�'�l�w���{����;��)�}��6n��y����-��$K1���n�(�P��h��:����s�$�hW,9��R��WՒ^wث��@2`�~�uᕓ��j��Nzb��R[p�͏��s�E�
DՑ��X�.HTMU>��
��&����	8�uc�W���2�d[�3ԔH	�t����	ia��'3�F9A1�h��\Jx�r�Y�kZM��m��~z�{����޸7	���?� ;�$�
plw�� p|PSi���^�Ae��Z��V�g�'ʾ�@��`�O|'3a�n� �1�x�]��4C��
3�'�y���x�`����7��.����ˉpZ_9�#�h~��o��[�ݞ�k���2�c'g?#����հ���v�?ݽ���*�Iz*2�%q�ZPy%+9�Y܎,��^�}�A�A:�����r89���n�i1׾����}��v��N������Zown˭����jY�U���d=�h�?ønS��'I�w�<=u;����k�y"9hb�H�'A�;�<]-F&�Ԛ3��p���.�Z�]����M6i�W���?��0�X^�Ic
��Rb)`�}ͼ��W��Dw��&�c�)����僯i�����Q��Q��q�F�3��[��&A��,ڷ'IIv Q�p�{Co�Do��]�w�<��)����y�o_���q���Y�Q-L��Y���?Lpv5>��^#�gg�S�r��)\L��U�X��ɼ8ؘ���;��Aݠq��r�|yҲl���g�$�冃�� �,����^Osf&����șm�Y_����,��;�S'O;�
#�3���p�$�6���	
���Ϳ���Sz��j �N)�۞����Ƭ�I:�b:MJ���UV�u�QW��}�^wۿ�=��[�W���Iә��*�4e>g�k�k�=	>Tqwm��;q�a�H0��3�8T��Ϡb��1�����?�K?y1ZBA��9N�M<�Xhg<ey
��#�yڀ�,p�
�|�`��f�恸��R.��5A�V�=�xJCuL�?��ޥs��[6OP��R�G��{�g~SD+&���J�~�����C�T�n�YB�Utj�jd��5��Й��Pͷ��&��\�~=Jm����K%�W.��������'�h�k,�*Q�93p`	���d6�H�{�犍�
�U�3K�G����C�<��9Q��r�yK$�[�|4t|iJ*�?����.�H�Ť�О�X�E�sxf	�~-���˙q�ԥ��Y���ø��6K$�ab Ab�x`ad�g�g���Վ5Z��i�t{7���V9�40������G�]k�e����+!Jl��oS)߶.��+m��>����1c�$_g��#±WbYM��oe�@�d[hV<L.%��*�o&�&���tۼ��؛Kt�/���H/~k���0�9TCY�r��ds�*�2������?r�]"I�Y����Qu*�x��hni���3��{��v�����|���#rhA������G��\�D(3r��q�r����L+���㢟C�FK��L֩�15)���c�DY)�<(o,@}�(�"�0�cgW,�C��3)B�
f�0y��:���)�_�~���dG'/���-���8 �ԣ(�%/á)��XK�J��2�e��rW �~�B��v����A獙!�����1g���3ˆ���	�0���io�F-�NZ.n���tO,��� ��2@Ĭ����S��ד~���"r�](E�y��}a�������s�F�ՕCIC[B�y~�R��M`��ªI�����#�F�h�	��X�l)�P/Hg/��а:�1�3�:��`v����d�$�A6�5��/U�q�$4��7h�+U���x�6�U��A��c>�A�)�ݝ��%�UAm1B#��m��)�|0Km�u�l'��R�V�b'&��m]�,{�Ԋ�:�7���1M�*�s)H�=�?���W����d�z3�aՖ�򷪇��7��#��v!p\z-��ų8wA���q�Q��44Y��z��ծ��HԻW�w��F"�2��Y�g4�b�<�wS!��]!>����Ӷ�V����@���>���/����(#5���/���m�7n��?��Ӽ���.@)pg���C铇4p�S"��˳}����w$�|+G���7���=�������C�~��{ӧ�|�������/y�$cS�����R���S�m��W�V��8���>�_��C���yϕ2�9!Q��}a���G(��@�|����@C�JU��ᕘP�6�� ��fn"L`B(������|�n��&����j&� ��C3���Y��F������5Zg�8-�r-kNz3X�`@�?��-:�5ʇ���� YV"t)H������9e��"!(� ��pӽ�΀�\b�c��ʘ��H��nQ4���E�}��J�7n%}f���:�ٺT�qa��/F�š}$�u"H��F���79k��#N�o`�Ic~&&4��̏e��%]�:Ϲʻ�Q��B���I��>Hf��9K��|������5`�ڪwpc��۱ڭ�������֜��.��qM��N�b���)}C�{����2��<�׾�3pL�l��pq24�è���jQ�t��5J��4a���(�0"_1�=�'~*��C�#�-����%�I�����W{���!8���h?r���$��U�׵f���پƑ|��+ͷ�S!@RCg�a�@���pLʻ8x��q���]_Ry�;嗷T����zgǜ�cgy���"":&�
�D�{K�>Ǝ����\���?����\�r�ߞ����.�ֹ�y:�>�3���<��Db�"䪛�Shx����F¨d�[P�Z�����!�m�	���G�,#��q��N���ݠ����Gm�l�5m�Xm�V.\��a2Y������Ϩ�*���<��"L�r��4����M$��B$�]`Q�ņ?_��Cw�^zy�Y%
�\�<��*jcA5�B�q�-/*;c��n������,��L�T���0ŀ�-�&�[|��+u�S���"J8����EBk�,��Y�`�%mT2�������ۻ��Zw�N����r�g��A���L�:�+��0����D�ϲQt0���+nXK�f)�m�|0S�mJ�S��	���m-	�\�:�S�·ړ� �����"ϊ�)U��Ҹ�ا��o�%_J����b�����T�̣�{c����	��bb��JS����$�s��u�;�F`�_qs@R���M�Y�	�\�/�F\~ou�Е����t��M)/2@w8 �^$�\$xQ��;�P�@X�2���bb��~-�q�T��-x^4Q���#C9#<��M����[`rr��^�Ic�����n+��u�sc�v�΋�H���^�����+��doKCT�gW�O���f��N��ƥ���ᧇB��L����V�����ck��֌۵���y��KϜX�����G��i*R�M��i�����^�@���_��.NT�&+�hb�x��-�Rk����×$���$s�r�d��)��v\�o��O��<��JN;\Ǒ�{hZ���_	�G�b�o3t�u�"��.+�E�]�w�]}K0�G���H{{��'õJ��Yۭ~��ub�0i(��Fy�lV��0[���ك�����A�]�DA����>�:��6��6�����B�H?�U�&Z4�Ω�m
p�����^�(�@I�0?��ō�y�K��\��%F�c�����t\QE��j;|��Owy���uI��a��}|%��@/��/x^�G.�07ѓ��#��e]ցm�zs}�J�����W �0M��m��Z;C�����Z9~R:J�C�#F�D��F�O�I,6+>�jD"jd��4�9r�)��kr�ɠyY`�Y��Ar���誫�k];��>���#!�+b�d%�,�
&�r�0NvI@�J�(�L�����*le�q_�qA���b�*��em��#>"�SJw0�yO��VO]:��Sv�����}A���ߠy����n��Ge�˷x�ܟ�m��[W+�% �1`�q�XEz�L����Sخ�8N�7��#v�/��ҎX�����sz�����:kq���W�.��$��������ؓ,�~ �F�����$��o����;U?+�B���}Ͳ�'�s�*��!��GB2z�C��2�8��7��$�6^��g�� ����S��ǖЀ����3:����8
_�I��v����T8��q @�N� ����=8���"R���J���v��'ҝ���Z�*���B�ٙ��{����ZF#����\i��s��EԤl�T(��L��	�h�%7X3���$Y�����Y*��1 �i\s�#�|�P\�Cك֜Z�z�
	��|F{��.Or�S[7�g�zQ����<v�42S@�A4Q�J�2��& �$Yw��B6N��:�B�?�?e�[�c��hx�E[!�+�K��h��VN���U�� ��FbbU�ғs�Z��,ҋG1n6N�]Q�}���%Ǳ?��c���ze�J�V0Z~{��SJ�� 1���~�>W���+"I�I��2Y�1�I�Ȫ�m).��h��ye����+�����}�hѻ�*�f�t�=��L�1�~z�L��ι.����6���M��T�o�_�������й��ٽ��]{g�G!�ÿ�=�7��)�RJr�ѱ�Q.�ÿ[*"���ʏ�$�p�������M�&����q�p��%� �GW�R�z�c�F�J2N�x�b��t�����(R�5���*�=������=z��9z���(�j�>���^&�jiR�x�l7Ʋ^��yF�
���f�s]���|�3�o(y��NY��H6uw��w�~2��\^����c�I��D���p=r��^���-��r/�^��wLؙ�3�X~�4�̄��	.�T
�O�"�XC�D���zX��-e�[��Z�Ң_�i��3���JJ�4c�p���)��n��r���~>��e_���	M�m�(>#1���«W�c�J\��p@<��	q��%[B����(t�f�d���a��*�dͅ��S��þ����Ho��K
<�kI��Y F	��,�8���6�}%��rh/%!�2_�ꚉ3������\iW��h@r�'P�T�C�c�^{�A�Z�����ܺ4�m�(5w(p�#�1P[��6�%T��OajEJ�G�������?�������&̈́Uv1�z�����6oq��Pk������_s >N�:��s�� �W��Lm�+��vٓ=M�d�*������e���EkoW����*������1��������V��Ju9�5?�� B��$�Se�	�B�B)��Ȧ��)ަ��qV^������,�/��g|m������HB�#uI%���Y5����4��\�Mط^���7��z[^\���Ȇ�C�D�\�2�ԸI~�*�Q�!_����;�J��|%�eHa�Z�Vd%|�	�LZ��Yr3z� ����1
��{�AN����TWب�͌��i��|�a�-�rlVM�y�"�<e�I�߿���1�ޯ�- �s�i�dsnAzz�)z�!�Fu��w�T��7�,�B�IZ͙Bdq��E|�y)4V���
ko�U�~1Z��`��_q�\A�[�Ve>����7G�d{�;���}x��Zn<NO9�u��1������AEsss���D6ss��ȡ��o��<���g���e�]^C��wwS��j�����Le�O�2�������шd�Ug�FԶkܵx��8	R�
ł-�����x[4�BqZ�)P���S��6��_��'9��L&�����Yk0*ٴ�uVx���Q�G��jyn;��:z���V9�'얥���Ȫ��"�Mγe7�7�+-��J��Pj)�;�7׽5���l~g洵v�&vΡ�`�8{��T�>:����Y����j�>���ڗ��+z��MP�����b�7hp���Qj����v��0cf����R-�g��ѕ�.�"���1��IY���^�;Rx�k9�O��OJ?�E�m��mƇ�j_��Y���ɨ����㤷��Of*��`+��o�b�i�u��TDq%�D��yϷ�K�����U�σs����-Ϗo�$����a>l�6݇���F�;��^��DX/�O�Ǽ��M|=j��Z�/��g��! /w]�E;��-��e�8ҽg�3Jw�7|����|v�z9wJO�u�������	0�^��t���{o�W���;1*�er�3�	�j�:��9�?G
����������F���A��B������X6��?�[���,��㸔��-��C\��R�,�� {)a��!갯�t�3"s��|���5WD6��O������`�D���^yF�6� ��2�V8��2:r8���_>v
,��`:�@�{�����X~jPw���z"�˽8`h�r\�|�,Rh>qJ�i3a���
�pn���\Iʋ����2ִ������8}��OLBU�LlxC�65,�
	3q��Z�l��$eo����H����^��d�X�����2U�+�~�*�w��g)\��K+��G��h����ɷ_hl
�Č�N{�u��[�5f��߫�=|��?^-bSN�A�?�ߟ,R���s��q{/��1F���nƨ�Ũ�{��s�r����f}cd��UAQ��q�3p^qB��U	6�6�5���?*X�f3�T�*�:�(`��Ɇ��s��b�Q�l�گ���L�d����rͰh1��t���yO�հ�0�'0�oOX�֥響��#��ϰ�w����N~%�F�t\&�-�=|�ő�?�t�����(����yf_2�^�zf!5_8��r��[�OB�b&��n�����2ؾ�9�靼�>N��r�^VQsY8ʬ��φ����+>��8��;Q�)�4��h��s!��%X7]4i@4��%��G1���B�)AϚA$P9�癞��kO�O.�*�hzn!Ѫ/�$��'H�\�0�ձ^�殉�VVI���P�i�ӐN\"#���+@$���-��X,� �J�a���e����������ܗ��bě_`�3j8�g�w�Bm�z�Ftkם��9�py:~`S �����y��e�����b�B���4��<-��p���O�Y��A�N�f��"��щ����w/��Wſ����J��o���INb.�m%OV���N��<!?H�b��0�3�hp1#^ڮ*u1�74r$u*u7��ҙ��y��m;%_7�6��*q��c��!p��-���٦|K���ȧ�s��s���H��p+��R�v��d�s=�G��,�q#�qz�[aq��Vr�a��s�]�*�,/����FQ�F�ў�U�(eaf���i�ZȞT��鱳���}�Z����Q��ݧه��I!�d��[w�[h�&���n�6
��*���;q��a�M��F;߸Ͼn\+��6N�I�,�$���O[��LX�$�1�7��h��ۍ��q9�_RH&�()k�+h �
���
�?4�[H�f�@�X��*% ��,H�ѫ�~@���� �"��	�~���lr�gV,�C���1�����f]�8�sq��.W/��mT	�P&�P��s�V����u֐�☾x�']�8	 Ȇ g �a���5Ϋ�n��8�R�wO��ݮK�bz�4�L��d�/>v9�5�~���,G�Fҽ
MI��� ��'g���S��F#ꉶ�^��Z~��ҽ=iF`b���!���4M�2���y7��0!3TT0[f������G��*�Gs�r�<���W�IBspX�ú7�:�Ѻx6�z�qp��n:l�$e�:\u����/�����J������Vկ�^��3K����^4�������H�u��! �� �O����Ȏ�@I|�i_���5��c!���kb(Vz�y��kP�Ao����R��	1����C�`��!��cT#�<�to]�o�ث�X�� �%�ƴd��e>�p��M��l<=jS�%�)5�s�Տ�UiA㫾$b2����ά�pK��c��2�??��\�dj��M,"�2!j�J-m��	�k�޺k��u�e�塶�c|���N��H楗ġ����4��p�"�/��Lz���?h$��6����	hs^��1xL�=�JG�y���X���VT-�t����yأ�:�:����nן�b9����$J?�Rgq3����~'�q^�.#���s��u��yd�V��e�j�Pͭ���p�)�O��>��D<���h�X��`�-�y����cnӝԔW��Y���79���ـJN�����������W|�BTnV��OrL�'�w�ږB�r�
�F���8�/�X�nZ.!3̉�fPR�:�����:|���<�Lf\����1�<�����0]i�!b֕���0���CF�� �V�E��Q�s���\�5U}���D3�j �_�=��
>E��ۻ���}���0{?^��9zA#��?:`\SDs\����ey��Hy�X�B�6I�r��U�?a��œ`���&(�Y�Z��ِBmfn�C?�E�aW�A�Md嗰�pKq��oޅi9П�ux�	�e˰+_O�B#C�.���w`��Oi���#W�����"��@5����2���~�&���!yP�mq�K��f�0;��zU ���mO����<��Ë���7g�q���t#�t|�1:�e{	r���Z?E	�t\�8���o&�$�!B�Br����%���|ѳ��ALiv�������3CB�A�wUU��wo��������S\���u����[�ʂ����p�e6ѹ�^��uJvvf7^�k)m���\C�ǩ�Yb���LM����%ZG�㚹%ö+��WV8x)���
O� ����
M�_���v�P�z�Z�Ln�9<�����@��w|j��Ǽ��w��X��`��ߌ7h4OR�O�p~�xg���e�4R����JI���o���coht�s�.��6��)�+�Ʀ���w�:���Ӏ��,O^�Ɔ���Ĥ����@&9����J:�N�Hyɲ\~3�H����A[&,S�101_HZ��c����`UӦY�]��F᫬~������y�֊o#�g-$梌PQ�NV�?�Z���5�p���?T��kon[�5=�M�'��č��2�}v���yh��Y4�?F��gtq�v���ɼ[��>�%N��������m8b;�@�	�_�M�_�]/�/���M�W����W'k��Ǐ�>N�q�?��?j�ܾۏS���X�x'E^T�|�6���Q��ػ�&��߯��[�˯��6*7��ϰ}s�ćeN�}�X�[��L��9�0��?aWK�R���.j�c�F6�}���q��4oC��ŕ��������$���ۓ��4�o�5uYh����ˋ�ƭW�⟸���7kKKP�R,��7�j�JF���e���;U1�$S��� �A4ճB_��Ub4c���'֒�qw�^���_�i�S���{�-�>?Zܫ�G�E�W �5d�Q��!5ɋE���a'��h�"XN���?�_�ͼ^tI��L/�?�;�?��Е_����9�,�_�+��9{��v�����6RMA�u�e�ī;�A��oA%I�A`~�{�N�;{B;����WGT�{g:a�Ua����<b�%���D(3�)+�(���^_�^o���"Kq�u�	�p
朣0�fk����߻� P��6�6�����9/_&����Kf��X���"�l@f��z|����6�u��u=���J�)��h8qK��3������$B=2���c�[�Md�J�O5�e �e��]�Q���!9�Gqd���*K(@`�%�������]qT��W���ׇު���;��[S���e������(��sn���jw��1tV}q��	�o�yr����i�:Ͽ��Er
t�u�k�t���<Q�:`��VB�=n�7��r�����-�ֈ��OfH�}�hbe=��i.���H���&,o��O��<�6tm��	��ɠ#���-	��E��������zb�g�Ő��Ñ��ONp2R����(�Te�Z�L��0a
��m�З��F������4�	��_�g1��:�MBm;��k�*����[f�\�Z+��;��`ڒ���!����`+�p�����yv�V@"^��D?�wۇ����R){�n�9��&�ˣrvA
K��5���3��|͍.5�)~c��^/?�D*���!��pv�y�܀��)�O5F�M\�h���Z���K���d^�H�Q��P�s=�M$�2�m��z1�v)�f>s�w;Gh�!j}�/��Q9p�1�b�|�:���L~]�֥���}���|L�c�n)�t�ȇ���]9��\8�s��t��8s+L�u����K����l�ht6����{]p1�'�lt���Y\�ϒp�>�,�9**ު���r��(&�ˉ�oK�4��bK���՟T�k}�)���i�z{��Ԯ���@���]ծ�3���������|�����P��d�s�g3�r~[��/�g��B�&	:�1��=�.�F_�S�\K��+�t���A/~*\�\��_��_�{���o�ԧ��B �"�v�HV�,>p2i|�ߡ�7�$�� >c)��	�AӖ��6 ���E=zG^�J�6�Ck��'���:��
a]�/}Zi7S%�n�A�}���E�ú�@�A3J�x��o'��-�r����2���;W�FN�w8�`���*��Y��i�
°�S��N&��j#������w]\I�<�t?�C/Y�Ŭ�z�R��Le�[G��
=u8�V֤�oi'}cn��.�5�M��A��F��9��4N�������QP���m>��HI��ǰLI��ԮB�Ga4�"��� kf��/��b����Qñ��%�ƚ���[�O�#����Ί��o99�v�Kߋ^y�D�W�� a�MwV/t$��wϗsm��� ���f��E�$����z6����^+z���������"=��Suө�ׅ�sZA�l�V�SS�B���?d,o=��/2^b����4[���%�!#��w�)�i���Z�E���L<2 (h���Z��n-L�1.4�$T�-��ۂGG؅#�͂@Hʸ��pӯ�RĚ�E��C�^9�߲>]���d�쫶Ο���Y1��W�FHwS���`7�n_��FU/�+��ʠ����,��8;T�|��[n��h-�=��K>��.������A=��-�ܾ�޾�Oձ���ۭ�Z7�ttu�2����Z����z��3H�����}�ծ�ut\��Y��5S:$ߚ��_�j�<�*�Z�o�$<T�rC�:w�8���r�x�����|������T�Ӭ��-�u�V�Yu?x<���C��1��|��v�S|�j#($7!�?/)羅~kp8��m鵋~+L����,����%�����{6q��s��\�ڢ��	��O@(2)�����Y�4p����a��໵S�|��%�~���H�0>,�O��@��j����@����vٰ!хj���h�,-�Z]�0�Lu:Me����7��Wm:��*�(0!d��e�F��0���L��q��m!;rg�La��y`ex�a: 	�`-�-���J!ԍ��
b�������c$��!���?��(�m>�B�B?����,�����<�h�G/2N
���C���)��I���c͠@�>��������0%o{�[�*5�H�������B�R�hz��T�np�s}��B;�U�^\�B�z�x������= ���|��3mA��k�W�r�]�Q�7l� 0%Յa:b��$��8�����%9�k�1/M���Ll���>U��&UO���k�<����������M9s�R���gC|x^�ps��JK%�j����S�I�m�o����z���M�=ۥV}���}��h}J[�<�~e��Gu���Do%I��M���D�%�(�����y�:୨��<H������_�ʐ�7W�a�d���"�UǄ'it!P��^&�)���_=}�;J*G� ��2�!12�g@��'��dS&���f�˴�ļ�v)��dW��z댈!Ƒy�?��gEf?��3��aT��sLbh�m�K���ȝq벐ҽ��4ص��b<�1Q7�2��'�z�
:���c�¾�j�ʛqZ�����<����]�&P0���/�P~P�=�0$,&�> ��ڲ�E'�8��+9�zp�-�i��C�L����ގFC�)�g0 :�ǭ�:�o�_D $w׃?/�/8���O�s����֟�D�Q溷��8zJ�#��l�S$@�����Cjmet�lKe�w6��-�ؑF���Z?{Y���Ow'�׉u�7pg���<���bA%����e�����?7Va�p�w��~���OL�`�l.�@����#����{�I�J1�P���
��ȑ/�@3F���gU-g.f�,Y��}��_�
W�m�9�S;k�U��A�ۙ����l7��< �W���qJ�f�唜��;�RA��Q
U���&�����^�B��ɭ���_�c�)b�}:h�?
)Yz�g7�o�ׅ����S�}$���k�[��:�a+v�t{|1{|�~g�׊ً`^ul]@F~!���W�w��;�o�<��}F n��^b�� ���k�ՓO��+/�+�����I��\���?�fo��NP�sk����qt6#��d����\�^� d�n�uj�T�R��U��V�:,���!������]�$3�Q0��@m1�k��6��Fl���tZ�ЋT�9E/�� -�\�W�) �S��H�P%b�r6���?����eχ���`�Q�״�Ѽ�'f���X&���K���DH*i�N�ϵ�x��2ϱ�@
���5$�x��`�[-R��j�gW�y��X�{��Dnj2!݌'4�n�'�8�mֱ���?��J�p%�q�&k�(m���1=��BI�ر�V����v6�(N?�I��L��$��`1�O�����!��;ߢ��?ͧ� p�M�H�E�g��>:����w��~=�-9�ϏU%������L!���(�ɾ�L�8���*|�#���y��d��wךdjFAY��ݷ��&��q�ꬉzo���^��ʜ$<+f������8���c�*��� O��gȂ��, �tD4P@�6⃉��Ëz5�'�@CԪ���`��N0�^+J4R���i��
-Н�t,\�[�A-:�#��ί�i�/ER
A�VB�6"��ɛ�ɖ3�6���|%|��<�r��a͕���N*�s�����a�Lޛ+3���P��^q��Hp�V��,��\)�+�-�u�������Ac0z�i���XG&�&�|.�:��Q��Z=��!���W�Bv�x,�L�	�GZoX;���x�q3�wj6�W���g*hK=,h1C�5ts���}�/��2p��2Y:@d=����"?��:�d°��h�$�.�l��fm����	����b6k+¥A�M��/�>NQ�<~�������Fx\��X!+�0X�U�|������:�2�|!FQ�N���E�X#o<nY�a�w���W��qz�&��1�L�����M�	�Y���C�����.�~�kn����m��K��4����O̺� _\j�/%�ܵ�<L�n��<js\�o���h��4<`��]�7Χ}�H�p�π��R�/$������_��9��K��z{C˼�������X��ĩI�j�.����a^�m��X����s�3#��f�(�I��ER�`�g��+-�G�
��D9w�'���us��6t���0�f��et\!9[)�+�^��Y��~��at���&	2T������2�k���I�{/�.;�.��(8HB>����FR-|�2�ĕ�p��-��'e�e��H�䜌�]�3����@_�kD����ʩV7��C�j���:��\�u�$�J�k'�
�H�����B �ڬ#\�*Q8�C���x\��D �����Pl�JN��Y@�{����&P.���U�f0�;H�r��^�� ����Sag��]�2�Q�rM�q:�L~�ah�]J��e�ۓ,?�4����'$H�K��$=al�$�[��6MǢ���"s|��X:'n�+`h�i�`�Y�Ñ�`@H���X��=B���̀��xwN�� ���,D59�7�
`�;�������tZ��a�2�y�r�/�jZ������Y�s 語%|]��,i�Ʊ�9���3~�f�Dgӷ��N�s�"������ӑ7��q�s |O!�'�߂�hb�d+�AR7�c�.��;G�ū��@�������le��Gԓ��%����k���Lfr�x֘�� ���� [&D�N��+��@�a`� ���HH6��pƁ� >�Y��j�SV�]x��g�N��Y�S{mP�Drd�+t���(<D��I��k����qR=Ѕ�jϬ���#ڌhZ�з���MA�'�ai�L/tM1�~g3$�VNs,�7@``���\GCH�����?�P=�:}��.��>���(x��)��!H0�d�%X �"����lu"��8)0�x�(��Ŋ,;���"��&d.�0��@r�;ϵ���)ں��W�L�s?��0��ѝ#���K�!N�͎�0��	�罥�m;��9z���/���x�~���x����\u_Ϋ�ꍨ��C�kvra�.����w��Ci�����й��zP�gz�l�߯�n֣�>a��p��G�+i7k����ir6Q����T��Dn��#Ue���BJ����뙫�GX�Ւ9�Q��!*�h� �2k�=R2Np��c{\�A7G�>W�;!����r�dqԖ���[ӨZ��'!	�@��ĬͶ�����u����I?��V;zq��q6�s���F�U�azl�i���4�0�t���3�����Q��s�y�~�r�9���*\�K[����
�y�w*�h�����^`U��f�2��^H��]耼]��YY����),����L���d$�a;�f���첄��:��f����Y�	M����)�Ԕ���6��e��MY�emw��l�-C������K��}n�'H]S��
����e}X�w#��d�7a�.�]\�ܫJܦ�^�+�tr�&�50iUB��c�Z�u���bb�j�n�˱��D�.�a�^F.
�7D�x�"���L8 ���'�*�7�\m	��VR#L2����m��zųP�<�gb�{+�eT�$xa��]�����jzq���	5J.(jP���0��@��;mu��!�XJ��Ν���LX}��.�WЏtp�]�j��sѕ��΁Aρ�&O���D���
�md�gF��\�Czk��_���2�Sy1S@�02+��dH7`}��',;�q�r�`�]�0Ɠ�f�Qj���Adi�_����ޙ�ڄF�f<�j����_v�X�؍@f`�,�_6D����5A$��X��`C� �L��*g���X/���N�-�=�{�x�P��{SoA ��U�c�y��:���@�B�B��\8+s4�*Ԛ��D���=܇�X����\��o�>�a���-R��MT	�G`B`o�p>b&��!MG�ڂ��b�^�ɌK	�(&Y�|��V3^�Y9t���T��Ҫ[�9_Vw�K����ud�1<uL�ͣ6c��Tn�l\��o�N��(0t�<�U��Gj$~ٵ��+�ے�|ZO��4���G9��u���&��>�˹����qo;k%����1^�k}�Q�����KᚫV~����x�k�65�GF<���g�Q!����#`�▯:�tX����!uI��w�w}��m{RUv��7�!�"Ui�|�L|簑��VK�.�?�c���%�ƒo��qj�}PBO����.�k�o�1SaJ-�x�8�_�i�T�ۥ�j~�7P�'Y��	�Q��ar��ި��$E�Q޽���\x�NA;�'�Кg��0�h��҅w{��cƇ6��v�׿Լ�<~C�֋���|9�_k�$#Ȗ�L�|eB�p^P�K�7$23�L�Ň�a�~2C0@�T������LX$��h�u�&-��g!�Y�P!�au�3r�^��vs��o،�r8Z!^�/1)�Xɇ���l�]ܾ�8�ᱥ�4}aO������M���ޒv��H����t�����VP�	�!�a�Gj.� RHT��������r��z���׻�y�g�iv�8�c$HI�8TGL�Ol�G;p ��6Wiw��4�#&u�4��
P�*��v~nq���m���v�j�L"6�yZU���*�{n�|o��Z��?��k����K�d�z�Tfdߟ�?,O�=`K8f��f���@�Z�~ۑ�S�A���W�~m�]�=A�đ6~G����^_z��tn���@]�u�.۔����0xpѸ�qJe�R:��k ݕr0x��G���V��qt)���+trL����+���-�G*d]�`��Z,����VҲ�w��aVw`Y�6w�t<�
���[�~�:������)�v��f���ls]Q|�W����ѼDh��XB��!^�(oPö;��)����m ��!���fUM�2�B,v�^1�]�<rB�
{j`a�Fv%�_9� ��|�0��a��@�qJ	�3��^a�w��Zc�%��[%*nL�����=�e�_o��|��>\j�;\N)�mG�
�~�B��]91*��4��]Ʈ׍-g�΍��Pd<�7j,{W��=��-�+9�&A���V_����^���D([�oS\��`J�]�z~a��B�1�b��p>��7
�k��w�ܢ]^�pJ���w�yp-�l9�����3h<lx��{�(!k�i��p��L�ü��b�P��mi ���Y�v��D�A�D�Z��璦��2��Ժ?�N��ds�J��7�u"�jd�U�#�.,�$��O�T����1�Wz������~	;x�YǊ�{��l���㩝ɾ�ULs�8D�0��X�y�E�[2Wo
�'�VNF����lDnā5����veB��o-���~�^H���S�U������!��oа��p���v�G�*D��ȧ� 0uV�Ip���� ��-�f�v�$ڝ��l=��W~A��@�?�'�()��M����<�逶,���d�@�͸��7�%=�����WX�ȃx?�S�k��h!|[Q�\J\*���Sf=�xǌPU��C@���m�E�I_G�������V���
�� ]�,�b���ޥ�yn����}ٲ�	����� ��	Q9��.��>Y���fgW��K�-��Ҳ������bw��/[�qJ��T�S�ٿWҥ����%-���'Cؙ��4l�;I���Oizu�<�X1�"k�>��D7T��D�7�A�$�rO5��?֏Z�7��@un�8r��E�7m�����8y��$����H�z��Y��2���Fٴ0��L�q�h�ǋWM�Fk��,�Q�Y��ML4h�r�$�'C͍-Q�-U�Њ!��H�r�>��@w�Xm՟+a?��F4}��ԋM�ٖF���~��W��.���h��A#�$�B�� WG5 MMJ34K��u@E�ױƁ\c�R�%l[�~��6���Q���W�Ƹ'm�V�Ę�V��rs[��*�ox��b�V�!&���z5Q��8?]를��Jj�����rt5�坡��7��P�(׸�RH��!�H;��Nq�EO����h,^��J	p�mإ�i���v����d�-�z��Jq�s�0=j�M��qǈ���另��<GH�ˉ��o���2.�;w��T-J�[N��oG��W��$G*��]ǈ���ص�C�mz��:�U��� �%Q��~�F�Z�g
Z�Iv#�q0�/L%�Y����X���d�1��w�����ʃ�L|�A��&<P!j�J��2��~<��^��܌O����S�����7�=��{&��Od(��.���&���<r'�L+�h}Dj���&��~d�|����{���B;S����z���W��Hu� ���y?țՌ��E0����V���y���"�υ���,���rܹe��l�}��:V��h�|����{u)�)o�ZA�ǪЩ�+EeI*�s0|k��<�(~-��B�ѷ4}�{ �*zI��F��;�V�u9��/��n�6�"�Y�@�_F�S�M����Dd�^z�!��01˜X�Fv�sb��?�.�V6��yz��/'js5U�3ZBw/�Ǹ����x{q����`�Qbm��'?x6��uc�5\��:y3:�/���Ɉ��<�~5���e�Å%t���Ӏh��$,G��4��(3����O����y^hW
��.h�G#8�_>H�R�>�C��M@���/���_���g���[	��Rw'��.fȠ��è�	9,���X}u�4L@�N,�MNh/F�ĿJY��_���n�8��C��d�]���=j۲VН;C��ãh��
����WV���@/��2w�W��h�x	�!aà!iTJ���L@�!����\v���[N?L�3廬� ��_��@�˗ƄiG֘3ڥG΃�*����*4T+�ڃ�s5��QSL�����k�뫝���\K���]*2P�ޏ�ad)��<�^y�J�	4�|�h5S�q{@u������d& �O=�og�s	��wi3����Av\tYv'8��OZK5�t+w��k��4/c�%�M�d����֩��I{�����!�M cʑ���`Nb1C��½1u@����Wӯ$��f�	�N�� �3��BV��>ݻ�"_���?��b�^�(�@dS!a!⢦�3����7�I�5�K�� �iruK(��{�@�r�������]+5]+���KSM��MN��|w*nŗ��?��SN����舎��!?S�p-B�o�Q��Cm"3.��>��ˊ*���ou�"�7�P4:�EcU������oP<N�@زk~���/���_��>�	(W�l`�#>�i�M+Î�q�ѿ�����6��
ρ%��%�<�B ����
��3�?�T�7�#UFQ@����ˤ:����ߘ �>�y1��}��KÞ�+!-��:R�q<I��J��s�� Ҕ�J�9.�E�g�;�4z��S�ZǑ�4E� =E4L"l�g�\�I숞4� ���	�W�q+��E����}�)���w�*V�i+ba�Q�hy��͸I\t�/�`�M�	ޝ\�[g;���l$z�7��%7袓*�q�Uf!���G�������3�閈̧���r����}xp#���^��7��D�0r�x5�O����mW��Wo�q�~�2��fô& "��`Z���Ciþf� P���ݠ�1$�p,U�����3�w��3���?v�����
_�T����p��KI�sk�۬�����H�����i�J7a��W��t��$��	����S���T«qz��+�	�ye���&:�P��aA-�s��,<l�x�	5���Lh���a8��i:�ʢ�Q-"����jJY�ʙ�؄L���@��A����]����}��	����)�E�o����x݁��n�m��f1�6�$?Vϯdº\EN.�)�^�����XkT4���q_�VB��M$q�q�ݯ�ïɫ���6�>�Iw��Ϸ1��L�j���a9+�-����Q{�$���~S�w�c5�u`(;3�^����н�l�}k��qfHz?���yC^��-z�""��r��S�%{��Mt�F�:sڗ%�JV9��g
�V��Է�O����U���Ͻ�>,]EJ	�H�_���HN7I�8�sJ�G��R9�u9���n�"N"dε��*�n�l��+5�oay�5&���>�R�D�
���i�#���rނ�g.��$<굦�4��l82�q�^OQ�4�h+uixQߞOi⥳x��p�aw�\8rs��8�>�U$:Ƞ��*`ᯒ`Z�.{LV��5�:���Ԫo���UHCdqA�7�nЫ/���q�=��R�3�C�pA�v}���4���8���8}��kx�����0�
��PQh�9֑��j�fx�7�ޖ��)������ �����E22Ye�*�`%;�p3����2�u�Ĵ_]C��4��x�F�V�e8s�q������xu1U�D⚣�MY���wbk��3Pl��D�k��g�(⟌`5�bx���� ���h�>}G���KDn%1�� �FtʝƖ�`�CfQ�;��i-������"�T�mO�� hJ<��]�,��m��e�f7��V�$+F��oBh�����7&T���2'��r¾��~�ա4xҰ�=/maǞ1�$T ��*�C��+^���=��q�ƥob�R���3^:�V�C_�r�oɦ�Sz�}�\���a���J�rFm�Xu��̡��o2�Q���$�MؙF����`��3�>��G��T��E[hՐI���1:������g�9$Pq�j��"JΛ�"t���4p���V!�G	s���k���y��Lk�{�l?���(�T���ZB� ��NV��5kn�{���~ֹ|;6X	5�I�'�A�xD�CFyS�\˱ ���?C��CIl���d�j4�\�<������I&0�q�DnP0i[��
,��w�%�b�}�a_�ox�& �Mq8�Y��w���Q~L6S�Å�ϰ���>�8�VD�Q��=J�����.�@'mk1F�Rn�Π��A-!�Dh#!�����������<�L�M<=�d����Ҥ�E�X�R�:�S��*�j	|&ϮqgWխ<>��"��֊KϾhӰ���P�d~E7nU�\��ҼK��������	]K�MgB�'���6w�wg�:��/�L$��sN8�mv{�]\.��
��ՠKpp��}w5��Y�`�t{߳uQ�Į����>�:S3u\��>�V���je�N�`'D>���璛�Y��S�wk3�A�	%�A�1�ӫ���Q:Bb����x5�*�w^>��g��>~�&k� 2���ұG�Pi��-�B��d��l�+��6~Fk�9�,��<H�V���H���$�S��X���3�k�u��h�'7�5L��ѝ5�Vzo�$�ڝ���u%[���+zԳ��� �����mR���"k2o�l_olx���8d.wK��+��Q���6J�x�V0k.�S�q�h�c��Q�C���|�D�懅U��D�;�Y_��,��C��hx ���e����U������P+����X]� ek�+Z�^��&��T���}kq���:^9.$_1�9M�.a��Nϳ-g���a;�w^�^��<F�p4n�B��4�+;�J�*�+^cE��A>orU��:�~��� ĚQ+�wS�������_yas�Vc�<;����%����sH�q���}J��C�/��>b�Yj��O����p;M��9�(�~0�;|Q�Շq��'�׮f��
C���Ç��[xC�lj/�EՑ��:�Nc8����?V��I�;���!�$�ʟt�/@\��e��TN��MK�'X�w2�a���K�!����5��UMLG�-���ee�{WF.�
���r͠;� �ء�*�Hy�e_����Z���l#�b�yYo5~���AuU�Z	o����4r�[�cw&�.����n.N���{��_f�6<�iw��TN��Jvܳ�zM�w��F㒹p�r�_S�����KM��%u�1=��Z���6��a�w�����{�7��&����؉20xc�VYX��܁��C��wBOr1��rǒ�X��b[�����#��^�.[�'~�z2�ʼ�Э���΅w&SKC�:�+ݟ��Ty�U�- �n!�b4�I�����\�8��E͋�$���G��	��LO��n��e�TE��\�����+tQ����@a�2�Y��GӍLr���m�:k�I	'��g�'����<@;�08�V=F{�DZ������W���e43T)�B.Z�-ȩ��[KV�PF�"?��n�F�+t*��U�Bo�D�k'���X����5��;��b�M��NÐa�;u�O7��(���3�*���Ժ�G"�w���M�b�ڗ����c��++�[�|f�����ִMNC�������i��#���S�q>�;�&u�����g;l��cŌQ;��R�GBU�-AE�����k�U5Z�c��أjo�����R������y���_��8���:���ϻ��f����G����Wi�g�Bu�^~*Z�C@i�z��Ev�V,>��-�8�zD%Y/�$B�$�k�=��b&���k��Z��������?�9�s�^�W��i)]�т/�T��C֒��l�!Gh�K�l�tU��Ro���,*����*�$3�E���y
�*0��Q`���sO<��a{���D;o}V��K�w���������YJ0tW�/���e��6<�'�mA;�	�`^gZj�!�������B�I�\�������l�Ay��݋�@/��-L��(φ��a�G��[l��j��ꇬ_���O�iH]�x��nR�%��63MA�S7�o��c�.�QZH���@�p��{ng��g��LԳ�ps�j�H���7�Y���K�0a[*�~�@ d����~p����DrI�����j��
�	<Ul�F���	֭�8(�Q���Q3�Σ�L�Rz4`�J gj�R�ףo�P�g�@��$����,;J��ŉ�?Q�t�]�f NKX�Mۺl0�X���H�w���"P���t��+X�-.�3J�!f8A�����TG ���#K_�nP�y��Ν�@�?�ExX#���9��5�7�ΗU�y;G:l�m`��RQ�1>�^����h�����⭴NsD�G
}�E���i��b�P�;o��~�%��!�`�P�d��9w��iι��������z毕�Q����#�Mz{L�I��f������:�2>�Ŧ#L�.�4�z�Af���0��)g�8��S$���,�z#l�4�!�/�,޵#eֽ�/O?���Z1���.�vX�9���Pcj���,�''ze�p��g��!G/:T/>�G��~ѼR�$KL素��'B�����/3�u=�#%pc̤0������I������MݤV-��{EhYE�ْ��>��@�����HC���5sil�!ծ��epg�4������-����v�_�G9}�O��9|'	.�� �|Il�c����� ���&��oD�U�̩̎�u�:��-��_�v��ya���|���:L5z�f��C�dK���>�7��[���{�|��Ƈҫ|7A��	�o�&�
����_~m�yY�Y��9�̰��ͻ�����Ť����#_�;h��n���v�U�M�!��ך�4P�l<��	�U�:>��Z�;�˭q�c>i����N��헟���R&^��*c�%�q�e��=���|Z�^U����?<V+�*�k�?�1%?=���*�ࡎpy!Pg�9�����Y=�����zvFa:�I��N�� f&�u��2�\en�+����a�Y���P%���`DR_\;N,5��S�����F=��+��MR(C�/;x�>�݄�Ӌ$mF ɜ?���bD-*2Yq8"�����S�@LMh�"�SK�H�ݴ�\��d�o���n%uw]+@���N$ޏ���B�������$�y/r12R��(�V��ЗY^�)�}�QVG��uo��9�����?4����E��� �G�ғ`:�E���ew�82Y��X8r�2i��rR�[�d��E~���@^�!��D*߶�r��UO��ٳq
o���r��%0�)Tg�8`���R��V��&�E��'�*�J~v$E"���R���ٱ!����Q�S�a�2п�2�o/8���"���k���p��U$�\:����[F��8z��_����F+r�]s8-A_����V�k�u9�J&�s�b �?0Cԉ˂G���i�x��{.�Ta~�R�I5����+�$X�C�^����.a���.���I��zWٸ'G9��z�)�T$}$tHs?�����?�8���_x� �����r�89(HSd�h��)�l���P�Z&O��r�I ��/0�xCDN7~��.���~wq��-�DƊ\��V~Nq`56�g�S�钦�Kt!H��I���R�u�-<�o��eQD�5erp���J
)G������Mdh<0��^�;j��x�v�kr���Ѭ�����ACC�����&�mNɍ�l[�	���&ga�_9K��x)���B�ꮟٯ�|�4�����9�L ����ߟ�$�e^q��Y�o��.رѾ,Fu�uwf~����������վ�e�h���[��|1[��6��=W�ٻ�'�w⩞ѷWtZ�d�@���jp�7[U���fY�<N�3�3FC���m\������`$cf<z����b��/�I�<i5�Nbc��x�T�6Oa.�����0���%O��z�~>��)��>��Α��HL�b�}��ٚ]��5z�5z-7�/��z�Q\t�Z~�=���B�{93KGZ�_.����`�qB9�-��qފ6{�&]�bRi��~�ޟ��$���1/�֏����:�������v+=3��5��C}w�nF�D�$酑�b�{��Q��Q�Լ��xx;��ڢJ��9���^)9����[���>";k�Qܟ��mz����}iu�w��T�*��~eO1DXV�C

�qA�0t�ˠ<����n��(���%��I���e���5G��n�Z��Mܴ���Z_�V�6|� �����?l q����6�������$�4f�Ä�)"&����}d�����B�����cl;��W�v�3���Fl���z�a�<_W�M�������3b#�x��=_@�T`����ݍ����w���p����5�S��?5t%^��zeаm��a�{֑��9���Q�IE��8l��
�aV3]Ha�E�����έ����{�K�x5� #�fy?#~��:�'�	���T�N�k�~t+���gf��wH�l
:P@�P�Gs��C����׊?Y��D�+��a����OC��SS����]�E{C�u�di6���
!Є�� **ZZ��m��t8�4<�]���Dvs�}�d�i�eq����$&�(�P�-vqF�Fh��)�O{U}-Ve��;��Z����鹵�ݳ��2#�Ϙvμ�N��N=ݒŠ�(�H��ec?��]}��ϋ��\�s?����oa����y�����OӾ�9�}BD�԰-�m�9�,�-����|�XIy~
c��͆�jA em����o�W����'|������-�l��"c^��BW��h����Δ����=y^�$�3��	�=�R��珑����G�_`�{Hu�U�8~p��qt"ڋ��I���ܒ��GݫM��N�J�}V�v9� >�$����a�������������%�.������\�����l�^_���9lxd2�:��w�u�;|���;�z�X�"���T�0�SM%�6R�u���j��f���.�J����:mb���}x,=�?Z�@�E���e�[$��|J|� N
�Fx�ʸ ��4c�c�'i�l�����;�3�V�EhyA�9��� �n�o9�p/.2��S����R�]����q"HD�bĠ�+�x��3�" �c�$�Nt���1�z�9U��&�w�;�Ȟ���D6�5ᾯ�V/�k*g��h�a'��j �14/���λ�D�0m{wC�[@vQN���̬l�ݧ�Iࢧy�t&1�8��8]�M� ���xz�I��#E�B5�w{<��)) �ۥ�Nx���������4;��0��j['5�
4�og��,�vU�/��7�lZ1UC����B�]`��R�&�*	q��}%�|.�P�D�VФ�-A\mz�](��/Y�6�/���=_�� (��Jz�/�;#���J��E�a���(u�
�}��ן�m�7Y��7�j?��%U�-�\�.��k�
�<���Y��N��rF+��#����W�[�Z�t-r����2��G)^oE�h����`��s:�	۸N}�$�������;af"�ַF9k��E��_?�5mi�w�Ⱥ1��6!�!`��ᠯ�c�7�|Ӂ�h�-cv�@�������mA���̜y@/Lux��o����HQ8qF�Ѳ��=��߸�h[�����d�;u���3�o(Oh�ch��kl����]�9�n������QCn�@��Վ�~�����D���8cÛn���-�c���K�i	�����1�k�O|ʉ:ֳ �-P�R���'����_�g-��ubNPj~*%\�󷞕�
��`�aY���Q��N��ejr(����~��$���U*˂<�-�+��Q��e�ڵ�S��l�l��t�AD0@I�tG'�-����Ã摒<�02�!Ey���7Mu�W��%���}�c��}���Gܪ�Q��M1G��P���O�d"w��Y��$�̆�R��S�=RU���r�d��Y�����H����v��J�B�}o�' �-?�SX}ƇC��(��d9��s(�+uR��	�D�|\�a�{� I�<Hz�p?U�	;���7q��c����UJR�ڞHH�YA�@�S�_�W�%��BD����Ra��'������1�o�W��_��M�m���p�\��iY!�d��6Y�����X2��~IW�ps����&v8~&���L	��y���(�"c�r���U��>}�HV�����V��b�1p��|��x?uL#	b��dL�;�IXK_�u0`{�!o[A��z�u��-I������j�$ԡ���S"7y�{)z ��"	����kː"�qA��BG!n\�ШpC�M��X# 9�u|-�p\s�=�b�����e�^C��d߼�:yӒ\<t�b���Y͈���������04#��]Ol((U3�s��F+��{��z~=���ۮ�%��%��� -����[cٞ�ͽ��"&E�+����,]�ݳ�� I{�Ȗ��٫d�7Y��פ��8 2[���uyہG;)=�����5���{'�A>]L&��Z�(|`�eY��t(�Ȑ���8>8��!�&�s���.Yҳ�)f ��`b�RC��[��	�M������-$���ӽ6]{w�b�s�T#m��l_���*��yo������;������c�:��q���^����mxt�p�~�'�qyd���� y��\�d<f%[8x�zp��']�7q%|URS�58�_�h����z��͡S��먒�Qa��fGo��Ns��3t,_�x)��s'�W5C~!��a�=���I�T:�
Ty���w�ʝX�s���w¼��O�ۤ-�k��}�q��ӑ����[=�5y��X��#p�<�5�{@3O35�^V��n������)�G���y�v����<3��E��L��˯~�R|���'�N<�z��}��}�6���(x�k��)�����T�a�S�L�������94�(Wo�8��_��E�P���s�9.���@�gn��\����JD���ym��$�oo&.0)W��D�Lx(d�M-�4G���R�5c�rlk?3Z<��Ћק��W�(��U<Cb@�(�/E�^�O���W��qN�A���OI�>�R�λ ��HI��/]�AQ&R�n�-�@8�d�B!�I�$���k,Y	_yd{Qk<��WQԂ5Ӯ��ˠ����`ʵo"�ْ�� P0�/�?�&���#����:5��g��^U_*/�,��M9c��b0�9��J���#���q�d�\Z����C:'D��G�� �B��BE|}%|�-0��� �����\���)w�ڮ�|_�1���j�󽥼�Ѿ��KA_I���'�G/�����3MGg��<a����ê<�6��<�c�Dћx&��p�h	�ܚ�S6���:�������$��|�\�j�����������oP���,_�ho�W�����̏{������x��]�H�}_��t=���Gjueo���}\V��\��ǡ��2�E�L��Ƴ���P����B39>�����[˙��N�X?-� S��Ǣ@V�h`*���麐���(��(���� e�޳x�f�{ՒvC3{�vǢ�5̡��)�g���9���Ǚ۪�W�=1F|k������Z�p���~�[�۵��`�ȥ��c�ś�J˞��ʒ��ZVZ���^ ��_ۡR�n�Za�����{��Vt�}ilY���nH�i\P��&�glpY�Xu����$uW?�����㼃���NK8�G�de���b�Cڨe������,���DNʡ����i�CÙ(�g�\�!H�*���� �[���.w��(�#7����.���zf�)u��5�l��ϝ�6�T�ӗZݕ���w�R�
��Hp���������z���\լ[�cV��h0T�� �Щ�j����?~n���[�݁����iVA*���t��s�N��؋�1�}��)���E����(`���-UT������p/���)R��9��E0AۅCс�h�-��	�&�KW��P�@�	�I�>TK�Z�8#���W5Ӣ�S�Vӓ���Ci �_S�Ͳ���b����e{b߰��(h������U���f�:/Of\��M,�r<��zP�;J^31s�I�{�O^�?o=����YHo��z*SX�z�]�����R=�-i���_]���$��n�g�%��	a>�@���I�I"դP���r���Tp,z��c#�$��߃@5���A�Gnn�76�b�WZ�F���vd66=��sgb��y�&V��4j.4���E�,z����'��p�>�8!�:u6=�?\~��OP�@��*�bӑ�O8�sv;�Q�3>%�T��o] ��o	�YS�LߨYT�}�v���(�N�� ^���ZL:m��MF�H�z�K5C��y�b�nV��YS8��)wLi��
"��e�`�ʎO�fb�)k5����-���1][0M׽�y���l*z�;f�ƹf�Ɩe6��}"̂��Cj�3�A�)YU��PԈ	3�G�z{��+�?	� ���}���,Qh6��bj\S^6�Ld��&r�_Vǌ	��?q�w"ȯ ��9U.��K�Y��Q�t��OY��ގ�IHPA�UZ��U��X�(Af.���J�����Ҵ��I�s�9�V1@��Q��92��K����y�U�\�7�å%���������nc����ִ��;8��c_S�]�$8�T5�g�g�w2\yQ6tk}\��΁��hߪ~e�y0e����Iiɓ���jU6fF�4N{?6p)�/��=7k����k/.�ÌǦ�=^�qάwpmBO̊yI����e����Ҿ��ӷ��\8�n,d�����y���Ae尩:?]�?eTX��m���pt����o�� �zA^϶��>A0�P0a��L�������o��s%�3�q2�WŖ�lw���}?zZ����".�- UO���'����ټ��@4�[���r2F�q�l��A��)'a��H_��L�V{�e������O�s�1���u��*�5������s_�g����#�:��X�n)�jNc>(JJt1c��
9�G8~d��S9�����ԯ���K6��������l�C�M��3�OEE+�K}~ ��2k��i~�� ��
��Y�FEf5��n3���u����s;:������r|M��jd3��Z}�-U��<��D���-�(tc�����_G>���Ej�n�)��� I��e�L˭T�=׻��D��%ȕ;��b���	�ᰛ;2`3^��(�w�Gt�ݽ��c��kJz�kx�&��o���s������S���j�bnoI×���ʁ����'��8�kr���z�a|M.A�\�%~��w����J[��/8��X]y&)�KDd"s8:?C�8��\���s�����m��EjI�H��Z=h_��	����f��	�k�7�I���L���+�@+����^��{�7S��:�-Z�7Mho&I�i�	�͠?��_bN*��tO(
{�N�e0ZPa[>/�.����_'_�ψ���o��X",��I<��=6����r���}���i��Zvl��t`~F3nD�˴^]e���⟹�/�	��!@*�e�X�j�����N��4f����]�q"6p0̷��'��N��2��Bv��հ>ݴ|��&�=0:���.<��OM �`�'p'�#�NT�x����K�9������@�����+�-� ���.vZ" ME�"�bm�-L����cl���݁���t�3��֚�����T��7Q�O�8�v�"}TQV�4Cw��&ׄ쏄����I�{��@x��$�D��;[���z8��b�>tC�}�}e��Hx�c%S|\�h�o��i{P�|�&,�N5�{3NM�.¹L��̇Ȝ����6�Cҏ�.��^7�#3Q�'H��B0�Kdh(����@���=xle=4�����~I�P��~���Sd��%�����Y���j�;�~tC�y�k��4Ϸf
�q�����^V{^�X�'�%n�;�#W�kuõ�-��K��	����������Cߓw�OU-�Jk�������~�G��p0�����W���w��q���7g���_���g��Ww��g��=�K'�7t��܋���\ûZ����s��xi�
o��o~�x��)+�����
��sOԞ.�<衿$[�4���p�s�?�soq�rK|d����b�k�*�m̵���/��u�@����xr�}�l���ӿ��]]�'׆�)�!i��A�M����sBK>��@?���j$6O��9A�٥����x����$|?�Ż�iV�ՇB2(,�����,Ɨ����C�P��<`z*؉g<V�(x*?�Q��k
7�$� F �(mdѽ�~���N����o�Q�h���%`��7�l7g��a�y^/F��h֌TZDi$��ӈ�QD-����z�7A�~�v��Gp�^��u���+oH`�ݝ����ǔT��ݳ�oK�W�ua/a����,w���x
X-?�̎�J����f\˪]̋^��q�غ���FR�;�c�&>�D4����A.�7��m៬�?I	z�(����x��Jg7Z^����=���(�y�c,��x��-�iZ�|�`M�7�{L�Uew��	A�΃;o?D�-�`x����[8�!��m���nΝZaՍI���@��w>�ةv�O�^��&=�{â�Qt����{ߝ�+\�]*� %V�p"�ն	�9��)m1(��3s$�_�,�p��͂M�P@S��M���3a���������Y�$��J��d�Ϸ�?)�NM���S�3q(�X�6n���F�F	����6+��#<ǋ=ӛe�e(������a�S��_�X�L�ה�!�S������P|M�I��j�;��
�N.�k���$<˷�2#H�H��(����h�xd����@�u�"���N��b�x��`C�1���r��M�z��a�5��8S�,�a�Ĝ�:(!daH�$�))�@o(���瓻�B����%e��C[�3��6�Qoox*y�0�&��3/��i_�eTXM�X��T��t����u�.zw��x���ǑA������2X���C{��f�1I)�Ǐb�]��+�KWP���xn�{��F��L��o�}��`sO��rU��p�=M��|�D��A�#�b�l�(���'�ndE�=c���'����Q�����} '(��U���]�����ux�`|q-Z�
S���Τ�v@mg �ԏ��#�۔�g�^4?��z�����#����;�������9�����?�w~__\?�u>��Y��H���8=�%C�N���d�����ϴ�.;2��~�p80^��bR���]bn�ǰ�'�{L�9��T�%w�h��n�#�&أ�ӟ\�xaѶ����bJ���m+`Hn)�I�����k�R�,��+2 �R�����|�LMVg�L�+)ȺOqcqJ�a"�*Yb�,8�&��f���х�����=,�V܄�g��|m�����n��J���1^P�س���A�Q}��	ZQ� ;+л�F��C�������$�[>���%���Y �c����0�bi�Q����O4��b'��z|�vy�E謬�b>SD�ɁB6'�y@�RtV����Nx؇{a
X���J��~|À�.܏�HMQɆz$2�
�T8��!��Tr�-J��pz!�Y*m��ia?�Y�Zx/^����ԎKd*�ތ��p>d��E9�BjU_�%|_p4/�O8' �bC퐎LWG�uBҰ����&������?_EOX��9v���~=Xy��]!��o�p7���;���� 0Ś�̞��T��B���	!�rkmϓ6�>+��R��W�5#*��o�)f�$Z!j<G5Y�7>銑��5��p�����]�%2�#�LB���`_�����H9G���p��A�&.��E3�c�6TBqn�il���9��3$��Ip��aO�Vr�S�7qiM���S����MiFkiD�-�#�~�Gg�{����5�M��3�12l���L�8�I ���*qG��sf��4�N6���q��|>z�SU�������b����m��uD���.=]�u��Bm�y��ߍ(�V�lCEW9�K ��Ң]�.F���B��/��~y�b!�a�;1�z���V����dZv�V�[S�I�󩇂��ߕ��.��߬��	~�Y�"-�[#��э��o���R��iK�?5�3�����[��q���n���~��"�*�\���e^�x�c���Ŀa�7������R���o�O<�jepx����9���J1FAgR�+�n%�{!?jt+L���Ǜ���SnϔҞ��֙�ӥxX4�t�'�k�<��məxqղ~��3|m�5��N�a�yl����p�Rk��#�[DF:����醬�n�S�xD�m���)Ӡ��g�����KfU��NTGO�ЩE���b
���^� Y�����??��"e��9OO˫L��rFG��_�W-	ǩ���$�}@��RKՂ��%ȫ���}L�^|��r-v<��w���9�/u��I�8_vw�r��8%�'!N���;2[& _��W���K�!P�p&�Q���U��h�N;ĝ~~\����d�uOj��a�P�i�k�v� ��H�@k;fh2��4�\ۑ�b��@/U�A&e�/�9�u��1(���.=W5���HZ�N�8���_�����/�jڱ���y)��#�����dV1-�a�PD�7d�.�X��:3��`��#u���*���[�bdT�n���u�{���lTs�M�W��9Q`����T/f�q@�e�8vAy�UG,���I?Sf�)+h���'�	PK��;���)��[��=� �j�;��lH�����H=�O�	� {�2�m��SB/<��i�1����yr2e��S�u��ě������ ��6������^���~�Đ�0|�{��y����m�llON�y�ͬ]�������8�R��H����(m1D�&if����J��h����9� ��#@]������G��ѣ�%��'��Я�bq��`���q*�)�F�SD�]�;���4?%+x?�/�\/�w�����&$�q,*p���S��(��ƅ"��BŠ2d7�v�����L�&�KrU֯����Z[���������D`��������p��!�5�x�zU�L=vq��x�g���~sĎϪjP�F\������BG6�ȤY�i[b6� �Z4�]����~�bW�K/W�0ȱ
{�j��d��f1�aB^*�tT͕-�d��2C!��.-�Ǐ��Za�5�x����[���4t��[���ɮ�GARwQ��+rn�'��Ǝg��	4��d5.)��f���|�[�բ��R��W"�;դ~������7�Qx�m���p����Q�����)�C�m�kLn"DR���n`pO���\�t,:��Xܭ4����ܮ�Q����+O�ɘ{�(�O�O'�h�F��Q=�#����"&{��2vOF�� �F#��vRds)D�J�B!�KB��a��ݷ�-��Q�!B�#a�7G���\]h[��/ހ1�rC�9��	rCnη��ϵ/xA���N:� A��C ó��(zd(�c|r0R��%|3�N���ւ����:�}g��2�bޑ= ��şC����A�a������-��k�In�-x��_�>+q��6��|�JJ�1ؕ����)d�1SȊ��t��g��8mH*�3IB����a�<'�焙&Qh�/���z�w}�ps#u�q �c����B�]�	a��vV�ύe�����AiM���s�:[î6���A�Pе�^����߶���M��xH�1�0A�������LV�Q"I&���gF�����c��_�������/��-���?ڠ�X�Fe�+���ބY/���;hࠀ��gX�}n��+��(�#�%��
~h0�?�b�8���N����4g�:B	z�������d@��Is_$	Ƶ��T�l�3���!y,3G�}��G�T�J7�eY����Z8r`����*�3)fuNv2>*�y��b�ڟ�VgBy��đ�Qu@�.�޸k�;i�մ�Y��M���72puPծ��`6�7���&8#��I����͋}F�m��`H*m��� 2�H]ߨ�>_
��X}�)��7ö�(Fc�	<vG����X-�d���hVJ�<����b�}�'�}����C���ӟ����&C�L�I��Z��Dʭ���F��<G����떄i�_B��>�c����ἵW���8-�~l�>�H���	毶(��	�I��_��h%^>��3p�H>Ai�e	nivO�E�f�d���|�;Li����R���Ӳ�E5x�/k賓Q�v涹2o�Ӓ_�(���o�$l�{�4�y1��{w��?�(s#(��L��yJ�������~��׊w焖ؕ������v�Mw��Ch��wG?R58ᾯ��Ѓ��`$U�\)����3>k�t�f�rJT�����L?M���qU�ޖ�rx5Zi���x��?�@�����uR(�S(�:�m!���NW��?x+Il?`H+
x�ϜF��G������ڂ�u�����x�ē*�(��CA^QBQ$:4_��B���PwQ�w�@VpјSԺI��Pz$��g�G�c{26La��9G^^�����M|g�/�usƋEC[齆%���U��R
�����M+{����]ϵ�����s�o��9��BYsG!��L1�%4��Xȴi
M�8�_� ��v @&+i57|I�Z��Ja g0����x��=9�v+�xD+v�V��N-��R�}hف�^tV��ްWM��7s.���BR�eN����|`�ı�E������]!��t��`1��w7�m�|��}'}nӮ��OOo�!�mƒw�Ї��=H�w=���G����,�q����+"QS3�0�A�Q�M��P���sn�4�PGu�i���r��<`���4Ȧ�r����D�H�D��)�����g��M{�k�FrQ��4˙��p
���_�i��_;=��|��CG�a��00�\�xؼ��v������/�?�d��M�e�����1������Y�8��R~Mu��D��,�M+u������P>����8Т8�2�g�סw�?�O7�M��`=P�`��D��E��|]��##A�,�f}1ub���x"��D˚���Q��}Gs�1��S�C=o����fR�S�tcV��r��1 ɾ~0�Na(4�42�[� $�G8���I���3�^�^ֺ�=��v���7�kn�G:�٭wl�&��R��a����WS�2ll:�8��Y�J:a����^� raJ�hv}}�E�������q~-�78��f������c�'َ%I���3�ؾxŦ~�ů$|#�e��_��8D���G��$�*��
�J^�clwnLDo��Q6��
r^̼�u�����Z�X\S�½���L2L�]�w���G�K�(�����E_Tk�݄��8�B��9f0KH��7�H��n�����%w���8� 89�x+/�|�ϲv�̞Mp�%s��-���g�X�)#TJ��-�b���nۓO����˷k��^L�JM�J��(����U|��F�߹W��%�nK������ܴӥ���4��~�ʚpB�N'�^[����n�M�v1��:�*��8k3��Qp×S�3��>�b2�p���X���D��TV&��a�j�E`Ř�N��0�Tu�}˓�P�V˗g$Xũ� {�4��_��rQx�C@�׀�(uO`��ͭ�	���ȭl�C.r���E���,�V���@�q�fHR.��5�gH|9�Y&n!	��+�u?q��'�l��ӹr3�(��Z�<��0�R��%>(�y+���C��:yk��{��Z�q�܎iN�����s����R��&U���-���@�C�2q�r�yH�3������gT����L�~�뿺���ݛwW?}zɊ���G�ڷ�{ђ��<^�$��=��"t`|�f�`d�����K�$�Ċ�!2�x��ĂII�K��ND�*�k��,i�{��H��9�V��$:#�Cgr���?̐�Cv��"��=t�y0{c���NH��/���u[�V�7����w��9 ���4>�+p���;��t��z�Pb݆���\��8�����dX��k��F_�i`��WO�}�B���u6N���]S���ѧ� x�kv�x�R����qe��iZ�u�<��:���L�a���ѝ����0ش�����F��&7��~_����C��t�5�p�����5�-��\�����2nl?�Y�5F���B-,^E4��Jyynr:-���E҄�@�R�fu�Ql�s	!m3�*���'A��\#x��Ϡ$���w%�ԚM"�@��ˏgt�zv��D��ʖ(��=(��sbݪ�۟o�kW�]�*�>�ˆ�%A�\��Z@"Ff%��rm����s'���M��s�yf�.�!��a�O���b���S����)�f䈕���R�����k���B�i6�j�R|�l��u�ɜc����X6q���@�t�����7L��Y��(�d��(8"�r��&�zʬ�I:��?�9s�8c��Y_}��ճ~^�.�mB�9� �n��Z�q�{1��ۼ�4c����m�i��a��o��U�0��	ʨ����|<�oQ���x�C�T���z���P ��_���~�M�kY���J�-�@3.Z����&����2�i�1ÿ�zp��sݬq�sj�Z���̴�j������Vw�f?����Q��ǻ�x�僨�g*�����3�m�αi1,�(6��-s^�����N�z9ې�ܭ�&�=X')1>�HD�����ИmQ�)��Jw�L��ݙ��k�;-�?jX��raUg�KF����ٚH��Km�0�E�<Ʒ5+:K=���ƞ�}�C�!h�d��FǩG#Us\v �vd/��`�7��Ƃߴ�����ȟk�ԏڏP���������4g�+De<��$^�{W��H6~�.D��M��g�Z�B��%�B������Y�̪��j;��?�-�BRu�T���$�y�J�R:O#{B�o��P�E�!Г���`�T��Z�3m�V���L©~b�I?XI����^I���C�����b�tm=.��O$o��0�%˩G�Y
��bft��o���X�t*))�p���cv���o�p��\�C�V7�� �iB���D5�����k�S�1�|Q<����;fyEM ��@�L�� �ceśV]OFƧ�{��+8<�pd�M��D���~ہ��d��0�C��3�;� ���c�t�c���Ω��տ�G=Y��-}�.�S�������$����R�8qnOv�2L��&�fH�G`B1�(��ma��[�Hn[�4�S{H�W�f9Y�q�KP�2ц��_�O�UA�d��Z�_��C9��>S��o/ s�Lc��Q��z4ʙ4)̀�~�O|�=�ŝ (�L�S�|�xƓCGJ��r1(T����c� !��#edȲ^�X��-�o4kH��K�ܑռ�/��	̯d.��}O�_'�&:�f���I�l��%��t^^O7�:v�Mz�c��uC��j��p�o���N�}�eY�,�J�[���¡X2c��4�q1��0�Қ>/x�3[T�;O�E��C�#^cQB`��]N��g�ɰb8N����J���$Wt�y�j��2B���au.0����h�̓�Y�d����ˡR�����J���5vn��ݸ=��`�Jʌ�=�U5���i+p��'A�Z��<繾�p��7Y�%De��PՄ���1�������f�֌�nБ|ܫ��`G�uF�7��W�!�U���m8s�8,2�cq]άi��!����MɌ� \����bj+>��osD��m�2\둶�F�̙�*L�(��� w�{G��,3��k��r`�	��X:˨8�(��NA��ep	$@p���2��[��0�3�ww��lp��������Ω�n�{��f��2���n�4���
��k�5�z\V��ej?���))�����9T�C!�i	�W����0��rd�?]

��_��OK��v�ft�G3���"�+IN���w֣����r+�V+�B��{��k^�<��G=���Û���7P��J��8��Ǎ�Ҕ��l�;:#Q
Ɯ�2-
!���
.�?}d��a|GѬA�z����GO,w�]r/�D뷬� �P^:�c��o�
`��Z��6�N"�2w�Qv�կ���9+��۶���ڰD��8�n�p��0��N_a�'���̎��ϫ�$_���c������G���9r)|.����g�$��ܺ�9�@�[�N$7%�����
���4�DG�a��]����*�h-�F�H�mg���k�iEY�Oۧ����HV\K��a��\9�hL��w������6wy[)�@Z���	�۶�A��a^<n�9��p˩-�u2�����\�魅K���6����*�B�M���ݵ�/�l�7X��d���g�͜m0X�ɔ����/�}	H�y� ���;~�ӊ���.���g��#u*�������J|K{L�Q�>����=��=�:!G�O��n���7s�TE@��B6���HD����`r�@�}S�^,���	b���N�|.#��D�#>��u��8��v'�G�rLx�d�*t$�y��*l�%��4z��Rj��?��C�s�}�v*ߍi�n��
�T��Lhc�	��-99Cʼ/��w�]��Ֆ��2h*�"u���z�4�|R.�Q�Y�H�4�8�7t}�r&{mR������ൊ�m#��`���0�Է�����Rj��ԕT<@h㏣��]��J!�t��jW�G�����+\9��
u1��,"z���ʞ&�?*���S�
����ϟ�U*ϩ�3�ș��'N�=0ԿqZ�}��؟��G�F��W�|g�V���C�]%?o�+b=E(E2j�O��∆�H��U����6� x|�5���p�]��&=hB��`g��~�����T����j=���������X�lr.����_	���"��C��\Z�(#���K�$UNФ�Xt��B*���tuL����?A�X ��)j@?{�od��=����V���l'��R�X�6/{-�,���+�2��D��l���Oǜ�/�BŹBU�Z��/�cP����4{�$�u�]�$�$j;R2���_�dq_��d��\�������"̓k.�i�&Lm��oF$�a7�`ï��H>���z3�j�I��Я,�<?m���}VJ�O�h�]��;‣>XR���S�
ꕡ�߷[�~z�G���x�iޕ�����םn�s%��B����'�$����Wc\�P@di��M}<���$��lO�fCF�xO-^��{��tnM8�#�qe���u
��[m��E3���m��q�pT�U�5�tc8?�xY���P��'k�I��<���I��v)FW��<�c���Z7&V�lyc��Ɣ<��',��S7�~iUe����9$��'�s� �ΰ��1՗)"�&,]�<'�%2�lڔh��{9��2&2@��/����ͪ�W�d����M��ɷ^ar�*��$8�;�5�曒�}��Ps�"�I���d{Ž��.�����߄��(4[;�6(�����%)GS+2�kz�u�'X(�%���u���Dk<�u�	������ĈW��Y�0��ʤ\�~�e?�0����ضY�k�����z��//���+��v\$Y��O��uz,�g��6u+��ѭ?��[R��&���G�9E����O�זk�#�٦6�u��s�DE���;c�n���)#����[���g�q旞����͌��6�f���&C{^���6 Ñ��l����18ʷs*���v�9sr���ph�fj� �6q�a�õa�h�����>��؇�l��i��ϋ�:�n�<��j�/P"����z޷��ü}]�}�o	�Y���,�����=�@��x<���|���(.�*Z�ZM}�ܗ�~=%� %rW52���M�fSgӣZd׌��
�*e}�03��K���ɣ��㙋�|�gp��*IDw3�H ��Z������?*�|l�Nn��.���{PD�{���5p(�_���1p�ڭ�W�[=΁@�5j������[��
%��>���	j�m��J�Z�9jsj�lOw�~.�S�$���d~���	�ȍ�u�z���#\�`/�5�U�(Z��h���$����ü���^U�c�I�0Z�dksD�/�貝���G��?h����	��p'6����c2�I�N�g���w=�7����-�iӕ-��f���md5��1�i�""tD�<������bWb|s��&s�p����Iȼ=���Wm8��a֭;����ӣ`��ETZ������d��p7��R(�o�ζH��E�]#\�N�d�[4Z��܇�&�ղp��	S��.W��,Qh���:Z��l�ȯf:ϥ�M�6JN���'��}��=5��8Rc����R�A����81�idwy�7K�\*��"�X�޿f
�g�w��RA��N���e������������WMG���ْB��	��S�u��1H����ޗq���,���o�g�
� &Cl8�_d�f�����h�!�t��	��/��u\�K���~��60�W^ާ��%��ߋD��>��(b9{$S{8�H:rI�t��ߛ���?��Q~��+�\
�~,�U��F�C7܉1��P��|E��,�;e5���#pH��R��� ���-��l�oE+�nd�/����Y��@���
#�?�;8�����Qf����kAI�M$
A*��2%&�@x8%��k ��(QG�&�+����o���� ���c��a�D��ad��l۽Jw�U�vK�[���c&�V��Sm~��-gc��e��<��`r�?���@�!�+�E���c�l}�.�	QL�7>j�7k����Sū$���ɕg#�,�����ȄU���$5�f��A��n��f
S��W߀A< F`����܉L�z&V�5a��n�g�n��H��e�h& �8i����Ik��B̗d��zW���ѯ�}���JhvJ��K���ݎT<�>J����o7J^�&,�G�Zn���A�,N,�M�-�}.d�6�A�(�����IqX�e�K-��ڞZ�j=���9��E�{�	�
�����7e��tï3ّ���=�&�W�Agk��ڸ�b(c	k�:������2&=oJg���١���`�YAC�bO���L��M�C��	0����b�Xr��h���_`�G�E��[�>[]q�V����j���V�����������՝}7l�f�K����mh饵��Nً��R�c�p���
6�Z�<�#�lz'�P!�d��Hm����f|�h����N^$�it��O���<U�9�\��.:�������m�n͇"8�9����}�p�(���]��4��7��?u��:��~�V��Z�x%�=��Z���ļ}46���Cx������)�$%��o@�M&�eҒ�5����n�.�Yﻧ(�-1��	���c�vU�!��]��54��^�J�6K�J��!,�@>Q�����(G�@�,�,�Pꐜ�q����~m"	�U-C�d�Ay�k�ܾ��j$�7�R�Ū��B9#�Bfzΰ�N̞�x�D�Ĳ�!B�b(�H�����L^�`�P����h ��SZf�!�[l�)qA���~1��b7�MT����4�̖�)����~MA8)y7����]op���l��^;���|��ʿ�*���eҠ{V���
�����oO8g*wN
Û�"gr���`�9�.� 8�k�YLqx�n�~B����ƻ�$xԔ�B�K�&�O��{������\+֒��꽊TO��H��h���NM*�!̤x"���w3-c�>*f�h�ŵ����K��Ùx#�lo�~��S#����v@����~tM��\�c�#ae xU(n��`�`�%��u��F^r��؏ż�N_����C¸������Jo+n:���6��oLi�\D(u���lcIEA�xڶh��V��9��C���}7����C�\̼�iػ�����X�W(������2D퍦����$74�`�r�r�혏��Z�:�Lm��_*���y z�^�DҲJ�ٿ
O�Ht��S������PĀ��%��/u9�����J��P{-��������!�P�k�����^��|�!^����0��Mpgl�l8 }:;>p��|�,�sc�v���h>�n�z�:��T�C�r7[h�s�q����{�.�zs�1:������[K��K��BC4�l�y΍0�g1�읊́�Yo/��Q�e|�̈́�zDU���΂܏JnZ�Cx�.x&�=2�������|_�濫��}����4��pU"'���R@D]?2b���`�v�q�V��5���l�a=]X�9蘲[�����G�L�\�fR�=Xy2��!��NV=�j���*���\G4���yy7�k�����~z�?�X5�N�j��j6o8�N�:��CB<`ϋ���O����evZJJz���
X�B��6�ey�� � 7Z��zgm���Jd����/^�9���u�75�ٟ7�@���%�)xɭh��m�$b�}��$X�vT{,`s��:@�J����F���C�����_}7g@InQ�PUr���"�+�*r	n@�ݟ��0��5�����0s�108�e�����Q4v���AgO��/�p&
�����+�SL�V4t���!���	�*h�(㝨����$Z�C0U�;..>�7m�'���+��ӯⵦ.'b�GLԹ�T���4}�`�����*�q�zwثf��k��KJ��K��v��O����q��'Z��Y�G^�c=��Cyjl����b,��p����)?�l��lq)OkF?�Ib�L��%�g�-��F{��;(wS�m=����P����lѹ�D�r?���jy�I�����U5�wZL�2ً�/��G@��<��Y�z����j�>����p|[#��s��gcP�}%�����#��"����c2d�/���w�m}}qr��}���Ҳ��؎g҄��$���aD���5*���~'��a��r[|wa|�
����+n�O�X5#�sϗ)�q�)�j���8��u�m��,�3���N�=~��ܩJ	��2%�P��"�4_ql2��/h�Urˤ8pM'��p����ϟ�c+���N%Un+��]��`g��:���*���D�^'��Y�)� [N0H^>aG��k�Imsp��(����S,�N�{*o�� wD��?w�K8_��ij�)�2|����r�).�)u9su�]1�` 
Wt�u���{]L'����W)�o�-F��낾y:3yz�,��g�g����g������仂*,�E|��Ou�ـ�0ν��I>Ԓ��7w�~џߩ���'L)�c�J�y����˸[�]�"j6c޸�P��aޢe�o���21tTG�n
��Xn�J��$GCv�T��8F����9 ���6����u0x�G1����JA���#Ra�MD��8+���B ��|w��E��y�l���xL��MM*X�R�m2�W]:�;G�[[4U,�^���}���R��,lN���[B�]�%$ܙ�>�4܎�U�g�v��V��i�e�:8��2�{�;E[F����>!���g@���c<����l�K+�]C�c��1c�:q� !�������<��aE�˛�6���T�_.m���p����"4u����l�K xh[a6.�J��0�D�Ul<�$�B�T5DvɁfr㱓�ǯ���v�o>U�� ��O��Щ��D��{ЮT�z���i%�;��/&��A�.J~L�1<^ ��'[S���]�08�9�K����_��=������ l}�XAJ������Hq8�??�+]'y�v���f@A��%�I�=��}vM\A~����\o���`��_]˵��yl�}�U�׈\q�U��-��r}�Ϩ�~4�����^6�6�%:%���ۑ��zfE�Z��.J`���c�ncO���~�,��r�I�|Bkh:
2��,~ڞw�*��V ��E �U#�<����T��? ?K�Kk���V��������3���r��o������T-�,�p`��;��X�x�#Ȣ���"Ytf8m&mR7N'�o�{��O|��F�rī���)�!v����o��#�(��=���>6�����h��Y���B���J�;���D�MAfc�
�u�+z��D�RK�k��Ӥ3��9�T�k�3����|���`�ۋ)[�u:K������d^�t�sK��A)�Nq>�C���ryIo�0��)����p����L���b������`U�U��L�n�u���e�x��h\u[�_��w���������W�0���yDҺ���,���S�pR�^(�8���a�FN�eY�1@���S�L�͇E��0����R+7'$���}
�_Q7zg��{�߷�J�t�����$�<>��ߨ |�� J�����x�۩����S�NxY5����g���)��ߞ�C�q�Z}t�Z,Y��[��L/��׉��m(l-�Z-p>У�XN���?���G*7s��K;���yHO�D�}��@�N@ba�M�r�Cda����"����Cյ�l(B�@~�����ܚ?��� �0�R��-�w���B<t��7l [Ɗ��y���������Ujx��#�DT�Ԇ���I�Q��d�I��T}lS�Aꆆ|���c�j@H�J�p"W�D��I��ݲ�����n���B��wy_m��5tB��L?�!.��Kqp��9��X\k�=���i5_su6o(<S���*�e�QŇ@��7n��	J��ηT��Z�&Vb�s����P��j�:�0r����|���lc{����D�6��'�͈m�\o>L�$3u��*Y4�u��$�1ߑ��<�X��*G:�3��	�:�O &\.����`;ÊEoE_�����s�+���0I�	�G��|H��QPDC�
,�r8á�}��`T�q��."�G��0�>[�RT��^��g��f�<�T�E߫���'��q�^#�Sʺ~�v��ju��ׄ�Ml�Q��&2�&��&0�5\�\t�Ax�:9=;�h�{�%o"�R�@�=��A�j��y�ٳx��׏zi4�/Y'h��=��f�y�W��	�b��K��j��2_�ƭ��!�JY���m��4�X�ck��$�����k���NY���7s��rCT�=��l�c�X~�=��h���M� ���\��:}_/曹�D�EU�ݵ�a���$f�a}ѭM��c�(��,I��,�1�<�� ��\q�
��E(V��{�%�tAa�h�ى�B$�5$S&U	��mzOk������Or�ᰡN�/@J	���V���Sqhk�0�;��#�]R�m�g�5Uq�����|���22�&��1놘l ��V�e�;eF�����'����[�h�V�ؔʻr����6�u��J+�F�7(h΍�E	S�c�EЙ��oT�>;Q�(rm�<�R��F��'�b��2*�!m������k�9��9��9���ڤ�x�:��I�9�mH�ݍ%8�^�|TM�f��r�a�t�����ުP}�1�g�Ě�]�ͤUr�r!�=�^@���bb���j�{;�W4~�j"��^��7�m��"q4P����l�C>V���K纬��?�����	~��5�?� X�2p�u��<�d2�K�t$��ɔ�[���Oh�`�pS!���g"�((3F�#;�bZ�m���	�E�&��TQ�J�����o'&�/�f�� �?�~	��w���[��:�EWL1;���:�6ٔQT���Z�m>����,P�f�r�\-Z�-�$��̼��yv��K���byVڴWy�!�#0����J�f�]&$3\��t\ԣx�Z�+�WlW��P�V�3Z�uN��WV��`gΡ�z~����Ep�7���{�N�6;&������~��22����85����=|�����&U��uq�sq�ys�u�v��8�y_������ꠀv�q�GK������R�9�ʍ��v�f���X�@I��82d��6���^����ϧ�Y+)�l.�+{��Q�����ӻ��=;�q��ȿ�{�>$U+npc�N/����~�T�}���]uʌHv�87�?�0��_����g�4�~ǦM���Z��-��G���sa�,\Oc������e�z���i�;�Li��,}���]�glTq�r/�+���dZ�HH1��R�2L~%x����<��͒+�h�?����&�Ռ\>�E�ib�Z#YC(�'�W�{����4� H9�T���QB��^�j6j;��V�oȸ.�$�;���P�}���&�_��mK�z5��t��P0���'�F�	�ݚt_Ď���5��)�	f�W��>�h&	&D6��i�ҧ�d��Ξ�3�i�˳�=w��v�gd�'���j��s7�����q���A_�տ���^F�#`�Y�j�Wq7n�{�&�?�&��MA@E��r�5���D�UsnY�i�[��f6�E_Ům�m�f1����[m��c�׋���[��F�׋j�p"S�H��FU *;H�報I3��+�����B����9��}�o'Z���<��Q����cPCW���_Yqq軨�q����?�����us���Ͼ�AB������&��
L�cV9�3�l�����	&�%�vt��V���^;�r��p5�!T,}P{~@4�9���؎�x����=C}��Q��B�1���bT\M���v�i4V��u�?�4f�ܚ~9�m�š����v
�J�d�x���\E(�-�C�$8N�N�lտz���YM�n���"���Ϋ�Pk���kd��������=�S���sA��P����__i������/ڭ��〣L�6ra���(��9�	Uo�[֭�s��.���܆��z���������8��lv�>(���<��U�F��!v�w;Y�[gX���8��$ʆh9嚎�ɧ�9�;IN'�^t�=����4�.��S��~�c��'�c�����R.vxH����B�ݐ����G��Nz�>Ia*%����j�>ߟ���ʵ�bi���<GӦ�#����(e�}s]O�hd���U,§o��y�B6G�q�}NkI����n"�r���鍁��d�ia�O���;Q�O�c����;/��y(~~�!�,/��yU����M�_�o3�+�.����SC�\���`���!�v8�qj�� �����@?a�W�=UK3(��������i?q����$���g!항g�M��2���;Y=���UWG��C���N_��3���l���K�,��ƺ�Wv���=�F�ͅ�=Qm+[�ۨ��ܔ����!p��.�G:�.���E�|�b%^!c�v�y�4*����R�:׽�ٲ���ﾽ_c�`o-&�|ujJA���t�Ӝ�®E`�qv���V&����i�����9�.qE;Sd�U��Ut�B�[U'��JU�PŹ��%�걹�*�ѩ8�8��H�gp�:�qŅ2�I�U��Rъ&l�G���8�U��&h�R�M`�Y+�t�/7�;���8���:j3���h�U@�A,k��Gڗsu�!o'K>��V���d,v/d��$����gLaML3�ȱ�����Z9'��{(�37�7l��p/�G2��ߐ�ǬSL�J���Fo��;n �Տ���F�<�J�%�>���b%\�s�T�>,��m�8$�6jB/���p���C��S=�&���d_d�x�Fڔ�u�2��kv{����5��v-���Y���Ҧ��O�Rf��ڶ`w�&V-˒�p��`U8�>�>�����?	;�9;�9v�?����V�^k��ZcZc��#b��ck����#��`)4!c~HJ��No^J���n�]Ǖ�y͔9l�9\F.�t>j���
���O'qn��g�F�l����v��s,��Z����A�T��b��AŌ���5���������c�A�+s�/P������O���������B؟�y$Y�x�/+�V��4���̟U�Y0�X���@����	7�7	�А�э�?Ä*��^]�t��	��jP����>^���[�28B>���|4�:�����%T?��.�p�y�)\.�달<�Jѭyz�2�YD}������-�@Ͱ�����ת�go����L��,�5�e��և�y.ΰ�e�d"�1�i�x���y��8��xe����� k��?E�z�$�����C-D�tŧ����Y ��+k�g�w��J-�t�X��N���y,�A�y����N���H.��v�r�+o>[��8 ����������:��ֶK�VRV�6,X�r�SEI��j��2i��]Ч�|��e�ח������S���7;�֗�s��E(���ms�֑�C�d�D �oT�����"
���9՘8���4d�8C8�]��a=R��~6��:p<��m!���rw�гms�:~�B̡��k���Z�]ǻ�\�v���h�?��t��gR���WkUʇ���� 5<&Pf�x�]�H^6C��c�J���'t<|��W�|m[���q (aK�i�C�^��;�\�����J��˪��rSI��g��k:v�eΟ�̵W�P�/7z��l�i�HU��-�� �+�Ғ/�iH�:���Zg*�o?Zc���Y)�Ǖ3�+&O0i���_��]�b��z��(�f�Q?EF��3+�E��k�	'%L�*��Ă���?_��MA�Ank��w�+W>r�5����|��]�	��}HG�5Ǖp�[�!�V����Z	��c)#�mRI�LmӋ�P�J�؜��c�L��\�Y�3��d+��"k�9���ܙ�50"~h'�~�$1�X$vn�ח��$��
��'�ޙ�Hh�X��_�t�����D�x��:�U=��fdx�}���`q�?���R���⓸�@F3s�^S��Җ^y��p�4;''���oz�����d�<x�ĽuZ�	�nd���_���&�&F現X����*j��"�R�#�l��+�����m�����1�=r��Gfxmu���Q/lK	.'BS��z�$QUF#��KA��4��X(���GL�'y�pc\�?��.��f�	s+D������v���1��� �yS�fS�aW�f[?�qӣQ(�;Õ�㈹�4��s�8s��!�F�� �r�9X12��{��!FU:8	.Y�#� ��Lj������H�����Rʳ����1��4���;�o�����t0$��g W��e|��4j*x�y�i�'N���'1�������">(�B���"~�
~�B��e-Ja}"���HT3&)&%Ct���
�/i����OӲ��Ie2�	�}"I�\���it�)^�t��h�� �4p�N�W��c:�G�O��f�*�R
ưQ����,�Y�cz��$VR���+"dl��0��cG�\;�������٠%+��"Z^����}��H(�}K���X3����T������M+���G&���������mm}h*ޟ��+ϣ�d�I��n����������'hHC�py�ɸ�w�P�s��N�o���0LS<�eU�d�A��74��ŷc�+yc�?\�(!�o:6@I�3��3\=n��kG��bYԅ�hܭ!{�'��#/	R��(�m�j��_��,L�<�P�],���jS4�eg�/�S�1%
��Ҁ�i��,��l�#i�!�3_v>'��K���.ڱ�z6[3��JVb��֌�z�$% l��������j2W߉��UElX}p�Ɔ���~�hW.����{T�N��u��ȯ� �2�����68Φ����}	�&�on�՘69�Ztq��Y�r�*[��(#g>��PGn�g�OF WIN��˷�U���~��h7�[��P$8�I~D�_d��^)j�p5�{�U�ѿ��u����8���)����:����if�h�h��q��alwŉ���м�p�H�MCfR;bB�b�� a���9d�.9�)�y�����,>�N�k� x6�����{| ��;);I��It�'M�ݿb=m�}�C��qT���N��u+��pa�r{~V���!tm���e����f�"���Ϡc�|n��w��1^,vk{{��|�,Y��c����Fʋ~ҁ��w5��Y:��î��E?ΞH��@5�$<T���0��W=��7�vFc��'?U��d������CB�w�����x�=�Q�3y�h��柿ki8���W��^�f�<��2ݔ�*3uښR _�Ǟo	�D}Mfa�1&	'N�S���
t=�X�S��	?��c�q�;�M�2̭���\�tj宯��o<]��r/��\/�NɣKΩfF������߰��m�n�ө�b�����?�̸d� ���������x�dǪ0m<��,Vj�3V�w�Ӝ �r�Z��,|Rw'��H�ɥ�t�wm�J3i��5����*廟b"�o�s_�p�oGN���d��$�S���?�d�q1T��c��P�G�Ա�\M��(���Z����e�Q�h34)e����n$B��!
������`��/�ʵ�44�,ҭY>_ly~X`u��/�La�>���[���&|��<�&<�K�RR�_��;IH� �� ��9���c�~�Ϗcc���k�3�_�߻s	��vG���Ezw�:N�s޼!?�a�aFg�[wl�SGe�+��Dp�΍c '��ז��΍c �u�=�J-�aIu��q+�	ﯼ��̣脨&M��Br"��z�|��~�t���ޝm4��&� Yh�܃��9�j���Ɵ�Y˖��}��S����G��d��'8*�or���c��V�9[�)N	Y����͂N����O��F/2p�ߩ�U	�4�.�rRNFz�ȴ��|G�k;�q#�oN�M�2U쫑2��r
�H^��F��Ib�������h��?'`L�0���AA�n,)b�
���u��_�����,�)��*�b���	���槐�򋘨F{P1�y^
�F�C����tr��"��dڱ���'?~E^�*QVѐ,����pp)��Q&|�H*(��dЙ@4��
z#��0(O3��S�U�����^F���c_��h�?���9�/3�g�[��ps�	�Q&����.�y������_�7~Gv|���$&��|8]膯��(�=���5��HX�A�g�%�ƒ�5W��!��EEl�":d|j�`��e���
������A£�1��,�u�K�T�(���E�	Q�j�r��oD�[S�B��Y�.�GN����&�����Ml��/�2��?�%"���~��ړ}p��%��7"a��Z����1�J:P��0&4�:
�։��2�Ƭ7H�c+T����E�]r���\b� ]7�V'��ד�n>����(z~&O�t����O��U�"N�y�ix����� K��l������hɢ��'}�ODA�c�N�kx����<-�N~�#�P���G��|W��G�=�H����'|�P�|Sb���k��'�F����p��;��V�Ǒ���	��
��V�{���������Q\�ũ�O�$O��>�'�H4#��[Ay'��p�M�?RB�/���a�)q0�O�(��v7���#{�����=;u��pv�B���)�wk���A�k;ۄ��jm��ڂ�!$��"����Zϥ[��3�,�o����<[Vl��A<Jν���..?�hX�p������Z<yAk~�t��״ֹOӭv�7	��/靯WA��w;\Dj�՜z���u����l����J��
��D�oee&�q(���Ʈ^�ٟ:�s7���=ͭ�r����
��FH#��	ZA��L�
��O��6�Z�'Q�F���8s��Mһ�A�i+���kZ����"���%�]��띰�����IR�$p׵��&��{\�`+��|hW�$��gĻf���1Q�]���l4)z�/�;.�p �s�ka��Z�c�y"{��eif��5�LȮCT�A�\��t��U�I���ɯ���I����~����ދ��y�Y��3���Z��$xL*E�;�s<+EKM�����(Y8�S�cU���,���4�O������C'脧�Tw�y��3e��t���XY�W7���������p�ra[mS2M��6�6,������V�6���$f�Y��a
��Ͷ�.ñ�r�_�O�A�B��A�^��(���q)o.��H��H��$<��_�n�;��B1"�F`�Ko�Рl#Ϣpʳ��n��Д\�.�P߾�M1o��\��tcb�Wի��\M���&�=���M: �&Ӌ�<x��rљgSD�uR��?�5K��	�fs����?�.x�Ix������\�8ǔy�c\��襞��I?i9�9sJ�tֺpѼpջr��@PҸq�<w	9)�^G���Q?x��e.�` J��F����^�ou�F��}Zx�}�"j� ����Hc�!��_V��)�s�,9|�h�&?�6
����-��Z�9��4:�t���S���AYp�ܮ�\�y4�1�k�b�h��'�h��֏���r�|e��:s��n�&�.�N��</Z��\���5S?I����$�Y�b	�$����A[�&@�*���/o��%�aN��H �W�X7�Y�آB��������*�y�z��c���_7��}_T�H�'�t:4	oh��Ce���[H��o��ټ�0Qͺt�-G��7��AD��K���;���E�^!2O=4"�F�Jq꿦�46p��P헆\ �:��t,�?ǝ�L�R"�P�_�!���g�*/S
7��S�֧�Փ#���4����V-��]���J�����3 ��ϯ���6$!�N��jC!�f�']���	�>�.wj���_�Q�/��W-�XRx^�"E�ְ���Ȱ;�;añ�\�J�/dY���$�Xt|6m ����8y��	z�P��g**΁������Կ�
����P2��ٗfDA�Bm��q�\D�LU�{?�a�^�lP��e��7�$��������J�*��a[y_xz�V(�5w,#��y�6�7g�(Ӽ/�ӲE8.
7S\��,�D5ۦS����n��f�E��Y@?���J���P���(a��؅�$�| �>����(��HO�v�)5麅ڷ�9�aͩ��.##y�B��l���G�P�+<3��(�;��m+�S���6�{R!,@K���1׹O	lH?nKʇ?(F�w�,��x��T���uZn�7\w���k�Ҭ}C��f���^=D1����8?u&�ޣ����OV���2����+v������r��6���2���rv�����,5�- �ȣ�(�Y#�^c� h�"ڨ��P�_��W�Ӗ�Vr����P�/�j�R�Y�a��^��P(��l�n6Pxћ��(E�D>��FC��|3VPv!T~M�*(�
_��'������YIr ~���l���tlq%Re�����{Z��r���ʡ�}ń�Y��uK����u�?�P�l�eh��X�i�Mt��/Y/m�r<�V��a�j\3��*!�U�zewu�Z�����rOJK޾vo�QtB���vi
���(�ܡ���W*�d��X%1��ɴ��Ϩ��.�B�e�תu������c��ex&�}%��L7���M!�XL�����O�<�=H"�A�.��M?�402GӇ"�X�e���	��E�U�1�Z�=��z������,>������wb ��z�v%u-ڊ6�"�hQ䯧n����(_~�����-�/q�Rn���Ưn�y�~�b�$td�x�C�@��ǁ��a��[/�+��0� ��ׯ�� 	֢�e�|V�ܥ�7[Z����1����Ǧ�����$��t
2��)+$Pw�|�<���.�u�=��F�Tľ�FbX�Rn/�*��5�ܟ���'ȼ�
�L���:@�j8=�ҿ�H�u�vB����lisj��Sc2mH���or4X� aQ�^��`����t�{'�Xb�.dl��z�hޔj���3��3[
�v�t��8>�0�nk�^�}89R�-i�]�z�OG�d�}-��@Sd'��`E��8!@��},�=�M���LJ���|�s���?\�eT[��w��8šX�;��E)P�H�b�]�K��PB�K��;����.��~x�{�8���1���}�oε��u�N����_����9d	�n��@2�9�k���,����fE]$��)z�٨�V�w��tg�F����f���I\��R�X;� �`�R�Ex��� ���.!c��HK�,xd������~h��'�Rv|s@���&��l�ޫ�)�O��Ս���cצ��U}�X2�F�'�|�7��}�S:z��#c	�[���.��X�εvi��'��G���#���Ƙ�nC«���Ƨ�.�'�D�۳F��9C����Ov�B��t�t�^���ǲO���^.M�-z�З��|���m��?
�5�3�ā�J�߃cG���mk��W��)\�M��?�@�s*��[K�SZ���KkKV\�-��)hyK�x���dƌ>�F��(�
�r�I��n�1��k�/-�r�&��f~V��Հ3�
~v���{v�v��N���>H�0����.ʕc�h�_"CC�ə��>c�+�� ��~󵽱+4��{(���f�oP�f�"���A���"��lB�����˷
�;y��}vV��2��������~�g������g;�)�q;��2`ʧ�v�|fJ��7n|w-��cr���6�ؿ=yɬr&�� AN=U ���g�0�!��V]�zj��<����<�#SF�����>*|�wľ[�)/��&m+� �	)�+����Ω�9/�97g�6󯖖�@�-W;�GO��W~W;l����z�k���7K�hg�G�3�V.�C�Q��Y�W�q�!���� ��ߣ�{��|��`���ǒ.�u����ѸT�`����|�<E�e�v;vu�G��%k���T �Fo������0��Y=F�/ob�QJkJ$m�=�,2·`���o����c����~�L�-m7�d���%%o�56�&o�^"�^O6@ɝPP���+�jƬ�%HJ�PH��w��M����f��T���B.��6	�/����}E�v%�:�����&���:J}�����t\l�۬	��27�1B`v��*�ʥ	�.o�u'�����qb��h�3؉^��}@"���$���1� >L���9�Ҝ�$ߺw(<Y�k���:��R��R`�9&<#j�Yj*����z(�%��\�P[��������_�\\>�[X�̴CeG��|�g� P%�;E<�&W	:�yG��\WÂBs]�����~dۑf�lga��A�M�VK
QV�?�$��ɤ�L�{�[���u��+?z4�s6�;E��z��y���2E@`�?��;%m����۩�R��HE���^��	�z08���twu^�K��&�z�d��d�~3�E##���'^�n5��S*J�(g��E�����A ��x��=ԥ�i�4 �m�Èu,��Zd��y�-��C�s�
?��*8��l�a���������K��#j�[����T��Ԑ����.�B��t��'�-z}{3�4��yv�Oz#Zz9�x-�#�\L*��\r�=�|0��P\�?��.�����;øQ�Y��ӎ����@�����DV���T���?o��{�Xu�;f7
z��Q[Q�d{��,=d�?��w\�M�j��١ �Y& nߴ�J�z��\�g��!H�-�
{`n����UmŘ��
�����<�|���D)U��?��<���=��]�ѴN/���n�y��5d����G�H��;H��m�-;yۇa��8,�]�dK\Sb������܀WZ���Fp�o�d��V]�*%[~�:�:���o�	mԺ73}�T���������O��q!fa\�3H]�j�_T"�(dhb`e`��:<��W�ݭ����H�[��V�L���(V�����Z	/x��s��۔?��X@B#�
�)1��Cg,jܓ��s�p�<��Z��~&S?A~�$�!sW/K�O�}�c�RU\ڔ��Nh�M��[�����׫'��	�3K8S��AnjF ����tI5׌��T�⯊��VNd������j�x�����}5C�w�E`mX�3sn�}���lnN ��Vg��a���H�۫&W��jC�'��x�Ҟޛ�ji��޷����nR:����S?���fH��b�H���AW�YK�����}����4����E���\I�C[l��*8���!���2�)�
p~�cD<N
�S�i�g�b�����C�A�k%u;I�e+�s��ׄ���^�S
˔��5O?}����*���-AԖ����y��AGH4Ϫ��o����a�����2�~�����/˥:6J#���J�:߈�%��6�5n

|4�@�N��:�LLI�*(��23�)�r�����|v��+��m/�r�^ә�]^׫+.�ؗ�'*�Ƽ�* ���RC��ڂ��A�x쒷�u�� D憛�x+���o�ÐV��1naQ"�Kųʡ�[����:YR�̟˟��F�V֣�>n�����g�����[?�B:a
��g�|�xE�ٳ�O�JƄ����x"���'�$��Z׋�&��oz�ł���W�_�8�5�E�|�T ��aq�" ��Z"|u	������`�|U��H-,�
�$��꽁U��t�rb�����w��*�7���2R�:�A���4@_NR0ꕨ�eʥ�׾�	�~1Í����Yː+Z`�*�f&=.�\�ː2O���%Ŀ�y7Ԇ�����k������� ѳ1� l[��Z�9�(�Ek��
;Brrֈ_�!]U�Kd�5фx�\��4���"R{�+Ҡ��\���Z{��<|�3����^y�'���Nؙ���yWI\F�rтy�@�5|��g�{k>Ҵ/o߻M7�Is�2�̴�������7��8W����42�z���N�!61��=��<�÷4?���_�m��u��{=��$�c�4�୤����oY̲�V��J�{W�=-��l��X~����hF�W���Z��E�̑��:d[4	�./�%'����{�!loi�q3�C1+BIl�,@��D�>X�A��Ky����u���5�%f����W�f������7<�B�GK��6���Q���C� �ܫ�>��w�?��ֵ�K���۠�[�{#c'Hv�;5Cgz��:�/�጖ふ���O��.�� 0�M����6U`������o&V��n4*t�� n�3L`�rklN�ux��MJ�&d�T���P�轃Rm���9�{�Қ�w���9J�T�c��T�$݇nZ�hZ|�;�ĳ��:gۧ;�6HV��\�`P�.��_�8�8K�"hb%�G�y��x��=F����_-l�y߭?/B�7���HɦC��f�HɆe���p�7���kt��N�{m����y���[]������Ixʄ���N� g0� b����Ǝ��tl�gu�������)����)��
��q�%��C8f��ƚfP2��qMb9=g�����9���8�~�ǡ�dǿk�K^I�$䉰���L�ָ��w
SoG�8N�&�Rc]���[]g�]��9���w�
��Γ�x5
��rm뀪S�Q�Ta�i�XvxB����� c� `'��C�m;V�9��+��$Z�0��>HnZǲG;�Rla�?@��7�\OZ��0o�O��U�-w��Z���Kk��?����O�}d&�/����Gd�f\,!7TMѐ�J�N����M:�N\���|��eO.�j���������|�Q��ӧ�T`��h�s��j��/�t��=[��$��:�2�:�~��?�M}�zò���9n��n�O.^�]�����h��4�k���'(�'�-��^�^�F��=���.Y��b�;�)$&K�A��0H���z;�ė�V�{k��]�#�nq�+#0mfY����jS����(	`v`���!�܇�[�z�пm��0ݷ�Aso��;5���4�S"����v��~}j��'�do�c	��m�8}���Q�|Q�	��F{?�p�~4���x[�\�gï��o�_�^v4>�"~�"�G���޶e��!��I���ɍ	��i��33�v|��L��pRm��tA�c����o�+^��$�ƚ�)�w��O2e:YO��M��4�� ����ʢ6�G���u���<O�=�н<ݎ��s���9�JB[��A@i��,'�'[�/��i-��-6I����c�S��Qze��`FN" �d�hg������LF%r<]�i����D5�#xY����F4Z'j�����r��#6����u\6������	D�����`I�.��S}6"�+�5Iҽa|��Г߽�q�����y��F�l�~�:'�{�N#�X2�{�i��>fDD�DLy��|��u���ə.�|b�>�U�p꣤�D�q���OM�6e&�/�v:x�O���j�\M6U��=Rz�ȏ!ErdK��TR9��0��������D��ړ����Xj!�F����.������J�e]Ol�B�ʻ���Y��OL�J����7���Um�a�Aw\��'�]�M"�jW,P����1V�^R�/�鵌Pg	; q+����<N۞5�ֵ8�C�fׯ�+|(�3Yl��1�:��S��1�6��n�Y�:S�zrF�������`�ZxӉ¡����0��ؙ%�D���AO�.�%ل:�`��A=iɠ"����)�][H8�iL
e}�L����)�VRZF�&*� u��7Vt�h�6.rG'̬7S5���������2�������	�-//LII����"�1N"�؁�|��ml��ƀ�FBUē��X±��q�go&�����	ٕ�]ע����߽�G'�+��)kǸ*�1�
��9��q��)��Kt�s@;;���8s�w� ��͙�,���}�!m�}�7�Ƅ���:�?=�DR��S��K���g����4J:u`/W�F���òK��*{)w�Qv����ERX�pυŷh��4x���Ӈ�dh�j�M�ʗˉ��k'��:�*):�Θ,�α�����h�o3�-_W�߱@��%�=�$�H��؛]o+���=��m�����D�'x�5%x���@YˠJH�j�|H{+���Hd��k��&Yi�C��׬��³dk�YB����0���-<0�w�����,2K�4�A�s͠�}�+*B`�.��y��<)��R`�8�e��:��^��e�ee��� �4�'9�#�o���W�s�4���id�﷯��R�a�����r���p57����D_����{;<�t��{{�|7��C���i-�8^#�����4^�fuשϞ�����Sx`�4�+cJ�:v�,/0���6.���"Q�=r	�:���+1�d�A����b~��S3K�S���(�3G�r �:4L]�.+�����D%��>-���,BL��|.(����s�]���%c�i�b��P-�86��7�Cf�ԥaµ,��2�tb��Y]��N֣䗘엗��Q�/���O޴�L�:�\�C���h�������!8W_a��|�;Ec� ��X��p�v�E��G� ���x��p^�Ťc^ ��j*�`*�z����9l���S�Lvk\�ҋ�{ת��ԱD� ��g��������ck�W\�_� ^��}�mP���G.����=� ��tQ"L���/}��>��_�(�G�i��B��W6�Ml��{��;�ѼB0�D��� w�%s�l�����th����?7�F���g��s,��\GƟ��;�9���.ly�x0PP���jwd��6�����.3���UR踱>ͨV����1m�'�Я{z,=�Nu���U���{������������*��)�����������-�9�?n�w�ѓʱ1�ƭS�|^�\Kw^�����^{��y��/���O<�裸�~�Y�9���3\H0�KsPJ�U�ؼ���ěZ�D[& 7Q��nʋ�.N�*�(Q��%�>�������z��!��>a���c�7��ۥ��Z��Z���%b'�Pp+��כ;k,��L!�4� ��O��ݽ�=׿�&�{K|_��}蚉�N>��I�����Q�gQ�'��/�t�
�
W�8.�ms�w�N�K7gd��"�Ī ��c��,T��t��,��k�g���L�0>��[J�j�ե�ai�Z�����;E��L|�����M�]��QUHW:OO�%V�ݗ�ɮ2]�G�7�S"�S��S***RRR������IKK������k�����IHH,,H,6e4�J�fH���g;������݉4zh�;����>}���.���0ß�֛�J��"���_�'O� ���tU���+0��P�sEnR��Y�b_v�g6��iPV��2��8�N�z���z����������!<�H���fQ4 �Y5C(��R
����vp��a�\R����+��)�v&��n`B����g�ް���_����y�����nf�H6 �g�&:��O�
���*�q��>�-=�b<cf%�'���!pQh�̙l4���o�8�E�C44C���a�=l�N'���He�G�*��E��C	��+���Q�01vn���(���~�3]�ݩ*�Ϙ�Bw�L�*)=˾�>�m�g�VNX�F��z�5��<?�	�rL�� }옪��}%�g��֍ܿ�f���Ŀ3I�h`��9`�R�����P�y1O�r�xR�H҆�Fz�������|[n�4�-KȲ� �"t���?����|k�<�CS�~�#�u}փ\���.y��b�
�]Nd��/?^�,{��ӷzn�Fo��θ�׾�o�.�'L��)��jAP��A�c�P�E�T����Xx �j_�&�r�ȅ$���r�|�|�F"�ޭ�+#6emg�L	a�כz6n/Z��;�K7q��u�wԁ�ܱe�A�5�f5��e���[�,��.
��/�����#��Ve��X�JG&�)����k�����_�fz)0�U�W����x���ǭ�Azpַ�T���!��PЋ���'a��۲��H�b���}��GRI@�(���6��8 ^{����:jyqO�$Y�_�@�޾ANZ�9�ej�B��L���fQ-n�/�/�U�չ@,�N�L�.�A���@�V![g9w����Ư�|�c>�H�l\z1\ϫ��>k��以�X��uF���[L���V̢�ɡ�mk륦٨A����h�T$Ꙋ�q.˶U	�B���$Y����FL�.���k?Fbɉro�h���,Z|%��ֱ�DH �
زE�@!W�(��0�|M�8H�T@~������/��H���
q3ꃱ�Cw
r������C��~T^���(X*_Q��u<m�B�ZnN'��<��ɺ7v�)t�� ���}�t��T�r�){	rxq��~�t�}b�Ӭ����{�81�g~j�y�&F��	3��Ey���f�{��8�L�G��� M��uy�3�x��v�F=tj�l8�i�����_%/��e��'�89٦�kt$Nى�ٟ��$�?5��6��������9�z�'u��F9��]��C������C�IQZ6��s�J7 
�ۀٵ�f^$��#��=_��C�c���/�ՃN,՝.赩t�����%�����z�L,ny�.�F�K����l6�_-'U�~���q�0h�������%��/�-:�IS��;=ʔ�r�c����P\�J�E0��\�,�Cj�Z�9HШ( ���POH"Ԧ��X9 bd�dw񈦦4�j\�j�����T���2-�*ѝ���~����aB���_AR��?�/m�	�5?������1v"���S/��e�!i`����L���f��?(b��A��V��.�����7��׍^7����f|rbղ�Y����	�4Ck������#���������,�K��,��fh�X��~�Σy=���O�n��o&$�O{�iko��!�Ѭ�v]��4����#Ɩ3����X�D�CoE�3��E�d���O$���>��h
���6��s��f�t���ylɻ��N�����x����Q�������"��_�s�L�DT�rtl�}Ĉ����F��Mh��vAK��fQor��r�4�ND�S8U>*`f���V!�\/�a�K�a���I���>��D!{�Z����|���P�c(T@��g:k��q��1�����˙è��X�W��r8c�Ѓ�o&֌%��6���9O��t�t|��lKBF��G�n�1X�P��<C� �h��'�(����Xe�
qb//�X� S�>��S�v�MV�f{���c�g��E#�k�4�?�mJ�Y[����
0 ��꘨QxA.���N�������G������S�A�D�e�˶��|�?�;5-	6��G(/b�G͠%���JX}��]�$~�6Wp_E$'�qf��q�A����[�T~0V�tv�t�����`z�`d����SC��?xo�PI2	#F���{�;��}:[�򻨎}��ʾ?�y��t���n78^/d�60�G���k�F]ǩ}@��N	�SE*Tp9Q�ai�0�L�9�u��_�̵aud�>	u �W�:�[����kr$��b��n �����zˊ�ڟ|��כ��^�&z�@�_�Ęm��^Y,ً��K��&��1�Z�˒��>&�+8#OM��7���Hwj���X9������a0�q�A�y�\(�UD9Cw��.��b�@6�"��ϕ�ȼrE��,v:Л�y�4^�ah�JB�m���7���2���`��'�7Kv�Ra�sZҲ���|{�܁A�^�L&(��G���B��Ǡ��!�|�������$oʕV�_pb)i忘��|Ъ1����;��ҕ@�&�KS+�=0F
^0Q�ޮ��b�il�X��0Ǖ���n���T
^T�Mƣ�5��%+��@��U�*��n���f�$�?ɫM�*�1�E�i�YF�O�9�E�)r�/����ZR��=�QX�ǣF �}�u�X�1b�M��lBq~��F�6���-�L+�-�d}�<,�k�9N^;J���.��'���^�J1�,.��؁��VV3��s�4��;�@Ëπ�G�}*yt��GM���a�E�v���Kl*�vT��N�9&��R�Z���n(6{R�uY7ڒhS}3���޴���$,���H��T���^�i�Q�$wR��~)��Ո���=��f�EN՟����4Y3������;�7S8��z�=�)GZ~&�5J�f���@![�Df��Tw���}SF=F�j���"X�A9�P�L������]����F�Ҿ5�RK5��!���ڼ`dh�a�����{�����X=;x�QꈥlE��hZr�/X4}Rz�=Iu�-�h�x�K�$� ��@\�[��Z���u�r��9}�z}���3Q�(����Ε@˒Dӟ,{�Z��p�R��D1EC��_[�[\&�ɹ9�u�F��U��f�w#���<�#�L@��O����Z5��M��G�h))P"_G/UD��R����*�;o�̓Ld+,���"���D7m�U9�}٬����8l��V�{:��e[_zW���e��e*�%��L�`_���������Oagb���ט��W�:|B��ocmz��В��d�����)�O-�<&>6�Y=*���Ɛ�v����w5��Y�)�$���w��B��l8id��w2�����4�`ܦQ��;��\ Dq%9��G�֦�,
�t���.�I+x=�a~c+Z>��mN����r-(b��E��"�}�C���*7����%�����gU��A��A�DF��m&�0���%����K�A�pº��-���P@��.�ge�pc�`@����#,̦(\�s��N��h���B�[�'#�BuGpq�����S��F*Uf�񊩽����.��?��m�3��o�I� �(���7�R�sH�0��e*|}BF�Z2�����;J�w�����"8'���I�+F��uX��{�9�OεV�2��{�.a�<ސD���~�(����q���	Y`ʩ�5�)' a+c�����fԿ�x���0G������#�%�L*n2�9a�k�?���T\��0-�����=@�,��,�\4�����AͩqE�{E]&WPq*��~$��\�w�y#>7:��fs;���J�g��D�z��E��NkL��"sG��Q�
Q�y=r�r���>\K����9g��[��%�%��C�մ������Z]M����*�½�eџ�m���}ѯ��K��Md�0q����Wr3"�Kuh|����T1A���Z \��b��y�A�s�Hln˲��L�g��S@�!�q3�w)Y�,���#!���(~d�÷Zr��4
�� 
d����C���6����� {�!;z�vj��p�Eo= �p5�w���qî=�.�q��Fcӂ!϶�Y�+o�3_��L�_-`������w/v�|i�fa�R^Gg>;/��7&?/	� �L�R7jmᇿ0ο�Z�ZD���]�Y��٢�Y��ك~m*���^�nz�D\i���X�7��ͱd�怍��q"�i7�m��A\�niF{1�~���q�9�ǥ�L  ^O�:��� 32G�>iV�����X���jf���=��)y��x��t��L���M0�	����s����V������ۈW]�P�Z�M� D�q�Sq��e�B�r��䯪����S	;�3�n}��-�J����3��s�1x�d�MH4��Xہ��[�qU��C���ҫ^�W1:a.�֜dݕ�����¼Q�4<%�q�W�f��QM�ʙ�1���b�䩸�З�u,�<�1){l�����2��G��Á9��pN2>=�`h��V�!�f�#�,X�G�s��	}L�W.("O;0dT��G>L^�+ԫE͈~v��[�b��t���Ŭ�i
꾒?ˊ+	8p�S/5c@���^�#0}�85��<L���A �����"�T����f��X
|��]���x<=ݵ�?pB��?C�?��@��rWvoa1oaq�{�yL��P���T����E/�F�Y�|�ѭ)o�>���;8(��q �� ��T!����cg�'���b<�FR;��G�ʭI���-_*�|���]2F�۪���9��x.�����O�V�)d��"&_���n�@��ѽ�YE��i7=+��O�F��~~��ˢ����-��H��T�7���O`�❅i��	�NJa�8��t�Y��m}9��$��$u9`���s+6����+�<��%�j����h�\kj7mƽ�c[�]|r4ʮ�/KWeӡQ-�)󬷿���N�86ʿ)���Aw�G9���ly�b����Qf�n$��j&�Dc|	X<C8/!�n~r�|MZ7�|
Lt~�7�6oo{]1x�������1[t�f�5��_=�M���]������d���'�����,�Q�@�B���Gw��ߝA/��ni_x>���?��O��m���P)��)2��~�P��V�Y�U�&+1YP�+*��4h��wn��:%r�t�4鐒A79]����a���=�G�W!1�l:6������)ś�����-'���0��g���r�L�B"�6�eOE��5K�Gz�����V55Seѵ��]�%V!���_őc���e����+��
�����f��Q�1E�ݏg|�h�.��Uw-��h��`�a^'04�;
���L�����U�i�h�5��ˬWu��:��N�rP)D�����اRfKtVN���i|^����n�S�����o���/��K/Xx/^egqz�ڵ2�.�K/��C���T4A�E�N�0{`�*_~q�%G`�)LrTA�<̴�s�+���?�\Tl�;y�{��Е>`P�g�X��ږ�zA�9pjn�}����KJ��V���2�h<K�m����ʌ�Ϻ�ٹ�wv��Ԉ!~���L1F@G��T����sކ��)��+:��$�1�͠�z'l����Y��SȦ4��t�naY����6)��4	@��.:H���O碭�M�1�О��/Kc�;:�D'q]�O\	Z��tf��ZA)��u��TYlqYA�l�U����6Un��G��*�#Z�5��<��֘0ƒ C|Lo�D�5S���u<D�S�r��T�v�!�������?w7�X���SK�L�!h��$�1�� ��8�6e�Ћ���Ǚ���\����A��Ug��f��>��'��4��zwY�2A�L������v��i=iə�S�����ӇG�����o���VO�� ����5n1#(��G���4��^^��N]�x��}����|�x�Z�46�lvD���C�5�]+Qd`�%,a�RgBʈ�wC@V'���
�9[�u��6�A�D�P��(���w"s��������Q�"��}�2�<�b,U�06	~-#y�y=���&z[���5�/e��	Jw�q܏�-m�1�C�,�/�8;T�͏�{�i��䯡�NSɅ����E�.��9����?H`�RR�l6a�UA�K�H�2@�d��q�y#ʘq�`��$��F:g鏵dL�`���Ӡ�A��]�4�����������m��)#鹍���D��zaթs���w���=޹U�yt�R���U<����^�զ�A�}�R�i׆��-(�yp��- �J}��q�!s�j}�9&�&��Ƶ������-�����&ڂ��V?����$��߶�����N[��?�cƶ� �ߠ�ѹ�TJ(�� ���Bm!�� ��P=�}Л��hL���*�\*�6<�{BS�N[�f�F��Y!v�砕��W4����R=�B�y�3��GK��3hl���\�ҠeS2h6�$#;��o�;Se�8��u� ����y��n�l��3�\�oO�j�
�~+K��#r���L�[��򵥓�&�Z��<m��� <���Ժ���v�j(�|*�~���,jw��!�]~��O�ɧ��:��rK�S�h���n���TQ�>>��D�5����:��ғ7*��6��~�op�A�e�V���S�*�H�<e�)*������i~����O������D JU�, 
}	&���N���R��Ms�^��Ϛ��5�Y\j�ʾ��k� =M�n���b��`�G�ث���-4�����]�zII�Z�(٩���Zq3����H���o��М��5�y]{#x�7�q�����"�:c�X�kDa�+�݉G�EѪz���3H��S�
vJ�SlH�U�Trv���+��+�(��k���5_�4^J��)/t���7ChDw����N�wsҩ���?�.}qQs����M�N)��X�>�<{�C�E�^�X-f��i��vv�mO�H���u�ޣ��𻖝5O�U�`LV��2���Н���.]���=���=��K�9��ބ>d�(�KP~�� ���l�p���
#�fL
� vLRѥο�QU����r� ��	U
��%+�X��S漏�"I�\���D�
�p�E<V�2F��޾�n����bQ�$�d�IKF�6��7�䕮6Mfi)��ī�iaM�C�`����gn%�`��i���T��I0t
����ZOuU?�V��,�U�|#�2;W�m�o��,&��}����?�����]^�/��st��������F�Ȫ�S���C\������վ��r�r����GBз����:R����cƵ-@�ӷ�h��Wrbag��s�3,�ᲅ���˶��]uK����߉�m�O�Q�0���;���w��?C�=˷K62T�$Nq�{�e��9:�,��|Z�_kh�̢���K�ѫT�v �L!R�ku�T`�=Y����Q�����Xᷧ���2����ٍvD1����L�:�Lڢ�02r�=K�;�ꨎ|7��Y���6�
B��B�袒N�b�y�}B���Q�y���OPf}m�����cT�6��Ѝg��X���J���X���۬��7������n��hЏ@7<�o�
��+��ȟ<'d�PSH����DH�N-r�>�d���̨��0���������TH������e��~�p�Ij�>��bA$��"��O�9�����)b�&Wg�
���Aq�iB�X8�E#H���a�R�߁�yw
���>S�4H$�)tH�dR���*�0K�nzn��֫�Lz���?)����xr��*;�����Z�7�V�ÕHoA��jKE}��ĭ]�0����V��ma6����@g�_s�|���?��
l���@(�m:`w=wm���Р���K��P�ه��/���T�pҀ�L\�%�G��`R2���lz�0�J`���\�h2��t���&�ൂ�1��w�4y�>��T�ݔ� �@��r+Ě�;*��,U �zt��Gw�o�B��IځCP%T�q�ϊ➓������K2I�ֳ��l��+�/��ҳ �e���y�N�#]��	���u����m��5���O�ǎla�_�~%>E~����~��*`��XAQ�T*OE���r'\��[r�#,j/���ǅ�ǧ뚶�вrn�����e��M�]gQ��U �ֵhT���m�l�_��x߇*�1;�W	R���S���[�Q��d쎪>cqw���v��;��i6:�@�F���
�\n/Z})��Q���8����Gs��Noy�[Z̢�&r+N���EC8�|ݸ}�dU�9MN�
VFh������Q2]'��{�1~�V������DxB���V�Z�a��MI���YR2ZR�C�n�V�!�$�6u|dn0V9'���D`¥BRMbs��2z��tl^e��fU��'��N3�D$1�d���y}�G�ߢ_��Qe9v�Jw�xX�k�:,*o�C���� �k���Ն��.����'{#a���r�T���-�u�b��t�pI��6*�����V�ݽ�s�k�i�� ��X���n�/?	�6��Q�h�L�*��D���Ld��S#U:��X����|�̾1=%�@``w�G��\Q����[�O�)Ftufm�Y��ɾj	ա�������j|�7�"[gv7xz*6~������g���CnF��l^>�L<X��'� �Z�{8�)�X��(�� 7�si���*��lRb�r�,��D�
�7G���z�+��9��@�{{5I� L����ySlz{_H;w��*�n��sK���o��鰶��(���;(�(���䩼M�2`���A~�����<�!�h�������l(F������g���E��I�ns��_���$����{�A�:�	nk
�!�%:N�t�n^*h�/|ր#�4�b������������kZ֣�ѹC�U�B@A�l��y��r�`�	��Di���|���f�a:��y�WV|n�n(�6��R��݉�&WH�����\k�\��X���i�9y�������B�4�C�Q��.����B��܀"��0�:ա��9֧%�_||�ǋa�#� ��!L���Ϧ]&&��������UL^/6� !kO�0@�d*��c�ƝZ`&u��R���^9B~��,��k�Φ�D�}g�p��"oY �̐6ϑ��e6�'�A��۩���%w�?eRxN�ز߫�x�g4i�5I�R��>�hwa$���Q���������򷘼�[�]�(9�����JC&�&<=��;	������iU� �e���NN-�Gp�Zk�T����G���B+��+<��*z!��D���32�h�����!��\})��哦|_>0�^�����2nh���p)����W������Ï�r�i�h�H�f0�̈́<M���P�K��ɷpH3؉18Į&���q��Tʨ0 <��R��Ǎ��C�I�?�;!�*�:6���gP�c�F�?�;�6�?�GϠ`��S�56��Eϣ�v����	u��Zъ��D|߮�9Zsxp�N��eOU#���IF���53f��m,���2�{����|Z�e��c�r��f�e}��w�mx<Lы�Uz��s]:K�>�����ʛ������uQ�-ZԻ��o
M�쯞������@
�ɜV �7����|�Oc�I��>3��~����K^D�1�����֩��s�?o5u�5e�Pu����>����55JSb�C
]���2��K�K��T�z��]!b��O�a����QՃ����5���~���o	朣7�/^ن��֗�_���4G�7�Gl~�Y��@�_�dW��s{��J.l-"��Τ�R�V��sJ�k']�7�4گ�=��-��?ȹ��P�$S岨J��f���S�2�DLă��o�Y�Ax!��l��B³�ͳES��ȭ]o_-��(�GV����5�n�z�+���W����<�Z���;Nɭ���W���zKR�j���������ȿ��)����?���"��H`=˗����vqv�7~�]H�r��L��y������`���؜�����j�}�&��%F	HJ�@�a�����%)�1�a0���K�A��������η�������l�+�羯�(��~�_��DOq�h}��,^c̭B�f���?��;<�B 2�'ύ:�*�j�9,������U��@g�d��Y���M�"���)�����
nڭ��r�26Ur�_)�uk#��M�5�]��I�]�@i3U~�6�2N�t�e��M�l#^�G��"V�u�����P�g��dT,�x�e{����^糃Oi������]���j`٫�)���������$��Ɛ�If�@|��E���t���yÉ}�5e�v5k\r����q��?@��˯
�.
m]��f�-��Q��jV%|!@��.8��Ļ
�+i�����6��t!co�U��;�DjA"L��Ѫf}T%o���s�Hd�ޡ�$��%��?���$�9c�Qo��G��U?~�.\S�3��aߌ����#��e��[�
[J�YI�[��-d,
���ɀ��m��~�c���vR;$y��ۋE�+u��O	����94��*�;T���~��4+s��&FBƬ����%2A1B���Z[z����m��jA5�� �	�##I<�}_.gwnĎ$�9x�� ?7��0�}�64�6E�*D03��C���c�#�x�PJ�m�-H'�>NBJ�d#��=������EdVc�F�S��$��虠���Qx�)�!�U})��W���}W�!�7)��qh��:��y��R�iV�\�Y0��wV����﬉=5G��2���2�]�ʷ$���3@,q�1K��#������R�hde�>n�[muyGYo?��m j���Q�`�{v��7P��9���0B�T-*�  Ѐ�/o^	+��Y��ס(r�jV�����m��/$���X����vҽ����\�Y*��`.`
x���2�gF���Z{�G�/�4I������t~��X���28M�T���HD'� -���흽G�姌��|N�XՂ`�*��4DS�f=d
�.�	��4�<�v��t+�o��kMS����~�z�ւ(ޤQ$k�E�~��epm��r������gG�0����wґ�v�]��!�u��x����.~�|��ѿ�?�z������ܤ����(ܰ8ۜ�h����~ւv�B���#��A��D�濖p��J!J�65ڎh��E�{I��){��t�I�8@��-�H�����+��(-j@5�i����x��pD �R�_���*1��ܙhH�$���}G�ei7�P���o>c��.�����D�y黅��#ҟ_>��e�����m��1��>���鹎�M�����@L�اY����3��3i#F���Q/���ф��?Cd��!��7�7z�h�,>3���7���^�tx����Q��8�Y�!���ML�m�I
4+��ԩmʟg��Fgg�����M3�?�MI#B��glbU��!���n @� hEJms�e*S�|��C��m�:��ϯό\�Z&�|�P��#��N��y�3�\D�]�p-�lټM���*Y�-�>�ab��(��s�]{�`���`O �A�;�}\&i�J|�~�˰���s�#��������Y��)�`d�?��|�4n��N%I��Gn�G��&���g�ؙC(���h��
����|(�ɳA|��Ǣ��3�Jq��^νG{h��菮����HP+./XR3�)����=���#�?��D�@�.�k���B��٣�﬿~	<�}�:��T��gQ��٤Tq�C�S���_#��WCn�n��Y����aA�y�w�P�oZ�œZ�6ޛ�|�w��D;ީ�ϐ	������_��'#-��bX��s�"I�?�G��5�rb[4�#czM�?�����L2ש��i� �n�	�m⢰1�]N�����Ȍ +J��`�l��ilo;3�N��5��9��~��[��[Ӄ�_G}39��'pw��c]��s���G�����.!�	[�9J��3?fk=��ݒRR;2K��D�W���h�?���1��o*�U�>�������s����j[>pQ�1�$���I:l)33����hY
����1�WY���q@��x�&�ZP��ծ'>:��W
�)>�_�(�
�ǔ�bzj�����x;�� ��w$�@�h[��\IB~����&i� �|ց:��T;2���`݌|R�1��nu�a��x����N֖���c��y��_ĈB�RZY�Z���J���>�Ec��f�+pX:W{���dt�"�ju�h��ԘM�)x�
�c�jc��-4��&�M���їS[�2�f'N�o�հ����)-kZ�n�����jE��TC_F��Ο�M"IL����3�D�֘�r,�eT���Fo�vϰ#�Aתg}A"%C+|m��Tܭ}��]ղ�\7��[vU�Iꖻ6�'j��1:��:�xe],s#�3�evk{�>��ZjKh}���^� H(D5���LX�O��aҢ������d�N�l����PX\c�l���i_���fꘝ�?��D��F��J��yZ�F�nj�)�/ރ�fToG
��y�U�f��t,��՘x���a��V������"����$�ng.���]h�q͚e���Ǎ���E�����T�8?���3ۑ���l�_jWJ�ۢ���삟��:����j�|Qx���3i�s����e�w�Hs`DS=:�Jj&���YD]ֻ��#K���u�%s���-�C��DOa��5�J��9����;�Er[ۨo�:c��O���e�,������3W�b��\����c1�c=4�|�ǳ},��ÿ�3��xF�������&M[)p��ڻoPH�.�́%��4�8�b�(�069j����Z�O$��K����ݸ�(Y1{�~H��B�!�����^;�:��l�#9=
<�9Mk�]�9M���̿r��;�:��!�w���{p�]�S�F�'���ĩ$b𣏔Ln��Z}��?�Ug�W|�;Ϊ����y��]{^����ޥMB6��u�@�[j��"�[��$���]h�����'�3_��;+M(\�CLFTM:M���ґ��~:͙�-��أ�� ���W��"$����E���Z�j�,p�FY���W,�$�؅��_`z|�d�4�K�+�����DX�����}mےf�|uFVE����ò�o�krF2�8�I�� ^�����N�^9���l����5kT<�h�x�V)/�T[���bbZ���

��R.ѽB:�X �\g1���v&}�ݍVB|��?ezB�8uLp*UO�a��%�����0�r�h�Q2��I�}��	��HAP���쳅5�aUp~w`��Oj�$c(ɗZ'���lic�Os��I�ҙFy���:���_��x�+�Ec��MI��r�	ʅ>�v�T�#|�Pr�mP��K�T-����gxe�� o�O��l:H=�ΰ�k�-K5M+�%[A�WN³��@mI��V��9�T���<�s�<#�V?�<G���+cV�S�e:�����o��Jq����
=��*��m�jO���nű�d�Z��fc{?�X-A�U�F/RG	K�@����~#ۜy���QSC���^�A�ja��4qS�Z�Jah��7�ז���U^���p���@�<t
��X#?�.���B ce�9T𥔳k���И`�w�\:%�t�Sji_]��U�#�����kg�(��qo`�/�Ȣ\H��U�|��ᦜ��Uٽ�߭�.=^u�@ާy*+IH�K~�z�-��V�M���Er�ej�GY<���}�{��z�vB����IB��6I�dݏ��7�E�����;�)�(���D$�7���8O`�1OȐ",�B�k;t��#��ܭ�D?/��)�<E�Ķ�8��1�p��s��ڱ�(��\�Un�����7�$�b�DFv�U.ou[LR[6
c���,I�j���b?�E�XE~��dַi�.�K�BP�l�v���d2�k�~�����VڿFl���&��fH�� 
�Q�ANs[J�OH�l A����e�D�pT=z�`n���%\���6���AZ�0�?��u[��7�OH����զ.w2@���~zs
�i�[��Y��|��C�e����ث�wY�k�UP#O0�n��b>ݏ6�~+��ξ��߄ՃZ��#�%��<��y�K������f�p���o�$���/�=�ު����~�V�x!�d{�F�x�cyj)��U����%����ҳG��r��%��p}��i�S;,�I�oV���-�����j��(�o��X�~P�W���b�������/RuxN+�3�?�8~��Yj�4���h���}�Q�Χ_��O����M����5���f3��ӥ��(/C��ڧ>��zD�Aģ�ߕT�nCjW���uˁI�H f����^D!��E���;��t���^��˩����w�*�^'�Z��7R&�.���Q��g�!=wu�ůl��FXL
��K�
�B�z����8?�ԛ������9�D�XM�Pg��y/fF�%Ĳi�Ʋ@���Řy�OקF���-��2����C��8k2+[�^K�슚�
9.8=�"b��Ψd�J���ud"����G<�cY�T����&A�l��x�*�7�GZ��U����\���%Yr�C��s�U ؠ��S1)yGRmڠ��}���\*cq�`$�RPnΠ����n��l�H<����;E�y"��e= C0u�e�ųԬ�x����G�`���hLR��hb��Snlf����k47���HM@�=�
�3Ǐ���eL<6������;���<���6��e1��m�U�w��]��'AQ�%�y|����r����KL�Ĳ�[���/
�6�;|���C若x��#�֊OV	�U	����:z��;��k���T;
��f��_����t����b�~���{큃o;�+R��e�����*���tb⹢`��������j2��i�]�.|o �?�u\J�������-*_`����R��R~%f0���@%��
��UQ�;����4������Jl.O����g�!B ��ȈL��/�$cԤ�#��6����C�k�7���GP���1h$Iy�\����^�HԍFj[�ЗJ��N�E������9cU�L�
�̘w"��2����I��95�5 oW#D`,�&�)D5+��1J)2��>3����f����2t�N��R�J�����R손b��_X�$r�sL�`3A�2;u:1��Vh�Fι���.��2�!��I��Q�F��G��c���vX�I=}�� ��jx.�z���+Y_�+����某�)4������
�з	fy�]O�5�3�m=���������T�X�Qɂ�^g�6L/�����Py&��v�*�Pr���AԷdܣ�o7 �}����9
#r+�꥔� ?��,�X�[�v��)������������4�$�ѧ��}k+��w����Y�]~����7*0K�˙�k_K��Ț��	���H�O7<϶�̴��e��&<�?���t!(/��Vx�}<s�~�}��S|y�0v�x9�6�0؇����O�ߩ���i�Bju(��I=+�Zα3��ENS�a߷ު��jr���x�&fU��{ª�>��T���k�R��&U��v����2���t4D��D� �4藲Y7o���y�k��o����Y���,C!	�_K�����ݎ��TN6�N9ղZ���W/ʋ]�:���ib�+�?��.�&�������1P8��J�rSr���Z���?7�q��V����A��^���[�O6��C�үh���A��u��}��X��/G��Dٞ)�c��5Vz�4�=��ƞ��m(,�O�qv-�py-�QU���r=�&Ä���_��Q�b��K�~"螞w�W��uO_F����
@d�
�h���DY�f�Y��m���yhG��[��?�&�ܭ��˵ȣ��֤��zn�i��Q,#햄>��y>���u�R_Q���4�w���Ԏ�`��}�K�O���
L��	$�&+�v�����������y1�T`���T�dW�ޘ�}��z�4�+&��ɱj3ʌ�mO�5J�$��:R|E���O��1���gd`�gd�������1ğ��s����Bނ%t�����q�x��wz�DH@��� ~S���ЀNs��Q-��m�3Ӹx�'��qt1ц�V���9K5�������j������ǧV&a_��5�V�ͪaܰ�%+<w��Z~zq+�xP+��7��Y�L+y�- ���G;����!F}��_��e.���{�R��ߓ����53J��?j2�)��4j��0zj�)w%�EU�s���"�����ˋ��H�j�R���n
	�s9�.K&7/��bl��tx�K~��\����D�q"9?%ف�6�����x뺃�2�4�%���.(�V=���]��f���$벱�T&��O��E�D�e�R�(�`������YAm���0�?�ĉs�»���A�~$ʏ[�@ �@zi)����b�"��|}���&��[�|������WcԨc�K��K��k4�R�-2�o�1gȿ��ȶ������-�4��QbZ]+�n&�M�%�r�([���f��%*��)�҆�����ɿ���	Lz��xV�y�z�JÙ'�8"/.h�Wy��%��4cz�T��"U���2�� 0�d�E ��!�C+#�2{��!��9f$L�H��z#j2�3m�6\Q�w[]����^&ٷOn)d��lû��f���~�/b�����e��g�JouM��º�oXI�>��S9�+k�d.�K��Eqd��d뭆��")%�0��ҿ~5��D�9��>� \�<ړb��)$���+kg�|�BT^�Ƣ
�9�!POt��� ����=h9g���]]�MCH�kW|���P��NG@��V��p@#��&E8x:�?u�ܩG��H�C��!)������$YRy����3�����q�"�$y~�8ߋ���P?}��/�_�[j �hU �`����L!�&?��@U��"�e�T�_�+��ˡ���Gl�1`��)��H�k�ܼa-3������Y�$�9����QH)��$ai�U�jƚu�.��&N�v��)��*L����	[�H�c�O�G�J�P�`S?�,����BQ�W���T�T/�I~���a&�.��+5�,ET'�zE�Tp*�g5Kp-�w.�{�Jb�\D�VL�rր�G�b-��e���w��O*�!/'���2�.z�e��������hOx� �ۢ�K:k �At.%0��R�t,�|�+����|yxEk"���5E:Ȅ���̜_Y�P*����9]��ɥ�r�@p��L8����Pe���S��7N�4���]�ſ��
�g9=�j,:'�f����h��׊R��[¤Inǟ�zor��W)ؿ�yW%z���7�?�O��G���"�r�\�3�i� ���S�H�aeaw!��G�;�/״���S�:�Mz7|����g��}��{���f��<�~��A}c��[I	hY�Q��%z
�"D6"ݙ�~n�������������9|��h(j�l}�w�J!���g0�wg�+VR����Vnn��{�W�]X�����O�h1���8���M�%��Ǚ<7թ+ä����G����VΫ����f��
��Ǭ�]()"�ٷ]���1!�X����/��*�3Z�ua� '
+�a=g�^AuR��"�~�@����MBT�:�F�N����ʏ��_�# j�j��yp|���_��Ua��S�����su���p��cS��>��4��bC}1������ٴ�����) ��.�ކ�Ґ�#�ٸ_	�%T߻�� �A�fcFD�X/7������M<?��s<�jpb�}@+MP7s��V0z��Y�k6Y�p���hR8;��\׉`�P�)3�V���?�\��F� (�Q���8`�o&�$^�O�T��ũx�Y�)L%����<��g8����ns��*��g�R�n,�S,��i�'Ǫ�͈7�=�F�$��Ve^Ә�/�/�T��Y0e�Lz��(@<������[~U^���m
6�O{\�-<�vU}nz��qXm��͵�s-�P!�P.<k��$ �(��.x?�?�����I��_b;A�h��Z�,���p�X�y��d�#La�C$���mƜ�����oA.f"�����E�W��jX�l
�q�:�  f$~���}Nƕ%�W��~���v<�0w�_�Ѷ�m݌!�����D��s	#B�ȝ� @�D(D#&�]j0&Q�~�M�����Ggl�ۺ3�h���qP`R�DR�jRJ/�mz��r"����������k�WQ�M�x���������zD���Rm,g!�R(3�o�ю�=U�\3�#�S�9�*����:��K�ﳠ�R\�d/S��t2�R���kS�V����!�V��W��V&n�����N��D��|F��O$�w! �y�dF�J&hHՂ�g.�^���|��п3U;S�t�6�ֳ02�/��N0��r2�_m�Гq�JQ����JM�æ�|�ہ i�:��~{C��ir�`��{�ox��i�x�<v`�Nh����^sZ��u:�w1E�������[�ҵ��^_3Ӭl��S	/=#�hj���*I��\�↢y�gB6�	��z��1"9^�vq��R��<��{�[1<�C+8�
��Դ�#
�Ԕ�7t[�љ�Q�Y�-(+�(+"(�#��Q4�8��]����
���PR?_ά^��̰�?��qm=�i>���iW��"0��D������^�x�!��0�I�����u�]PS�UG��ߣ1�r�u�U���/��;���{���Xu>:�Y�oL>� k7e�I5�D�і����)JMM{��N�|g�̄>���z.:�wLA�W\7���r˷�ò�f}�uRwx�z�Y��	����S	և%��/{~X&u�F�����<�6��$Zd6>�"���p[Э�w�K�+���_<�C��H�ָSx����� g�[m:` 
x���f^��~/�~_&�ۺwz׍I���p�RN��������l���a�����!������U����٢Ӷ�Rv�S�3dF��>&�s<?��(��Q��Й�V��g\�R0h�5��1N�v��R�ܫa�W��,$R����G����ul#��a��m���=H�#)��
%�Ç5 �#�{h}�\�4��;Ɨ>��R�n=,���ci�+������8���KL��	[a�.�U(��_7BP3��Nͮo��-���%�\aݵ���������������=%����f�P�R��)��nz���/yz:�y���\2+���#�Sx�ɏ'�"�\�;���Ŵj�_ռf&��?D�d�g^X�^y���$"�Y)��\h�Um��$�O�L`��l@��9�:�ȳu\��N9Z�/^�F�{4��շU�Kq��&�H���D�U���<b��.������QA��W	����%~SKJ^����3�
K~��$&���Pp2��y�ZA^��]�1�٦6�,�x;�4�a�}ʜ?y��Iaw5k��Nx�ԇS�f:�z���R�3��jV��J��Ι�9�C�޺�[H�W:qW�I��)ݲ��MK�����M�d�fEA%��5AKm�TJ��������UR�Z�iS��C3�`���Zc��:-#�ޒ��a�,�����z��,DP�ʭ0���Dm��Q}�P��P}��r�{���4*�f�S�R���e,f�&͇���k�d*�dlǥ�#��+	:7�FX����Q��{���Y_�k�����_�����,q���,�j�^%����-9��A
�M38$?e�ʠJx��AU�ऍ[7w�����IC�zf�W�������֋z�1�Կ�֋Dؕ�rᆃs��9c�㘁KO�: �I��p�S1�\�ʫ+���P/�(p
Á�^`���M:N䪘�dM]K�!rQ�ߴ�]�v�r>��wB>H��ʣ��,��5������;�2ȅ>������ȿ�&���}�����_-�=�@g;�Tg�������%��.bSA�%�T����������Vϰ��a��;ʊ�ߥQ�ݰ��(��)*b.�p{��0�e.aNZ�|nz���Q\�7O1Y� �Z㵭�V��̇����xp�<)��7��}s�J��MB��t��f9�m�5<�u�|o$8��^=S�06�������+�����nn>����]�ߎ�'�ل����k���e:ph.=v����Ҏ�߬1�A,Gލ��T�oQib�C�\��ЄNF^i����t2^��QΧ�-k�g�Rިd�j��keMhRM��d��T��x����*dM�6���h���� (�"����T]^�6����̰ࠌ��D��Z�}��^��DC���k�?ӟ��@-�ڑ{_�\�y�{vŌ.�-����$�ᤔ����u�+z"_-�3�g�Q� ޳�s�1�=r
��>ϳ�����3��q��e�RV�9�lfK��gOe]�Ʒ˃?0��*�J���TN���%O8����	�^s����it`�nD���5 G�V(某 ����i5M<w�|!;J2-)�)�e��B��F�k.P�w��K
��CRE_Y�D �^���3��\;s��Ѵ��ig�}�}}O�מ����ĩlG�)M��*ހ�>@L/�N�_��c����D"Eu�Z�{��y�c���18��2?�gϊC���Q?2��y���2le���DX#<��bl0�U��1}S����d�PRxu1���ZV(e�X[�L���4��g�p�K��cʗ��0���;�Xc��v?\.��T��e|�?WE�77���^�-��MDO#GeA���WVW������,���la>�zb���_m���~8'j}��0��R ����V'��CzԭZ�0ΰבsz��Қ��r �<q;b��g��H/r����Ra,	D>�1�yE>Ӟ�,9⚾L>�q+\:6�qnȥ�	� S�f�g��/���F���L'=��]ι��Qi�+��{20[g*�T���Dd��!Z0����ơM]Ӏ��A"u
֟g�ܘ����"��'v�4O�c�F`HIa��u�_!�jyi�~*߆ja}ݔ���B�W�wD.�X�:ʪ��>� j��TD�����~ww�#-���FN��j�_�Y6�F�2�vЦ×�?�b:'�q���x�7c("��L-(
7 ���)%W�Ai�yr�{���G��PMf�
w�z��C����2�ҿi��)�aL*�����_R.�����}��=�a��1f���?#?|��d�_���D���.k2�n�M���aG P��s��@}����-Ua�譎}������`}��}�b�k5���4���3�#*�g�A��0���_�_�&���$�W߷FH�6��XT��]���'ɹ1OӅ �����_<��-��V��],�_�]�w��}E0h�0�E�Ղ��8Z�����擽�pd�Ф�溦��䇩µ���F���͹W����G�5W�_���Jఏvhf�\�D�p�O>�Y����)��3uzۋI�B�վIjLBWd�����ؔ5Kɪ�	>��ID.���c�/.�5�>�v�`-Z5AnQ/�Ȳϲ��!/��D�Cx
1��fl�5 ��ޙ'����x�;\����g��v'{m��u����_��̯4���׾�x�^��A�I�-��A�玖�'�b���+���[�o~�������[��[~��n���ÔӢD񉭢C�;��@�:�n�4_X�7��&�	K�t� fJ��H�rPH�/�u��r�#��.ʣ.��\�h���0X\�Z��0���)4���[�uθ)7o!��8H���d�A,�# ���8��U�*�##i��a�ȑ�󐏀"Lb{&��R+r�|�NB�gI�%�lP�v�S����c�����w��K�k�?6I�,W>M)����P>׿8_��?ڼ���l��TiΦ@��1< �?�'��n����
7	8�?�f�O�lLr:�?�����Q�<�䯣F�w�?�9]ղ�����:�ߒ�xG��v(^J�j�ޖ�F��	t�w=���@�@�d�����훛M�67^�ޜD���j��&4��+���i�}׳j���mWۃ[�]��H|����4�ȗ=��GPC��7����ݓ5����8�vj�+�E�m;i��b��ڳ���y(��� +�I��gS����ӿ��-H�@Kq�6Ε�����18�!�A��rm�k�k��ե��p�����>G�4H�)º&
ڣ��U�B�i�A���z]�4��j����������������%��)�셂�y��u�
�������ӧ��v~��=i��/
�q��	)ԣJ�^ �S�� �?P ��ݒ�Z5>]�Ax:\��Ԃ��a��Cc�L�_��� �\I�S��?�~�m$��rn^��v�0��_KJ>��R�9�zV/l�/�^:T��`�˽�~\p�jH�P-�f�<�%��q0N�f~�<�h��*0ϡyipvH5&n�����Xaz=]ep�b�4��ic?ek�x�sn�$v�.o��y���T.[@<>�'

�~��w�5�~*��H�����%W����""��ľ�/GVP]q��Q��k�D�щsE���E#ПV� A�G���$`�����Cm��8ۑ1ɘ�C���ʘ"K�G>��#܀ת��`�N�lg�J����F��g�2W`��끭G�r]�6#�=�p�[�w��f����3}	i4�!���D�)����ߜ���|�x8�W�4ѭ;��0py�)�3�<Aϟ�E ������8���=�Q|?�M���B��ϴ]hSX�k��RJ3����ȯ���]+�?n6���r����5Q���<RW�:������4�C���Pv���m~�2om�Щ3��#V�*��&�gPR@���<�լ$Z��B3�a��(�R�eH`F�Ÿ 3\��*�����G�"��(�,{^B���sB�v@��ц��V������sy���Șt���J�ܶq5�볅���ڸ�({��&ɏ��/�J����d�\�`�!��A�+Z�Q'7����g ���6w��{ 8����%םy���Ţ�/c4�.�hc�y��������_=����j���c}y�����5�3� �|���PO�S����S?���<V�K).��������������Y��)���-�іѕ?���w�=�p�������z��8��۵�x�� 9���j�߱NhX�a��9�=D�u)�:*7���kF鲙	�@�>ac���5|�5���(}��珶ӂ�T{:qx���UvR
<8���).?�>���z!1:��Gі�v?f\�1.z���5�[�st�PǾ#�~��0U4���	zk}�]�nު?�u��aҌH�z�i/�i���ë+��[�޴���������e�����g�No�w�>PB�c�YS�l����bFZ�-�b���B{,�3��,^���:����-�Wb#W�N�����Z��ě�������*��~𱡰��%��(F���\c�D�8*\g���$���=i���>B;�Ao����o�]���pz�dv�wm�j�f+g�zɻ���o�U�'h��%���H���aS�[T�00f���k�����IM�����p���XO)����Ѳ-4W3㳪��O��	kB�hߨ�s�����>`�N�\�U�x97��h�?S��*�m��'\ޱ�Pf6���@�o@�wV4��cy�c��Q����"z'�[�<u8w�f"����Dg���3TS%���fddUVVvt�{��+_�lg�Q�d�o�����~��^] A�g�4�iA���1����1�]�`C�A#�bF�#��Gt�dD�L��{�s!(�"���{��an��f~[�R

C� �fu�ݙ�Д`9��n���� �/�4�S�Α�9Ղ��*�)�׺8mT�Ƥt������6ȵEb?b=, ���>Я�ͧA�
��C_�TK�(���mS.�@�1�8n���]@!ĭÆuM�r8�TH��U�h�pd��UL.���ްڮ1J�ܱFZP�,9��+�����K����2�~��4�z��G����]��9*ԧ����7������E�UmW��,!��=��,�'�}&*Ē���X���_Ĝ�aQ�?�	Z���J_A��<J'-��si�l��6	�:py��jW��i�����J`�oTwv���S����.��)b�y@j����� )rnP=�n<(�b$2x�]0��Y���ϟ�4j��q�..��\
�Hna�G��C%Q��y)�JX�\(�L�O^&��?�dЍF����	���pԽ���ʑ��V��a�3�
?������?���%�;��ňƳW���w���)_�U�" �ѐ1�̖�3n��=��+�����荳�����P\9ۚb:(���R{���]��G�_L��8��	dL%�өJԴN���uq*�y��J:�Z��z�>��O��"�G?��F����Qݖ�C7P�(��� ������d
&6���6�L�m���-�WQ��fxW^exT�����:�t�wySu\�J�1K�I��7W����x>��򧵇gۣ�e�+��Fu��lK-��(M�:85��sY��B}0���Z���(5;�[XdiXbdK~��;�?�1��߉ߋd��ى*s	�)�f\?�I��׵�.M���.�����������q���𱽂2|s�<3�AH!̹�p��ȟ�+(1X����Z��a��!n$jO��V�r��h#����OC�y��F!cya�wU,(<oM���Ǡ��׸�c7��W�o�_�t2�T���=+�j�L��ؽ��fηZ��=/{nu�d��~��2���C�٩ii��=}fB�'�|J�\s�����^��)}���6��u��}�����\���g�w�+q2�:�F�T�â�dIݩ���H?"+�g�VI�c��u'�ݮ?Y7T٭�O�Ծd��gŝм��tD笲������U�ho��>���"{ �R���]��^��F��>��Yn{ر��z���������N<�n�uK֨ߌ�L�2{��x������S�3�wC����J��#$R3��Z ����e�6�S���[K����M���߱~�]_�'L	��$U����Z�j;�m��~�����(T��W��'�"��݊?�V]�>��K��0t��ރ:�1n��]�����l���N�"T���92��'Q�\�w<ӁD%2܆}�����+�6�{dGw��c����{;f�g'n'w&�Q~��W�YHJ\�rrF
e����iz�#	��W�<yQ)� x��k���W9[g�]x��)E0���"'�@X� ���;!z�Ї!��$�Q"A����mǒ)r9�G�/Z0$Z�>���@�jE�#����i5�`J�*d� �@Z�33��!��ʟcn���Mg���H
��M�F�xD�ʲ�U�3���K*��V���"~�]<�׸V��l�q�F�h:=���t�>�-�̫�1�9����;�θ䫦f)�>�{$��5��S�5���36K�86�6�RF`��C�AI2� �§�"zcqbE�^{�o��I�e'�b
���@�C�m�t��Ӻ	c7��;��WM`�u��cn�*:����ߝz�-y��b�;�z�H*��`Ab�Ա�����o����Cͽ���o��i﮽�[ﶬ���[V:���Zh�j���`�H�7�N0+��D���,aq�R���VU�Ŧ��QU�d����6�p:�M��lx���O� ��~�C,nl|=��k�f1/��^���_J��i3����azN0���)����m;E�w�!���it���-z�����-�ǉ\tu|�ʈ��$z�Cyv��J�j��t4�s���d��%�RR"��(�*"�d�	S�`d
��l̀�4��r~D�3.�d����z%�c����Ͻ������;�8�G^2�}+|��B�#��><Cը�GKH��\	X�@Oͮl]���4+�+\�ڋ<ZyJ��i��6��\�ԯ��;�W�{x���ݶ#D�e���٥�h��~�;�
��r����~��p֟���$Ц��S@̣n"�����I�� �5���Y��'@��-e����iv|f�1�ќHrTzđ��8��a�up�i��������G���Sr'�!��=�%���	�cq��5�(t#��í��]��,GW�s����+��S�S'w����Gy͆�Դ�J�iW����&$���Ű�mn������ҝ�������_��=n�(�A
E�(�
-N-,hq��-R4�bm���Kqw+�/�P�����3g朙�!����u�׵�JH*�Ҟ���DZ��}��
s�~,:��^i	z�ȭ�ՅK�~��n���L��ds ��8����XY(hb���UW��4^J�U��,8��~݂�|�SU!�u�k���>XH���#��ҌNfeF���g�{����%}�Zg����懤�>�v"1�<�[s�?�l����vD٣
V��E��5��K#�S��i&X����0U�����8~{g��r�Ϥ�xU�Eh�@�!V�;b��卑���� �_�Y-dxmd�����W.��I��Rl�/���=T^0��;�	HT�W6��i�v�Q�g�т +�;~��"f�Ţ�a*Ϯ2F��=��_�)�����m.�\,�P�,�.�}\�԰a����N8�]�; �T{6�� �|��?�ؘ�Z.O`}He¿�m\����6�^D��*a����W��ϱjP��Wйj�%#��q���#�v�y�cwe7_�����pW`ǰ�mg�b�}�q�l�mӃc��oȽ�T����ރ��Ń��M���}��iA��R|m����lZ����p⎉|͹o�j��uK9/]��<�*&�"��"<�T+1M0�ѿx�h�,��-gH�� q~��������ف�N�C�#�rzN��Q�8/@�S������ן��A���)^��A�슆VŸ�p_��`@&���n����E��g�L� �BQ�7z���u�P�oՇ��Q��>�M'P7���R���� D�70X��j���$�H���3r�q�δ<R�ĺbD�/�~�Xm��\�A�#Ld�t*=:�9G��FK{�-���KX\�N�j0�I �~\�|����15@��rq��b��LVt��u �A������*h�3u��M�J�CbA�Y�θZ�������� ��o�EU��h$���z,�g��$�-�<�dw�42�:��VT�B�R1Ω�:���U�Š�2��/81C(��G��
Y��-m�T�4 ��:	w�|��<r����"YU��*�G�&�%��h6ǓP_�mN	���*�7�&Op"�8�y L�diE�(�W#!y J�Y�C�^���^7�|B��X�+��+1�&���VCc�%�H��?��w�fV��m��|r�Ԃd!�e�%�}��6�n��ە�7��# =��,�݋��qp�B��#0��_)�� �-)�3Hj��޾6�E�&�I@r!�f��C��N���B�^�S��-�Z��� P�����zn[ta��+�n�6�������{%[�$�0�ʝ}��� 	S�j�=�xړ���L�ᾮ��oXy�մs��DilXM�pCc,j"��n�j��FI�l��uw]}�m��$�G�쓶u���Di�?�}�dDo��?�'	6�z��^�1{ND�����9	[�;^W�r�NU��\F�nY�|��D�vlO�n���qRש%ݮ��_iG{~-���?Wp��X)c�,sH�b����<I�K5Ry��e�^a���ri���=ˈQH���[ �g�i�ʇ�C%ӑ�}{A�x��irq���{M�d#��
&R��V��G�S��S�ci���q�cx ��TH�P�hl�y��p�Y�h)�jK�4;q�SHf>��ƘҷSۻ���ݕ.
�+�����B���gRJ�Fu=�>�͇���'���c��O�h������-�]f��U�rL�vQ!&.�$�O��<�ەT�4��V�����m�@���!��|��u�NCc1��T��>�I_����|W9�:��S��B*�O/!�O��Q�<$�e�E�ű��j��O΂$��E#DU?����T���bu��ϊ�4�]���JZ[9>_���tbƌ䧈ʷ�*Mm����G*+�+���9DWƌ� �5x.NO��KO��0�q����Z�č��3?H��-�h8P�}���`P�+0���$d�ɳK6��\�d`'�����>�d"$��A:zA@�?�0~!A��엟��TLmiM�b�D��9}B��E���J�h�5�2�N��� {��6��OK�>���A4Qz�(��TBTJ��3 �٪
+�aD��&��t��*��Ĺ�įTVˋU[�\��Z&��)YT����`�zhͲ`�����f��`=��P�W�{���%�i��l1��S�=-�p#�����Q��MT��v�?D�%��0i�=��ٺs[k��}�۹�1���v$���ҏ[G�y���A'#�HGy�tY(��wg��i6��5��!���!e^�'���B���ͥT�G�&��7
Ӥ���}����@��]���E��=쯣�3Vç���s�)®u#�����������m�O|���7kZ]x��5i�|�}���\�|��� ;�� 2�O�b�}���0b�j3,��c�2щ�MA���/N�M�I)~���$�v�h�=lqe���kQ�_o�D�('�_�/5,��%:��xzY�q,fN���ª�	i7�x#d�+�cPBdRD�h�s�4qʹ��})�\!�A��J��#�;������:��(ctΛx�����@W�G�=�{���b6��9p�AC�h����sp���ѱ�T�u"�椎��g �����;�;���6~��Tˋ�����#	�`C�o�~�������h�ZU�:�K�J*c� ��d�p��Q���^Q�.�5����k
wd_}��\?���~��u<u��5᳜�J|q��T��w�Ĩ�
�6�{�9���RâŢ�7�t�F@v���7+߾q��˫���-[ԕ1��0�G>�E;�K;gB��E9�-�TCW��f�w�N��"wqZ����=sd�6r���f�qR�v���r>�r����1���0�4<�!�mcB�Tb:OD�m%qi(��
c�'F��BW^�A t��e�́[�7rf#bf#rj];l�>��sp�/)�4���ZM_YM�1�ȩ��9ȥg�Į���囆��S�TOXW��3�'��c�$�(�K��?���P(��SІ��	��9�q��Nt/��H>�1*�a�>��1�J����}>N1P�h2i�|9���D�C^��,����#�1�S�����,���PHGiV��\�,ܝ� ��_S<�����6%}����n4��5,��/Y�_}��*����{���	9W�f��:��<�<����\�[���9~�PZ:~�2���pR|�Tߖכ�4}mc�rz(�	2��M,IsYB6ʜ9����c����u�Rsz��Bͱ-!j���4�x2�y�v91|�U�U:�x�nw��lP{.��3�̠k��Z��_a�XB���^�������B��A9��dY ��3D���o*F�K�g���E�~D1�7I?���?�Afe�]󗒼����6-������\
e\��]&MR� g����.F�	a�a�R	����(zX8����p������R/�<,ƽ��:�:��K�K��E�3�j�pjd�I-%�*da�%�Z��aC �����KzLO��m�
]�~���Y݈�ϯ�3FĦ5�ż`EE�੯3V����i�#j��1	�@.	�z5Y� '�`�CR� 0�,��ZnR��4&�~Ԉ����>j�i���dD���ʏ"P���m����H��BI��T���b&�G:��p`j0F<�� ��ق��N	sN\
�F2k-YS��ᯛ��J�y����D�S>�Ѥ���͞�6��>Ӭ���P8�X���SX�stw�׬!r� �'�kǗ����2���غI>W����y��h�>|�:��~~���U��w�FFNV�2E5��:�)�1�I�����ȋT�p�D$
P� �~��;�V�
�ƉO0��D�",Bd�~J�V8&q]�Ae��'7Xn]SCȠP�}wu�W��`�S�ǫ��ƽ;|�]��r@��I�5�fЖ�i���~{��;ᇜQ��|��K����P+�)�|�Q����,����?�^�yP���~�*Y_��]��� �[h�=Գ=�~?��I暯��6��g�_�6���o2Ru�
�B�${2�9M�.4�v�n��!J͛���`&�-��#�7����e���.)~L��&<m�����-;4��rK�×'�i��Y�׶��[����+!��:�W�\�.5p�{<����6��Ku���&�Y����!���_螾k��3�%��R�x�*c�x����彅�N��5��ɕY��m
����v���������C��!l���R����*C2J����ʪ�9�� qC���	e��+Y��`��QkԦ�ƉW"���Xߢ���[;.l,D�;�ħ�g�an�*�D
YW��~��ͼƀ��^v��HM�	KԘ��ЮQ��wa�1**�����yd,���i*U�K��6mNʛh� ��о�U��|�eM���GXN�辰�'n��~?���8Tn1���������U�h{qJzӗu�/��w��bu%;2�;ǈ��幗�N&��}�L&�[T�3��-r����x��v�%�\�n/3� ��^�o�EҪs_�g�����+2��EhS�UѺ���3p��$����y�;�M;i����w�Z�j^�g���}��iO/Ţ<]<1�@��S9^��l�D@���� �x��a����8 ��(S@wr!A9cB�b�"zPDQL
�����8�^ ��[؋*������Z�7bԯ�����wN;�=��0��� V�ܻ���ӟ�N���Q�	v솀bZ*W�
p��٠���G%�2G�0<Þ�0<-w��+֓oy�I�b��g�7aKy��W2���j����.v��G��hL�_����W��������%�R3�9̱��)���-�}��."�,��V��|?u���'��j9T|����:;DmAz��Ko[�<[eL�܍~4_���O�հ�Ǉ)f���C���j��f7���RG�Vo��*Q��ZS3��P�x�a�_(ޣ&�F<�[�x��)�����Zp�h
&nIG)�س�v����}m��FZ�Euh|�8߶[h�/q���H��+>#�l��T*����sr$�b� ZE�Wɠ�s�T�M׬JL�
����W�'F�hWü���|3V���{
�#��EyWH���-���T�[�ڬkg�D~��5�5���g46�I�Ԣu���43U�k~p�Ml1�F/�L��<
p��]l��U�Z�l�C�-��)/#D�""j>~�h�_	N�D��3����^E6/<Z&�֕�7��D�����{��e-�1�JR��&⻗�O���~Ü��k%�_��,D ?1W�ťD��wP��s�߰���;�Ƀ�:�_�mń5�r7��M|d/��.`��nW)7���S����J�aDJϟ䖄�jr��RW,�I��d�z8ϊ�ؘd�/zw�`meu߻c~��o-��&#ыC�k���_C����j�v��r���{?I���b��w��9!z�t��scs{%$ŁWk������]lE��l)m2�����`�ѱ�2�D�����@ a�	�d�@��2���с�F\M�é'ˋ�Y1'�d��,�߳&|��̊�3�Ss�@W�p�p��o�IV��)�`!n�9���.	v��N��~$��z3���w��ZQ3��t�vY��F�Z	�����S��G��c�rؐ�~�`I��x���|}w�/�y+���9eK�~��%������6�灌�W~:[�,�u��R��GQ��~3?d�YS#���<���?Í3�3}v�w֫{��7MĲ��dŤ���S�vFSn�@�g/O�7��5���e�>6�6|��z�?.dF��@������r�������3�L�ʿ�Gيr�E�K�*[F�q��j!lQ�bC��E��ʯ��^� ���\����P�y%K�m��G��OMF�)��p��ǲv`7�m酮�8E=�I�3�Du�ߊ{���~�<��'j��2e�{�}~!ly� 7�\�7b@ }�"D�%��z�o���E�&g����y'#����\b~��L� =�d���]NGlNGG�g�_���XK����OQ[H$?d<+�iTә�~5�k���j��!H��4�P%�:������ۥ���ٛ���ks?K��(vՙ�"��������S���q.��~X%����i��0SdGS�c���O|.D�\ν����g�i둓xR�}��ş*�S)u9Zɿ�2��
�JrOp��#��G��3	F�� 'Fh(�������	�i-p��i��Ow,����^�����ǘ"���r��/���h�rx��t�����¯�$�>c�!c��$�{pz� k��)M?WA/�È��f�I�}]�����v�g�mg���*�Pl���E�=ηNA��S9��l��T���e|�����zX�� ����n��j~%��(��ũ��mL�g3�x줉�|�hbK�1�k�g��WI��0�Y`���d�I�jsE�;�)��_-`0�=I����>	�����Q(8\X�6��M��'���W�9Y��e�-����mqX�s\��Xd�zjI�آ�!�Ni+�T�"]���t��L�g)o��֥�$A�nI�}����};�����'c#`e-{����xdݙtE�|�ȪWul`���8S"��NyU���y�-��[�	W���)�l�1�� �2E]��̌�?xд�ߔ��0	\�Ǌy���Gu%���ã2�UF�C�\�g51���a�e�Ʃ�kIL��Aw�w����]E�7ъ�*��'�@Q���KX�KQ`�
�ᥙkԨsJ��*e~M��I�ݢ%��:6i�����B. g��� Wd���,5���	%��,h�5�	��L��t��{BY:R����L��d�$㗣�����P�xB<'+|&G���$۪'�((0�6pՌ#��$��[ј��|2�}��}��9�?D�@���I��F�??��Y�.T/�>K���y�6��7�!X�7�#{�n-�⟷͠�ٜ�.Rڈ&��|�(��ieܩ���`,ka�k�ڪ�;�<��!l�6�A�Ȉ>:2�r��7T7�̈́����\b�4.�C�dyu�A<��K����c�����x^ێ�S�6�����5�|�����������x��E�d����H��Pz���p�gG�s���.)҂eM�F^����\��ّ'W٣����7Mٷ�����^��u��W��?�??�u�9e��s��!�`��y�)�z8�]�տ�(�hKe���Ls4?�y�``�󆌜���_�?%��N��p�>��"%���x�,a�6��H�1�'o�W:?���ǢTH��������.�~��Z��Z����X�+��C�Vۖ
x׊@�~�+�����!N�ǚЫ�I9���[�;3��\߄�XFe�r�C�Bc��ʔ
	�M�m�J�_����͵=�?)?�
Ĝ��1Y2�KcEdF��{�#Z\LG�����M~��+�5u���{V@h1i�Y�$�$��C7S2���V��y�.�nh��U� (�E��+��4���- >(~K�Jsd.~��#��{~z��p���g���|Q����|���A���E�E�l��J��{B�6�*�'_���xݾ����S.��$�2�
Qv�v|�qwRu��i�ZX;ʿ6
�52}�aa����B2 �1�Ť�)�2�����c�D��ι��m�������y����0�V+��yY���!ǋ�1����Hw��ǳ�R�A�T�~%3�$���J0 O�[�\[�\[�>������.�B{3��R�#����Q���Q���ɋ�@g��#�۔�}���.g�����w�1�Kj����f�"f�q�2( ��.?	1 Vn�!k$����v��zy��r���M;	��hx��c3���z�OŔiU��(|�a�=
��%`C�e�"���ÕH���ݾt;������/.�KO����i�ɚ���y���j�N����'l�6�`� R�~*���N�+u�����#�e��~�3�l�|�|c`@�e��#i⎋i2� � tE�������2ƻ~Џ�Ū�C�7�a�C��l^�O��	�B� Ƶ��W,�4+�>|�a�;���n��+Έ����1���������������F�*N^;�'�}H���$о��7%�-H]<nm?�^�����{ͪ0�ELDc��}d,q���~�,uzq�����X0`~2vs���[ٰ븾�;����ҩɃէ_����}�	ʀ��6�3i�E]�b0ZJ�3��6����άX,�{2��S����cx�V��b_fzF1)��oEn	��=�Gb��3�C�<�Ɗ���H����X?R�C�)��7�i��7u,�빗�,yI���n���~����U�x��5�>�J��n�g��������w�Q���g��?�U���-��爟�|'�S�-}Z���f��.��W����e������)��s�sJ��t\�E������N��0�H2��i�Im�"���_/�����L$k6/֡tY������IO�`����4���;�L��Cd�y]�����$s��93���}_�X��a_�(�Ojz�����7���g��8<Wk컆��w�8���^<4$�^(����$�/�d�oH�1x�*+�D4;?�N�f\�G)d�c�%�GaC�Q�w�&�H�J#mˤ�sO�ѳ�@N$�e� ��ؤ�̨�x����P��٨,6���p��H]� !�C�쭀ak��3��Ά���Ƃ�1��\�o(��/�����Ξ��l�=Nٻ�O��̯�;G��9���G�VW�o����*	��4�2u�& �f~��l̢�S��r��K���H�iZ������XL��C��U ;7�`U�>��Y�k���' Z8�D� SR;EtJ[hFOB+e\��2á݄fWe�But����� B�%�|U^���E�r(T����}m�n�s�Ў�^4�^OTX�&����޸{���������y3l��	�w���JE���G˟^Z���(���Y��2���8�9��&��P{������X���H�x1��{�c��R�1CrAr����O:vH[��/.PR��;���b�d u:5��A}8?����),!��G�~����~y��"񨩡����b3&��Z����dRn=�ⲷAy�|����5�X��:�NDj�GU���,Xۧߧ_����Q�����i���s��� ��8FN۹��%�	���y-��FUu�1�>��s6�쾣X@��lkP!s��*���
:5�")�*>�T��x�4���m.��=h��ʪ/
V�Z��v��I#�)��M5�;�������F�ƙ��;�:� ��J1��O9#�Wk=m��ߠv����#j�����-W��K䔹@�fr�$��0���>OQV�[����~u�z��jF��E�d�v�lː���l�l��'Z/Q������m�} ���6�g/�7;qK��Z�񨞋�}���9K;��`�͖�(���~Q"�ۉ�V#����h��Q��*�b���a��1k:֙wK�$�fNA��zR�*��T��<ăG�{�M$�Tf�>�(����{N��+�Gt[>�N&�×4�ڝtgՒl��U��N�m8�9�#�iAy*�L鄴佚`bxG�BZ�iF/V$�^TN�kg���������em��G(��AɃOɑpuXF���#G��(}`�1Y�Jy��a��q�AC?��>z&�����
T��v�=���A�q*�o�T��$�ؒ�Ҳ4��7�*U֑�/H���'b��u�X��!3K���(�Ic�j2��bK".ר���Y��}��7�f<��Ey��tE�7r[��/l�yg#�F��/���[6�j��,��~^e�g�lO�e��?����Y�d��n���9��ǅ�;����.�75nFČoɮd��=l���0�e��:'{�.3ףU���4cw&�_5�q��/G��I|�����M_�3G�F6�r���P��B�M���ess��@���E��C^b�T�j=J�4"�1^��A�XH�W��;P��ۚ�ѹ����`�@ֱ��d����Ћ�SY,;؞	�I=Q��Iܜ�1=�?��o����(q�%�/!a.&M+&K+A��]At�\�F(�b���"c�$V���N����p���)���afGSi.2��ʵU��4�� ��zATeB�5�Pl������չY�c�ԌE�#gb��Y1�,0�Y��%{�M��]�Gk�΃k�֖k��q��(Z$��+��LG�J��xB&��vxT��;|୊^�T�����GX�������m������񀎩��	����X0���B��ɡ���k�8� JZ�阅�qj�6���lbbm ����_t�
��O�[& b�e������mz� џ��K���ڮ"�env]e6�>�oߌ�z	U7MT�̢�Fè9��*<аVKB���:�G�]�y@�����>��*�j�9��\��5	G���[H CE�R�F�2!]�b8���8w<�I�GPH����*f��j;T�Su����3�I���д��!�j/���m�X}K�~�i� ���F���cC/6[�O{a�[~>���˥�MO��Æu�m��pޙT�d��c�>��ۘs��8�w�j��EL���ؗ�� %�ߝ��j�%<����1����;���X.�u�}�p��X�1
�\{�iP"�Pi��5.�f�h�o������Σ�5��_�̬DA���i,;w���1�Zj1���b�(xh}{������I����I��{��+S
�3�xJW�2�����c*���:P����%�@�
<�������������	���147|ܥGO�����z߸�RЫ��1�R�5�G�Bke}<��� V�	�"���/�=(�hSkb}���Sq���]�)�5����b�5�!�ǫ5{%�XQ�$�'��D�o*����%b�<��N?�~�r�Re�`���,��GfDѧfQ�FѺ�=3X�0���YG�Ui60�42<�Xd�9��ٱa���M3[@��v�x�c�fm�O������9#��Y�ل
���f���e���pO݁���@C|m����'Z��7Q9G��n��s)��*͏�������vn��D1wFf40e�q��I�o\����4�ө������Mn�<И�a|�i
X>,�m�Qf�qF�p>/�n��2�c����n����h�$ZU�<�T�\�Eqk��)�%7�_ߡ>�$�{������36�t'�o����	�f�-� fC�Cg�T�8�{�ߌ�����i5�JIi"���R�w�^�>pH��`|�%�7SmJ�|����8t��3u)Ɵ���=�i�G�%��{4�Q-0���m
f|�+`H�'R__��݌6մ>���m΄Y�R�ϣ(���'�(�eA�i�C�AG�c����-1�>�P'�#���J��Q٫'a?�E��{݋�#�^dD�
����Vѻ�i���JX�(�����U|JR`��rt������q\$$�[�ў���peS�1ac9������$
����I�|������$����5m|�Trl�_��\Ȥ�mn��Zݸ�n�����؈>>�tAD!%��B����{!T �T��I�T�'#���Ƹ�=�h����}{-�Fs>J��0����zs~�Bn:��(�M�_������9����{/�p*K�Ȝ����4m��K����G���-��Ž{��s㻉����U^�g�&a�[���-��C����Iԍ�����F�i�Jd�, �G����G��!B�a�g[�+B���3�MH\X�0��4�@�s�o��� �j!�"̷�n��Ki�B�66H��aY��Z��T���[0�9���20|k�.�����~28���6��OS\��{�_w��|�gC�l��r�0��쭶���70wU���S�����݁�#�"��B��a�(F�)�nt"��Y7�I?����`�����Z.-l��7r:�'���zH��Ąn������R�L��?I|��EcivG'��� Z3n������<��.��&Ὼ��6��,���.W�h*�Z���EܮC]_C֦��@+kk*��]�:a�o s֗ʪ+V&���B���J~��B��c�r����8��P��y8��O�uBQ5����2D�'�`�x�r���`�`~�VP��@��Trn�_-�m����s���SvG��Њꮯ(�	F{��t����T��X�ã�,�/sD"�lS4����WN��������ǩ2KϿE�y�&����C�^秓��0={ztry������S����Ji_+��dQ*��e��ٽ�0��밚/�ؚ�,��X� UҸ�.~��̥?����f�/Tn�@�\��5�G�����:�Y�G.��CWuw�}n��f�!v:y���&_9�UFZY6��z{�����;�R������wo�ս�#g�1'�@yvX�u^��a?�<oMnB>{���z��ggRge?1I=��Nl�U5)�mވ�e���Yt�K|E�f�~f6�.���CϜ��]��Y�$�c� s������:����%��6�y����%���P���}�m�'�e7����믦��]Y�KC]��µH��Mmca�AY�F��I�=$�>��[C�;H�,�0����9�G���!Xx,������� ;|7���(^����Xx�+JDҕ��A´U��������j6�9)��.P'B�2)�Fa A�sA �3�Ss#�'*Q���7�w�]����.u������h��XF�X��$ ��
�r؟>��@K��J�{|�byG>u�ݏ��T�
��ܭ��"�|����@
՗r�(`E��4IE���Tt��)Z*Y�������%,����l$�?�$YQ�_d>�����5��ݪ�;��woW&]ky$O2�ھy��}�:%�ʝ���DF�&"����	4�����q�z)�jw)�L��f)�8r)�^���D��������L��jBq1�k��k�T��8�fh��xz�8��L�F�{�2����u4ï��Hm.J2�'�vH[�g�Y�,�9i����uF?:�=F2E�OUb{��-Z7�q��P�):� _1�II�*�B�B��c#�04Ì��e��g�wn��\R�Y��y��Pl�Xt�q�
'e�nq0(mg�@4˜�������IqX�C�hAG*�xl��¡M����@*�2,����)J�����4��/F���JTj re�bz�Y�������s�A�=/����"ZR��?�-���~<�-H��y����{��]7�Pr�.�Ln"�{X�s�V��?YR��M 3'�
)��7:-��;9����n?}���$F�+��V������t������Ӥ�i��4�Y��؟��{~������z6�6�3d�r9��D뵇�;g4s�[L['�hc���`-�H������灲��.#	b��'���E�N�^��o*�Zo>k+v[�cՄ�{��e�\׫^�f���>�c�]Ǽ~�L��b0B9tiif	�V4�k����g�6������Q!��ɟ�Zi4+� HR�?:ɸ�����Oӑ���fA�� �����j����4]�j�P��%#V7w�
��s7v�6v�8yB9y�1�-�I���!a�K<��
�nQ�h�����������B1ҷgo�r��#(S8���p{&�:Q� �Y`�k|��2No��O����_Ǌ�OO%��q_G�
�|a��~���S��,D����ik�H�X�����}E5�c���)�B]�Q$[�l�Q���o%��3���}�b�m�}˰%��ҿ�\��'�>&����)�^p'�b�b�]ۻ�	���Μk�r'9�\:̪�X�ಇ����V�Jn�����w!/����2�ُ>�W�M�J?�/�Ae�^�ΜzO-�ܵ�%�8���\��v4ݗ<<lɱ�?��cٳ�t��.z?4n�C�Ԕ[L`ހ/πK|d.���eo��S�i�43G�f��� !
ڲg�dl�Mޠ��j@Y���b�n�@;9�����6�Ojdr�k�z̶r�z�l��k�po;J���[||�;ҵ.�P��4�]�~���e��2�I���o�N7�h׶��.$k5�NN��(�I�ȧg5�|�S�;쑨��:���#.	Yѷߞ+��Vm��j�C�q�������;�zX���>�y���0���%^/3���e�N���@�O���O�~��rX�d�g�Atf
�h-�P-G@�0U� ՟�ࢲ!�Wsm�*�u�&�e���|E;�������K���K�/�9��s���e�R�<$�j#�'Z#��c.�9Qj�%j�K�����FUKT�ȑ=p���G�-/V�\�:�)sr|��jm�q��ȑB�8��c\�5�1�a�%,�I+kz;M4!�����O�c�h!�ik�x�g�-��?7�)*�]��xuV�)��f���~���-��/R�_�2=��V,d-&6�ɏ�s���Pq�N!��)¼�/�e�Y:Ks��������7�����V,]�Wț�K�k�� 8�Ƴ��ō�7>f�"�p�*R�U�r���6?��1^���֭�w�CcOIc/Qb��L�b.��L�+X���J4���-i�s��aǟ���{l���f3�
M�M����PR~-ot&~t~t�M4��ՒgP���܈�x��z?��z���x-�`��
�5��٠�~��Q��k�1�!8���[B3��X�6t��iH�2��I@Nlx <��"��Z�OTG�����z��>�y������k���$���8dǞ]��a����������B�Y��o0`*:�k�������.�$k�$m2���K�Gu�P�Woe��5!�S��Q���dI2m�N�K�_d�8���Z���`����Ĺq���X�>�Y������Vz��0��|��2	�Q ���q��#9���phkpH��7z��o�v�v���7=)h|�3��|���~�����,���Χ��i��Y�Y�X��}�2���XT��]P���lL�n˰L�1�a���[ǭa��_2����xP�v8j���͇OB�b\�*,����Ē�ژ��6	dR�����o�(U��*3�� :��	�	�4NQ�WO�-B>��S�M�U|>�0�
��$��fv��J8�w@�Aֶx�[L��Ȏ{�t_��� ��;u|2���`�����(����r:·�k�c�&\v���C}�`�_J���ϼ>>{Z�V���A�m c�^����+����������N�j���wU�˞>y,�}�;���4M{I�����(;��=EE�
?�!�>����vu�9K�_T_UF�J߂���UG��:�����Ep쭄�Fqh���b���Zp=�A�9Z�mD�RH�o��0cتa�w�?�����2JS�����V��"�l�u�M]h@6��=2@���)�o���q�`/OQ�1�������lݚMh�������<cҗX��E�X��R�/S��D��#]�^�vm���'[�CN�v���1��ސ|)��f�%}�[p�ͤM�[�@�+�˃�����)=��^�w�z�����x���^c�w������� {A棯Ù�t��l��1~���"FP�E+B�VVB����n���C`@Ț�As��B}���>~����׵O��<
����׳hM�^qd��X3�������_�F���#�����L�k��-�ο�~�B� ��Љ�D*]��	c@��Q��$��I%d�N�/�I�Fj�ɜ��;7�@�Ŗ��`�bѿyQP`f���v�/���VK�1�Bl.p�X*�XF�.�N���--}��u��2=�#��X�<i�������-A�V�|CZ�a�l�\��>��������9��~�̟�^2��v�?>"��S�u��niy�bf��"sjn'������8����R�Y"��v�Bs��mG6�&����E!a����	a��Ly�����8�˚GL+1�DI��v*�æ��;�i[-�����l��CnO�s�L�y�q�r�ׄ
z�Pj�o�����3ٻ����ͥ���W��j���� k�z�c"�g�'ζe�x����%��r�z̝h�=�Lr(P�u
�B�\���o�dX� ��ɡ$g"�p���ܒ��Q��@�8�A�
.���["W�G��]��b�#���: |X'26o�^P�%��o1��z��`��IG�s���p��T��z$ �:��yu/�e�����R��s��T�rx^�Z,������k�{�>ݥ 1D�6�q�@@�a ��twH3d0:�����--����{��{���u��s�}���p�&�[�5�t���-�oC�l^f�'�>7k�\+nW�®eMw�-���?S�S��5B�1\d#�s��\�ͳIF��:�+��]�+2\!|�W�5�
֜�*�)�% I�7�����U����6��C1;\�7�RIL+��;7x�Q��������Q8�[s	��ז13��uV0l��Ta��a��t�k�#�J�g������Qv@���YBU�q���w2-��Nk�3@􂱷,Iӌ.������:ʅ{��g籈����ӳ���i��\wI�H���Rs�Ѳ~�)��Mα�1�b�25`�*B�ۂ�
a1c^�c���f���B>�k��⤡6��FF��	]٣X�t�Ɯ
��D�S@�;�h��}y��v�V�h������	k�5�Q�g�$47k��O���m��=��}�?_�Y[o��o>�����="D��w)��-��{3H�{���kH{�b��o�}�Z��z��`6�dp��B����J�B<և�M9c��y3���?�?n>E�6O�����6�Z X+��c�;�E�P��W��w����<���d������[d�;�$�����@. `\��bRE+�9�!���F�D��iv� �+$4(�M+�K-&�+�HG�FiI�C���2��?`�룚�U�"�4�QG������ʵ�4e;(���dO���R��YW���"x�!�"��f~�j��Z��1d]}}������W�'���r�F4/Ik��)�G6�b.j�v+d�+����V���"�~�c�����Q�
���k��]}$f��l���,*q��j�R*^ꂧ�>kD���Ȓz�t�{�y5�j{ �;B�� 
aE������0�@eu:�\�I6�-���� `ݺ�J	�첟��X�)��S9��C��fQZ�ƥv\��=g�~ŴNF��%��ۼh�j3��q�It����L����i��-nf �J��%������[`J)�]��ƒT��@��\D
��� r�:\S �b�n�3���7$����_��eXAUJbQ�!�|3_hD�I.����ꅲ��u��G�U���ߊ������D�~|q՝�қHj�r-=t�V$�^�l_�����g'a�#Ɂq��k/��G�6�#4�����	�\ފ?\��\s�j	�8qh~�L��`{�F��`۞u/p�=�J�9���9��p�Z:@��+�j��3����F.},�Q�%B)Zk,�d(��Pp6ݿ����8LͰl�t�fѮ��o�[�灶PJ�9�D:���τ�ϳX��
�m���`5��s�M\׭����+ޗ���Y-��ę��+��6�x�
�0��-��`�}Yf��W�⻥��
W�/~���o���/���o7��^{}�?1_�^9�݄���&����%�A����õ~��t�h��~T�e��h����j�.�5�W�x!w����[[����,jKD�L��[}j˳w��H_�$��E��':���Kp�}�c�����}F
���*��p�t3c�I�e�sd�����K�ƒ��"������,�s��:����X�c�BG�����Kn�P>�.�L�9�G���܎�'k9}+��e�j-��}i�������Y�/Ս�H���487��Cu�&A5�+�]�6���"5ĩ�Ku��P�c�}l�P� W��Ѫ�Vћ 9{?r��ʗ��Q��B�J��3�迩��a�I����S�p����F�ݔ$�f���m�I����RqGw�/�:�W��[�)��R|6~�2�p��9�E��N|l���3���DM���Ho�Hm��T5��K<�K��_kOU��(寰5���z�l�M;���00��M������L��Ɨ`~)��k��ۿ�2��Qd�n��,�nU[��/���`[R[���)�uG�����~��aX�f���T.B,x�_[���y��DT��z�ȌJ�y�)�7a�������fr���o�}(�(����%"�4r�
�Y�hz�Z�k|���i�WUV�d'�2����z���=�Ge�F�$���F��INl_�7�LB�	@��J��퀞sA^�k]�[���96���Y���Ǟ��_��#ۇu�{��B'_�giKY󧳌6�rۯ�	4I�A�K�;��AX��N@q�Q,q=�(!�e��>�Ǉnx�������o�R�𵲳It�Y`�vs�-q.z�������!���Gt��H�Oȇ�X9��#;Sa-�-h[���w�s"Q�!��G+	�{�����������mJ�mj]+��
�Kʙm*�kB�ǐ�&��d���L-G��b�¿��`N�G�`iɿ���ϲ4�a:h�y#d��%�9�-����&�2�3�
�v���X۳�X�X�[�&�3�Xe_]�����[��t���M��È�+S��P�C�'�t>���)00!�n`��p������q�8�=�h�ݟim������w����$��߹������5�Q|&�ѩ�fUN�8	$��f(�UD1GV=�o{X֡C�z�l>�
`8���ui(R6�nj����@Z{�)r�1�;R������:�FE�R��逢�y��/0t$D�B��IC�_����M��Ł&����(/���Q���K������'7�+b�@fE��/�x^����Ϻ__Z�ޝy(7��?�7� w�U�k�[�g�-Ղt��Y�ƭN^�~���YB{J��s���Z�D��!&�sԥ�=!\��A�v��>�A��v'������X�iN���oOu����#� �+�j�h�dR��h��M�>/k�����B+�·� ��o���v����e�3����zu:ξ�ߪ+�0�;<ik
W,�����W/"�)�7�ғ$�R�6F|�Ң�z�9o����e#Y(���{�3��m�M��왵ģ:}�	�/�]_��;qjy��oeXm�aU<��||V:K���

�E�>��������gWVI=��T�*-ӣQ�1��%spx�j�Q�Uh���dFi�{]������E-8O2=���`ɩF��#o��d���g�&��2hdAp�L�8�X����0�,�_�5\�b������ߡt���p�2���,����dbR߾�� ��S��"8��4M�����8�ВCƙE�YPޙE�m�����;G�v��o�7j�'0����<nÀ�4�I1���n���#1d_d��\#�A��u;���AE#1Ŝ�n�Z�v��U���d��<q��g�?,��]���99u��
�X�t��W�ˢ�թ*���S g�q�E��+��,ƾ{��"�Z�H���ɠ�NC�����@��t�X7R�3���h�Fx1��$}2�v\�#"zZ�(v1�4��\u��.�'��h��N݁0'N�ц���]��$Z.��1d��@E]��5�b������T����'��E.ف���]�ʍ�n-��&��c'�O����n�Ψ8I�i��8��I.p�&,k��I�qN�&39��Ύ��Q�SLa��oY$�A ��	yI��u<���Y����GK�L��q8�]%]io x��ݙ2���ϡ�hg�y�Q��~�=�P�Ӏ���-1�D+�����	�P0T��R���9�����Ь���YJ�ҧ�Ц�УD�	��X�TqR��D�V]yŤ<A��xL�Me�La�O��/B'�+zݏ0��[U�+$��~*R�q�f�l�r�Qf�T���wŒ����K����_L������3P�'�b���([�	��l�ed�5d�-�"m�
�q�(��O�EoFQ+�y=}��+���3>���}�t������9�5�˴kn��v���)����M@˔�H�7�����s�����-�Vپ�XSCJv���y�V���������&.���������c�]�[�&4C���9J3���X|���2�<E����\��Y�2<&���p��U{�m�C�X�q�5���>b-uA��ftꝩ�u\�k���m��W-��f2W��=O�ۏ�N�f���Qp0G�ko�9�Q~��=$͚F
ă�!~F��C~�A�"_4�[x�&5�	~��5E��z�|1���xu��h�����K��b�g^��䓼��ܡ�P�Ǩ66��_��El���~�?���lV��A�kȏD��*��?�ڟRD��#Ud
7�x�������q�*�+�s&�^�N����h2'�5�	$ J����w����BB���/��|ۡs��VDv�NFl���8�F�Q��O =��F���η�ݟ�h�P͘ �S�:U=�:;���_>������й}�N��u#k#�T�4��\��.���~蛟�yQo<��%z��9O�A���z�E	$����<U�ϡ��ϭJc��Kdx�y��>݋[B��*�T�����VB#��ۛ����v�l�j�ȏj���%\��wq��������|zY�q�Q�	��W�����8
��e%�W�z��+c
�KV�Є�������k��y�u�N�) ҁL���4�#4vYܙ�/qy݂4f1��xr�,פ0얻2"V9e�(�e.�;R�פrm��S��~��*#oo��(������Ж<��?o�L����3'aF-�30�x�{���d���94���r�����.Y�B#�D����_FI3��6Bg�l��m�b*�$s�H���m#�;8<���Ds��')"��И��"�l6:� �����NP�5�t���9H�����w���nYH���N����R\d� P�KCCm�l|9��a���g������/?��9�U�1���p`&̤���A<�#�Ѥ\�*6��.l�7�!��[!���d���������bV������Hl��S^���Ih��<d�"�Xqr��n����tk�*_��΅�P$�3%���e@:� �n��<�X�����H#�aU`��q�0�}u�r�uk�����Ͳ֑�������������3"����0������p7��A��$�8��Бozj>)녩oV��?��m�n�C�gyN� �s�V���n�|�CN���%��VTPf����n�L �{��O	��1��B���0HXa���k��b`aɡ�W�n~���������W�y��"�@G}���𖬹���{����29k_,p�=L&g+s�xo_��B̥��>������y��x���6��\��ت��{z'V��aD�n�	N��T	"Ǭ�87�H��t?�v��h�7nk�i=0±&-�c@��VgYUE�3cf�=N�ق�p)a=�Vc��%�e�uV1o��	�����ދ%�������%4��/s�>1C �9{�������Vϝml��oT?H��u��O���S]���Y�~�Pc��[��R��$���K�C޵� ����,2%�O��*���r,��F~�'EJ�r��ɢ���՚���|��������;C�W�'��-&���g�#��5:�yt��FK�(\�����:`���4�%?޾Ϥy�aB!W}���Y�u:����m&���=b�]bs#J~���4X���7G�3�&�K-��<��n�&�ˮ��H1:�\8��l�mm�Hh*�5&s�wZTb�������j�k��X����#iުnz���J~ۮ6t]©�MNX��_~LbPd"fL��|!5sq�>�F�Mv$.�ٽ�]�'�*���ʈt6��­q�[��}����4�DԺ�
>R%���g�N��-�Շ�d`զ$K}'���MŶ�:&0؍��p�z ��:�9�*�p�[ɚ��!}�^� nR"%�I����}���7f��y'+�qȟ���BQw8�-��b�ʈ=N�M���Hg��"4lT1�ь�����)�A�ۢF���#2(�e�+R^냿������1�T��b�H=H5Y�IV%��|HeR(X��믪N������q�?�NCd�s��,���f��hR'�+�N�hȐ��#���*-������1GP�%���0z
>Ю-�
6� �O�6T�.,AtЧ���e���|�+#*,�C^!x�I�I������P?���L`g�=�C������aP��Ұ�����{-2b0�������s�srH��fO׮�����aL~��=��=���C�`��&���S=��o��%d�
f���s��}V��1�e��m\uc$���	(�jϷk
�3 )������e�j����+��1S���Ӊ��j/��T�b���t����_�����a���Y��Y�Xy��j�TU�_���B��F��H�Wǩ�1�	�|� ���l^P�RУ�r%�%�s7e���̿�������҄�nY��;CY��ojb�'a
a��p�F<���KtYI��~�Iu��:�eÛ�ǿB7V�"U鰨����2�(u��p��C�@Q�L{z�	wAp!֍�|�2�1���x�/�Ϸֽ��5�mͻ�]5��}FGt�|#��n�t��$��CaFh�)nA���R��N=�w�+y���͚_�HC���ƍ����7�u��J��w�j\�p�c�'U�����P�)�G����oW����Cz�ٮ�%����!�\�f*-F8XB�iT��`l�g(dWwk�~<O�7�	j/����5�Y9�@�ƪ� ��@0	��}���n^W��ew��Ҭ�+�F��*ޚ�`�p1���  0ǜҳ��WѠ��V�c�@S��oN�tz<�(�����׾���9 �L�Ĭԋ�������-�LxU�bT�ӑ��K��LX0�z6 �Z)���Vv�%�k�����,�t9.���|?b�����f�_�" �O~�_م�?��E�Ç.�BՈgJfлB�_m��c���b�V#Q#��Dl� �,q_�Ĉђ
����[Op����<�7�s��p8B3i���I���r��C�f��n�A������.�n��<�+&Ĉ���~���W�(z����ŮR|,��z^F��T��m���j���^}���X���T�ɘ���ʛ�I�o�����*n��(B �d��R~��̤+ �?���G���*O���B�
z#��4yϳt�w���M""�zK^����]�O�7�fP2ϲ�]�z�e���h�Qp��h��(�s"�߶��_��lxg[��+ � bLH����Y��Yj����m�_��Z�+����@0�XV�� ����ׯ�bq�b�*Ļy�WUƞ/�����ג�@��|��+�HC�:��+}�xRC(�a_JԮ��]߅n�2�$锞�gZ�{��H2`p5��H�Mz���n$��Vw��A�{��J����)-���$�Eli��J��3�9j�
!2�WJ	�m�'��q��ݯb��]��̑2!`�S�W\�?&�;)�2t�8f��'O��{CAL�:|���	Jpfs�
'BE�� �N�h�w:���:ܐ=�IٻT��&�v�b|%��)1�,��[xp�Q=�~����M�g_)TO}/�c�N(|�g}5��Ş��5>�����$������lz�nw��cG7��h��C���%��BA���Y{T�$�@���H�/-��:!~��B#4���n���.����н/#�����T݇��y:%���#R"�g�O�Ѫ��K'����cd	@�>������6���^*t4�y�n��W�zM��V��L�w�K���/�� �F�c�ʰ�8Y��8�-�ܻ����4��a�_�ʫ�a�i���093h�J�����7�_|�l�]N��>M~�)�rI�xs4B�(���wi �z{i�4jGt�<=�kә"����v��b'���A�)%���D% ����� �C�@[\��-D�~U��jW"Mi�W=[v7/�DM����dG`�f,w�I m�k5��U�xYNg/��N��G5W�7�1�Z*���j�o� $�[zUž����q���i�G����<X1�HB���1���:r���j?Ρ��;)+�}Gh�g	��5�<���>fI�h������&�.�����K�ߣm����@�j'����e�z��X�4�${Ѯֿw{��O:h�1��/�j��:���x�P��植]��]����f�sݏp�)J�w���֪������ZC^=�S�ҭXB��hz_�$]у2�n��d�_I��i��ePC)�t��P5��)^��XF�Eb}��=�z��w�:��&���찒4��H%Tw�B΄��U�NZ��cU���"��j�F8��_~��1N�]�Dbkz���oub�1�ē'�P�It��ɋV��I��{�4Q:U�?&�D�C�� ��K�s8��(waq��|�p�S�*�߹�<��4�X5�i�K��o�w�M�����{��Vtʪe�z��:�1 5E �����GC�k->�W�-M5�f�F�sb�&0YD܂ �#��9���a#tH�y���)��L v��!��V�]��C�z�XK��rn�qGv�?�bd	��I�^��m����jbA˟ө��ڬ�Sŵb>�Ӊ��?c��zi�h��L*;"ʦ����g�+��P�����s�3��q�a�aj���N����^��|��2�*΍M���
��f��-���k�.�%�X�P��4�m��~�>�'��m�z�4�u���Qy��B"ѝA[[G����""s4����~�}��C��f�gM��cJ&��"�N��Y�q�l����r��������'��f��w�e�q1<�0@o���K�1H-��ؔ�����|a=��6�!�ɒ�X��fx��ݵ�IE(�!���ق������8�0�bJ�lP	0�U(���Y��q�+>��/ų�L =[l`�����&��z}:�	��q����IC|��,�.s��oA�����6]��/�~���z6���8<�{W)��a0dB�du�����L�uܴ[>��RQ-���I���*���5�~�&K��H3�r���{�x^CV��,���[6����X��4�^x?pK�-eXm��z�m���{C>�H�(D�9D�\:�6�Ȩ���
��J �۳�Y���?5�&�B:��g�?�µ�0��-�f0��B�Jɞ�*�fN1�Ee=��o�꿹ս"�9�6޽��Tj�t��s���Wm$��[�򩴡�����w,����!�Q����T�ѦC���^�~���ǕYY�V���Y%�%ay�ʄ�}Wd/�9z���H�܂��]��P�3ĭ�������׵�Z�0Y�®l�t�
j c�SawF�M���Q�H�(=攽Sw�9�";�bPC�&q���Yi�-9��uk�l�\*F��N�Q��0�6�o�-�o�U�˷*�^�la������M���2��޵����2H$�)ۢ��D!�
��զ����ӱ����]���2�ݒ�ۡ[#��v��.k�F���E	��+��b��%�:	�>{gN`'Q1��&��r��㵷n����&:40Z�p���xV�cH���ԃ銏��}�{[�L�k�E��]r��!F�+���uf��Ĭ�ʣ��ҹ��e.���D��-��הS+��\zt3�e4��f���%G���c$�q�&8�^��pUHF�[�Ř�� ��i�N��X�7ab�@�N23s�/#z�e"d[�
Z��;�Ncb�n�٠���+�y��m5�kW�	ʆ�i�������.����\4�h��Xom�Qg��_}D�OT0�8�I�#r�^�p5�j8~i9���[���RϛSϗR�;������k��3�F��3����ך�U]�=]����d�k����Î�2�1TL젅�YcHϫ㌂�2��֖�z!�eva-vQ�*}���/�_�]��U �>v���t v�<D��r�����\����p ��M�팡(@�̴���L#H4��Y��`ס�L��=D�����z�u=7�b�5��s#�z��m��3�~�o^"�ҷ�Xx���0}01|��?���n�,�w��x;e�����A��~k�[�~+Z��mr�G�@&��:.N[�grxq�s>���C%��a�_��`�8�4�u?ਮT�r���rd\���x�@������=m���2��]sz����p9�a�崎q��VꚈS���r���w�����f���ԄP�:�2 AW��sw�L����(�w�����)E77ie(\x>oBx�AxR=ό{Ăw�I@���;��e�iY��z�s���y4*���1�TƬk���b<��kZ�D���-y��`+�W�w�o�bdWL���@Gݰ������7���D}�3?0�z����h�
b�8>�aK
�4~����Æ����F�S��Sj���^��l) 2lr�����#����S�zR�����#-׋�����ʨOy�Ÿ\}ص{削*���-
������٪�72څ_�57���CK�@��*���(�����d�,�� ��r:�j�1{�t�_��\C�(�hV7��=C�_<	���r:���1��BKa��*�)����Z�g�Z���� ��$e���/�\���z�*�a=��!nP��s�����[{Eㇾa�������
x(x&,�*|߷Ob��g�$'�Lh�Es��|~�� ��`�K"��wT!�u���D�9u׊�D��
p:�������Y��.�p���.���0���>��__O)����%��xo��%D#��&�t�_A��#��Z}�����vV�STLu��n����N���H`E�Z�P_��c|kb��ɟ��\�tR�lF@Wi�X�����V�J�#K�6Cķ6(o���ڻ^jۯ���|aX�a��Ȍ��'1 �]��	v@{}�
�	��]�;� ��c���%����IZ]�o�N����g��3�_-���vM1"��j8Tݙ2�|� �����qO�'@"���W��(��̿�f��ut�wN�.�����?��g\ە���~9�c ����}�Rh��u W"IO�P��x��:���������̆1:�_3��gG�'�L:�_$�g&�����s.�ڎ��n�P�|���8�1��P�%�.c�
�k����Y���2�n�f���Wy���#h�4$�@PEX
���p�T�
�����`u�֗�vS�o�O��	͠�s����_��_�_5V	Wgx\4{��G4*J7FЫ�2��c���o�� n'wh��x�=^(��.q�-�-�N�N�N.�L�L�x[��>���Y�Es$ "����(7-���{zHb:�.{+�8(Ee����gg���IZ�����V�P�>���ޡQ�3�n �o�$��猥�1����꧉z�6@�wɱ�؁xK v��r(sHPP��m&3N�et����/	C0��:��U��?�\��y�V�?Ji���Z�����:K]��%�P��H N��(�H )�I��2��y���rZj�#f���ܯ��kV�Y�,i�7]�����h{ږ���ԡ�/R� (,Lv��_���
��(�'Ƨ���x�"��h�n&����?RA��5.UE�T@�JdR�dV�R-��%v��Z�������v�������j�E�?�AL��;]��/��I�Ⱥw�wO�*{��$DvA�z,��X��Y��+Zm;�E͟��]�"s���گr�
]�9��V����Id����>H�&S,����կ6��t9&�ձ��@��؊t������H��8!Yz�j]>� �������6%|Ɇ�Z�
7��Y��q�!���0Z/�$wi	Ea� -�W^J.�����?	��V��S��	K	�H�)U8�uߧ��*�tWi�jN�_??��3�l��g�VN����⥰Kh0����[}'k]3�R�C��,��������x�~�,^��M�G����A�R���M���l�hۦ�b�"Ѫb���˙�1�L�B�1_�1�T��z��+��8�v�t�W, _b�;��A�?��|߸qB�e��M�E���;�1�"�L�-����E�!tlD�)S�	�S�s%9~�����M�9��V*�)_�����Q<T�LH�K�i bJ��f��3�4C���IÑ�G`�	A&V(yt����FR�c�/U)s�`w��M,J��#bȦa7SF��J�̵��7�gw�>�;��㹾�[�������s�H5���a�N�����̱��Q�K|��������ѣS��ã���V��n�C����YK7�W=�lN_�`J~D�aG 2 /��x��0�{b��O��H�������J~�>1��v ��rl����>�a��g|��_�T���Qj��>�+����LC9�J�K )m( k�Oh�N����@Wg�?y��j�5x����}��w��gc�����+(t)��.��D�$��[�@�/S����4����t��rO�X�%������<���4���~F��naK����^R�
t���b�#��ID���P��R��R��R0rrE��0lǴ>ne��m����ȑv����-��u��?��{QflP@���0=��MH"]�՚R*P⫑/^��?d�R"� �	yuX�^�6��YL}�����p�Q������/!	��H(�4s���i�P�$<:�IQ,���0�{8/�-������I&E���X廬P��:��L��*�6�g�'�s�cm#�ܱ���_��fZ1�~Os�ü��'
X�:�?i����@}T�0�ix�O�Rh�RX�"s0h�)�=�^� ��_C-���zۅ���j�����
�h(�I؅U�R����!m�V�9-�����ہ�(W������Q���撦�u1���F�f�ȟn��Eݴ/�y���A�)�����6}E-w7;+��5J����z������D�U]��<�B4L����,Z�[	�|�����I)��O3������\)� �m�������L��Q�y�6�˺4�|(_��O,���9t6���4����!�
�cf^�,�B�*v-<�Wpвⲳգ��TR�[q��YZ.��g�F��5_��rW�6D��L�0�����ޤ@:QX޸]eN��n�oD&��I����&ƴ(r���R��{5��W/���k�N�Tq��Qm�T&���v�]
����)�(��s�a�) ÜC���<�m,����s@�����Q��t*�����(W�1�(�e{����l�2f�\Ov~�Z'�2����ňJx׻��q�b{O�%d����Uc{���4v7-���?�|;��a�Ge��h]��pg���fʖT�pi�/v�|��L�`y��9�^jBOt�]�]V/�ܮ�g�'�q^>�pqh�@���y>�Ҳ���h�8ǩ�"�6-,>sl���i|h/���*s�,|��qT,�_N�>a/����8�@����'��d�&N���Eۈg�Ȫe���$L���V���|s3�h���"�i[0�.6���֊�F<E�1��冑�_�}+?L��ۃ�B��H��eb	)����|�I5�QK�Y_veHU0Jqڒ����࿮�%۱v�������cy����A2
�$��$����QR{b�����#�W=�#c"��Q��i֡C_� �=�bJD�+q����9Q��|�!�G�/��$��B�B;ڦ�G쯎��e�ˢ�Y�����k���$h9�+Ο������(��l��鎾�?����=�̧�� ��M��C���n���d>�p��A�t�TQ�sk���O%�����ON�&��/�	'���H��/��Y`�>����(ܦ�H�#Z�U�@-�����C�������D!h���q��*�P��?�p�lv��%Mp�+��Hc�|q�>���i��B�{vmM�0fW�M[r���9�L������kϡ�FH���R̆;/�����2�f�ط���̗��4M�kv�W�^*�� c�6�=�tO<��Q���v4�NtI@�
ydq�o�QxrG���l��XְF�A?o��9����5��H�P2�I,?"����3m|vF��>��i}��;�������em����m�Y��Bq)C�Y������Kx� S��>[�aM�/���s�,�g��
U��/_oU�p~x���e"��D��&���to�Yq�rc��cwI�q�8B��hR ��H<)���ק8��e[>�>�g�V��97�Z��A���Pa�G�o�=��.�_�:�e:�R�M���{e���fn5u��Fs<5ߴ�����i���3Qo��a҃�@`�:b	
���d(�6$��o��:����L��1b ��<��;�,tp�#��@u󉯏�.�� ��V�V��,���0Gc(#/�t���E%Ǯe�Db�^[\2' ����C
}R��!Ɉ$��/}�,I��k&`im�4D*�%�P������i2I£AūM%�XN�aS۔+|�{BӀik�^��N����.&B?��w��R�6��0��$/�]��Yt�Qa���G���鴖~�Ǜ�������}aI��>X�|�Ej�@�t��(��x��[�vf	p����>U�j�:��9��o���a��c*�%���I��?�	g��vy����`.���5ѵh�3�E�zB7.(���+ϑV�tT��BA����>u�Z�{fl!�]&���+5���r>����þ+kyr��3�:�Y�����n귋�Ń����S
ךe�o�՚_�git�X��c9x	��6�b��;�A�Tm�����V>�K�؟O�)b8��!Eۉ�@��`�0�]w�:�L��ڽk���!�������Q&����ͩ�5��	���y�os�>R��ݗ��m�p�H�J����6�����ݝlW*
���T��6整{�t���}�%o�f!�I�R�uʺ��_�Lˏ<I��ڈ�5�%��kZנ��e��u�J|ŻbL��]�����t�=���L9�N�""������+��M:����2��= �N��՘��(/�00(n��t���e���o:Ln�~;����������^�'J��[�q����0�#TE9�Q�+~�p�Ɔ�kN������*���_��4Mh;},�#-�vZ
 ���R q[kR�C��V3A3��.���^�YY^������<�k|N�.X��if���2�������4����+{��C�������+�@����=K�V���eeW�p蜀)!�k��΁��%�nC�{T���[���|ٚ���=�\�����I�c�p��ڻ���#�ɽ6�_��x�UE�� @+���(�4�nxLUp�Q�,�W*�n6�~�b�����V�O����)F�(,}��^�o�v_���������#�?3>��>w��g�l��>�#:��6������Jz���i��E	��>�`xVڝ���.e�o}�>��=z?I�ךu�H�/��[41(�3yx�۽��Jm: ��[��9qDH�A�R�KdKL�CMA�U����eB�7����a���п�n>�O�(�����ۃ~�!�V�]�^�҄���9��&Ա=�G���`��˲���T��D�����<�@ov6ݥV����+���� ���U��"B�;d���Ii���Tv�/Ds�w��~u�a�\�2卽��!x���z����o����a9V�ETB����aG�%���b�ea#)�����A �Y�o愥א]5�M�S{+{eU{px���"����{M��((+�H�{�C�^�e�\�L�:��:�{����SS ��[�EV���~"�1��b��/29w6=i�HK6�n_�Z�'���4�fz��@5��2�w�ξI�4�Ut����Cc�N$�����V¤����,	CQ�z�C�� y���������Fq�������MqOǍ����K�`�/�Fg���q�
f%OF�p݌�IwZ����1�u���'9�e/�\C2��i
s��[�z.�V��.&5�����-�8=�O��MkYUtqkQK��9T�b
�>@�-�?j`��%!V ��g��#�kr쿨	�ł�`��뫧1��$����uRK��)���Va��C��؁�
�IOvx��Ӫ��ͤΦ�ƌ���D�l���@��v�����5�R��_��&X������'��kߎ|sKT�/�r�P`�l���_���S�js��8E��i�r0s_������+�6,�'vt/?�}��\ -D��\�$[�qG��gA.F}n�O�ByA�����}���Ԣ(Ą�h�kyy����eR׀�ɋ]ȿ'��fQ��b��}���;�%���Co�uu��~#,������y�>Te���"y�O�`��`l[�����NO��c�Ú��6>R�	�A@��n�C����ݩҌ�P@����!�tKI��{�?�V�s]۳�����y�}�#�8���������w�iG�����m7�x�`D�q��n>�	�袳Eʉ���o��]9���v]O�{�����ǧ�
�N�2��.`F��_ ����X1d�T����zH^yV<�FdڕG_C%��S8*xEkkf��7�l��n����s�{ւ��ȁ������ �As���O�j�p�77B��_�:�?��F��'��ݮ�&�Rl��`�UHz���CRSc�.#$jp�q4�C쓇Q(?��	��� uctv�����y���fm�ϳ!?P\	��o��0��I���}����#�e���M{��q��e�Y�*2�kN/b��W?Z��j=^"{0a��o�q�/U��>��g����'aő3hQg?��3m	yE|����i�vb��p��ԍ�ZL�xh���a/�8�w%�u��ֈ�E��Ú���H���e]�&_�2�[�G��eǿ}
^���"s�u�ݴs��!�w#J@��w�\0I���R��S��}�I
Gl��������PazQ�PQ�.�����EU�:Ë�}�d4d�,�d���ս
��]�mNM0V!l2��d~���O5��%��J��А/��Kl�D�sgsٗH��E:A�\�� ���/ts���r�j� 労xq���s��C-�P<a�|�Cژ<�aE���2�iH��N���b츉Y�-SX��ޛ�<n�,��4�~o��a�f2�wnZ�]���W�OnL�]����N���Ϸi�eyxx��ih)���gp�S+ۥ�R&�����$6��~�\��H*K��
�a�}OV��1�|]�Y�x²�k��e�G2f?(�C��b�6�K	N���$k�\�m�@0��Boe��I��IQHarV	�����s��ݟ�ִُ4�\��|�ҽ^�Lw��%*����o��ߙt����|��� ���.(��;w�N�@�
$Gh�6
q��^�i[�p5���q��O��u���䴞µ�kd���'nA��^ma�W1Ϩ;c	�7����a��z�9(-�X]K|���/*��<�2�+7T�d��Gc�h�,�ZPH֖����W�v��UD����YB~&�>���3�r���8G|4��=G���)�./��.�0��/�ߓu�d? �|�ݽ���:�S�F�v���1������`�)��O��J$���($���=l�S.a˄��1�*�Y�G��&=�ѱB���ރ�m#}�{c���}r����5hq�v7��;�P;�Q�>�������T�-��cODy���r���_�/���aI�P���qL"�j�Gn@GK$P[�F�vj#������P:ٱ䤇}c��;�,jË�q�����ɖ���
ΆQ�-��nG�F��MW�P�B����;I��Cf1���!�p�]�,L�\��-K�<+C��!p�XP��\�]i��\�I��R�5ȟH��rt3���w6=IS��r:�_f���yW�LiPWY+6�d�9;��44�}<^�Ryuf���ջy�߶i�c��z��%	�@h��ϛ�>Uodn��rA��2o0���["0�q��8{�n����f/��f������i���z�ϻ���Ƴ�������N�蹌�xz6h4��'�@Է���~�Ǎ�D�d3\�Wԕ&�H)�9�R2��t��W<&Q�0�=D�?}��ظ��8LCvO�5�6���QZAx�j���L��Eo�K�rLcurf�T�@/�2�(2#?(M{�=rd#%��>�� �%�}�fGR���i1��,<�a��;g�B���S���E�C�#p����eOޏ�5+Y	�Ls4�~����X�{ 3節}B��(�Lx��|��(>v�񥕹�h�I�ye����v�-�yK���8�*�R �ӓ^����ȴ�@l�U�l�����>C�ۣc�;ͤ�ow���KE%�Wh�6����0�Xx786�	�p%
_ܷ���#4���S�F� �L5�^W�/���ޱ%���˥/z����g�v����<Ae����<���,-F����{���Cb�m�P�ɖW�v�:k�`����UKx�CG����E�y��yթ��`�%��?���=N�h5���яJ����(Ď�PZ��������s�ۭ"���σk�Z�h�vx�!�7�s��7N��g�p�)�9{��o�H4�8������R������Ͼ��q�[�;����7�XrP�a��<
P'U�hɰ�S�ۆ�,-��t��'c�f�f'K�{�r��E�{F!���0g������2�%�:��=ӭT:�߰a�B����?ªk����vw��k�$�N������}Qj�Æ=y��`�R\R�L̈Oω>��~���LWkg�`k!mw!kɀz��قhA��gF�|ڂU���d�"�X�$}T�v�2�n�D������t���8:%���Q|��G�^H�ѵ�j���p��C�Y�/k�n�(T��&���v�fe@wz���΅-@"��`˼~���`ˋ#i<Г�>G%B�u�>bi���Z����ؗ6uw����yD^t+C�b�焌�Ϻ��"��#9-�Fl��Vٞ�O=���b�9՟Y@���mm[��yI���:<r\.̰�`y!�p�g�Sv%����A:����p�T�έlI��WU ���W o�"DYd6�9�z�9�#z#���%&��$�R�	h!aX��C��w�3���9D+�`qK{�'VF&��;����2VP�=�{M��^e-���=�ZvF3j'~�qw¥�����l �ZQ1��f����`^����RB��+�B����@A���FHT�Ƃ��2I���u���=�%9�Y��8��Lr~�(�#�B���$���#�6���F����n�M����N�'	�_s����g���-B���񺉴��ף���o��(���'Ê���q�i�l��HJ}����Հe#[���ˬ���} �@������w�I�`Gz{�����198m��K�_=�:���+T�l�y���R�����f�'�M!�*m)��Q����y�`)�dF��M�JL�ŏ�&<�(����F����S��k�$��u&��1�S9��e�r��{y:I��/߶�rpK��*o3Q�/,�P�X�>8W�W�矊�=�1w�rX�kS�.�i���u�ɚP�gO���:��|F:u��-�1��-�y0�	А��M�O����ڰd�\O�z����Nh��0E��P^Y\�l{�{ʫF�<-ds� �pi)�*�Ќ�O�lZ�:9�]��0�ߏ�o
��\Rkq{A�\��&-ƭc
؈�=��ʦ���#5x� ��9�il�s��p��W!/X����{�g����p�T����2K8��#|0�ߵ�ʯ�K�#�@6e񊵬�������Hc}�ő���9�A���� ���Jy�{N`�H���)Ⱥ����y��نYrdP˿8C<c>	�p���e�+�Pr���}q]�;�{ߣ���l�k�)��N�n1ֈ!���c�5U��'\:���p[�]�lk �;
�6�26��u�N.��W��ew}W����B�.�F�Fਅ��O���Y_�n^�#R�e�7�T#p=4?vV�xK�?�*�owe-���ԫ,}�l@�%�Ka���<�zL�W�UN��x�e�mQ������GK��^,�n�<������>K+�&��+w�D4�/O(�t�ڛ�LnՅ{�}�Fu���:G�[��3�g�t=�z:j��=�+<����x1��W���Y�@�� ��q�Ǝ�c"���>,���<��E�VEsX�j������,c@�!qo��>�t��o��vp�0f�6){������.�u�T�OkwN/tl����˟��t��A��_v
��_�շn?��E]�͢u�%7��4~"�*fzMm�M<C�1G��E�/- Ր^���X�a��jĬ�A��T?Szʜ�3,��c�Ьc=Y�RnVQZ�7� �Q�N;k��-�俽��Ȅ���7�b�=ȃ��p{�� �Cײ���/8�� |�ܛ ��a���L��\�o�:��r�G:��HC������?�~��T�z�]2��5�a�"��ܸҞ:�rʸƃ���W��W�1�����K����1(Pr��%�^�N�������/Uvxln7��1��5D#/��74}O�r��є�y8�߂K��[����e�H�۠��X�1��8�Yp��a2w��'P Y��!9[8�%�:�K�j�?��hy=|%�#���@�!�dTqfZ��{)P���pc)���^���|���a��uI
3|������-��/M�d��q�'Jd�V��:�|01k=مd[��?�Ҷpټ�5�@��p���B{j����rn��M���7H��}���o���t���ﾦ�߈LYn�ی�mZ� gf$~��3x���@e�P��kM��7�46zux+I	�W������x���r�����6I����g�
-zި�}��O e��6���{��,9�FA�S�/i��.�E-OЕ����)��բ���6Y�D��$�M��Y��g�U�z&y�7�g��P2N0���	�����VS�P3������?����!���QrM�tp+�6.�W�

+�o��	Y q%a���y�!���kI%�*i;",��م^ak��� �'H:�~#�B)x����8c2��&}C\B����*<\�b�ˉ(5��i(5:��	F�w���*�"2��"��!tLJ8�&��)���������(�߃x��f����K�S�K��?����n�Ap,
��]^���of9�Q���a�76�Q��G�:F���L�`�f�)A��ph�3JN�L�#������~���/әI��Œ	��I%7w#ZH�lh�l�s�O��Op����&�b��f �bqK,�qH2�_3L�P>����<����`ϰݳU\�Z�ԅ��<QՆ%���N�+�M�k�@O�ƚ���d�3��Qʫ���kѤQXg��=��H�b>�y��\����<��gN;���[ˠ�~�8�K��A��z:w�яZ=/��9\G���>�e0뵻qS�>]���?���ƴY�d��&���_# @v[�r���_q�I��"Z��:��ۜ�(��|���pМ��[R�c�8f�5���eW*�%�`��
����z��.���j�U_8�o������j�=��,}Ei:G��7Uo�bSRi��Ź�G1�|�����E})�����6D
s_L�܏GttΞ�9��7X���a2m	��m����l����V�˹���2���t֋�[TH<d�IC����т!�Ni�0dn:�-	�G��8�����g�5����t� �0��c?��.��ę~��9�o�_t���9�q/peJ�d:g��&t2ɰ��̅���٫�����oA:��87	<"����fDS5�l�f5|�B �f]ۀ�l��%��Y�?�vK�z��j��<����{�ٽ�]��;��N�����΋�󮝍2��Q�Q=D�uu�&I~�)��@�[���_�z���F���}噣�VD�A��Wg�P;}�-���
d!y��`cI��3i�J�QQz���>�����l=Ž&��dIC�r���e����6e�PgQO���j���N�T�����K���)"..��+�1�f8ǥ)�ΗQk�NQ)}���[��B�*�2J�($�Dg�sc�음^��|�v!���cR���v6t��eQ
����H�@�P2�s�2���������|�}�}�	�ۇgt������7@8�Py%��"�	��ͷA"ۺj{��.����f@y-��a�sڔ�����0�@VԉH):���߅�;�M8啝$��V�䆫�Rdx��S���@ K#ce@ȅ���@yر���P��d�wΥ��5�t��J$p�a�X�B+�ɏ�aH/��!��ȗ��!����υt������XU� M��k^)]�Dj*h'��!�{�8 K=�-�"�Ҽ���9��1p8�5�J�ci�/��;��P7!*:I�4�X�'d6�!t��qt�ؑ��k��i�y�ٕB��?Ռ��L!PNf�׶m�4y�%��h`��6�㳆��}� ��u��,oF9�yO����:��10�|��K.�)h~hFH��{.�0��A��k�O�[�˟���S�07�����~���%�A֨�b7�%����,p�F*��3���o��kx����U(<�V�����i�o2�A���E��*!H��9�Z1V���./�R�2ܢb���;�ۋ�f��ÿ��ʡ3�o��z-�q��C�dy��O�z	�5�V��]����a�C�j�j[���:p]�䭥3|o�0js �������@p�� 7�$��;��Im�۬"/��6�W��+�R���+����bw0x�1�x�!��m��P� ҏ���i�*�m��d̪8[�SQ���=�π�w[:�}�K*Wv��;d�z\*��V��^�Q:WwȾDx�!���������\����߼��;�z��������e��_/����k��y�4�]�je�,l��l&~�#=RݭK��o1tZ�`�����oO.R�*N��[�N5�x�=�op���h�N������fB:I0����2���?t����B�gEQ�1������&�,��H),C�7�Ml!K��#�𱈖UxL�!||' ��C�/�����|dMu�&�pHe�l3���́��|ku�W]�߮?��ܾ���V�=;{4��;	1�e㉙T>%n�yg=�N:�HV�G����N����ٖ*��9���b�_��s��Ck��i��'�fdg����,�+��j{�-�0��IoG���$�*_՘H�G�q�˺�˥�M:�'�֜�IN��N`��'��t�2���2����n�˲�&�e�f�( �i��Z�#��@)K�R!>7�q0��4G�YN=G�����3�A��D��?폚�.�O�㠱��R��,�4.�㞛���C��&�<a�I,���t V�q_�T�;:��u����<��b�90�-�%|�9¯��x~�R}��q@ԃ�d$��U?�I���r�B��+�F��"��q0�"��F��?��V�)z{�W(#�e6�*I-I����b����џ^Q�˵�N�6��qÂ�e ��Hdܿ����}�:D����!ط"m��a���O�6Q:����+�W��F!9BQ<8��/�:+1G���6̤�zOZ%�^l�[)��G2O����S������e���h ���InјѐDa���ߏ��[^��������5Utcd��ӄ�zӋS���+Y}[�p��,��^���b7������-�]�j�!?������W�y�ዖ��ł�
�1��f�<L��5�RT�I���2�G�Jð�UK���-؅U������n�40�p,�
��"Px�Nݨh�������V���I����l��zq���V���,���_��ɱ��ɉ_�����P�נ�X2c�%r2@�kF�OwH�ƕ1��Rld��x��ί�.�<�%5�,��:�6,�B=�>�.�S��<b��5�.)!$�ٕ�ߩǧc�2�{������&���|H�	�֢2�NnK�bʥ�&AZ��J�Qpfh����'A"�l{��0g�&��|�o���,,�@�a��Ӣ��O��4Z�mc� K�<�r�npr��7E���R�k����,�¿�ʤ�t@a=i���D}%4�ص6Cʊs$���
�//�}�k�w��.�x�������*.�|Af���n	��_Zn�l�t糞��<��챉;&���eq@�%\u���ph����E�sLd���J�Ϊ�l��N���i@��D��?�j���n��S����ʱ{��'۱���u��4j���n���P�/���p_��v���iXh�U[�%Y)&�t�������NB
"+{ء�QM<s�w��
���l:�m����vΕ��./���44�/h������^m�Ł�(��<�����>����`Hc�>�|.
|�Lz��m?H�|�Fc�f.����:�xnr=��7t����翡"g�(fAA�.l3��`��gn�`Nr|�)"���"2�߮�S���8z�~�,���wJ��ls&*<eb���h،�yU����z�qsh�W����T�
s�x��x%V��w����/_n�s��r�V��	\�?��> s���<�y\^z]zc�%�Y#F���zi+L�"$.A��w�A"��{�.Ǔ?�b��/8�j���z��0X�f��d�Xuڐ 6��h�9N&��M���B��w�����&~���$$����ʰ4���
��^2��q�,�a-�x���c�a�U�dn^1�1��Ջ<�$��'�0^�0�nF�q�	X=�K�"N��%IaGbf�k�d.�^U�x|����
�W���l$/9��7��S�A_fZ��>`��A��'G�Ͱ I�⍥��)�lʏ��Ay>I����8�i��W�}��֦�^���ϻ���U����7�}1N�f᢮�������|P z��̦xF�j�᜚�Ȯ��th%�3�8ʑ��c��z	/W�C�{GC�@�ɕ�8w1p�#L��^���6�u�bP�Ţ�Z
��H_̇�i��@��vsDs~�˔@2*0��U�3	�~.�^���d�\,��/6�{��ꚸygՈ��w���᪽.�1!NdٝhCe����{K�ˮ�ugy�>��H������#y���؅����|ׯ�������ɉ�
M3)I�5xH�������0Ț��~�=O���$	��6к � ����n��^����w�q�L��(�� �P���t�k�N���bfܖ�k�tϰ��L҈�;0G>��lkV�X�r}j4�,��uT��c�b�	G�D�u����$�>uԆ��]`6>*�x��t��6����{��w������H$CIK=�a'���[͵��Z'�:�^������}Ǘ2Q��X?lO,j������,�7�m�\�y؏�@��Y}siCK�����"_*��Z�	\'�3~��h�Y1���©bw��$�Hu+�e�||?��&�d��a�)�~yI��F����=z~�]�O�>kԙB۞�c�J�~C�VB,Wi��!6�"�* ��s�89u���im �s^%r���J&�\n��W�:&��e��ӂ W(�
r��s�ɭ~�0��0qs}��d�+FWS\������������ύ���zх�=��l|6��md�I�OT�N'�����N��~G��v������ɧ�2Wi����\(%G����kw����8�M/K���}\ט��/��l0�pe�7�v�Vкwy��VyΗ���T���Y~$�UZ�d��c����Tѧ��.֮J��碂��@O||��+��Q�Ԡd�8�nv����Dou��\�)��;F&P���K�Hѐ�ub&�bϬ=�b�@��H7"z+7>g �$%�稐��t��ƀn3���x��"{���OoJ��Vq)�i��%��k�`�Nue?��5���G�C��������k$�#L ���L�^᧚��싔���j	g˲;%���n���uסa"<(4C�
d-@ڦ��L"�rG�;��+C�8���6x��~�:I?���ご�fR`]7��Q��w�%���/FP��JZ2� �9p�GGe�a�kRD�,�&)-C���ߩZ�e�Ѧ�t�|��)�n��*����+��\
�Vco�5~P�:�kDWn��-<��=d�I�R,�j�|����<]��E��<�D���21;:k+�'�	h��Jr(c�{Q���8��=��C�'�a0?�A8g��j��%q�;��+`�^�����}ғ,K����|��f
��
WId�� 3�X:
�<n�\n�?�hl��_>�MD�y�涳���R�	��QB;[� ;cA�y�)�`H��ڭ~�5���� <ݧ�vg|�w���͔N��u����E��Q>����Y��匹tx���Ȃ!5[lp�]�<����c�T�� *�[4e���V��%$�NvH���Q ��
�-��V��-�`����>�c�B�pN9�ӆ�A |��8�'��Gq9������u�g��%��8ּ�U���4�xpf�����)ð�r�d��a�+u�h�_���h݆�J��i��9�`��l���f-U������ �����7w" 5K�ɤA�ŏ\j��{S���yAd��5��3Ǐ½�k��ă�dC����]炙���9��I�S$j.}h1�o�Cu�:\0);��L0���:iC؋��stՀ���
��(2�V���s��˶�Æ��J����B}�e����D:C2>o[�)3�0�|"4b16�:���pw���Rc���&鈭L��Fp�kK����{L��<�rm��QR��� ��v9yM$�D�����Du�(�(��U����O�۴�/�܊����Bk�Gu9a�L{=�)A>Uך�p>��Q�9��$�&�藋c`�A:g����8+��Ap%��@0�1�Y�u�H�qu�d3��EC���HMҁ�������L��B���6�>��V����&��;j��\o�Ӓx]����z�:�
�^�Sp�W;�\xx߸�&�����c_9��`��i���k��ch������d��a W/ъ�,�0C\��,�S�j�����a��M�yv�9�2>�^܇�
�G8O��XF��Ǵ�(p����i�x����~e�9~�����ZY�#�N����x&�pr�h;�E��C�ZU�+R��<x�}B|�-Xv�3栌���]��Cц:��C�)��C�%�DN|&����`V��9t�FL�i�m�^�V�u�Sفӈ4D3�Ĕ]^A	��ܒx�+y��	�mV��jT1�?@���֔���̱e��o�Ƌ���H6�룶-GhK��u�,&�2�x'EͰ�2O^~�o�[���� {"z"���@��ɩ4L��{� �f����>WA�#�+�TK��7��/*y�����|�_��k�= �T֫7��l~����o��2(&��&S
��c�YT���c�9qF�ZHT�\�.*W���i�G�YVj#T]���7�-|����N��8<� Cސ\��[XT�/��kk��zW�jX���W����?H^�vww�����kW\�@�DBW8�'W��>� ��aq���힤!�@�J�m5�8��%E�>�
4�Y_�i|����?&�ߘ����V���jd��u������vV�����J1y�)�:�0��Z<�qW��Yf��y����K�	]����~�E\��daQ���}���
p�Z���٠/T���h�CM�ႇ��Q��r��X�}������ݚ�ԓ~���cb�C����!�U��_6I���W���1�F�vҎ
�	�ֿ���o�'�B�M����CG���J(�Xa||�<2����I��8����J��l��OT��z%����Ӛ�x����>xX5��|�ò�{ Owt��/}aΞ-�>	X�h��E�u�3�������~�V�mүl�#��6����'p�+����٫�0�^1���i�%VS��CPDF�ʳ�ZV�����@�Gi�&��L&c��-�d��>+"l.���f��E�DR�˞$����T��|�/������*�
�؛�|C��f�V.'w�/�G���@͐����shp��)�m_x�\T�ۯ��vԤ�ށU�ȗ�ť�&?���R�+s�V�m����	���UNk���5_����}&j��y�V|*����@�O|G�D�+��3B�IӹBq�*q�:֯�$�>�����xN�;�s�����R�Gy"|�90�þ���׈��)�Ő%���9HT��ׯ�W�n�G�2k�{�~;
�s��ڑ������5���&+QV�Q�2+|U��t,+W�Y!?�㭟�@�}�:6�S�/�h�MsS.�/��|��s���X�L�_��[A��$ ~�؏ qr���>Ֆ߃|����G'�9�k��i%7��:��x�$�ګ�" �� 
�Xb�8,=:Ow<?Ü���~�k��tH�ɗ��=-����Q�5D�f*We�P��]N~��
y�SzM޲t�C|sɅ1²�Љ��mopR( 3T�)m��4�j&�S�OT����	A��9ű9ú�{^����']=�h��ӡ��|�y�6���$��J.irOc���f�a�$��h��`����@ߔ�6iH$�1�|%`Z�97$����s����.t�e��h�DB��i^,ͧ�.�����Â9q!ò�n�޿��G5k>}��2(THl۞��3+��_��������q�4;��j���k���B�x���NM�W�o7s<<<�N�1��TU�U��-��8��E�V�ђ�n�m	!��+�,�FG&0�Oѿ�h�̣#�
�_�?{ag�xXN.Aj��6�~{�F�c)*�$�<u�����H`B�.,l�������?,kBk�~�Z��؁N3�3Q �����ڂ3Ua&_�����*�j�վ:�ɖB�Nu�t�p�w�'���g�3�.���-ξw����g�(v}՜'��~q�0�o�.0F�x_߇�.�""�/��zZ��h=uZ�v�/>e��;�i��?�]�}�o�|ս��OzX������>u�6+-;��ۊ���H�*Yau6�o����5<����@lL�s�ύ��y�|s�SE��tKU~8�krx>��Nҭ¬�#�P���r.�kW�
�-���r�?�#2 c8�wf��-�tCL�Ш X�2r]�Ep˚X)!�N��m/�cC�/20�]%P��'�(�C<A�W�fӌ�j!�gJ@!4���� T��#�S�p6]Ls�m���\�q ���Q� C:��Ga�������;r� ��́r�X��Y �W�!fO���
4Y%T�a�)f"��B��2�B
�,a&�P(�-|��	�"��X!�	���qvʟl�2�������!��� 2晛_��'����������s���è��h��8�T�b}�9��?����R@�`5�@��-��m�R�:f�4� ��k!�xF�S����j���td�:#��m������N����N������Ռ���r38���xM��tnP��[���D�ک7ҍu3�(�d�L ���hB����]���i#�C0&�s[�Gh�!L�7y��'NE�W'��-�/����)�:�&�ͮ��� ~MӀ_wֽ��}�|l���{ѽJ�]Jc1Xg(�u�XE�b��m�n�������A"�&%�D]���;2���2f��eDc�8��#K���9�LR����MQ {��6w"�K�9X�륊c��j0�S��շ��=��� ��]1`�L����I}��bQ�^Q�^ѹ�;��
UXr���:S��l�Gj�8cѱ���v%�o�b��e�{�/�;IsoOuX O��HDt-+{�����[��]��Wk�<��rq����2�,.��ahf�Z����.k�'v`DU��Z���f�.�0m5_D9'$��Ě ��D<[Bpڪ$�~e8��T��V����dpF3y�yCj�$d����YD{o*���u6�by�ߊ�ퟰ6+Z�E��`��&ȼ�Ԯ��o*?�ùtH�8���G�>t��wO�<�Ի�!:����hp���ży���NL��1���8l���X���~#�%��z�{�%��r�ϒ]��z�фђ��uQ�s���ψEʟ#��ǧ�G��㟟<9;�;9�u�M���F7��[J�5�
�9���=���Dg�v���VQ�m���	�P�/eZ/��\6�s7��z�V�?�mc�2���I��S�G�q��.g���˸���?"s�|ߙ����XL|�i�[��ܱ��թׯ$g�_V�0�	�)���i=t'm� �F�'Yzt��Lԭ8�Y�L�]�|
y�f�I���9U�d���l3΃.��Ʊ���a���i��9Jk���	�b�"�D�,R�l�������n�ڤ����ZdH��c��� �7B&>f|�`��~�w�Ļ��J{�el�N��#\Wu}�����/��� �S4@�H�|��hɱ�f�5d[�����6���k���n8��R�Q`2rǵ��H��n�[�j��A-	�l��L�wz6�}�����Z��z;CV5�E�����˥~�M�K�����ͦ��E8�޹^�SZ�%��3�T�wz�)�k�I��^LT������}�-T}m�`{��W����з�����QF�9��~[,�
�Q��w�x�K�����	\$6.w���q�;j0�$�Ԫ��}\�W!8쏢eK|
��<��m/��7����G���X&@�k�S��i�}e�9�+�P���Q����ɯo�>��Ի'E-����/�`��9�嵻\@�����,tƎ�璠Ȕƴ���۔�t�(�e���"�ǐw� �X�v��x��Q�W&p5����cM}.#;h����u)���{ڠ=�o�闷�����Q-w7�(�5�%��Ns��a��������k����ݍ�g��7���7��~��Ô����z�>5�V�j"�_�8�>��������?��lT�cfP��^@vlU�K*��0؆2x��9�"����Ơ�Br��?پ{yΑ���������'�J]�>a�J��e#���a���F�O7����2�A!�AJj�<q��\�4��@\Nf >��!lqe�m,a��F�r�����\��}l��~����x�S�TFb�Qn��Y�~���SH��_iZ�XO���B%���#�:l�Z�ț	m�Wʕ��L*�����W�1%�{�s�v��r�
U;Y�2B�+��t;q��C{NĵD�]_�g�[N[@cCPG;]�r^�*a�(!Hɤ8;�v��{xEI�w����b�y��Y$�3=a����l�ӫ�i�iШ�IC�ɴ�'
@L�^X�͔� �Vo��i�������b,�.B�	<�M�lJa,�IL�D.��`m84�)�!Yi�I���#��g@��C�;g�����W��jB8O�M�e�͛��?�4j��j�0����VR�G �`|Z饪J�t=�(�&ه"��I�G2}p�g���,�C��O�9��������T�T}�I:�|�a�0�!ك�FS���z��nc�8�������%�!"xx�_6��W.�j��K���φI�r�u���y��4'�b��^V�����$�Lr�m?j���MF㬨���s����fuR��s-]���o�:�V���/8��'j���v�)���˅��y���l�q�S놏7d���T$��ؽ[�E*�L�[M ��z��Q��1�0���L~r��h{k}YE?=?%Ϭ��T�uԿhkg�OeNy0�:�下�ڋ�Z�����ŗ��^��i���Ү;�Z�� ��ŕZ�DNZ�\�	��ݗ��X%�Fb�߉V���j��xp�";ݶ��S�яb-�%�-���6�Р��_���[���X�k���X�84B��c���<%`� c_��3x�g(+&�D=��l���O�C�jx�Xm�j-�������k|�2��;J�ѐ�ف����T�y���,A	�����i:�g�YCI�}�:���)q��'��d�VOPʏ�K��6������R%2"��
��>��(!Ş:�PH�Y|�2�����*��YM/��AK�������zϙi�_b�;���o^��\"$��â{c���*���v*Y��0Z����۠C�������^�@d�ƃ�ޗ��l�A�!��N�5�A�8���Yke�3��j��[4�
� ����^Q
����l���5/Ϝ!��E�3J~nq���!�R�wF>�q�SG�?hc�[���4�5XvYg��;�f������(�'�剁�����p��!�J�5{�����98z���e���!+	�_H�'�An|������x���qz*�:��^+�n�}-KdA���F�Pߴ/X��u�X�RΒ/!毢�ښ"(��>E��K�#>�$�x$}�OG<�G;X�H�΢�|JԤ ��Z=gq�I���B�ί�/8���דң��G��j.d4�

�>KDη>�� �"�����*�{��a$B�N�,�}����j��a������Y�\x��T́0>U#�f3��.��4����_�����ݯޟ�ތ��L�]��l�q�����~k6��
�0^z�?D}u\�o�7�)]�Gw3�ި��1@$%�{tF��H��� 	��[��<��}���ǽ�^����\%>��2��R�pIkZ����%RִUFV�q�|r�~&�3��,�Zv�\�CSgA�'x�H~��ZϨ�E-����av�(Y�)gQ�a�L]О��ݿ�M)�\�����#����qk����*x�B�> (�ɭK��=hC;�rl�>��E�)����֠Χ�b@ξ?�=f�hD�G�����d�ۛ+�!��Ll��,�Pd'�.4I���O-ZD>z��j|>Y���`4��GV�R)�C�U#7/D�i�T�p�#4��^ \F��b���0�ߨ���i����o�nrzp�G;�-�
����^`��!����"^��Z���p$�:0���c�]�QA�0�{o̎ˋm�J��
%�|�o7�~Wũ'���*$���A�SI*��-���<�NM�syC���CMU+��wclkd�oP6q��p,��J���s��.���4���\����}2m�^����aʩ �N�͌�̢ۢ*.�!1���㉁�+�6~��sP�{)E
#���ZK�����r�W��3ɖ��r�4�,�h2�_}q6V1�_�z?P�2D((U)�T	�Dc��@3���H��s0Lg&�+�K��Q����p����C�������/nS<��ԏk�<��5�}�V���Z��	�	�@3���!ԭVH%5��cg�>E�E)�F���i7��)4����~C%����/��	��ԛW2Sʃ��A����k��o� ���]B& 77x-����ƪ��ⷀ�I�RI�o95<3�9	��A���4�]��9��A��~�K��{fпP�Q͐=}��궰��l���5-��Q��;�:�ymq �7w�"�J\��#4��ۛ|����#�:�!A��ud.P�� ��(M��jT��D��� p����"�<�Q�
O'9�t��d|c=�_E~{�Ĭi��9�
�#�I�\�Uq�Ղ����ѹ��L�;vw����04�-����ot1@��f8��;|�����=Jc���+H܉+�Lv=����t��ϩaj�[jG�~���Y�쮭��0���l��{KB�"Ke���#���S�.U�k�[��b*\���������7�!pl[)�M��TH&�<DɁ�]BQ�@��XV�-�9	����p�\��r��V�GFW7����u.^e����ѽ�t��oz8ȭ�
/N��u:4��0����#|���v\�~a�Yu�XN��J�M��r����py)�A���s4��{����Yq�k������cGh1z���;��4�ķ}2|b�R'Ƿ�y�����Ri�U���U�q"�+�C�2LS��Ժ�)nQ��Ǡ%�V±���Jl�8\����}̇6P����W�Ƃ�����IA��ɫ��''�-��� �V�Q��A�h̰��+p��<�?��wI=�	X��r
�lNj�1{J;�7��[}���C��Ͼ�߰׿��cVo`��w��߭{��=�x8?}�0�x� �x5U�p}R!2���~aܹ�o��<&�#0�N 6m�U�I](�׹n���Ͱ� l��E���wω�հ�'��v��l�<��@ǖ *�;��W]�G��Kg�ag��yf��*�Dq����FFĸ ��\�1c���N�c�wUTTCH�$Ȁ�`�Hu�<	;<;6�YN36���U�Ui�����g�߇(i�q����aR.�%1F~���D�ȁU�ٝ�ǲIzm���N��b�X�o�?����;�n���e~�m��x�h���ھ��_�Tv&��6
QkK �)�@s���Z奥 px���02�i�Q?=��|~�{>��vV&���0�@��qpK@�8�!lAU��d�q�:����Dۑ�O5%$NT���`�bs�u��N��8�!��4�E}2-3k���1�7�5�zw{�v�;��n�]k���`�~��+˶=֏|��n%���!�gM��9o}�s�n�b-�yנ�F:m$�C��J-fA�2�Q�mEWLM�G7�A�8�f�,����NAg<��ԵZ��ԡ%v�� �`;VQ��	�}���c"�iql�@C/��G�bW�vXs�Cەf� �"M3���������\ *jse6*[SEe6������h��o��|�r�8MkO��ZU����9�9� #�A����><f�T5@�.���<��C�T���I���U��QP����������-`f��􊔇���+sm�e��eҩ)��e�i�8�`>�hx�,m�H�s$�6��31!�xdH����6C����Z,��hҘ�\�{h�8�De
���v$���tk�!�g� hoė�\��;;g���N�:�P��A��#R��5)�3d?�!��G�ђ�A���`��+�����˃Ct;0���_yb�Ku��-x�]�	8��٤��Z� ��!$/R�_�b�M���j�n	)�=�5y�|��*6lVe�X�d�N$]�P� _Tϑh��ŀᬕp�F�%�<=�x���x܎[�����l��^��ۺ ����$�����:�tzi��C�6�,�h;�-^�b��ڙB�y����;�܀V���l�T�C�¼a��~�+���Y]E5���M|��:�(?2ap50���
�h���@��b���'�'iRPPh��\_]x��+c'��nk?hn~{H���>|$����W��q213�h��}�B�	<�-����/�柅��*Ԥ�!!�w� �f���Q������~j�if��������`V�&�!�E����4��k
�`]��_�0��?�@pQ���,JW@��뇞`׃D�5�����Kc�+)q9�UCh�f�.�?(��m�@w��zr`�g�B�nE���K�������<fQT�C�2�����/aޑo�ъ��e�ZC�;���غ��~�>|{h�|��x���g=�n���v~���g� �րR��R!���`���)N�C"��W�
�-3��&�R�C�F@S:^�~8�K��ƯQ��+�+G�^1�p��E���F�'|�"�<��r�1;�|X$��L2_f�I����?�/����(6ֶ)�ێ��昡�ez��-\�w\n���ƒ@��Rє�s�s4Ї��~��������M)N= 3�0�:*w��$�$����
�����\f�"Cn��s ���k�������7;�\?�2+Di���M#W�k©*a�,�;%Vw,{�=�Qҥ=ɕա�F�hR���d����﯐V�`tQ �4+8n���^6"zxe�2;	D8�������_)��HE�N�J��m^Ӯ���d���T��U��8�1t[UX�|0��7E�V����O�����gi������o9�'}(����K8�p"@�ÙY�#J虾�^9����JV�VSd��[��-�?	��'��Zd����Z"��Ϡ�����
d�`�"���
ȵ��YD�Yڲ�ܥq���/3�!ŕ�����!���*�]M��l���K�hi���Ju�+� ����!t�p��a���H]����B|��E�嫸jP|�F9�M�[p�^��"��[ZZ��&�B�(��Y�14�g6�/5K�O�r����I/�공�LX@4zۊ�+[y[��*]���im��+�yɸ���F~��}ct]@P�r����)��N!˂I�g�I�]��z܉>���Y�X���!�n����pAN5 �1Z��Oϋ,x`�q<3�����k��-M��A����d5�'Xŷ��>����Ɔ7�WK�[���;���O��o���o쇝5R?Q^0�`	d�!�Kg�.��b
�nr��� �t��L���6�~M�-�sg�k�8��j�W�5׷G�4�]$�Y��a=��&y������1�����e���"��3.�ؑ�!�z�MY"ֽB̩�7�:c��(�ѯ��]�@�zk��)	Ȃ+�,��t���,�R�����=T�ȥ6��7��k�0t�i@�&S?��rR	tV�h�n{vZ��G�����-�m�
����2����7m��f��6R�Ƥ���g�%�ZV� ��S�½�>�U�	���D���_P��pI����n�?�������2R6�/[�6+ �I�F�(�,���0e_�5$��Aq3��󜔍J�������er�׌��������#�WQ[g ��D.��:k	�?nN�e����}����t4|�zz*C����5L�-�H��ϛ�U���>�\d��k!������6�`��hT��X�S���� �D҄FĠ��k��ɠ�LY��{P�	J5����~/|Ev�����x���_�琽�����=�2�<Z,��� ӆÌi�Ȳ"�ʘ���tj��O̺�9�V����-��~��.������T~��`�(��yDYQ~�\,�`0*SX�0`Q3�E��C�(���Ct�8	� :�T:;�����̤%���4���E�b�l�[E@9�q��b}eZ��K%��$ȡ:�$i���z��t�Z�򖮭�Ce����Q�v��Cy1��3�����1�v�oQ��<c��槚�n-:r����|@%ld�W%�M3�!�0��(^�u�����R"�|��>��t���P���K��|��h|��h�)0(d��� _ၧ@	��D���wW��̑(�t��	1a$6��;U-K͈�-h��~����5�pv���UF�_Mv�?�X@��+aj��.m �;�o7ߐ�N� H�*�����L��\RY�T4�恿"���?4�N��Eܺ�bC�pj�(\?�3�]���	�[�m��Rc&+9�#����n�K�C���c�is���Rtu/ٻxx	�ВU`*��U��ɭT	NY��o�C�:�Φl��i��l]kd��4�4;9�SL�s�PeÁ����d�g�V2@u��i�� �L^m*�y)�w�=�祩�c��J���]�dT�rm ��b�v%�'Id�`��`��e�=��߈v��v���b(,+#)ڹ=������"C3�ǒҚ�F¹�(��j���{CZ��2^,� �-��?fQ�/�����̌nJSP��Q\���.|S|SC&O��3A�RH�R�����b�?;IC�HS��t�J��[�EE�T����a �-�-!�yy�	z�AO������F�J�(b�t��U�p���~rX
�&��o��F�_2e���b7���/g�����nƷw����o��;^����+��p*w/�Pt�����D�c}���9���V��� � FU ��{�k�(ej�.�JLȇ�D�d '��Ru�(�:4+#�KC�A�%{~l��V���{S/�
�s0 �j��4�6�W���7�(��j嗋X��3�4�U�OCg#��Ji�b/{&h��U�&c}x>\�Og	�XH�����^V�m좪�Ѐ�LT-Cc��/*�rKӔC�b�S0'nBm�>Xq|Z��*����=��-n��V.�5$00���L��%���3b�RWG�>�!�k���߉{ڡ�t%��!�-2��z�z��jZb����W(��n����z���V]�3���|�+�DYq�̫��j]�P�3�C'G��~��,v0œ�����4�\H�a7ߏ�� b�v�������b;� Q�"� )JtЩ��z^�W��!(�X�����s"�2��?qw5�U-fS�'���CN�Xu]��X?��������xn�/0�vz�qa�����g	� ��K�r�VR�.��F�kt�m� Q�@N����Y���\��mm����%*`w#����f��|qs�B��<����w<ԩΜ��\�sH�����^׭>�!;�oW���%א���� Io�>Pv`z�dJ��DjP�TH&��������	E�7�5�0��|_L��X5�6	�utqR���)
so��f�U�2�RQ�G��*@�Kb��rzwr`���������=lTʅl��;D���!���3�g\��a�$�鎺?ωRx�NQ��Za?���*�KS8�t�Y9��jv��@Iw?���n?@D��0��}©���)���x�M"*�dU�$_�<�:�&�VU�v�#��Ѕ��|YY"�/�~�.F�VFn�`�3��ܸ>�O��YA[W�(�<(*�mK��Z���[8h����t��[��+�pMP8�_� �Z����e��+�FBI"��wW;+K���
T�ʣ���t�P�0-��<:W����T�3�UZrw�`��V�=2cw�DV�C��FKz���O���F.t��5�r\�_���W��x����vii�ml�s��q��xvo\{�&yk	~1q0!�2^[uJV��B��wbX� �^��*Z����+�ug�.�K��TA�lpfK��e���|��ȼABK�Y3����7pri�����oY��<ѥ�fVo�,����@nY���m�Qv����,��� ��L/_�~'� I�����
eIL1pU���q�?`��Z�~������-�v�P�:5�C���[��g���Tx�Z	�FoV�[���������B�݃l>��x�����
hȮ�TlqJ,�ŉ�V�(V6��^�c!������g���Jf}� CD��P��l�F�_��ǘ�c9eٿ�
oQϏIw����r���;��07�uur �Ŗ�h5��v�� ��F�1Cm"w3��T�� ;�trS�-}�.9A��8�'Ե�]*NR��Ea,�y��Gp�J��+��p>n*�zKkw�梹�=�1�}��f=O�Mo����ǋ(5y�_�d�,7���ڶ��zZ�V8��6A��������	���N*����+$e�p�����)0�Wzv^�j�h��C�Ed
�>J*#���vܪw��:��,Y�Z*�YR
Y۱}��"8��o.���$阗f�ja��s���D�jy?��$��E�a-����D���#�&���D-�}�u��.��Ϳ�L���ח?*_~�;15l~X)�;��¥2�O���i�5���/
Ll?C��f?q�:l�.E��������I 4���c$��(��]����ދ�u��5K���������a��<�~����9t/�ca���O��吿��2������헭n�F3�_e�2Aw5}��"��y�em��G[�Ɛe3=�\�/FG��l6�9y�`��Hce�	�j+Ʊm����q��EID�t[,�y�����y�M�$�/�|��mJ!�/�hg�����)���إ�&��%s-_�o6�؄��K���dJ�/Z����h���pTz2Tv69�.�g�=�Sn�1�GFHAar�]���������ތ��]�����4jn<mj*	�V3����Ca�F��+�z#�p9ޠ�t��]R=�G(�(t��ĳJr' �k
�Z�i��hTymnu1S�E�23U��?9��Ԋ�#�:U�E���i:Hށ��r}1V�bN�kB��Fy�h**f�/t&(՝�����3	�1�Щ�94�K���R"�1�����r4E"�-/&�h'�g�)K7�2{�-p�poͥ;:�++6��p�tp5T�HT���.X1/��"<�"�-_t�Nz��H�H�[���db����G��+{O_w��Znc�B.��qr�}U�j�L�ReޖhE9���I3��}��|��Et�"ӓ,�5Vs;��<BߗS%D�(��y��,�u]�F�ϙŷ�Y�6-h���x��-���\�\3�o!�О�v��d*]� �q����URL�7c�V�W�Oh'�߱Y
I�#�L��_����r��3u9ɕc��0��l�c�8�$�� ��dƍ�dv��E��oH�3�#�� �{;�D�R�]xV���{K�{����)��)�qX�O�ð�&�������<u�8 ��{�h$=8��7���a��y5�F_���C7�&?[��Ư�V�@��xgϫ'I��L�ۻ���Sp窸i��2�������o{�����!�����c��_��GRn�D�g��20ؤ3��[�h�]�L�+�ID̻\����x��^��@	u�
��h�R����sn>"�PmJNm�|~��0[ls�)��!4	6ٱ[�0LJ��B�
J4u����Z��9���7�|��p�a�l@��/�F⬨xe�S=�]�T�-��vƛh�b)���=$3�j���]uOO<�s���AF�x=SV�U[K� GV �Dz]�/}]ݎ�[�\A��~�~�� ���Sm�>9>NLF��*>�Y#7��ߗ��A7�n��n�z�=>~��U*Xh���T�.*w_�Θ3�F
&b�8wE�C|<���7��Wu�76�4ط=\C�E�M�-w�d��|�w�t&n�v��`��S�ۿ�[�7�B���v7�5�:��P�؅N�s ��S\j����k�'�6?�llA:I��P3��vBS��:�N�?_��Y��"�Co����z��>�?ܚ���8���5���}��a0����Rk�/�g�Ss8�Vo�y$�,�,��X&e�c6E���>�
a�L5\r���8`�!xLH/� �D!q��/*.6���r�����T�Ù^a�v��%�@|K@�Qؒd-|��J8��.rF"�t�[������%&��_���x�Χ�A[����')��+��ۺj
��ű
���09;�z~���n�Y��(������ݼ�\��S���糍�����ۻ�}x��ʧ��O�_|)��xx,��{z,z����V
�����=�h��	����ڷ� ��>+x�"��l.��n��v�VTxF]ߕ��i��Yrm�7е��v"�����$�a�0�I���l� H/���+g��F�5��f��C�Y6Hn�&���2�2$�yF�s��_��V���.����O�^�*�9`�����)��|�Y-�XJ����u�d���hZ��!�a0Z�5lU�h��3�\����08�h�5�K
�C
��so�]��U)��Q~�^=ϿTCEǕ0H�n���1�nVn2������b戜����Y��r���V
�SA�j:�:Y�<�,C(�CјAtW��;��c��Sg7�j3ֿ��*'��9Q���P�.�_ jy�;��b�2ä�W2iVܟ{|Tn3u<FT߱�ZW��E��6�&��WR�zz�~TA�h+W��U�kȮ�04�M�v��y�����5��\,����ƕ1�E�i�^����U����k��r.�'���~��Z�9�;\��-���㰐��>�b~ѳ#��\Tc|y�0�ǁIxh����˅3m @>���f� ��Kcna�HOw���D�� z���V������7ZY�*/�5/��"��]8N�: �"u7����:�E��\:�D������I���}:�B�՘H�½L�!K�R���#��3x���hB@��֪����3�0y����/_�Н9מc?�@G��|D*a�m钕��p�ϟ��7�Ai$a�.�xY�G�S�Y^�*,t�F-�^[���&�)4̊1��5�\�*Y�g��͙�~4K���Ó
�G�U���,�nG��T ahܭݛ�n�(���T�mֲ�-���Rg��L��������S~@�>[ĕ#X����~j2�{����%��1�Ǉ54��]Ht�o��׬��v��y�&����^4�Ar�`e��DA�H����"7.t���]�Q��b_>��
�!_I��Ƨ��J��E'�� �"h+�[6� �	A���\_�I{FH�'���z�/	�i��b�JJt��gN�0��r�
�yQ=�]Ի�̥�-���kѢ��������(�6��BI��^�^�r�͕�-�������H�?���C5ש�W/F�
�|˚ݴ;d�r�OF���&3��t���m��EA�7*�ٗ�c���5c0��R�|i�����n���0c�����w7��Z.t��k���8�Z!)N��H�M�WϹ����d{��@'e��0A�d�;�_��]TUZ�8�2�6�/(n���F]׋��_ok��:� �Q�y���q���J��=�2�{���x�H`����]�Rj��|EZ�;aK�N.�PFC6̅�K|��8��f���p�z��d�6�K1�)�jX�6R8z��p�����#� �b�E���H�Pǿ��!C:�N�E�L�1���&+ټ�T/f�J��B�6��5����#�����=���R��-��~등��~�*]%���sG)�R�=�p<��X��aW����� T͈&`��@�v zn{�`�2DS=9�mp�θU��I�VY��s�%+iGP6k��1.ٵ}�E����;�� =p����"pv��n�('�s�i�]9)+)D�l*��ʓ>�?�hI��0���H�u~��e['��D����Hh ��R�D�o����iG�ld�
A
՚�-���$�����^����$��ZI��C�q��-:����>z�h6�����oصDz���I�Ry����U�@������/W�k��!$�,��+�N��X�ڢ� �I�+4��Kr����޿eE=�[�ܴ�?����a��&p'Ϧ����� "�y�m:�$�q|(�v���2��/�>C	�ƹ:_"//Q\�y���aR��بI��� ���e����%���F��$!N��ۤƁ�*6��p�{�� �%��M\G��6���Ų+W�د&�ZkU2��WV��>io�]���3�����9�թ���I��7�j�G�TC(^�h�	4Ǌ�|s��JƝ}��f�N`_�}b�Ieǟ]�'�p, ��P�3%$7�;��s�qlL�;�[$A�?��a�õX]����t���B�J< /DD�a����ݴ!��Qa,����|WD��;1 ���#�Y^#�P�0s�s�e�:����s:o�b�P|�\�xx��oݥ=�<��������e���ן�S�:��c�i����o���9�r=r���O=JPʭ|3��R���_1�l�I�����OQ�*8M���-)�)秘�_;��W�\�b�D&��� �z�d�7
�Wϫ5qc��E[�Q����%���
1�.e��ʲO��5\�*�ym��&�V)�R�R���i'D�2:*�Ti4��e��Ѭ�ka9x���W�L��_��J���!ձ-.�{xw��m��#���b�'�srЇ�wh��҈ib
�kx�%��)+�)���Z�A�8��&�����~��a���o��1YP�!M�tI\�q���rhEG�W�g��|��.��2��-��.h��I���B����֙�! D�@ ���I�m�#W��8��ӕ��޶�.Y��J�9��l m
{>p�!�������m��F�s_�ĳI����;��}v��q1jn�Wq����������q�R25���R�;`qE�a�ܭ#� B���P�mcz�Ƃ�~ %*��xO�S�Y�~�﷪�_nZ7��[�of!ag�����p�0��v8_&d>�^���yf��0B���Җ�ք{�c�Q#�nO�fC�,��haߡB	����(ڐ��oh�K�FkJz�J�l-��NB��>}�/��DJQяM�(�V0�f�n�1r�5�=9������٫��������ZE%���z~�NI.R�H������"�zs��%C�xf�+��ͅ��ܼn0�4cr3rw�&����ֿ�����n��������礮�Vx;�d���@�ѯ�LU�q���R�t����dŒ�6�=��!���:��l��h��=�]�o����ۂ=�Ͼ���yܡ~�	{��_�, ����V�߬��.� d��箃[��������@� c8��Ӣ�[��gvs�K#���;q!�h�")R����P.j7���W��~Hw���cv��Q����,_�BQ�&��ю��o�p�"�Qp<����-pS:"L(� ,�h��Q{!/��@]��*�5HϴĊ��ܠ��'9�I޳I�F��GJ��\f�wG:Oo1bY&}{�)3��C��v��E!�j����r��t�'V�E'V��u���H���b�}�i8�SEs�.2%�EH�@���gv�iA����ᚴq�0��$�lpW�P��Fci͐X��n�4}�K���~�w�x�T�UI��ըV�2��g�^v��E< Hњ]3��İ�f�S�����o�'�֞:=�ν�^�Wz����,x��t��d�Y�w5�!�]y�i��[TN͆q�%;���#S�;נa�v��&}vs�)w�fk?A�=1М��>�� QbCf��w��
�3pe�9P�Ïg����>�<m��;U�:�\�����H3�S:��U�-T�&[�i�I�|& {=mu��u��������5#�XS�<�Jl�7���*z��3'�~�x�8ij��\2��C[�
��V��]ͺ�A���Nw�
w���9����]��]��]�)��v�G�G.�<~�����:[nE*��+��v�~�[rk��� �Y�_��K�9F�����	ziN�Ò�1�ro\���쥏�"y�D�q�~&������Ƙ��`_�6��+�$n!��mJZ'�j�Tݼ4�)�7���N��������ߦ���oڋ��[''`�
0yZ���hs����H}5�Aa�^@_�}*'���kbJ�-3�$*b�;��[Ba�)�lD��M�0����I�ۅ(���1���G��y��;ӣ�9�ҏ6���[���������!>?'�y���,"M(;"²���A�zD-���m����xw��K�c?��ӄ!�Ei%L"�+WB���|Y��Q���<"�Z�
���e��� ����y��_�L��Nv���?�6��nry
��ON���׋��\1�XA��/���o��B���kupqe� �t1���^+*l 9�gӑ���,��p�>v�r��� P�,��`�8�8	B=(�L1���P�f~\�%���NG����6������E�ˢ����F-��݉�F��EگF��(gp^�e��:���"Ykn89Y���$yEK��C=�������Z"(?M�!�����0��S�+���lAB���g�d����u�t������}� ہ�yﶥ�>N�i�/U$��X8qRG<ۢ���p�L%�gߌg(�6���K.�?�T՜G˔
3[��ؾ�Af�r%����k9Tڐ�a�n[�Ԥ��4�����Y:��Yc(b����V=t�#�q��	�<*1���N�>�������`�ިiɌ����4IE�Y��+�o�3���gx�����1�X!�(����������קɡg�<�����A��v��~�:R���[��+�*53���S���N��t��u3">�ޮ| �dHb`N�'a�W&d�Udd~�ݯA�`.p�fK{� �b����*bdZ���y+��IN��i��R�ؿg��b�~*�� �s�\ �	{�˟g��"�H�<��N��.�	 �Y���n�%�/�d
�U�d:�sI&�9�O�(ZB�����HW��_%��k�j@����(�mAW����e���~������xr4Z�{}��e'��K�B�sM���%���Pd>��/^v���/?���~���.�ь=p�j�����g[ҡ���ԈIN����PN;$_��k'���l��f��׀��M'�@ڬUD�[8a���^��^��<�г��cU�mZ�mX՛^֕Z�M?bS;6Sn�d��ܑ���Dj�][|�1�e=stp�-ڿz�� {e�P�(��}���������^���]w����`�n6����lC?�o��;oV]�آ�c����)c]�¤�ޤ�B4	�-�v�"�Ya����g���D�&�;�H	�9g1���Yx.iuɧt�F(�Ge+b�Y"PN�ia�啳�>[���p�Enz����W��/?J��=�i�=�U�oݶ쬶\�CO��?r{X�"z��ۺ-;?Z�t[u|��*�9`+޸����m݉�Xn�"���O���2���,z�7���/f�/7�k4��t(�	Ye���T��j�,����S�����;r�u
�db������[ ��d�j�x9��ô�P<E�p?���~""ZCl�?��Aݼ�QW��W7o�<,�{�.�S�K��[����
���u���㧔���R\��W�j���պ�2��܂�k₱�;
_q�do�\~�W�v+5�p���EyM\�/���lX�Q�:�.2���3�\�OS�tr"�����1��{;�diI7(����hi(����0��n���o^EP�Xb�<�ΥLF����F���z1��#�|�kEA�Kֿ�8�p���u�o�bԫ9֪$�v���.V�
����=.E�2�}=��FuJw�p�����F�ęF��x�x�g:p��x�|X�5�C�}��g�+�#��m	A\�^���J��F�f����~�<��(�[-��������%u��<MT�1z$(��]%f��P0a|]�%ś���R<=� e����ֿ��D�2��֤MC��W���Z�.�d��c�蹧N2�[?��fd�m��9����A��������ל�ۘ޳L�!��9�_�|M�r(��s|��b���xFE�ٷ"ϷGm�e�P�fy�sz�B������>'��'a(/ʟK��{�f�xs�,���K����U�B�Ǒ���o�6��ύ����,�3^�f=��n`r{�U���Tw���|tgr���?�<����w��]�a�;�9>��`"��3���Zo��;]�Y��a��6�׻>_?��\O�e{�����[��&�ܑ��7���H-Ѓ�#��60 �B��[,��	L���"�IRYG��ݘ���덋{��톧������?�ġ�?jNC�kĝ@����I�$����@p�(����Ȥ)���-V\*J�9-7�N����Y�H��,GK�2�0��1�&��\p�H\�ר
���L\n:���<�~/B$� pJ��C\aO����0�g|�Ry����Voy>��8��?��~�	�dLbg�{V��m�3��х=5���	?����?KM����:����(�
t�-������)\�{���s82��u?�58�������V�"7>H��M!:C�"��ޡ���#���Tpi�4�,�CB>�1n��g�UO�
;"�h�j�`M���k�ߎ�O������c?/�zU�mjG���Ƚ{w`;y]�����/u)�4��V�`��[q�I�����j���D�qF���Y�͛q����oal�o3�|Xܤ'<u�^��e����� s���,U� (����T�t���}=q�!��RO��]M�=�?���Xi�n�:�.�;�m�&P|R�u�`S�y`�'
���{�
�J5��a��n�/��X�,�R+�P�GH��Zq%� ��J{lZ.�R�z��֬ڟ2B�%h��P�jwUw�݄��qn���h�F��0�]kW��Dq�Kam^���8Գ��d�b�x��4�z�fm�o}�o�;o��ׁ��5����ny��_�E�w�~o��C�	v����/�����O4�]Č���"@S.o������d���~b(]b�"ӣ|���1�Ŷ���JOXPAq�L=�t��>�Q,\��"̕F4���=$ª(?�ĤH_:^2w�c�"�hF��6+:庒�p���Xk�]��KD����g~�ش: ^�O.�@m@�gG��֎]ҫ^<I1�I����5���9{�.�0s���o�⏑��|�젂#M6���E�{>�[<J�}�G�<���|AlĖx�B%8�}e������)c��ŐE�Ga��[�H�0�s4&�C�lD�a=�|���}��#&.�bq(�j�����KX/�L�!�M�s`aE��$& Ucn��J4�z{�p�J�`���{�"e����y3�ܸ�*������u��m�Y%��4Ƀ�cCZ�B%��Y�ڄG@ʕ������}�;z ��6)j>��T4���H�Nv������;X�ԖBdq���щԅc.�r��I�߳�\V�[���>y�����>�QŞ1-su�YK?S���L
�;(�J�qnD�]��!��,؊}X��r��K�<����"�|�b�T�#J�Ny�|��U�:��6�w+�/
9d�_\�.�p�Aژe4� ��I �d�Ϛ"��F*��J���ѻ�א6ډ�K�w�-ݼ�Z��CF:��I9~/��ƾ27�]/�g���*���[/o��[+z�I�	����g�f��A���8��/�g9��N��8x�D�)��鰻�C����'����P�*���[�����!�t�����U��!�������� 2�	��Y"ʚ��s� �H֊���qI	���qw��ss�*;]�ۯ���T�{�nx��|�e��'���u�Am~���Kq--��	)n������J�/�-�ݵ�%����C�yf��~�3��9�~6�׶_oh��xY��h�:)ex�H��|����)8��pT3أ��`��!��2��N�nb�c����a��I�����a	���SI��$�C��c�53cK�J��9/�U���Ț���GW�+GwH"�ǀ�}1Sxw�%ź�G̰�d3�����xЃY�mc�bY57��HLQ� D��\J�o�8��8�d1��qE�<�=77E��e ���~ ��E�<��3x��z;%��.�S��d���4��ﱏŽ��y� ���rq-;��a�@Z1���\��.��=�O�Q�.�����%ƞ$�F�!Ģ���&o���l_t �5�}0���d��)�`�7�$9�Z����|��͟1f�����m�+V�"� �"�2��ʟm�-���K�6,��ς&/l�'����@�
�j���ޛŷ7���}�u���;�n���[L��h��\I��	\�	{Ib�k�i�?m%'w����3�[8�E��z��q��!ϑ��yȅ�m�z�d���`�H�o'�.䒦YA`�\��r�LQ�mʲ��2c� �Ix�D�Ng�Wt�-Oy��;{����:��)���c��
 %9�W��#g�O��C���{��i��\�Z�[T��=DhRHd�F@��R��^�ٹy�^zz9���`-}0��搏=Yo���E��^��^��S�e�6��֢��u缋�t#�4�.�4�4w�����$P���W��f�V131mY��s�چ���5H�a�k�G �M��R�����K������z+��W�^�=A�Y��Ve�˳H��\3e�	�ZU\1;���qO��FOg�Ĥ?��Lq�o�%oOK���H@�-Keid��,w�MF> ��V�&g��^�h�����DiH�=��u7��K��Co��������9p?H�}Vf�[X�M�;���YVPs�ocpEo�/#�!��ɱN�O)oP��\r����nZiAQ����?3Ik����w��a�����1��e�U&�(:v)Ly܈̀E/y�ּ2�4k2X���gp�S�88-���'0���.��d�N�$K��$�@�(:(�!�~�&����P���V�ȑ	��w��Gc����MD�|� v���Ԫ�ͬc��Q�>"Ey�.R4OO�!��[��	V����D&'�i��g��,FzA���d�V�%��.�R�K���&O4a�����@����ňV�n�p�����X2@��{����������JD�����(�L�\|�z(L ۠/�#�T�Aۧ�G)���<��V����$�Çc�=|�~\L3���� )��I_��N���@���NwP��N����_1�{�GH؇5I�~��c���c�G��h���롈���R�@���W�ա-�S&T�-u7��4W����J���'+�PB8���0?\8�4��f˱�����CR�jT�� 
kf���U���lX�1l�_s?i��e�"���Dt���u$��W	p
����0��1�� ��	sA�BU��7�# ���xG	EEB���#��K_;����0�L5g�T�v|C�zw�dp�-�2%�����pp3oy6zZ����~�Ȁ=��v�;��.bʷ�j9����]$d��:��U�P��s7���Ѭ���ǺO���:�����ś�h�^~o6h;�UQb���p�A� ��u�1CSU��]U��p�2#+��@#���S��M"���B(�A̯F����s�$������I'l���"N��̡����J��������x/Z����#�O�~IXj��ʨ]�m�O�EW$qk ��l���^yޞT�9�Xi�:Z��[C�&�7�B����;���H��h��()� �t2ڙ�T�0�V�o�Q1��X��Ut�^��tL���w`�T �t&� �d��H+��}8'�.P�
�).��&Y2h�p�Ǩ����B�{�RS�5	��{�m�����V��?N��?_dG�	�@Z�����v�W��Ɩ��(n�'s��'��6}�a��c�ʓ@������%e�
����4�@� �^�Ϫ�����'��܇����ie�@�-|W:/��D��<���:"��8mo �-����{'�oF�t��Ԫ}��hʓi�&��A
�<r�U�AG&o�d��D��؈\�G$�8Vա��w�5�,0�SV��f�HiY�e���1��ݽ�HE%	$�+b���ز����/5z7n^��o%>6޹_cڝ/7��;6^�'�(&�.n�Ԭw.��긾��*-)N%���s;���t�;�-����IDyXO�c����|����&�Tu�3q���MF�j��{��5�e�=�j���!�}�b�>��} ��ޅ��}Wi���H���r��7�U �YX��Yq�φI	t�����<mr��_���Zh����믠'���:׷uUPO���?iO1}�e-�#�� ["����@Za w);.6�x���p�s�-��׶"��"T�2֒���Sm�Wۑ�����Yw�_�Dy�I��s�ZD�r%'o���2\@ղ�?���m����8��fŌ$5lv���|~�/�a��琵b%fIa�t\=+2������C�>�3���լm���N��%Nb��=�+W�c!�v=�"�5¸P�>��@b2^�hÅ@�c9~�?ʤ������M<EUXyW_c������.��>�!��K�aƖ��I������ 1��C&�v��C?�v�r�C(��}��M�(��i�m ��lM�̈�qu	�ߐ�� ����IU����S�\-�D�N,�]G��Ub��E�8� �5��"S�X��A]!��lX�fx�������؞�܂W��g���Y��8t��Sg)a�6�xzٱ�
?��q���Vȟ����3����z��P��p���q�~���J���l�9������EgwoB`E�_ �,s�9wP�f 9�A�?�[�m�����������[�F�S�(%!�Z������ﱫ�|�y����|Jӎ]x�}&U�-�XRֿVh�:E�T���PM 
%g��.c ����/��&^���|e}m 0�����emF�y���i���w������ �q{������g�p�����ފ(̳fHH��=�2��`�f�W�\�ŀ���7\.��9���4���\v3�{�W�HĜ��<�7!M�7��_��j�(-K�|�r��n�+$�,����D�#x�s�a#��I� ��,��^�/�e>
�+ G�Q͐f�w��%|�|�LB�C�IQ��L�g)����5BK��y0�a\rƇ����$C�}A��O��6��¡��c!��JkR����=�TS��&��J�F��}>���=��ԗقl�o�k�Ap�T��:ew�@HA7�9�9_���57��`��1�4p}���m|�x����1�����N��.p�4Ӡ-��+k]!	�~�ٷ�,G��:�����	��ݢ��׉��C���͗���c��7�e�s�����q�C�\��x�rI+<�u´i2͡�nO�[W��Si׬nJ���D��Y�؛�����7m�����Ng�V�S�����ѼQ<ߞ/ox�x�g�յ/,3ԵĜx��^8�z����g��/[�5�^}U�����v���z����$�G��R�1��ނ7�+��-&�����*C/0N/�"MA�J'ߒL\K���>�u�FΩI�Δ��&�b2W�/Ɇ2�����l��e�ӶʥęOQ���T��ft��A"&�v�Ɔ��Oؿ�!s;�W�%�(��X
������E�0N�:kB�m,�w��G��r��xSLD�Hc���ΰ���t�ao]��A�w��(3��ev$��z7��b����6����Tb�rҕ$�FM��r�m���f�;�YЊ���6K���>�ź��[��o��-�����OJ�������́�����d� �N�x���Y2	V߇"H��~�]3��$��YeH�ޑ&�b�ز�2�%f��+W9 Q��7��񵭕�9�Or��i5C���M|WK����=Ԕ����j�4��FY���Ս������ؚ��W�V#j�y>E�� $�*GH�=�t�T��ОH��f����)Ls
��GB�����h�k��k�[��$~;�F��+��Dx^��� �PĐڂ�b�<�P&��d����n�a��]M�P9���H��aDbU����^=�P4�1����s��N~��|��E�n��Q9Pߛ�O���,�jk����\�'��=�26�����^�$��B�L��!���k��&Z���U�/Ej��o��)�^'��g�弒�枛8�A�}H�̔VIB�[�|�������>��0���c��DA�<i��J�WпVD�R�?J�i�����@i�ڏ9d�lS���Jk)l��^�7�s������_��:E�a�	�w�W�[�r$��ػ��I�h�Q���Ѷ,��pCx��"�Ҳ��s}��l�� N� xht�Ұ�bSQX�W�s`���B+�~JUF��Řf����������C���T��W�LIO��C���
Y���.[c�:�=��}�%�_��^|�xU[���mf�a�r`$��`���1E^�hx�Jzf��4Q�� �8��K:O����|T~��2"�w���TG�l1�u�ࣰ1�|������ �H�)�J�!�R+� �x.�"�����[�%I����ON`lkc�o��1%xHݿ��Es�?�A��^��2c޷������{�w�~�t�w�k���������vP�6"����̽+B��o�НȬ)?�r�S��O�@p�*tr�`�Z��t�"4���uz|ZB/�P�c�qf��ץ&	���s��m��Q����ai���+����A��s��������G�4%C`u��� Hr�Dx����sS 4E��ym��cs�L������:����(�]����L�X�;z1�(BI��y�o��e�/�H*��
��S���d0�S�<L=��!�J���Z�%ͬ��5G���_R 0��aN����,�!���n���c>Mٵ�L(�cU�؂���6�a�*m���=�o������۬��`��m���Ǌ�Mx��Ԃ��r�;A�,ߋ>z���A`��X����#�5�f��~��x��Dz�H|����`�U`o������y��[�lG��Z+ �� 0&윛#Y�0�J�pCn��y��E���NA�5YZ�,~�X���B^�r���*&!�P5_y⛅�\h��@����]G����XfZ�]�l��ۤ�pH]�� ��*J.}���3�\|�Zm\-�����*�(�%9J��u�,��㸀�lx�f�Mاz�-�Z'2����R�4��5��ݚ֓��Ĵ�l؄xۅ{�6��d4����<,���<�Lu�YDi���ԁ��]Ů��SKٽ�!�i�]���[�z��c�7�g�pŃ>���J��%�	d;G�@�����
y�X�
 E	�Gk�^m!�?�5^��I�^�jI»7�)�(��N.]K��z�8>��+�W�ʹ�*O|��F�zD�%�>ʸ3
��%ʥI�� Go���O�@*�@�;��d�A�m�(S� c/[���O�h%VC\�d��`d ;S��oz��Д8q��n<��)Ƚm��!5���Ȳ>a,��X���.T����5��ē#8����SDH#O��N*VP�cQ�mUSy��}�bx���էz�-��絖�3�@7Ñ�ܦ�v�4R���'w���s}��;��΀�ݻt��i�W�ˢ���n��h� 5��-Ӳ�%���W�Pz맔�O�@Wხ������E���ڗ.���`�6���ڀ4�0Z��y#��D��'a
/6C1
��
���jA�v�c^ΊR)6�],��g��DN����&rL�ZN���� ��H?�f4���V��.s^�@��¯�d���݈��'�͖���$M�C*m�U����=�)�d;����37Q?\\�f'��3#7�*#�&i*�DODJ�Sg���l�!�"�G
d� "� �N��Q�"����#�s)��ۂ�o�A�N�`�s&�s�r��P9a�p���b���3�s�_BU�C�7q�d?�X�L��T�wZ�����_iC�u���
+jI><[AP���_�"k�L|*� �fk��.*U~�@T��2��䋸���]W$v�{M�8r�z��/H��L&����&��!��.�UP����J�e�B�}�Cw;��f��-i�������;.���f�i��&�#MRe�:��W�*��y]C�	���k�o`�fIj�X��@�� ɛ'���2�{�pδz���tN|.ŏ�={=3��-���ȹ�qQP�9�q���7�х~��!�.���kM9_���;�r����j�)��'O�ы�]H���"N�W��:uOj��u�2��d�ς�8�s���c��L��RTE�?���":�~y�T���T��q��F`�>x��>8��=�Aû��O��v�9R��<����z���'�z�:@�����V&$d�[=>~�:r�M�܏/̾����P��?r(�ڧ�];4�L8�s`=�{a=�s$�!�|��|(��-��"l���1nю�d�p�tm߶����@o-|���;_kW�i�U{l�z�Z�2v�fV�D�R�N�N7���3�{$��^�b�u=�uw5��*��,h�~NG�3v�S�O[���/��|����fU�6]:yXŜ���?U��|,]Mdq�sd�5<S�> �/��5��*�e��$u@���1�\���$M`6�X
�T"��8�X7F"&Qp(�73�@�]�����M�8��� p\IF�T�M]���[X! ��.~j{O��Y��f��v���e��qذ������i�f������d �̀j�P#��t
�s&�w̅�D�H%T��$e2�(WA���B�}�X�P�5���H���
�Casս#lS�$��;�7�DH�,��Q,$������X���p3�{�D+���f�k(Vۗ`�`E
Y_���4��.�!�E�@B��p2�P`��L���M�K-�����ȋ��Bа<�<
PU��g��a(�U��K�"�����i�Ѥ�b2Jc���H��f����H��� A�C�|�&��O�m.V�,'J�1��=�r�#Y����
I�@��W,�� �tu��:�tAfWl�;�o�]w�e�$������������"Y��[� 5VBXma�el��mFRe���Ȥ�H��(87�� ��nR��'>�A��&j��5|�s��\7Bjg�8�¸�κ�θBαТU��s%���������[��s��s��|�����xR�F��-�  3@��ڟ7[��O����O[����3ՈH�#�ߨ��A���<v~Z�+Y4Ơ@�o��7�{	��/S�{�l}���|�'�z�օޞX3�Q�D^���x��.�(�����o�1�0UhY�����J(�pn
����I}�E��¨��v������7Npo��d9[����s��r�B�nѤ�д!�����3���p�.Яq��(]<��64vZ���q�5[>_�q<x�]��8�u�xeQ9o�ǿCX��l�X�ئ��X|�Õ��	o�������w��x����/�`F�U����A_�!�U:�U���P�6|�ۥ����7m��M��E��5ٸ����'y����K���[��=X)*X�qwHs.��&D��#�v�ZvSw�0Z0;�1;��}�Ѝ ��4t�?c�๵nm�\�Je�>����B��
>�)��N�l�C(�gpA�.X؈E�����5 A��4����k��־^����n�z������_�cI���ծ�ʔ_[�oQ��q�՝�V~b�`3��|f������5�`��n����R��ժ�U� �:�Ţ�������Zܲi�&��Vi���A��<�Le�Q��*�י��۶x���`r4�,��_�wC�������U�.Tka���iё�p�hL�8n!m:Y��.NlRCE�l�)�(	)���w���I)��Y̌����.{��[��f�����:�7������-�d�k��^s�̻FgYe O�Zv��^�
Nݾt��p%ž^�����GB���H����>����5ӽps�������RE"���z��(N��f46���gʪ�;��K�]+p�{TA��Z�R�9���SǕ��ͧYxȝ'�cK���w��v�ŕ�0����}bT��e��bׄLӆõ���:��͵*@�?�-~+C��2*%8H����8h��hH(E��L�(�m2�����$��ΪK���-������9���9 ,�6�%�_[B���9�Q�;��B��$S!� ����`�i�M����n�	5��\E�gTʿ���A�rz&[�v����l���*"���ѝ����:�_��N�e�L�q��H�ɺ���@�/�����S�s�V9��_2X&DG�?K�Œ�����ŭ:�e^S����ъ��a|I83�~�F�Bj�o3hˀGuen;��0�gQ��V��NZ�b�9O�c^�����(�92l�y^�����V�|����||�0|x9�a��d��>V��$K�c'���{k�e�7߁Q����+N%�'�0P����WE\`�ɼ�����
�4��|�C���銌��<B�����5_�f쟮��o�XNZ����E�*Z��TSt
1� ܽ��-rβ_},A��L� ��O� ����:���Z�6�j�0'��^-Z�_���l���.9fr(�f2 H:�hi�I�g�}�Y�M�5���3��V�u�T���U����f.��Ŋ���)�ˑ��v�OC��#�;E�&?�-��ֱN�r�ho�Y�-ðL±L����p�$� �_�rQW�Z�ޣE�XF輷�+�ފ�ێ�'5�"��וS�����ҙ�(C.�1���`�{���>I*vx�9IW����ǵ�>6��{-�� 2�Z�L�����8�zł�ء�D(:����gn���6O�ʝj7A�Ս^(���lH���k;}F�Dl3q� R7roT�<#�F������.��CQ{�ұ�ì�>�6�b�z�zE��_�1���G@�Z��NjeޅS�#&�>����́W\�K��Zo�)�l޸��+n[
7,�
<���gVI��*;ҽ5H5���,@%4E(4R�7�F�f���$���O�)f8�J~֏C���N�x���%�(��
�j�<��%��oz��{ݎ��*�]�{xh�,=iu��~�֛9��;o<_�+t&��L�n�:�g!�Z��\��\�Ag�0(����Gwc�U�io�0}8Ã-�UN���OS�D��ݖNg���%�<
hC��mf��lx��Ac�m_��2
R���bx1��Ű��;��c�ü1��H6]�\S|9�ܨT�\t�g�Z���q8���yt�"~G��l�q�8F��m��_���(��BD މ%�0��&a$��#�#"�ē��??`u���$ه��$Z�ES�� �l�Bt�Ӏ�E��sS��vQg �9�ז$��4��4����?$�����
�S�$��噺\��+��ʟ,�Ϛϴ� �H�1��1�L��T�*{���\���
s��ƴj��&�$�G���W�j��YK����N�:5N
�%g��O��.u3�o˰�#�ϟ7��'}�/��/
I
��� ���O�Gu�Fw�vWWK�w޵���V�U���A��zk;���Jm�⧵��iO�,����"M��^G���ĩX��<f���{]�;�����T���@��:�j�C�!Z�&�R}��Z�."ۼ)<3.t6�6:vZ)B���ٚ5&�X&N��*��"��y����+����To�h����������5�/4��As�N�T��8����w��1b�H����[Q�/u�i˓���~(z17Hٴ�^v�KL�n��C�)�-�l[���	
V�j1Y�_�Q�dPA(ҕH,0�U�����Ԫ�����&<��xzCt�-�غ�)����k�4�B}����},�.1H(��1��5��p�M����adU[}����w��l-�d�̌���@N5"��~�E*[���:�/Q�3aLӷ�jS�p�|X������=ɖ��ΰq�!�[OE�-pv]�G���ژ����1ME�s�����8|�3��	Fs�
n�v�9�7�uC��X>z�~xo�Lo��i���N2�F�G��G���F�t��ǅ���tm$��͓�t�}��Ǭ��;���]<�N��������:A��B�K�-K-�J+��BM��,G�y��P�Bzs)��������&Q���9p^A�RTa8Y]����]��Q���_g����3����q�!�2��⎥(������r
���p����B�3:�j.R �<Ц�Q!:0�^�a}�"&��#�?��2����R'0}/��{����y���w����X<h��p7�8����'����W.N�
|,��Ub���)}�Y�&�����别���SY%s�2{�˝A4L"K� fN�y��u�I���z3�!r�mN�u�K�����ش��j�����r���v���E�?��\�<�r_�|ޒ��Yf�'�9ePxȪ\c�#�+M(�Τ2Ԝ1R��Q�z�X�~��5G~Ϭ;�ve#&�T�4@ȿO0��`Tac�5*}�5"򥀚Im�y�D����Μ�%�{I���a��^��о^�{:�ڎ��a��Tςޚ�E+�k�j�Yؤ~Ѵʹ%/X�J��f�%��6��Y�#�~��zѼح�K�^y�Q���!�DV�:i����9/9�V���.sp��3��.�D�dԆ��,d@����
a��+r�N��.�ܮ�1�N��v='��Xk�r]lzc2J�џjZx�H�9Vo�9N�����h<F
��C��D���rr�s!2Zg��Y�� �e�Dn�jjM>eN[zlЩ}��߻���~����S������{D~=��i������K�������I݋֋�����4���8��
-	Ĭi� t����uj���m����_7<e��G���S-̀�$NrI�\h�9|�r�2Yl��5
9puĹ_ ������]a��S���տ�}j�����+��g)�A�u]-��-�i��w�����'(*o�B�D�^!sC\��S����Z�,�y�C�&5�A4Q��Ƿ��bc9����i��K��������3_ន^�v��GC�뗷���w�ܒw�D&vP�'fի�!�0��Ek��&�f�7u��\�T� ����=�᨝�U��ji��C�i��&����~j�PC��� ��@��Ѣ��Y�{r�tUP>��?���1
�ɸ�7:��*sY��
hHVRϘ���sU���us��\|q�}���3i��t�:��6��O��P���r�}|3�:]��Sf㶼x���{�ߜ[�H�}��7�)rՇ�g�=��t�e���k���J�a�kC�b���:u��̷����ז��P��0�� R��Vb����f��A�Ǳ��qo`�[Jߖ�L��2/�$!O�Y<�//T�p�!ү�K/!�;�V���� �5����Ct]ȥ��$u=�%~�)�O��q�[��7ِ�����CS�����p���������te���nt�2�ځ��`P�紪���c�/�%�
���Sy�L8�#8�і8�암D8� E��h_Q]���;�𫳴���w%����XK.�=�ݭ�6�=�ŅɎ��BD�>B�6�� �������(�O�=���?N
~bw|	�1y��� �
q5�H�F;�l�i%��yE�X��;�W5�W p^�jz���id�'y� �K�f�#�G��l�h��qY���B" ��7���(p<5��q{�O`E��������bt.TLfc �ih&~�����t�X8��*���1$���d��d��W!|�Mv>�}�!�_W)�� ���M�OE��4Z�eހ��0���L�EC�l��i��ސë�az�S���n.�ךKb�P"0-���V�i�(��^\A����g��!���U{����l��TH�x����<��"!�p(Mw�ޕn���=Ή>��|>9|q���O�&1+5��_-B��N��꜒rk#^�,d���BP��V��Z�p`��]�~6qΤ<Jv���!V�\\�o_cY:l�J��^��Ӱ����6��ئ��~ipR����p�&���%7�~�
��s5�5*��e��}��@iI`�W�B�����q���s�G�eQw��"pѣ�	g�jm�mm��m\C���g�[�%]�*�?qr�T��Ztp�~�Nl���ݍn���9�S����.��0�Zi��S���_��D�֤%�y~�d�
�ײXjw@e���0�6MψՖxU��lf�?Y��)��Q��;`?��u�zI�kb �[j���S@���R�&k��<�����P2�_�gɷ_��#�nVƛ�^�Q�2�K\��4e�H1��T��6XH"S'�c�Ĥ9���%Y2?r�5��h�(�*��0��5ϗ�T�A��7�8Hd����zR� x��:�A�#r<O��*>����*�^C�NN(�_��w9��+��_Ǡ�X�)4�	�}�5A���U����)�B@7�p�r��qm����E��������x��/�b^*sk���g�j�k�{�Y��{��K�t
_�Y��owmZ�@��_��E�ws��nR�����j՚�XH���O����UqX�����W�\S⢌��寢�����H?bo.��)~4���~����S&i���R�Z�M�iX�ծU�^�ؽ��s/�A�+��ybs���~0�J�;�����,m'Mk��6�n���,�~��=	�"��"V~Ր/^�7�##�f�i)��Pr ����W�^|�U�q�Al5�!&�'�'dB���2�o楍j�����˫�i=lܵ~ؼy�qb�wB�������߆�BqC�c�g�xy��G~o���F�x;z;��=)#iU!-�/��dV*�P2�P*��p<�>�}x�rM+	!� \��s�a$Mƙ�A8�d�rQ����d1�J#:E�}���n)��cg��ķ��I�Pêd[|b���P�ӵ�Y+|3?7��jM:���f���(|�:�Yoa�[�=�N��w}�ްU��>v"�v;�}6C��s�|[|�����n?�6��bg�
)U��۞7�h��v"�E�p��]��;=�2���{{<=[>U_>2zcõ@i*��1/�<�T�J�U#~�dºǑkMǳP8��Fu��u��J��o(1�OJ(�����64XRd]rBYv�o8!�o�⬉z�o��Kx�F���{�;�g��߭�r+�	{�<�[5;���%	� �7��Gu4F����7$ݖ�u��T#��N$����2xwmlb��xzɠc^�*�e����V���%>Y�#�u�g�AQ����13������Bn���	�3G�s�@�+Q��|��c
�vJ��B��+3��3˶�A���H�ܱj��l�D��y�$�n�Vi�1���:J6싚��^s~�u	;n�ԅ*��oԶ�����	ɶ�HTr2�f�N�U�f�L�\������m#&C��;�-�O[fv�%��~��Y�<���>�HDI��w*vJ&�C�#�Z���/qay�����)��o�~�5z'm~RT}���/��Hɟ�K��0���ȱ��eK9mM&7p�(��I�c�E��_�J��A^�>��̂~�7�^��'��H�w�SځW�<����˔^�D�-�a��h#���cHL���#��b���a�]���"�R����'�Ln�G[-��<�@�r�	���`��?� �UCYժ����^=;D�}E��0(��Hl�S�ģ&j%<=w�5Gn^n�S۽w�E<���W^.�9�����Kq��߅�6Up�@*�<�\��D( �`4��oH���(�@�`�UF���|=���(�#B\HY��?�Ĭ�e�!I�/��j�z����F��J�&��n6�>��Ϭ��Fg>�ά4�����,,��)�g��g.&ѽg�n��H9�L�٭���Lg�K�H�q��.�%;n��o��	����;Te��X�`V���Ho}�V��|5,5�a���������Nk�����0�R��I����˅��%���=��=p��t�t�U�V�n��������^Mg��*�;���HGSC?�l�nY�Aq�Q�Jy�޻z��e���T��oѷ�oŌ��A�@�1�[-+�vW�@,��Ak�Ǔ>	�8��e�� ���u��"�v����}��d$����
Ӆ�U���I�Ҵ���؅��4�3�Ŧ	>�3S�ਕ7Y&��Y]S�.?����(4�V|  v�B�m��R̪Jd�JO��BF��`���F`��BD��vDEP�,�������!�|g�|��g�XY�u>06�ѽ�q�2 �vLQ{S��.Y�꟩Y�e�4AS\�,��g/n��)��[�&j+ʘk�$�~�M�|񶘭�V�[ ��T��Y��+��Y��|����J7�r��$ģŻ9]o���a�O��\u)��^��Xu�0t�4T(
��?�6��f*E
�p�G���[N �^�B8饏%�)#�m�UR		��8O��/`�O�r�d7�-��~�?��PU�۞/�-�H����4��8���_�,B'���2��o}��_8�hNU����Q�zO���\:�ya2ÝCZ�[�\XC�*PU4#�Ri#�"���%�F�>�J1���6���;Nb�C�9�G	�B�tx��?�̆��)��͓[*�����0@�~�s�n+m�� ���a&�h^+��f}���#;�&�J����v�bm����&CY��Ⓘ����a�s������o��}ko����P���}h1!��₰��D�`s��7��|�i�`2}sRAS2���Ap�_�`��F���j��r��������!��=��5��u��U�M3�ː��REO��%c������zN���c��>ѯlR����󜨼����yh�u'd�'qi��יNº�����"���ӣ��en�]�NR�R�#x��	�q���h��9uz:�S�\S��c�N5>�Տl���D�w�HlR(��V*�}�c'�I@<�]��KU�8�#�u���:ԙ��¹\١��)�=;h�wCk��_�cA����/�vߐ[�kȆe��m<x !�,DP"�a��d���q�>F�w8{����������ʍ�̇�U=!��;i�#c�c���	���Đ�#�Hs���feV��bd�y�\���,5�k�+�:�Q?mFm�yg����("�/���~�S���4N���W��  �D�<gd���'p8L���9R��Y�&����_G/;�+�j�q�H�r��i a)e&��YeY5e5�MM 0w��U��V�V��Vck:�d)�_*�QO����'d��4�O�{���{�4�?-9�N:�����S�z�C�08o��5��GG��I���TаVVv�{&���3���&yZ>��Z(ᣵ1������sn��ȡ	H�����*�̅N���Ζy*s�J!2+b��]P������Y��fj�ȽПs���<P<�m��=����-���O������n��}aG8+W�����k$\�4
@L� q�v���݋�`��.� �/!��͆��}��kljj&$B�Yn�ɩI��bszp#X�C�&�F�Bv�?�~����F�l�s3���W�${��lo��_F�ں�v�Y
b���9:v�pbF�B���4H�N�;	�3Љ��=4�i�1�!?�C:�A��Pz����B>q��`\~>�ȥ��E~-b{�o����^��-�������&��s�F�.����r+`zi�?���_�kڭG�g���Ӕ�v����nق؇l�{��
��?�0�9#\ހ�^u�Td$H>����'S;�h:ѱ�����`U�՛�Tzt�GE��Z	�z�"171����������,5�1%�(�|�$�E!]�t�j����C���^��@O�њ�|�S�ZVďD�)p��K-r��nԄ`�IX,&��b1It�I��pm����V���o�V�m�U���0.�Q͡bF�����zYG!X�Xj9��uժ㡈����F�jo�8-������=F�Ptl��F�����~�4�.���� ��.�'��wc�n�A������S���5@GH�Q��F��J��R��� �iE~`��`����O=�Y��Ig~��c�,��h��h��E�CpX��!,�uqK� ��C��,,n�=��Bp�@РA.�������꩚��9�yN�Ȧ7���&����r}��y��x~���7GX/�ɥ��)��H׺$�@6�z?lP�|%@�(e�K� ��4�M!���0�S-}6����;��,����D#�9��U��*��u��&�j&ǽ�^Lbo���V%�}�ߔ�����А�L&�*S��FOln�/^��mt*|���R�f5	+�	���)m��I0�$�[�QX������<\9x�b�M*r�F�˔}S�X�ڼ��[�J�
���T��p���H��I9�q0�U ӕ,�y��ۘ���X��1f�7��Ѭ��c�({�Y/L�N��Y��~R�`�ԣ��:�_}���]�J��a2���������ۀq_.:�7	�lB�n����_�ʛt�_�pd��\���=ރg	Ɲ�kzH�� ��旉�;�3.�_�xj�-�z�KH_O���]��.�}��#�fqLd�?o�&�ܖ�e���B���H8'M�?ﮄ\ˆG����Y��/Y;B��R�I��s���k��6��b=�����!K3�
g߭�յg|g׬����:��ұ|<�
�.a!�2W��X�����33u�k���>�.�����Tf�%2Q�7J0����!mg�j���?�9_roƸWP<*a�۾�4�Y���Y��]��]V��U{Ns��#|`������è�-+�pgY4Etl<��yS�r����o;�e>z��J��~[�h�����}�1#{��#��i�@��u(��ըH���O�v!�M|X��ky��O��ߜ	Kw��<
]Fp+c�[���eX�cw��e���"ty�ѩ���D���8��D���.zYzǰ�R7~0��`{p��:8tBenl4��2�h�g,U���}�!;��@$������(�	 jW1,˾(���d��a̎�Z��EpiX�R��(�ވ�T�T��˄z(4�%���F���j{
4�y�*a�F��>��m������?ę%���{��#^���m��Sy,��vh2q ύy^Ab]<��L.�wָ4P�lf３�Q<��.��l�%z��GE%%��&B,�ta�*	ET��*{����wI�zV�/���ǔ���2��憸g�Ho�9!��r�W�x}���<��P�u���?�O� �j��i,�Z�qd���������r�/ALd�ne�s��l �#�4�	x'1��2��L�َ��-7��Y񜛇��r�~2�X!����f����V��Wx�\Ε��J���3w����)V�ĢwŜ��Yf'�,���pVo�G9�:9�4L �k�	�y�QS���j�rDd��b�����V��jk���#*����l�(�(�5��J��������ɠ����f���"�o7����V�)�`e����a�ڂ���w������;2�������})�mI;\�T��K��/������m�W�� �H~9k��f��0�9��Π�U/#����N�eRs�:g�֩��ޱ�I����."\�P&�],�?7��j��s�o�z['�J�.,�N�*�nM:a�[���`�N�a%r_��@�u��74 ���u��MgϺaK�k��7^U��(�)�Y�Æ�L��p��5� ���O+�|0cO�Z`��6����12��')o䬎vxH��T��))\!T`>'z`0`���Z{-d&���"�M�:����V�>�H�4-��Oa��θ�S�ۿr�5�icsը%s��|K/�hA����ca:�1��mK6t㪥�:$�ey�W�u?�A�~y�a�i<3��j��R�HY�鳑F\�'D�p	�ν`��FȢ��0�~>|�E������QCh�뀢�N�=���_	�-?H ��n.q̹$�.�[���f5�ڌg-ݖ�"���t�Uܮ��1Jь����QszS�jGB# �X]+�mF�V��bN�	=9��*�!���c`'8���4��D� �3la%�|�&������zD�7xgZ��S ԖXg�,������k)a3�WKF���ڗ����K�i�Y�av���<��}����
�(�������oV?�ʱ��"�Q.���}� ����7	Ik�_IC��Ԙ�4��K���_=L�$@@׍I�M$<�75��Fu��2��Iӑ�N41 �4���0���H�cp@�91�GEs���x*��]z--s�{�������/��k�n��Nz�H�z�V�?��{��f�k]^��֐���ۨa�p�m�0-�Υ�_��6;GA����Γ7�N��ȯ]�"��u���g�fG�v���I9��<}�m�~��\�[� �!Gy6��, (!�J���-6,�cA2U8�T�����[�^���$����b�e#^��
�Zj'�.���w�A)������nmU�]�Z��8��?��ǉ�\
q����p��{keGHO�N;�y�q���S�`-�[�T�2&��f C�N�[�2��lhw����]��%~�;
M�܆�>f$�ƙ�*a��=?AV{���E�m��&$UF���i�[
�/o���~~�ƕt{,\��M3Ao��$��_dd�w,��P/����N��T�&�4ƎiXA�c� �)�w��l/�׀��_�7oÊ�§���~� �'208��m\��?E��ӫO�߅zB�	 "�c��М`SF��3m�.��(�V���z��z�S.�E6g��\��mKo;絖����Ê��	�����('���EgL�rچg��/�L*��AQ~5eq|FQ��N��EOm�+����S�� +,�+�6�����g'����'�L�x��ɒad�@Zj/��X����������b-��?e�;n�O~=E�*����Ù�s��;�$��*�d�����Q�A��K4��Jn*����~觗fm!�#W���Է��E������N�~��'r���p	\h�:K{��Zd��#�Ŷ*�F�$`�b�>>�ċ"~=P��+a���n��It�[eR*R)�;7؎[�[g�[#�$��,Lȗ`�*�~%���	�ß����꠻�I�ǭ��_�b������W�U�?�G���U��m�ϥ�_��k�h��N�m��zB��{Ң9 ��TOP�t��7�A�ˇt�ԙ��gt���M��g�-�ά�"
R��F��#К	
����1r0ai�L3J}3�r|y�T��ǣ�#�AGbivL�Dkج�Z{����f�a��R���R[��Ll6���?�yTK�+�~.`� jy�X�j�����K���f��[->wuN]��1��$j���W7����;ȏC�T���)��#�ُ�m*s9�l����N� $��� ���F����p��}�����eP�<��'V�ȳ��q��8A $��pr��Bp�rSٷT�@�DwL���W!h��r/Y�z v�t�ğl0�_إ�jԤw��Tb[Ӷ]�w݋�y����#�{�]����n��n����*�d
<��?Q��^�my�{��{"�^��7���}�<�x�b�0fp&�9�h4'C�Ki��a�PJ��������cT����1Ã?��c>x��i�(��S�jj��āDfCs0��{�����BCͨ}�-����m��Q��h ��y�{����u�uNW�ߤ��a��Dy�Ơz�{ac�\|�t�� �N�zP�O��ߌ�����Q�H�~�ze����ʹ���)��`l��W�5̻���-�i���NR�i���S�ϼ���T��ui��׼,��Kk��?�{z�G���i�����# ����YI|n	b^I|�<w���؛���z��S�I�E7�b3�B�>�Xt��Ԓi�t��~+� /%�{?�+����k�2�'0�-���Gy�e.�fx0�~u�A�ݍ���)Ry�����D7�?�Sa�!�K�՛�"V��FD�$ǖMY��?� �פH?{����ޓ��̒����O�fAO�y���7��.������ɯ?��w^S?Uv V�\Pd������.qy�e(�遌8��3�l�T�^``����D��dq[#���|b��fb�y���_}�C�i��uV�ǎ��6�?~�VM\�`�r�{	Ⓨ|�F�����ܽ��������U�Ԑm5I߮M+�b�JY�қ�1	ʇ���x$-~��fe�H�c$\`�	�٠sX�`�##W@G�B���(��7�����6�iI4��:C�#�źϗ�t�j�yl�%^rU�m%"䤯�������]�����S�;)'�Dt���q�|q���3�����9�zx���}�*a��TA�@3R�k0}2ֶ�����D�&ib/�1��ᱶ����u9+Ȃ%��c��ؔrR������c���MүpPj�'�`�1t:��AN�5�&7���9�3�Edf9l��{r�w+O{h{�M��;�I�E�o�9�+��Iv���������;ne@K������{>����V%)u/K'	�^!a���Nc�2���7b�5��4��	Z���ۋ�{)$D�ȯ�wS2�(6��ooU�0��к䤐��[����bީ$>i�F�g.Jk�qN�D̮ɞ\��~cm[g�P ���:����MM�E�n�ݛ��[��?�ڱuDz�_�Z9G�x��0�����;�X�������
��$�0�J0yQ�r��w%8�$uz�t���P����?���f�T1�?{/��q�~�H,)LF�y���V�����`�C@:�͗:t���W���S���k*+h�)(Ϙ��1Ԅh��x�P	]O��������!���$:�K���h2?�&��K���2}=BdEI]y>6�^R4�8j�d�*V��yAKC�ϩ��fQ����x��aa��]z��L���z�~����r�Bpt[�:�5�-C�j���H��w� R�	Yf��+K@� (KG���yU��ȋ��Ac�y >;(y�(_8f��Jo �����0���L��]�M۽�x��q��޷췵�l|� �eŦ1+�I�谇r%�?���u����Sףf������b=��Ŷ�	��I������_�C�.f%�D���jY�\���i$	Ƞ-d�O��a�He��)�H-��1�Txm���W��d鐝 K��b 
��x{e�HI�]C��zm��FT����=�^SF�L4^+���>n�ùˢfi�,R�Jh�٬ �(���7e�+���L��$w�������%C0¾K�o�����v��<mO�C��m���`�nрo	Fߴ���q�;��$S9�7�H���x�2��H����P�Q�������Ps�$}���n��q�T����4n`���V�"�&�M��"��fH���ަʬy�E�ܲQE��)��[��bA]r��6�mW�/���|-��ث��o��"��E��s�X�Xg���ҩ� {��T)$��/\g�v}@0r@f�FsL��G���4x�k5-0
ŋ��|	!Eb�΋���\�r�\��}�q���Sh�[��� ��B�!���;CZ&��N�ԡC�ӄ�V̄�$�_��(��H�%�5��rP�wj���v3L��0N넜Q�d��t��o�y]�ۖL������C��AI�{�y��<�D0�!�=.K��f �'l���i�Y��.�������j	/��#õ�i�$������@b����W�q��#�d�Os@���]����F'��	��O<�PL�.7W����?3F��W��Sk4����V�y�UW���	��ܪ���*�a��W�Q|U��_�|2�u��L�X.�w�v�np�	�����	+ד�iv
���j6��,�j�yc4��߸_���Q��d��}�	"$e�l�C�*�ݧ�U�g}F>3Tt���I��XQ�%�Μ�y>}��ܹ3�4�4�y5�yn�fۡ��1Oo#���B2.����1'�~AJG&�P�5��b��p$?@+�g�����D	���G<sMB}�5�k]n�[G�=o�����1�J}d�+��i����R6�J�?��IT��/X�}c�2���Y�S�M,�wޤ�>�]?J�������^�/��(�
�2L�mH�0�A_C�@���]� SK��D��*T�����L�B�����D������х����Q=V�hb9��o0
���oڟ&(���DO;ϯ���O(6��߆��2��*��RP&���Ѕ��R~���~�>�Ȭ`�+(�������~����yk�F�F��ܴ����̟���+���o=�\*i)��X-v�ذ(���M��Zz�,�d=���tP��o�� ���/'x�*�ZQH��;����q���Ҧ������&�jo*�Ƨ��R��bT�h���P#Os�xAD��7Y@c2l��3|��0��"E�-jIXF�]QV�o�:8�����Z=8�|_����A�R��F�Y���U���Ю�qc�W�QfQ:ի}��6����P���b#g���*�B8A���9��xGɻ,��!?>9���
�?xlA���|H���
���qP �4��j��n�
<kpخ��~�4���i�[��o�H���ǥ*��0�����5S��(��_�G9�-�ش7��K���ъ$���a��b{12�ͳ����|k��.�j4(�'c7 ��)X������ma&�9���|S��,����CHĝ�$���������f'��OF' ��G@��j��A2�:#����mØ���y�pIZO�򴭃k�.��?��C�9�YLpJ�"Α�(|/�O*h��d�Z��¦V�A��^�rjmm�@����\d+,��Gẑ���M���6n��y,�ިɈ3$^�>ХN��)S�.����^7ĸ�Z���A]G���4��2�(��Ƹ���Ϥ~�-p�Jȴ�
�zp��&��e�V#Ҋ�.��0]��f

S�[8�s%o�w�'O�z��$LZ�������B�&hX�s<��W�t��t�ɡ��n"Zg��7���,��"#�Om�a@E�9�A�cDp]P��8*JV�������\B���a�(�V�01��
�YY����C�������W�Safy]�|�6��]D*�#��Q�G
KV>G����!(�z�͘�<����꽲Yʬ�}K�?�d��Wl�JqK(��h�Xm-��A���yC����L/Siث�if�,���P*s+�mG��[E%O��d��Э�.�>��iˡ�g��$V���1�cV>�;^\8}U(��#3.��ڤ5.�ͩ�M��E� ��)}�	��7�*& @�wAg'&F�S���J�Ȧ�P���'�8�Hj<o !5���YfJ�L�G��Q}�N.���Z����uV?k�M���ʅN��-gB��������}I�e��㒠�Q���Ѽ�=A����<��n��.�m��/<�?�������8J�|�(�H�~؂�u��SvR�X�$�b5�|ܸ�@ ��L��R�גK�4� .�oU�AY���c	����b�~�&���@#�<F�7�6^�׬�/�}�9o�%��D����\{�oh�T��LB�1{9!k1:K61��A��kN^d{H���8�va�s�z#8K(��'�k�È3�^�}�J������w����:r$��Wu����#	�c	�N,��,w7?��N�������n1�bnu�X|��ϧ����/�?�?��V��S��Uۡ��������U`CI��5�@5�������&���U?�]Ck6?ޖYEj%��/-X�;�%�P����Gedt"#�}�t���]��ď�Z�I�V��<� c3�@P(��;��z~CmMk}�Y��?�b�и��Æ���l�8V��x��d����[�&@�\qo
Sk��r-c=.*�����7B�k���[R�Ǯ��]���9�
��8
�=��5��U�]v��(Z-�!Z9˅���/J��p��<n�G����v�lK���KO�.Ck�R��n&���@��!����j��@���XD�O=�E,	�D�jT
�n1V����2;S�
��!0�!�F�#�lQ" y'����! ��H:t<��iD���ݬ-T*W���lu?����H1?��V6�Z"V�_� �>��������ּ�P)HFŨ�{zPVS��A�҂Fj��
�߈�wͳ�w�l|�|��*��g�[���r�a�|XZ�dX�=?.�=&(7��f;�m2��ڗ�³�@�Ţ����dlf���+;�}U�}l�؞e��T>�ʕʯw���\C���f}��kq�����l�k޾���DRb=Ы���~kz[q`��X\۷��Q���PbY;��Y�=�P��}w�2�����P���6ڰ��#���A9�vtLu�ܒ_�D���E*rc�2|&'�@Bz���x�l�j}y.}#�bv��"���Q�z��vQ���;iS_��#n���T�iG�b�����L�l����N�E��^ j�������%�rEg� �^Zxg�L!��l� p��(�p�3V��N>���_�fe�xY9�:L �t_�({��-跓^����Hg����!z���Aѿ�����CmҖ������兝e^P$_J����|8E�O>8��m]���TIh�zu3��G͐���3��e ��W�DNR7�͉�I�>����k�>��D
�>����d^E��RX}���8^x��I|�����|���k��F��5�,��,��{����������~v�U/�O��WRE��k�Q��%k@qo@�2Y��R_@����Kp<��4;I�|4Ǩ�Ҝ����r�?���5Nۜ����n&�I�$�y$e%4'!G�%��1&��پV�va�cd=!��(3�)�^ts��^�K��b	������ |g5#-���craOm��i&�
�d�E�,����ٙ%Ytw�uiՒ4�&��`6����+e-Z�CJ��X���E{��U��QW��h(���Y�¨[�����-�mG�T��Z�V�Hp�.#�ݴ6h)��;���>����KJ#�U��z�$�G�S�'��~��cf�1��]��\O�M��~�$��P�#�}
 �*?_�E�b���ԔHQ��v��Q�ѱ��������Ȃ��_,p$B �&��:NV�������d�#ĝɀg_m٧^a�k"?�w��fAD���8}�a����`�*s�>i�v�ɯlne��3���l��W��P��T�j[����u]ǧ�z�>���K�����h�\X� n��5�d��b�F��<Q�]�a���J��O}�:x6�6��g��_��W*B��V�EzԓϠ���~}�ԛZ��면����g ;��`Ϩ�Y��d�
+�����F���_b�ۚ5�Q��r��ǗrK�)�sb:9~��9����Go�(^:n�j/��g9�"x��Ɋ�Y��J�b���GJ��˴&*jI�5�Ti��)���b�f�����U��^g�-b ������N�#�A�u?�Y�Tͱ��%����pn{�+(��t ����4�� �-��E�����U�u��c��|U=w��u翉��������g����̶����Q���":�����Nҧ��mӠ��	ӁN���*��K*E���+"X��POdv�\X��9`�g� �����B6Қ�1 &2
1匕;"��%Sg�*�:#o.X��2{��tнߝ�I���ݜ��X��P�saxc�e���@�X�G��d�������[Fo�؋7�bexQ�{@�W5�z�.��V�]����t��'+���%���Z��N*�*���?��DJ-
 ��ɧ�1(�6�S��TV~������������Ƥ�,��S	������!憸�ԫx  ��2�e�>|��`��wM�,�����9�:ی�C�\z��8�o@#��?�I������G���+���՜�V��N�Ϗ��jL���=`�2�=�}?�y���Q2�p������WUeg /��z���E�a�^���Tt�B�#)�Q0W��G���h����@9��V���):-A��(+2��	������2F��j����w����9��n�Y��������A�IFG�-Q�z�f�;ϕh��R�>�1i�Q��M���mP�G��FR�Zn6e��V�Ʒ�v�:�5�9��ř�����M���L�ôX�`�)�?1a�K�Ą�T����5�RfI���ǔ]�e�)��$�/����{A��ĭ�,�%�����wPK�+R^��E]T��KG����E${?��MO���j��~�(�I�z<{��Q;��l�����@����y��f?VO3���$0��.�
kV�'f�g��+�DPiu�Ů�E'��u�}�+�! `�
�1k:����M�I���;�x2�j�(�L�B��ɻ-?W�<�d:Ԭ����Ħ��t��hѾHr��Д78/��L�k{�Wa� e���IkZ�{��.�U���%~�-1�{�j��|���R@M��OB��!�rv���+G��,T[��K�|�cd)$~���ojϸQ�ݩt�y�P���^��%���S�M��ܯ�r>����8v&�t����lFy�*���S������_��^L�(V=hO{~AG�eF�g�M��Vǽ5��J���ۜ�:aTY& �	���r��+ U���	������K�6�֞�����q��&��$�^�.,��T��3��D?sn����C� ���r���6�du��>}:I�|�(d���`'�J����Y���_�}��+���]*`�- �4�����՗E7$C�lp��_��6#����P��a�NW�eNbV���ɼ�S�Y�M��f6$�I�7e._e>&-^ȕ���9�D�y�]LuNm��M�H��ׯ�Z��X[�'~�S:V�g1`w���&;���5�.�W�O�������K�΍��bS�[g�$��f�b�Z��tfy3�^d��"�	3�S�嚝�Z	�� �b�|�؞�1�Zͨ]��8A=5K�'�v���|�5�*��S~�'ajU����'g.��$Rv�]�W�������u{n섭9�c������ᰱ�������������%D�=h�S��0�G�5��;�"VH]R�������������H�Sl擸"�)9���|U}vb3'���*���������U��t�����	�2x��z�S,<����,;( �vW9�)°5R��<����9�o�5}>�<;e:�J�IO�I.���ZU�����K����;~u6�[�������ΐIy����#t���)�~ML���Qe5ܜ]�ܔn"�o�>���,"t���ɇ���-���a�M���7'`	0�����1,��3p�XL� ��2��e��`�"w!~��	Kn}�8�G�q��/������Ko^��+��R�����C�G�,�Sc�t. ��TV]�J_y8��P�d�����w�dw�z��@-����ǐ�BZ?KPo6P�u���MU��{�:��˒2p�F�����-;�[z/�آjbN��ւ�9��VR�Z*�.{^6t�;T�+2Ӕ
S��n}��N�]\����UCt�J�o��<�8?˺k#��	�w�������3&�iR���h �eU���J;��R�p���ɪ;�k��^ߝa�<�d��C�L�������U��e�zIn5C��.�3?l!xv������4g��P�K}�+5[�b7�v�+�"�y�L�*�W��:2Դ[�L�$\z�ۙ�O �yl }�N݉���7#mfm�,<�,F��$��Z�j�ߔP���v2^����3��ik�ɧ�ى�����}v�)g�Ͻ|Q���5t)I_be�Ӝ}�1֧���SM�O;�@TM���PHx��Mgh�a�c��n���`�Ֆx-&�&�B�E��J<jǰ�zT����pΖI��ǉ���z\�J�ܵ��	W&��V�My�0��W�T>3g��Moj ������m|����j%��S ������|_/B�'V��ٌ���kwF��z �g?G�.1&hq^63B�
��o�цG��5�3e�4�q�U�|�@���C��S�-=�K{X���E���[LkѮ��f�SF�.�:�����-5kSlZ�c�;��9��Z�ɚ�S��=�ޣ�=���X���&ɉ՘Q�����f��q�f��z,��8���9��<�Q�J4�Ʀ�l#�X0��j�C��ќ�H�V�͞�8l�x�������+�Q�����'�[��!a6�\e��� ��Y��lh��m�0������2�Łe��p�?^���SJ~O���n�򝉑_�'ʗ����YǑ�C� ��j���5���)�E���p�Py���� ?5�~�C��}��'	��d�-Dz��A�򫯘S�&rU��x--,�����Mu�^0w��N���z82{~�|���dvy+��/"v���ѹeF[b{Ɯq��4
�4���	��O�L	���?s��>�pQ�� '̏�,�G?�,�'�����L���Ow������k��;4I��4~�`��!��WL���Z�"�=��"��)!͂����'K��\NL8|4Qy�?5Nc2�%h�M�&��'�#e�H/�I���!;�0t�_�;"��ve��tC�f���5B�-�s��s��V�?9��[��g��G�nt)������� vk	���ᅦ��,�'hT��椁/=��&;@��mϺ�k+�yb�7�Oc|�����6�0Ǔ�G���Z;�h5�C��LR7��H����V���\�7���mE5h1Jat��)�/����I��]�_9ÚI"���oh9�K}"�<y�.�`�E%d
�m�\�C�C�*���_��~r3;n��o�Cc��sit5��W��ʱ��ԯ��ϝ?�4bI��q:�����3^aljߜ;$ѡ�`�Z��#�����k��Ͽ��~����u�G�u��S��?��?��S�1�D�
�b�UxSi���	R"��jkk����"��5��oPR_���2���������
mN�2�x+5J��!������oCG��pB��f���U�u�h�akXyދL�鋬�h|>�㎏Ұ���$��W�v5G!�"
؉�پ+���ܕ;ٵ�f��.a���SY�x�9�m���ܝׇ(�]��'��hicp���`���6��i�a�ޔ���Q����S6��`�/�׷N%ʐ�U@2��)-%��, �K���_����RR(f}�!b�OGSWW̬,�u�]Xy�dυ�_�����/�A͑QqU��]z^�¸;�]��;��;�\L�'�_^�"�3ê�G�vU	���m�nOJ���N����{�׹U���B������l�pa�)#�%�]�0���-G�W�qQ{D��aUjZ�"�
��c�sr^�TM��!}��_�0�I�q���մ�E�YB�l�ph�������?KI�C�&��6'j�a���,���Ǣ򯾝����.�X۾Ţ�+��_)���?���`Ғch[�j8��<Nt���*g��1g�۾�Ms���W�˖&�= ��*��r��t�TX^�/j{7p�(�كId6��u6�q�Y�uy���
�2y2�B.Y�r���V��l�'sEB����WJ�?ܦY�*�O�pV��y~��[��(�|� /.dj��4�p�~�.�*�i5�4R4���q���f(A���ލ@ ����ۊq�{5@i�b�J' V3֐1/.����&G)�Vj6��M��c�
r�@��|2�+�<+�:M�&+�>�Sb���b���r��"��fp9�D��zz׊���)����:�߮�j��g��S����A�ul����gN�|�f��2�G�>�����?��rW����4�����&w*�TͰl[������WB�#R���r�&*~�!,���m�G��-���q�����>��9��r�+�d�bX�z��sD䒈
m����A�x࿥�)b�%C7,�A�@���( ����N�a	^u�D<�zB�!SF����u�uo�8����0"�I���ZU��܇�'��W1fO�����?7�
�I~��^���r]����a���Q��XGt{p#�=�>��T���%{�7����2R5�X$g��H:�:�U�^f��S�z�T����n�?ڑ���Y����\��U����	G)���d�v���W������������������x���~�ѯu�Mf+�����0p[�p>˄�~U�w�@��ͫ��PhV�ϐ8��b�b�
���Da�ZO�i-y�m�k���"��
~�yE˓A<@�@�4 x��,'�C�eg< ��N
>��m-�X��>�-WX��$j��w������Y~;K|uO�_v��^A��[�N����{"5ڗ)�����׭[Yt#���X�.Lc�!Pt(D0��#
����55���!����l��T�x���~��P�	����(t9�1R�G'B;C�ۧ�����̤�ٟ�����+;s��������%~U�W��W~�~�M��~��Ez�Z���L��G�� d�~��`�'�>�"g�K٤�mU�	�aTu�����1M�X.��������q��<���|�w��#��R���M5���'�H�Hμ��۷>�0�p|̴2:n\��8����~6*�҂(��/}��B��a��bF;_�8L*�T�Z�
��R�Z����A��V)# �((=*�2k̠]]K�);S����hDF�C��S@�M�Sgp':���j732.��j8R�������7���@^N��ֵ�vLmw\8m�R(�<!��kz�剉O�������L�5�������LP&�i��!uu���\�2.�I���v�������E�>� â
ՅLLs7���%/"֋�

�������z�a�,��\�rk�f�o�ţ��[�-��!~��m.G�{u�v��w��,��%/��Г��-��|u>�X���f%�R��jެg��}���t�5�S|����=�Je	�{%�@��۳�����Tb�D����-��h#O~�vur�3���eV�1)%Rj���������Ͽ�>b���9Eg���O��M�|��Y�gR�����>&`b��~-l�U�}�u����憚Q����\���G'8�
&/��K�PW!�s��U�s���S��%�	H��"�B�׽$�g��p�J���
9�eMB?�O��nz��ē%PA�կ�����di
u�*�	�ob���{.A�T[]�]97C�a�'!:��e5L�9l��<�-h�I�s�'�ǒ:�=��.Ε���q�eJ�-�s��ZT:�oO݆����y��%M�7��{�>�,!F�Te�K�'ʘ���h�D3���W'���sr(�������q�d���r�jN���?lQ�vΫ8<�8Ai[ϟ���¢�Y!,��_�(���"zYlM�$�iWnz�+�+�v��	��i��]��#;��Y:m:��t'�57Ja�3&�����2�f�Sn�&��e�{o&�eS;��4t�(��	E/~^Gv����>�Y�$W?"A�?[',W������9�C�;'�M��踱�V�%i�3:\��?�����������)*�$)�h6TV��+J:k#U���Ů�m\9��y��F�RឪA%t�D��C��bBRK�1� � 0�G����wrf���w��!O)����oc�YT�(:	Gz��oF�k�z�#��9J>�W�w�y�ܮx�k>��t`�ki�oI��
y0�� *=��p�B|��z�Ӟ`�_�f?�6~�y��HjY˚�@B��?��{T���\8�w�p�����dCAo�8�2?�FO&[}�F�쫲�|�)V���I�vҨ�	���y�0�2�(�����)�)&�k̼�H�.K&NT�6.[�>c}�LVv�'k��@��gk���
Fه����HI��MN���|rG���m"F"u>Σ֩sJTj��b Kܠ����f_"%<�3n��I��F��&O?�Pb��H�;}��i��&"M�u��'ݪŤvE�6;^��?��1�h7��ZK@]�h�vˌ��A����B�J	)���0�_���q��{7���5�Wǟ� �!�q�H��J/\$�V2�IRO�����f�/�pf�8�k�b-���/D��ss��]o�.O���&3v�Xֿ�Ñ	���A�$�IG�����O�<���d^lR��I��%�����,��袭=xp2@�ஃ	\�w\Bp�����;��%H�`��{�Wߏ��U]u�t����{�҂�I/|�?S���"U����-��!��C�Ъ�M�+4S�ս�	�	g�xNdI_ů�;_�.�5���Ƶ�m"kw�n�~{�(����?��}Sӆ*ꡥ��d1�^���om[h9�=z5����hr�%*zL)x���/ȥ�bmF�QA�U�W&�+fϐ�]0a(�%U�4�M/1��UdǤ&U0�# ���e�L�u�)&�j2+9�3�.q�l1����D��v��y�F���c��#�69���j���W�X�� ���^��+��c&���t2�F��cH�@�n\]{_9�W<+cs�6Ɔ�<�c��E��`H�:>F���D����gn8���E�ՠЬb8S9Bh{"�3���8z%����]Y�4�caᾶ������$\�>���!�̠O�]pdFv�e14rwFH�\�T�)b�q���в�kFnS#�0q�;�9k�T�+)��08��^��q1��oV$��,>�L��M7�#�&��� ���Í�wY i��A���Ղ���W���P��7|0�yқc=P`����B�Ӂ#g����r+=4�M]�E�����`�7�oKUN��w⪀RRݯ�r�����p�����B�c� ���M�
T��Xp��~i,��E޽�X_M3^����;*G�*c�#:v\�gK~b���(��k<"���bA���a�:����������/�'����-�ffSHHtto�f���$*�+r��(�v��_�_d9�N[/}��K�e�&Y�.g[h�_hWx�)��q֍�CT����~��̨)���ю�	r�u��^���'Nh�Py�(r�)ق�T�#����޺�g�����/��G���4�&q�/e�ێz1�H��23z��@�+C��<��t�@?�����aJ׏4,f��JU2�k֘����`����WO��@:a�ՆbU�>n��.!ٺ�t���.����Y���z����@Nh\R��P�O�z�~���A�PC:�̖���B��^N�2X�lL�A��X6Q9셄; uf�Z���L��J���
�49x�������zyC:n��Ճ�=|�4�F���U5���io=hKddv.Hk�#��XLf8V�r�;Ѣ�^?r���(]Y�sm�.u`T8B�2�,U��4g(t�d� a�uE��Ҝ���	{��h_���o�Y��hv܆7���H[��S6v���
���%ݔC�C����p�UBp�J�B�
}꩗5�0��])��.Y�$!��!�%�4e� �HmI���<����������~R��ؘ�Ĕ��=j����m2{� Ղ�D������ _[�h
��j,}��[�Q���%���Z|k�[)����6�ʞ���[�	:e�7Kc�VE�b,C�I�°�%��^�&����j<��W�ɍ�)��DZ'ls(<�(0̴.^�C�&/�q���V�b?x�]���; ��l��Pb/]Vs=�|G�� ��W�~��]A��ꌃ��S� � {_K;�:[:9{P[iEmaS���h��\����2�oSr�[�I}I�J+F�]"!�0Y �*�x�sTkb��D�T0ψ=ؓXg��� H��7��4���Y �拀^|� o�w�Ύ��?���X�]��.��L]�����&����o�0�3�ͷ�_��U2�T�����pXx�4��F�w&.wǼ��>ک��5O۷���~���j�W
W�_y�Ӎ�S؎���J5����EwCw1����;�;/�m,ݴ c#Y�}�IL�(g�a�7�]����|yG���?�QWmXj����X��.��Ɯ��5��S���BB�m��W�TwP��/g�%��&��7�a�}�}n9���̑�*H0�_@מ�|�}E.i�n
�?�X���r�/	�ʌM���W��D�~�݄[��	1�L�w֍{hQ)}��n�{J�S���g���)�����]m��)���$R�@a*r�,�$�������Cv��^�h�$AG��Aw`OmҬ҃����'y(�I��"��3C#�������n�?<�A�x%�`�p�u�]s�h��!D�oT3pOzkrmo:��1ɯ^���x+��L3��K٢λ;X���e3�*ϝ��VnT��n!��ASY�j4�1ή�o?�����n�M44BN�����O^��=s���`�������čD#�kKmZ�*��A�!����ƨp"�5�<����w�=sы��;�@I�k��3�����QSC�>�Ϙ�T��6�����+/j�qg�\s����V<����;`ۓ_c�#�������.��R�A��W��^�Hx��pԟ '���5��������������L��>����? �ϵ�ۂ~k��箝�#��q5%�"1�Rņ��i~����c���Ϻ͟����[�*Ӕ�E1�Ucʪ�cN�η|Id�T���|�D�v�I��b8�N��з;~�{�~����_�(��7����%�"󬐥����'#'Vf�Aq~��j�� �*o�����<|�J���C`6�c�Kց��B9
_�jѧ(U�aHh��h����sq��QQ��PZ,�;c`$���8mxq}2AA��F!᧮�§X�>+�&���	U��b���P�t��$.�%����(K������ɮ�		�u9�W�C��F?�xާ(�l���.*hإ�(�j�-MNݐ����t��lg��8��(���Z2��*�$����g�}e`A�Ũ���б2�Z��������õֵ���}�g�U��\4�YS�|�E8�q�;p���`f.�p�a��Q�:%/#�BE�<6��[��^1�$�GW��O�.ކ�%K
�'�RP%�Tt��}����5Χ��� sº���!6���IڕO��jE�`&��zp�s
����l{��;�x6Vsþ��6~J�z�S��^2�E���2o���va�!�v�e�!���'�v��U��ɟ�-���ߨ���+:����Km,0�������!�ɚB�M0(��p�f�[IhKE�E��,���;^�|7�u�V�o�UR
�������9������]���˹@�w�]�$�ũ���s�T�p<Uۯ=<u��8���q�6��՛�&��-��Բ������,�l�]���Ɗ��P�Ձ8k�\t!^�E�JY�9�\N���%�Lg���C�a��`"_Z�^L���MlI���AoV����*�؅ΛַX��A1L�a�%¡�2z5��Y/���EY`(������vɏ���9߬P뎍~����i�eo��Lp��� �MnY��kR��#�}դH�.6�'��]З����%aj��ާ��Z�Ac��<IQ�����-W�Bc�σ@٦T�M� �t��?i9:/�*��3n�]]k���3Rھ�� T*i�r7���)aЛKf���pP��-�a��8~�vk����:�~�1�g����++�@�L��$���,��KNbf3Ǔ1;�[#�����J�\	�������o��W?|l��U2tQ�3�WPV�#�{|�gV fA:�k��G��G��ky��MÝn�Z��I(��B��'� /��"T/l�m|��M�ޮ�vP��F�h�Gwք����\�ut<��`�TR��n�]0��Dz��<6��er���eT��'n�q=�F<	u-��i�fu�ұ�3��.��s�3���R�^��.&��Zo�O��>	�Ix��`�'&��(v��}MuՉ�H��2����K�L���{�ht(��´�R�+��I^�D�y�fz�v�"4`&8ɿ������&��k:O:�\:1���S���0V���c�^�Wǲ��3z������R10�᭸&��v}}=C�z�X�Uq�Ѱ��Q8&��L�Ƞ�͑J(Z�x¥�Y��rp�>�g[����{� �A4t|��E��l� �p����\�B\��F��p1�@d+u#=�kc*�ۏ��1I'��Bt ��e�) ov�W��G6Z�
�v*'7j	^�:h���I�L'�:�%�N���a} ��U���whU�b���h�ȥ=%7#�,���Ӄ5ۛE�/R5�r5�$R����?��F�%Z�@r{qQKN�KG���tM���%r�H��|`G�����^��x��o�L�wD:��P�y�󫧛�������:� ��+�\v�c���7�N�^�c^�o�á����r��" F�pL*���)�>��Ǭ���l�S��*r�"�I�1	k-G�&X<���a�������rH����ƢQ:��Z�l���P���5D�x���.D� �SESKx�lz��
Ѡ9�K^^D>b��#��k�Oo�dp���>��\�z#��=�a1�w�o{ww}+E־�W�&��vW��

:=i���q0�pw[Pr��{vi�߻Us��s7��lN=5���À5�J'�3���鄄�ՌAR�h���{�-C�=��%c�6��5�o��O�NV�S�!�9ɝ��S�lM��R�9S1'剬��R�Q~�ɞ�s>	�Q�Ww�?f���m�+���b=z�D�-h�rL&P�D�xJu	k�l�Xb�`0�Նd%Ъ��}��� ��pVMH7�ed�.:�4�h� a��d�����Z�ٚ��x�;�q�k�h���uw���ݏ-�Ƥ�� ߠ"?�6G˦`�ݳi��<c
�u�O.k�ө��O�U�D�W֛�5�՝�_������+BAf��b����΃���ձ���,2pq���i6>�a��e���Ah�e9��gLN96��,-W�H�w�+��EB�1��V�V����/<D�լ��L$��K=�m#:kH�ȿ��*����K�x6�a�z9&KFity����խ?D�ė2\�}�;�B'�_.�ZQk:S@��m~\�E0b.�L�=ܬ�Rr�E��ჟ����k;��D(��93t�|W��2�(�Kp�N
`/�茋���GJ��މ�d�#p�5x�k�sh�B�EZ�H�˪�Oۃ�e��%�E��@v�����..�_O��{�\Ю��h��b�D=����G����g��RP�ޑtڃϨXd`��"��P HLYYM���e���ƻ��ԭt$-�����#8ֺ?��{��"��jL��0>�:s��V߼���k%�W��2� �[�0����6f��p�K�hb2M�amSb|��k���9ң��r�b���t��L	�e�َH~ݣj���/SFm�	q��P�}M!"[�,ۂU���ݾ�_��ь�g�p��YM�r�4w=zcT�?uu������w.r�C�b{ٓ���*Ir���Q@t&��Hiv�K�ʏ��eTѬ�J?�ǫCR?�!�gk�� �e��M4BY��5XF��"�PjVw��|�����׳2`�R�eL� :�0 �����+����\͌W� !;�A��(FtY{�s%���m�toz��� ��!ߊ[�i�H&�Or�y{�厺M ����o�]������0����J2	���>�%�ߺ˴�;�]����JeE�͔~�D+�kʄ�o���xr�\<��Z�c�_��4ը��Uy��򲥯��2"N���WT��
�{̑{���K��ӷ��'&U��*�I,Z5vW�� ��Z�c%���RP�}2�CF�V=��m ��r�� �!6.���\��!!&��_�x�zju���A�ّ�c[�P�*!5�YMB�����m�!U�O�������vN{0ѷlFHΘ���8�Iv��R'�Q&��k;i�9h�;�o;$�����ӌ���q�H��m'�.JМ,c�Pj����慕�s���IoX+�'�p`����Z�l�Ӎb�V�X>k�6kйcs���Zc]�JT}X�� 6�r�q���1�d	9�|�Z��,)P��`�3Л�f5Zd,�iWs7�na�^yY}zn�I,^Bm�[|G8隆��-&�p^�g�Z������g)Z(����	 ��)�m)�O�Lz� G��t��P'�鏒TՇ��J�#  �6� �RA���B�A���춟��)^-=�*��]7�E�zs$�"s=FF;r`?S���&y��<m2��(�� �M�'�
�)$�m˥�fC�N5ٲ�]��[���32��%{���o*��X%�Y@�a�b��2���ӓ/���ik�M�����>�	��ZYG���>����(2S�e�K���e�	w��^ U�dJ�S�4~Q���C��8�AV��˂�d�����ܩ��L �4Lب�̅����&o����b� *�6ě�i�$���24#�D�`�c���x<d}�r?���q�n}x�<�Cj+�y�8��E�;7ux#:�-a�U���)��`�3��z��5K�.!��7��zC��D���+����,�<ꊁP��ˬ�"w#@� �x3��=�bF5d��&"J�D�J�酥4Bol��B�A�#Wol�8�3�9�M��`D�L�W��	M6���ʷ���W�)_)�H��ߋ2��d�j�����	�M�R(�"�=�
��VW�ڗo�-����w�Y�0C��F}����j��Y��A�6����
?%D֏F��y�2~���&��!��6~��ԯQ��AK���˿b���6�P��~���h����U`�8�ݯ�"��j��彚%+/\ﰟ}�,�&�@l0���sᕷVP��8�nL�wƦdT�n�R�b�4��O!�� ��/VQ�f� 9���õ/�E[Z� �`h)Ĵ���[�)�L��R`�h\��"��;w���ߟa����"����݄x��.0�,��m_hn��M��~<f-��ο�Ģ���0Pt�=���>l���!���+���ٳ��Yk᥵,�u�p��ҋ~8n?��;�a�p��^2�!X��f��#[(<V��>��ۘ/�숻�{�$�R�1<�"X�?�f<�ٴR��M��)@�ZU��-S≓0��c?NÒ���ㅲg�`������!��sk�<���]:h�t��v���H���8�#�7(������x����Ŵ�R��9&���ZAR�@�n&���O]��vq�8�D%�h�j�l�\#�W��E��b��l��J2YU�ҝ�n���kW��`2̭K�י *Ag�5
Wඈ�q���q���߲�ML�A/O�0���Ρ��:��QT�/����k}=gF;�[����x�굱۩�bt13�z�2v���jl\�Y�۩��T��	���zaW�w�o�ON��a���1XK�J���_�|�
G�F�|��z�9Ư�^���y�T_̀��H#���=^Y���`�A�%��Yo��C�X_�H�����(�K�W�vf�S��7FU)t��;{`t:+��i�N�ح���(M����ot��mM�;�KE����\�>��ux6o*�wv���v���)M!\,%�E1�X���� (aOyY4;����2�bjP^�@1-�q�b�9��^<������:��ŗ�T�e�K^��u|��(�0n�(,c56a���q8��ȅ8��F����n����o�swU�z�o�*����>��V�iV����dQ|s�=��v	j�Ze�*��)��bě�.�D��}JcS*�p��O�,�Kb"� ����҃��l}���6	s��1���d5�M�c~�+M��GUn��Q��d�Ds,����V��6C�d��z���˒Y�K�祿�MleP�74,(^)(�ҘNg�j�f+G�����ν���+�|��	/�z��T�0Փ{��Z�g�ƞ����ǯ~���৻��$��2��9��W:��O4�l���Q3�.��ͤ�3T�ه3���MJ½ْWS�c�5�`"C4Q�J��hZ:^��������X�9�6�æ�zGn��C��p&���*ܫ}��[%����?P��A4��u"�
��li��	>tR��x���r���~7B�.��l:*�kw���'X3�\�_���{;��:ImJv�_���.��A�G�z�쭎WԻ&Ţ5�ɓ���-j�B�F��]���(�_Z��@�:^�jJ �!N䴳����)G�p�gÀzDx�_�	��^�������ewme���j��k����ro�z����F�u�R�8���i����=��:[}�t�?)�--����%���q
�u�_h����P���p@�����j�j|q-�>��N���.� bq�r� ��K�?�@:�Ϝ"Tzt��L�wК��¸x�ᇡ�F;�����hHn@;R�8)wxe��ǩ�	V�m�aEa\��0���1�,�O��~�<=�?�$I�~z�C���w.BcT?�RS�d�^���BKB�D�f�'=���E�'M��x�P!��IL��"4

��E��?��douv��v�PL������D\NUB���@�,CR<o!D#fY6���ǿk�2ba�7P�Ic0%��f�9�
��Iz��	���;)ח�mU�P�e�Q]���̌TLR8t7e(P�h5yh���h���,R���4sݟ��~m��澻R��(�Y+l�F���ti2@��U�]�"��̭s!�~�~���=�{�-v��VȽ(��w�tG�sX�n��ӂ^�>�R�om��ڻ7����CXܟ�85=�c>����˓�d�������b4L����uy�*������:������u�-�>u䷍�������΁����J�q+K�}ٶQ�9߽T$�/(k���7��Tw�[U[68~,��+��������{Bz�G�I=�>�,�<�N<.�<.>=|��w��Q�-��#��/��6xsT��[�z��'0R�!,�����
A�D���lZ-l^�Z��������S��J�(H�NY�y�n����ڂ�ֆ&�R6��u"D�v�L�%���Ɇ ���j1^�@�shP�#��:ε)�+���W�O�$s�����G���J��������������S}���}�6=�+{�����˴�oRR&���.�'���?��9�mq**_�&f���K�D��\�%2y�@����5d�BÛ��L��) J͗�'���<)��V�s�����q'o�<mj����Y�^�WO��S��n}皨�|J��|�$�Ӟ��V�����@b��_id��ScTT����aA�_�KyZ��ъ��F�3I�ٙfO���ZO�Z�mBD���s��+~��Q�3ڠF�g׫�j ��9(�F� >S��{�)��o;Y%�9Z���FH�B*C�v�>�n�E|46��K�g�O����ǲIf$#1�I�@W�Ӈ����x������� _�]}���"�o��RO�LH5	^�Z?�O��ġM������2(��bR=����"��)���{3ձ�m����w���P�B�?\ē4��xdK�$D���f[�r '[j�Tx�%}���2�x2���](�p��c]��A��$@�؇�@LYf��ЊP��<7��qo�	K�C�s j�h:��+��hZV%FeM�*����f�|S<1�J��f�:#/UbT8�bl?vG�<qASoM�(�䇾M��(�S����&6�0"�����5�3��ӿӣa�M��A�B�w\4{���M��	Ћ�����Ok{�cb��9�"R���<
��	���׏Q0!���+4��29�n�a��ʫ�V�-f�'%���J�Fw{�MA��b�Jh�]������ruL�-̧|<�޽m���_���1�"�Mcb*�
�\b��6��P��8�F���X��R!~�����;��`�C�pF���Wꙅt V�Yw<��L�p5�����EE�������No��_(2�3ƿ!���R2j	\�L�KZ�済;U����w�:h���o;?br:3�P��߲	'�S�����#h��#���h8�=c��eo$&�u����,�/K�p������y�w��!]���dt�@c�8u����Lv�VR\��L�v惗kA^=���n\ⲟ�`�j�H��"@}6nB6v��L�����p��� ϻ�픨�u<b�����)N^��Q� ����6�7B�뢶딼�FrF�紋���߭��at#�v#<��D::��:�b;hd㻪�{�K^(�M�'[�Ep�L�``���3�9g'����@ 4Y(#��T�+o�򝱕;N�1i�>�=8� ��gv��Ey�W0��L�c~`��T�����/̏���M�x�jJg�wLyRFצ%6k�7mpo��i��E����ft��f��x8��q��2�I����{�u���u"�v{�m[Rz�|(#ڋ�D?�P�8�"�7	�3�q��%�Ш2�Ϣ΃3\�E��k����/����)�cK��H���_��%XzѾ�n�:Ϻ�E9��IDh���L�+n��>�(��E0�5'��������٫����:�Hɢiw);i�)�?5����W/�?��0>�NչST�z�Vȋ����HN�Fsc��;3����}���lJ\FXG��h�RR>Yu���s��Tgdt�m�l��7:.�i�1��^N��7�Ӣ��a'2�*#���Q�N���CB�����S����]Zn��Z�+�c�&;�ޛ�'��jjH�E�?�^~�zz�s�t�h����u.��q/�Io��������ʰ ��z�"��S�c�z���!�]�Ȯ�ܚ����tNZ
�R���Ec�{����J5[�ܕ]26$K�Z�T�7G�;fA<�$�_��d$"��n�e��,)L*Fy
��?���p4���si܎Sv,��Y/p&u��=�1Rө�<m��5�����(�Y7��:.L�g�K�J�o�D�
�� ����5k���{7��"�Lأ��k1h�)<������J!P0�*�\��PQ��B�:!-��}_G��H� 0Y����'|�0�i18��_��X�0���� ��"��&>ڴ����U��|R��%ЅE��v��Ӎݥ�[���(�Tq��*�@W˨,dB�Ũ冑02*�� ���)|S⧭8���.8t�;pj�t�f#�-����j�ά�6�LI�Z�O&21�L1��Ն�����X�<6W�}�u;������MTc�O���NU��d��N?W��TG>᝶�P��Ӧ�G+�m��|
-�t�گ��57��}'��A��I���'a��c2�[4i�jA������`яM͓���R�V��[�:|�*���=�_��J6	�yy�u?oβn�\�d�����rQ"�Q�ujj+�X��4� �9m�����u��H�|}�'�ʙ%K�
�p�S*�D�z~�F�J�fܨ�>ŪR��3��`�Io��18���"Z��"�y��F��"�p�s6W7�+;Oŀ��-i�vN�-�6��1?BB]�;��*B�f��H����Ky\�E��!�&�y�m�lm���L�1+,�?�qD�w6oh�Q������~HZڝ���иJl��ח5�Ui���	ǚ,�2�\_�c%W��م�, B�GB�}���Օ?8��ׄn&j��{! ����zs������Vm�f�4Y|Q�5��_�莆��lf�Y�C*�p�C�-�[��r�Y���O��A�����z!��k*�3��Q��{hTP��Dc������F:k&_�O�Ǽ���J3�i�>f �z&�gH�J��Z�X�-yy�ǨM�sŜ��夷V�#,Y3y]���`�c�	I��b���X+ܧ���yU�q;`�]�MiH�
����
g��˕�S�>o��R*�����/-�Ҵu�m������3���l����H����J���q�f�OT��	{i�S��I�JaP��W�F˄�Z���4e#{���!fJ`�Ls"k��{E�'����';��P _+ц�����*��:�UH|�I)�{\~K5w��s�pu��.�	���[�qUr����q��]�Z��-���g��޴�k��ֻ0gf��/�C�{�H/d�n�H=+N� n�E���?�����R~�;���'�0�1�g�\��C�a���l���c{�P�l�!n�<�0�P��_��Q�0r;�0~kw� @Y�Q)��07�ɂRl#��b�F����ȇÊ��ى����utRmm��_�76�ܞ,-�i�"as"����/��/�+��|d�L"��b�W}/g3t��P���l��Kd��+���f��_`^��,3ӉN%I�ި����?�7}iT���~bUB>}0#��6��"ű)��m2�Ui��AG����e��"<��(��⊋�����t�գC�W�^�p���c��i��t&������N㈩��:�Q�։�-�
� e��d�^�ϋ�&�V�����o�s�r]*�a���St��t��t�e���	�(���ok!X�K�I�rj�p��N��Ql�����r`m�}�����]�n��@]�:[j ���(�:�Sp�W&��ɧ}��n���c8�z߲�ǹ�T���V�j}���U_ٚ*_�|-l�5�y�r���������ˇ4���_o�Z�~� �������_@��H�㯣���{Or�?��>�I����}�
��Q�t��6��6�6>l2��?�ɒ�,�,�c���t�3�4<+{:[X�n����C��XN.��\E_��'�ޤ-�=㋣3Nv�a����HL�&����5�H�ɓ{�&;����ëWNR>���}S�-v�t~7M��?V�l�4�ߗ�O?UI��������ͩ�4�RA�n�we4�������|p���E�|��w��A!�4�S/Ȓ�T�󦬱JM7�H*��[�$��sta����g�@z�a� �����C����B���D���|��D�D����u���l�h� S��Sn�d[�,X���\����f�ٖ��6	[���lm/�a�U$��h̢�zv��8�U�[��awqw��@584���F�߼�ݞ�ꫮ@���5�:pq%�n�3!��
\-J��Y�u4'&�~��A����?�.^���1\� �Hd�9N�6���S$	��qhB �C�o���2��P(D���O*ld�k5n�,{�D6�f?u	H$�2��9���M�<�����G�����F�V��&�>��TL"�
h�L�?��y󸴯�tp�`?�u���b��eh��)t���K~-���#WKX��M�[���yA��]A?�;�MN1d.�'�1��ٗ'�Re���<�A��f%q�ʔ�F��
���i�DB��w�jx��a�A�Θ���BQ"p%)�<t�����H��׳�"�-��q���bS������b�^1�����5����0̝e��χ�<S�CJCr���J�;��z��0W������`1G�kJv�J���/�U���O�,)�H��!fA	�O��N��	��w=7�x��p<�f`�����IR�(#���pn4Ǐ:U���	���R[\V�j��"3#��r���J:s;�Kd��?�M2�ybI_��xY���o(h��u:�a�_�G������o3&`K�v�v,M��x��?�"f����C����Q��1X��e�F��i֜ci���w��-���g2����D�rRiLR)v���b[7����w�Μ��!i����SS�=x)���?��I�KN� �}�pN���fω8�3�;�r�=�vpa-�x53�Cn���w�x�~wS&�����U%R�.��_tG·�(�"��Gx�\���_�:)چ)�^C�����s���g�?B��(�� Z(Ԙl���Е�L�Ä�-qE59D��ɘ�C�!�u�@luuH�lt�a)�?����D�`��bԯ� �c�C)7�Z\_��Ix�N�g�	�_�@V$��E��J9/�M�>�T�\C#:NR�T����{^��.U�e�;��t؄����HmɪC�L�}�PL@HR�.@�+TV���_,���q�,��-���y2 |@�?� 8�Ɗ	��u#�rz���l�/}��x:���bs^>�nkF~C
O�^�j�7!nW��\��?�(t��s�k���u"�ޮ�K�����m��H>��2�v�)	�c��PLjA�DB��?�n����=�<X���3�a��i��!�r�?JV��x]A��|�m�����&"ޢ�DV���Ӫ8L�_��h���1GV�E��μEx5u6Am�5kL�D̒��|�EV�j������Ф�����������E�c��-����Gm��<+5P3�Y+�l�B�)CP%u�`�Iפ�U�5�wP�^T�Hb��ݽם#%��oȱl1�_X�1�Pp �λ�\�:,�g��mE+�ZnqԞ��aR�	lCh*��F�ŽB���F�E1H�!��1�Xi��=��/�2�2�406 g
�^����ђؚ�#<�eJ).=�Fu�v@��1zv��/�j���
J��p��.��믋�;����y���9l׏�`͈�g�\�y~F�4���x�����0$������ƳnV��<Pu�B}:�K7f�0�6�2ʹ�Qg��K ��#����%$d! ����ռ	:9t���_7�_) �ah�ut�%3k-�0��"i,6�pL���O��Ɩ����OouSf�}�7��;��o>Y>��/��7=.{]t���]X�HW�z�Y���;'<T,���=݇y�m�������y��;uw�UϚ��������Őҍ��M'i��� K�nϻ��ϑ<N�uRM�`M����)^����z�e�6���1x;���rd2�&%B�c��wZ`(�اak�a������}��c��=唐��aH�5]��,�l#�����#2�f����p�}�����u#�X���J�Z0�`�5��;��tĮ ����I��SNk���۞�>;���G���jq��_�u_f���p�m-l����f�H��2f�
Y��'�Uw��N�V�W��,��o&h�;<s������^xE�,2���v�f,Y��j�je�r<����P����u�ܠ��\.a:�Z��9�կ7{�6c׹?�?���`�nE�U=�_�+f�y\�.��Nz�u�Y�x���]F�K��H�f���]���B��	G5b�Xx,q�{��Z��E����;�4��Ieg���:��$<y����T0"�ny����SC��7v���I���b�l�P0uF�lK���R��3�Q����n"`�	�O�B�o2r�϶�_�Em^�S~�h���q�ߓ���ѐ��7lR&��U��M��,zW�=l�Y"_��/��^��g6�p�y��V�['\� ������s72!PL�!�Ռ�*�7����;vP7���S��)�c!䩭Kf��j"z�-�x����v�U,
��'m�7<W'Gd�_��:6 D풐_�>�BAzd�F��K1�l.5�xl��u�PMl��������!/�������������\�uHĖ������yC��t"����B�O�o5u�\��>�X�(���t֐�5����رiL�\%P�g�.�I:HR6��+q<)q4�B��<E��]���֬X]��dR�EF��٭��T�{4xǪX[�-�-0RR��m�}Ӥ�teI�kyM��-��t柳�!��5�~���ť���v���:�L�$���Pc�r	�>Ӝ�*Y_�����S�,c,r@���5��v�E;��� >@��E��;PGAf��$mc0hPŗ�F�ˊ]����vl��)�тjV��2噥���H��5�v�Ӆ� z�y�8wJ!�I��/���&�g�Fs���>m?X=�|�Y��M�7]?¾}���kd�7���.Q"���闁x��r��ˠ���N��Eq�W�^]1m���ڔU�0����]�*�1*��މ���<��L5DFCbj������&c�� L�b0ө*k�/�Y�S�`�P�"���ɹ,�V��΅� N�3��:��k$�ͧ>}�T��h�Ω:-�!W;n��M�O�M�G4�6<����]�R���q�$p������?��V4��A�m�9���į����[z�c�@���!^>��f�s��oS=��e��#��e��*�1�ZBȜ�>�|��X� `���Q�8��L�UgĀ�H��ؿ�h;�a�ɷ=����D!���!����u��R�?zỔgdvX�B����9��C!��v'��&K�aOu����(Y�n͈��NѫEn��B�m΢�6	"|
�b�(�; 9.��o?G�B텄�@����K�j�e�Qk������&��R�
���{�'���0�t����/�S5�:"7���,�%�o�8��CPz�WF�����c"���^	H�|�O��_Ř޻i]�R�+D*�x��vsb�W��l��lp9�X��X,7����I���u�Aq5�<���w��N�K�w����	�0lp�`��e� �!��\��ϭ:���N�^��:�Ou�^o�=+	惐s5T!�r6�84\2t^S��m$
�y��6���ye��e+�y����tS�c��u�
��
YR���KO�K�jadyC�嶵�M^��)ڃ�5(X^�
���hH��:�_�{U]Z����ixx��}���+��*F(ἲ��9]NJK GuG�O���s����w���(���;��<����ӿm�(�/���/�(�b�/��k��#8��~e~��k��/���ة�?���_}���`V��.~}�-����ȯ�d���D�g���S�)S���Hξ!�������'N�0���Jb!�;��(��{� UH��[�O9H	�ݫ$o�PS�ؗ�b���/�+kh�/��7�qo�)�@�n2�ٙ�;�½)����<��֪��0Y0������4<[���-P�ʜ_�Q}���~��s>X�BQS翶ql�r�i�6·V���ݻS�tȾ��Rs�����13I�l���x'P- �lZ��!zjoY�dTC���n4g��/c(c�|U��r���@������T6��o�:ޱ���%��;�����oq�q�^zq|>�2�):`3q8!���UYE�E�%S�l�W�cCP8ro&	-9c��u?;�4}.��/�v�!�?RT(W����W�Y��]��CLo^�� �U��7r��U'c�w�PtE(_^�`�wd\r�Lkt��R�.��6Q>���g�v�ƾǔ��Ͱ�������H-�LM�Vo$�u��u6��|u�/&:l��_4"��5�=mpu�,JE�
3K�����D�z-�l����|��У��*��&�v�)�'�~���a�<�4(�t_��AS&&�����
CH�S�=t��!�u��[0�Fx��ʕg]
.�H��������3��|5H��TJ�f�!0c>���%zy#�%����V�z��^�۔�-�lg��]�h;�e?��B�(�K�o!a��]�����D�z?]~�x	Y�>�G'�F19��dڌ*O�x�F��٘����ۖ6�RV �]�#��pZn=��-��2R1ۚ��6	�'���f�b>yK�����oў.f�Y:��(�)�^�H)��� �´�%���;��M�͌�vYޜr��>f�^&*���^��d՘DF�gS�܀�����q#nʚ���rF� " ՛ۓ�&(%�)Ӎ��!I]i�`�%�C�1�P	��|ϱ��Fbl��2�,�Uo+ӝ�V���"���\K���xS-�Z���F<�d��/���H�j�����d��Ķ?�M
W�{�4�=�c�E�Z����&ґ��:?T��.�w���!d&e�}R+����]�d�����"����m�,Y�㿃����?���lLsl��gĵ�k�j�׸�~���*�"�K>Лpn�Y���� (��l}Sw��aFa/<o���נ������y���}��󿞁_��m^�n�M��ŋ,*��(����q�`!��Y�����T������͑��cR���L֪a	�VA�ƦX�i$�~A���Z�nH���nf6x��yL�P���I��P�B�6��,XHv�ge������܅z��ef�f��^+��n�b�M#��w�L�Wth}k�)4�ӷ<���x�MdX���'l������)or�E�G���FL��5Q
�T�.y�@�M���ɛD�T!4jkE�@��qT]�ckE�Θ0�I�P����|c|��%[��y#Ak@�D���aM�ͭn�m�)p����H�?�8�)��_�kk�{B`��<����Y-" �t����o�N���ǀ��*!�}i�~H������v/��O��r�{��B<p�xb��ŀI��t�1��(dOf��jיr�pd����ɫ6L���4���'����D��m�8HR����C�5_~"z�eh��yК�SlUkΉ����@U���a�Wml�cnu7�v&���|��J�y��v��١��������P��������6<�F���������������TE��v��l��lsth�VIBoM�fY����Y���hڷ�q�����&VB�R���f
�I�Nܴ�?���x~��\pkѦt:m_�,KSl~ӬL��	�^a�k�\��*;x�ĝnS8�G^;z~��R�<^��K�e�>�!���o����r�����)���������ee���?��]�.�d��`|0�;/j�o�ǡ��A �so�jPq|�Vw��{b:y ���:y>�H��]��� !$T"��
dY�Le�:���k��ko��p���1/[%:W�.ل�����K]��h)X��)rR����	  ��@H����[WC<��A2^�e�^�?��ǣ"ֆ�O��	A�]pjN�=�0r^�)d3�| !���<�9?�QY��'I��J�B�x���}�l���(9�1��&�	R���&u��\l�Jm���.ͦ`e|�h�-���F��' ���=K^]ۈY�,��	.1)8���s��7	�&��6�_��@�m�
��/�j���l�s���ƅ��>o�%P��%h�ba<��R�SN8��9V�:�:�|طjv�Ł@xS���E-��q������^��9�7��b�wCI����+Z�����c;��&>��S8�"�2f�D�9fh��.L�F��;���,�� ��I�B�ՑZ��K}�F<�!l�cK_:��Øiٵ�v$�|�G�+���?G�����cF��|fn,��H�n�L����?��]�cm�$�с�>��3�v(l�Q=q� ��UL��a+h���X��'�.9)쀀��n:�Oa�����
�|g�`�p1�Gw�_���4�XLɶ��yp+D~��!J�����ٜ~�gٱ2.�O8����g[d�k`�� I3��U!T�'��P3L��������#̖��~�D���;����(��[�F�S���y+U2�3nG�9��}v}I��M9H �$��/G#^�����;=�$�Zj���y�����Xy�̢�I[��"-�YZ��U���t�/@�
�\V2��V̳IO&��@ ��Af�E���^
�l� bw�]�����bM!_�f�@�u�
T)=�=G,�"}�\��e�5����z�6�Pd�\�R�%C2C�v_��PR[�%�b�z�}�p�/�D��r������T�hj���$�
�R)��@�H���vT0�CR�5r+�Z�]QU�a�.�i#�}n�S�:�Ja��i�_������Dc��mդ�dj�c��%�w�|���s��͢�P�{?hiRxAy�v�i>���I/��E�:�����J��|�>��m"f^��[��$Hu�4q+һ�EGz�Ʒ/�q��$���s����3���P=8;�f�Jn�I �)՝vF&�y�8<����Cl��k��'��]��4�9�a[Y��Y��![�����e�^�?���u�֠��ǿ�YSoe�n�q��Y�:]�u=� ��S�䮵�����]*��T*��c��#�� ����!�ё!w��� ��v�1�-g�s����$�!�U��Z�sU	ޚ��m�1��r��$�bֳ/mpja{a�`���L��M1�*jzs��;"�x佬<!�~�e���{��7"����,���r2=� !5.9_ɍ�~�2����*΂e	��䖐���LAO���iS�Z�,��l�d�L��Bhb����m6$a5�G����̦��\�����i��q�)��RQevջ�j���>�&S��y͕y��y�����\��ZT�V�y�y�D�� ;_m�R�����9"�m
����`��ŃBAϗsGM@~>t\\�j���2��Uü�q}v���F:U��h�e�6�ZhUZ��{��EP�+/�}9���4��iw ��D֛R��}��q@�>	9y��N�C������:y<�5���2f#& �٨1tWoҬo����oD�1�b�):��2R���1=Vkc����L�Rk50R��(��o�P������`���~���K�1[���ǃ 2an]>���~l>//�N#�H*�vcz��P��E�@��� �I;��b���}�JV��_﫟GU---_a�-���Q�0����qr[�_���wHw����Wl�"��r�+����� 0��ju23z!�TsX�a�%ෆBCDI��\"��_��1�̪:J~�|��^�a*@�k�Ե��[N��i���
jKxJx�@/�EşL������m/MEC���������������M�	ûY�������'��9��i�q)JX��,%�ٟ\2��D�y���_�M�,��-:�k��j�nMJL�j]N�vA+Ur�Q'L��q�D�2u�I:VOn�:~7�ߖF�I��tJ0&����Dj��0�����ҋ�o![��l�3V�H�LeD�C��IX���I�\u��"����r����R�ԩ��/Z�\�����eZp<���պ�&OLi��k�Б�6��_i���]���s�Y�	J{�C�r<R��?�{�5d2�˘4d��h��	��L�8ܖ���!�y[l-��.�����ILR���i�'N�t�WG��W�伟����*�ؗ�hw��֋M��9���<S�����P�Q��*-9�B�Z쭌w=�8�5����
Q��@W`�tK��G��r5䘮m0�%	�:�$�s����x�(�)H}g����k��~��mH1�f�λ���rW���P]+`��eR��� ��j)��Y��1 ��l�^����Z��4|��}L���}v<��{Y��h���|�۬�^��:h���n���XN�X��cgƌ@tm��F<B�i82F� 
�~�B7�Ee��B\��Δ)�i,����Zj�W��U	М�-[��`��x/�'�����D{jx1&�Ո�XT����A�ғݏx��.��p��aO"������mC/�%�N��������n)�d��:͙��ٶ�|	��!�&g���B�d�b�bLy�.�Q�\�O[
ɞ\ ��q�
׫��wcb��Tq C��*a����^�HB�E���d��h��4��i�x�ޒѰH�3����b^ꎊF�,w�-���f�ND�MN�����N��J�����c�ZHͮ�ɉ��+��{xSR�w�w��Ǝ��^b��
������)\�W�ZܖD���g5�1�cZ5��@W�M3��#�`��*3��	nRj��"�ǾgD	kj�1�~Jٹ,�ܝ����ǣ���(I� W�سO˰	�3l��
�D�?0y{u����Ͷ��]c&�l?��Uֺ�;���v�Z[����өȵAOzC��1�t���8�=�R��p�������	7��Uo�
��)�M���P^J�t\m�N�8)^��~��2�W��Up�H�#"<CK��m�����p[�_E��@x��㰍4*f��t�����ϭ�ߝ���u�p,aj�O+�ț���ӫ�4�x[|w'�/5��S�t�������:P݊z&�����i.�kL.�QTo��N��N���2�xV�M��w�6ޱ-�Pa����Uc�S6R���PcJrhu�}�~ǖXײ�Jl� ����I=^K��!�caA5����&����G+ʖ�s���${�jjI`'��|v�Ӂ�0��9��<}�H�t���7������A��m� �r��77Ǧ��������������M�H�oC/?�!S��V���9iLVu�/V����!�Z�VjĂO|p�p��Ԩ=�D��ڪ��^d������3_Ţў�D3�q)��m|��bOW�u���l����̗&k���_^��gH�sj�Y��v��$���c{M�{L�Y������Kc�`D>PQ�#�x:�5�j�t��79:*KP W�Ԙ�m�H����Rk�M����"�K�M� ��C�5!hdY���{Ɠr�7�	��`;��q2�Ҥ:Ta�P.�D�8&�NS��4��ӔxŸg[�H"��qJ-�t��j�<̼v�L9F�@�5 =��7�?�2����=�\�i�n��o	�)��D��r�t5���5�˪o6j�H���ӌ����>[��*�^v��9P����ƯK4�&�3�7�+��x}}��ֶ�'VӒn��a����51�e`X�j��a���������u��u�?9��,��̦x��{�@o=ζ3��k�2�������[��i^���vL�𡐙�^0
�8cLt6v��w �� �NyU���6J(���GL�P&�Y��W@� F���%���Ӊ���V�tKA��TCRM�|7��a������ok�r��,�}�*�]Y�g��K��mI؞�����t�������U�����A]3���C��+�GF���ܜ�բ�Z�'P���gR�}���~tkW�y���_�)�_�O���<�� `j
e�OcL>���D� �q)��lh�.{���j��Z/_:\��[ $���������R�~o����n.U� �헆t�[��<��Z�U3���z��_r�Z�<'%'2gC���;�t�o��}g���
�ix逸������r��{�Z5�@�m�|F՝sp	N$
��P��>cPU"h���굪j��"��H�b����������.����^��x����/xx_͞���]0R��u�>���mr��nM�NFF>��������X&3�PrF�*92c�Xxr��[��$f��KE�ZT�(Y�L(7�i��Rs��_�6���IC��RZ��1�i�q�J��j�d[d2�Ā�gKJ�mU�4�L�BM��G��`��Z���q�F�41z;*�S&&(�����`:0oF�c�$����f�,�$"���rFMv����p����ɞ��
�*�	�_	"U�@��������L"Z6-�v�|�_b8?oG�x
F���3J�v�|>�:��n�L�xg����ek��QGq�1��"/��%�8{��_Ч��V��� ��C����5���0�V">�؛�"4V�4�F¹�A���cxk�����=�ҳss��~�䧖�Mv�|?��\4LZ��0�;
�KA�p���U�n�ov��n,�u��II�u������ֺt���d!8�g�|���ՠ��h,�Hփ���7ZXK(*��W'�� m�j>N�T� 6��x���i�Q��A>T8��4��+�L���� �c֣\����k	��I�"��T�|w��)����Ǩ�$�*B�OY�����
q%i4v��u����#�G7U�����}'�ƱMΰ�;K���O��'0GC���U�:�S�A�\�sQ��+\�9�K�AB����p��o(�I2-*�6�?9�L9��,�(v�,nǏ�ZG(�K��?k�-~=�f �`-2�Y{��٬�ڷ_��M�Ca5��;���}s}Q�si���Ct?��=Z�u;�vtLwv�,��?>8�/�-%��yKhI�9�t�T)�V���r��#a"f)�&��K��q'�t� ����t�ЯOUCPD�y������n�Q���8s�0e�f�!��N5%wk�����&k�P�$�zG+饡�"��x&Ie*�U%؆��>��sQuϵHsr�a�O����.�@iK-�'�z-N�X2|����i�]^��m,����u��V>՟|��e�!����<ĥ:f�l�j����^	�0�MZ�ڪ=%hG0�@{�Vb(����VHk�d^��ˮ42b�uNfT��4��GU�X7bYye3zp �i�~㩇�R����}?�1�a��Ř��9��ɜ��+�(P�s�"{�p��|���`��㌫�x�d�e7��প�z�O�|�['ˍ��"�E�Zh�����x
����xg�M>) I؍�`"cc��͌t�Y>j��������tVAXο�l�@�޿�Ǧ�-'ݽ��m����J��f�Ofc�<��j��r�2P���47?�q�#�=���f�l��4P�6�H�GS�g��`��/���'��C5������r1��r``|��.꯭����=����x�]z�ς�`�qf!��������d�B��ǅ1o�0bNq����F�*�-�.�����omh������D%����J㞈�Μ���u�_U��^u<no����,�_�ᎪX`g�j`�v3��&2H�l����Jmm�em�d�A]�����[[Ǜ�O�����:�����?��m��9�y#��\������nA%�TaX��Vg,Ek/F��V$�p��p�$Ɍ�h�Ĉ��t�N���Fx��t0�W}Trr�������D������'^�^�բ�����|��{��^=�ق�\��1Y˧4�!��G:�J��;7�}u�/g��v`j�ͮ4kd)�F"&��I�仹����H�2��s�!$��ɱ<�W�q"JvC[<�t �O�H��Q�DLF���Cƕ��^�I�����M���V�� �Z*�P�}ĜⒺ,�c��cR���0�m� =��Mj�����=���{+���o�����g0y%�����{d�y�זu��jI��j���It5������%���9���I�@<T���w���+��)8��k�M
y�Q�gJ%�DK���?-y�+���_.��;����������?���Mkɼ�����]�tbÞ"({�Y:�������t���JqJ�8<���fI0Oiu�I�S2+�HŚ�C$�C\]��^����Ӝ�0�l
:G��N"�/�ȏ=<��U\�SA f�J F������Zy�y$b�1�@ 
Q�g��SfX�ZS��ߛ?�[+�T�r31����`�O<�$����P���3C�/�����Bv|�P$U���g�����K�bm���L�u���@��Z@�7g[wxe��e��h����}n�<X�400[m'V��J����]�4�!2X��91s'�-)_�� ~�k�o�qWԆ!)c'�2�%^�� �%��|s�Iw��
t�1�E^;�]��yz�#��~����s�������wsZOW �AY��],*�*(獵=���+�+�X�o?��������t����"8&�:��ú9D��rtу&ӿ�f�ģ�*cM����|i6�Ѧ�iQ/ �w�(���9e�j���|��s��<:Q�Rj��>��f�3��\�D��h V	��D��3�`���_�1׭���[!d:�$���+��D���~�%�7�z�wf�rX7�×[Y�	SN���<a�Fj�3�$���Pq�Zqj�N#�l.�W�%o։M{�D/���Y��[˃��H�!��G��N��� �9		�a�բ�e���%��ͧ,�A�mel[�I�p���d�>@-��YL�z�3s��9�xW��9^��r���o4������(r�a\�M�M�ZM{V!{ �7:�� �����3�:Bk5n�@��>	@E
ط]c�iN���q7Bv�3���x���E%������{ϵ%�`0n]$	_l;�1�z��L�@3z
HNҷ�U�Mm���V;�)�[7�����u}Y?�H��G]�q�����̱��Uɜ�;b�|AS�.^[x�-d>�Dr��C 
펮��d�Qs:p����p�UxT�9�^�� N����&�o�E���}hG����a_aD��"A�������Yv�~syS.��K�A�ܯ��W	��=���[W.��@�_++��.wߞ�s����c�4uj�Y����(	%18��Y�qƃ��w��Ք�pŸ�N#x�.huOCx���A�S�Fg���23ku��|�J =G��Dh~�J�
�TU"�|$���K�;�u���?ˍ��2¨��(���h<��ȱO�}�E���#�Г�yDt�M���_�s[�c�s�����ų�a������AFbJL��VȪ(a�ɖ#=�'��s�eMY����ji+����/�2�6S�����`$^���U��ߤ��勚��������ŧ�����wḚ����Y�T�b�}|�o���N��0��﷞:��T;��ğ����{��>\\o�MP������/�KI�H�������+3Ǡ��t��G�u����`����)2���W��f.�-���SbR�����xnkx���U9~԰�:���������Nҿ�H�E�`�,\���%����l�Q���~ᝰL�A�
�a�7���1{��t���qײ���p~"�i�*{��~�')��E�%t5c(�ѳZ�$L�縣̸��pS�^-�C�+���߈оg��+!�,4�}sO�! w��1N�R$� �a��s�2塞�a;lZIhs�!m�7�6Qo6b�ۖW�|4�^���[�YV�ɑ`��Ýc|�b���x*5#C*�P���/������J����du�f<8�"%I?&\����
F�yY)a7�Z�$�i�d/·�V>}!�D"B�%���T�e���۳������'F��H@?�� �c��@}�'�$�T^�\enS
�~�{��~_��4���MG�ȿ��m�q��s�PE%���|������/4�2�>���7�ݬ��V�C �Лz���"Vܴ����sGk�t����D�5�,XfR�ITc��]d.�E���<5�W���"Q �Q�ça�\'	}����~����{��^��|����8JD
X=9�D�gh�^�no
�n�C��"cd���4ǰ)�,�
�3B�-���+�8^�'�#���	�Sfqڇ�2.�۱����{bod�F�D͈����#[5�l�72^�)�N�
�����}�Vm�B�һ�3:LB�?��0�K����y0?o����a#� �ھG�
}�l�^�ޙ����F[��x��7�ÌA�#@�Da�Řk�Nx@�I%��������y]P�AT&��\C��e�K��DE��[��l"�dr�d��L·Z���@OC3is;[egUp��厑������������������-|�z��ro5;�}����70��={�}|/{n/;5}U#`{��bc�V��퇘�z�QF��Դ�T��메���|[26紳����Ԟ�彆:[�l�o�!a�[;�	�R�Fc����F�10�E����w�6|��1� ��d��̴:��sC�a�q��.��ꠞ,�e�T��K\Se$���f��uW�]�%�3|�+��e ��u������t��?�%e)㦜"s�(�D����΂�^��qq��b���%<�e��ef>	��� ���Ub�w.�E7�bcb�V�ܗ��+w�!�hh�������ތ�)��-��J���J�<�3�j'X=]t��>�p��_�b�{!������
ْ+�J��#�����>ˢD�a��+�ޛF#�}R]aӑ.��6h,�Z�������g����B�剂��F�����@�Cw1Re[�ض�ϨI�GW��[ݍl䄺�}S7�2�6P�<f��1yV���</*�,���?��?l������u��ãA�J���0ՆBe��gw�T8_Q�m��k	�����&� �����W���K�L�ޙ^s=��u 4�ϒ��25�m$TR#,��I��̩ګ']��8
*���NT�nޓ�nƘ:qX�,[��s�6S_d��̏����_ʮt��|��8��Zvso5���d���e��]��"O"n;�H��eN�JF=�r�Xp>��Y>���6��y6�tfr?�*`/P��~r���*Ç�����1~�42 Jk���l��(�֌e�}�o�ד���K��� �Fpā� �����=�xL��U��Qω�Re�d�7�9APu���)��\Q����觲<�<�N��ȭz�Q?n�U�uX������J�l�?�9���W��Y��:��@�2e��:���4�b,�9�Yhx��ʋ�N�� ��λ_5�ƹE��R�>J�+�]�������w�?��2��w��r��rYgk(��7���E��M�۱���"�%#�'T^Ԗ(ا:U��������4��]}lp�u��s��w��׀L^ɽ��I�w� I�ϫh���'�=�V7��!e���'czLB��������p!d ��v���+6�ަ{�����W�>��f��}��%V�>�_��&�g��q���ӌ���b��������ѧ��!4��i�ݼw���w�� èo-@w�����:��I��4ߤ@i��?��}��Ub#��1a��ċ���0P$�a3�I!�^cp��rLũ/7�!�4T3��C�E�|}A�f��	A�=+x%�G��T.[!��˨���*C����$����H>���~.Ȥ��N [���R��6j9<�)����6㫵䢤_��+�	bB�H��&Y�$����+CQ����$}b��ţ���1J�~B5*��[�-�4����ڞ�❂�OvH�b�ܷ�`=(��d�!֍�Wd/����?Z]t��}�[�:<��x����@���������\����{v�_�Z�?:�;�h��ȏ�F�Ɋ�6-�\>T04�Nf�
Cغ����J��'��ބ9]�_��QƟO"�8')Թ�?�>��PW4����b@��~#����W���͝��J=Ѕa"��|��'*:#1Z��� Dv,ߡ ʠ�ݪ6%�Uc�L��]B�Y6�)e�~������4~P�X"�g@&�<B�S!�AR����0a�K�y3��u]-���n�[�K�/�ŕ�d@!�W]��컘� �-4�X;��[/Ä.Z�'�ި���f]��������r\�]屼j�{�w&6��@�}DmS[g�O�O١�#��������X�f�#3ADC ��?�ow���gBP>��ʐ��MĖGU,e.��L��O���'
Lfx�r>]�OM��.k���tG�4��$���j������Ctt�==5HOSO�SO�gE^�h�0�>\���Ct�oX�%8��$�U�kڨ}�-�t<t�t�-?`���a�|_��ճ����������\r����@�P���I��4��2�� ɏE�i���C����.����7����D�z��g\�fA���ᘭ�1�~���sR�[ׯ�#)�"��=q�ż
��w[���~�n����D�	\ʲ�1E���y �9X f1�S��S��ݜ�#@5�E�������L��#S�-�Qo`�ʨ&�+�B%���q�� ���j�u38�?����A��� D �B\m4�7!�D���*"�''�k=Zc]'�Y,ybɦ��T]�󛟏�L��}��qԎ�baVN��P.)p�AR�gO�KGli5�|�G�_�Y̛�SS �	_ƣh�*G%GY����m�Y�#������5Pf��N�;�_����
k<�%;6���~wf���O-��!��Һ@����0��	?�������l�S�H�B*3��i�ӻ
I~����M���O�uX�lk��d!.K<���c��=�Yqp�spc�t5�i7��DZ�X1�(�����I+�;��j<7��!�Ȃ�~c�Z�9�{�ȥ�
��g�����(��d����.�Až��/��/(mU�Z�[x2*7�RJ^�+)̼�Z�QvH�5���{��Ѿ�eٙ[���|����(����v��W�#���-�H�@�k�].��F�9��!@�1S�5���L��
��
g�sO�;Ą d���D�.زR���n�j�uyF�@+�cB|J���7�V6���0�)�$\�F�����=�M�oNOk�v�n��B�qC��PW?U�p������7
ζI�ou,>P!��W0�k����x��],%z���("ϗqE�M+��L�g��bAǯ	53n2=Hbz������^�A����*��r�*�J�,c��"�m5��ee�uU-�uy5y�����c���ݏ�ϋ�^�4�׋��Z�~7~���G�* �/�QQ��]W0ŕ����B=_�ƹ4�7-��s籜����M�)�o������--��2K����i@!!����f���ʔ��#U���J���������S���o��+��|@�q�H�$l��r��w8w׹��sq�R���T�?�Z�}y4�y���xx~0<�iJu�?ڊ��>\���߾Z�?i�Xr�����Lp隵�z0Kx�6aVc=,�U�w�i"��iR��Đ2r�
��MFI���j�}&�j����]l��-���t�
��T�����jw�DJ�Q�M𭠷U�J�0����F]� ��f��N�n�[��qX_��dV?����V�cǙ%�=�1�"����hP��z�D�	��D�@���Nre.��Č#cSQh�A� ��$���mj�_c�|�/���k�ndq�pN��O��6_К*;4��m�{(͆��/�pf������S��EW��Ӭ���i�ከ����Lo��>V���|���.I��B�L�X����gj*�] K���R���I}78�c��R���G3:�����ԁ���M+_�|ts�-pF9�ԧ���F��VvhΕn���^K�%T���n&)s�_sCU0�M6����'�m�|R���4Uo�,Y��»'3��tp-*�"�L5�����Pǭ��Lc�s�T�#"E6q�F��#�=���w��k��ໝ���"�%R�Y�T��bH��4�H	rЈ�R�0N?D���gᯛ:<:6��i��ܗݗ��]$0�;��)q�Ec����R�g�M�i�ž2\z�Rn����U�'{/��(	NF\h~�c��yK��'=y��;y���pE�%[�ָ�ﳅ��q�E�Ǌd��bY��	�nB��f���M�!uH$u�JEc�E*�f9�IBb" �^חj�V��[��.��$;����J��8�W7�n��|s)s_-�v�v
��?f�D��E3��%�'�y�:[�`�zLKt�M=s1�r`G'j�QX��_!vZ���=�*P֘n9�u�6��i��Y������Y������b���~c���wU������ɀv��J��:�Z�v�����nh9������&�w�}��� Ltc2Ǒ4�F0��I<�E,�G�z�*��͖��9��:�?vT����п��Ao�άߛ��E͢��+8�n�����H��xv�.nU�6FJcP76���� �p5��&�՜U��v*���Ƀe�hf�x��2GW`�����Z�*�����uU���h��E��OQ�'N��Aj�-򟣆8bC>R��I|�F�#[£�������]tE6�P����8!�]�?Q��SO�m�v��~��Y��6�QC��!*c�!څ�����SX;f�r�B�����My��ۈ\g���o�����E�`�����T�n��OnrM���<x�Z�ִ�_m�H��s�\Sİ���Q�xڞ��t��(�xL�d=�/{�gW2�W2>��@tg=c5U�6�h��m6����Z��@j�xFsQ���w-�ۼU���+׶��l����ucN�� ���"[s~hL�[��⣎�.�Zk&���`2��fH��դ�Hj�'��Hq:�!��_h�!j.)�͢M�Ht�����J�+8� �7w�s�\�"ׯ(I�4_�ʇ������W��F���3���6c��Ƀ���:�3��H6���`����Ki<��^&h���$��I�UL�#����d,3�u�'Z�x�[�3���+�^i=b$8�ob?޺�g11�����)ѬT`@3U��o��:�Bǀ�im *���!������@��y�Ԃs%�:�m)M�q��p���p�z�u����Y��WD}�7Z�U#�NrӬ��>;�����$���~( jr��ԓf����2~�����T�6>��֭�hb`lSAM�u#�����0��E#\dλ���#U��%n�1�+Ī�l���iV�������j�K�CQ��"k��hP��M���(cY7�c����f��+���g��\���Zq
sp{�#(
LCGU|s&��FVK� ���B�-��I)d4UQu�U�&� 	���	x���1��xא	d1���kND���a4��|<	At3M,��A�
��gg��#R/�cH!U���Xv���~�m�7�Ǻ��9(��^8��.pQ�r��ɽؙI�}��9-�o��������yKaj����#����,x	5���<QQ�<k�4�U��y>l����Q)A}��A7@�ިَ!�Oʈ��R��#�X�=F1g�m&�*Z��H����ePM�� ��s<8Aw'p�p�wwww8$��	��z�{p��U�����٪�~��鞠i6�)��+�4�� *��W��*<�}l[��f�M<ͫ�X^*ɋ�t�8�U&��3D�����+�~���@>(��!�("Ԑ;�J7e8~B�9����Kq _�ϣ�'�g!��
�چ�]s�g�	'�c@���Q^�fj�;j�r�e���S�mz��a��IX�\�אΧ�cD��P>n!��L"?8ɬ�6c���-�����S�t0���`K�M��@_=_jb��Q^����Op�>�;�:��	�� ���)�/���zS�8�ӳ�����gmŦ�R�|����+u�9� �[����K��g����Wg"�<W'KT/������;���Y�/f�|8�O'�8��>Iˠ"* -�AWf��L��|�'����6�{C#��/Y�M��H�ʝX푕��v���
T��'�*W�Ur~���!i�%J��@Jȝ�I��մ�ǫ@8���4w�����е�b�^�F����js�����	J�l

DRyFK�>���Z����d����8��a�e[/* �*��BMr��X��n�D�?��kw�}~�U�O�)�Ӎ��|��-�
��Y���Tu2��Z���D坅yP��(����%S�X��>n.�4/�/*=�.>�ZP7^W7�L����&�1����W&�}�?�����ͨ�F�
��m��8gir�������+S��ms#�[��C�N�I.h�5`F�2�i��c�H�Ǩ�x�c��\�����#��@�A��dZ�m��/�]�@���!���W��\���g�G�Q�K��S���|b�I�ܮ��>l;�^�K`f�o�ɽ���9�<ɾ�����_/��1��1�奨W�9<` `�O.f�.fpe�w�x�ݺ<��ii�Y���
ed}�#2L��^���T2��W� ��	#���**�Cn9}P'������[�n��-+oPő�>/��F���3�E��3��*8".xP=��O�^���0��HI��UD�� I���D�/�^�j����l�8*ozܔ0�]F�Q��%�ҧ��j�D���{1��X�3���35����g[&�A��Ml�����pQ�*��Q���{�nV�pM�N�:g���OnS�m}�x���c�x���Q�̷�,(/
Ɲ;#ĜZ� L�c���k���s6�,�B�ܤ�࿺?������\ҟ��zjx<���8C>L�fjy�غ�U�yiҵ�9��N�
��W
�ⴾ�m��'�̇�~q�شBI��ԠuL�XXzQ�A�1��׸��b�8xab� �B�n�#KQ7܆<�.y/>�&V�ONIOU�B�KXz���J��FѭF�;��"��o�xi��u��4�ABk	k�)�E���K#[�~�a��d�?I��ה2ʠ�@��86^�<=�#�A��
���n�q��l �@���_���S����T:�w/�4rf������ʹ�����5�(8�ȷ�Ƚ�˽�ƽL�Kj�� ��*��5Λ	͝#:w�5á�9ϟd����L&>�>!i��S�T�ƿ��(J�Ȅ6=Zz�~<85�9vTU���L^�U�LƩ�^|m�n���/V��**ꂫ���j�7�--m�Oi�;�O�ZQ��C���sIYFQNi�u��WE�X���+��˚Ƶ��{�ji�`t�y�+�l5>�8�V��%����һPZY� �EP)���0���**��]���#����u��� ��|�D�#
�4�V[��p�o�1�n�o�{�f�]߅ɇ����Q�"�4�(�Ʈ���87�7��<�>f�wv�������m���3��A!@��7�]��G��^Ml��v�K�r�L�F�����6=�g �w�w�0ڍʌ��o±��9�*���k���RGt�:�!��~��
g
Z歌���2��?pL��y�mg�!��V�v�+�רA�Q�8��v;)���43τ��Խ��yI����B]�xZ�9�ѵ�&�����υ!}��r��ڻ[����k�WW9��	��.�T�P�!�LG,�b�f���s�|W��C`v�V�����mF*Ȭ�\ۃ�/���EK'�sRFp����d���1��N��ՀgcG�������F�|��kǞ"<)-YCÕ��F�l���b����gcۯ�5�u��qO��_�����tj����diV�՘����W!���Ĳ�9֚.��\�1�eM���|�Odf�-M<	c4u2��yw.Cm��E�h��K�3�Fj@7]�.;�ǲ�-����P�3��M�wWqz����!����w�զ�͎��<��W'�N��c̑�.��y�0�R����y�w��q���� �{���v��l-*�u��j:��y�/�?GDM>|̓�g�6b :g��$w���!�  Iv!��j��+�F��hFl+�$�TF��$W=����㬔NĤ_����X~g`���@����`q*��N)F���G�߮E�Ȍtg��y�Aꛔ,�Qq��(�*���m�
L�+����y��O��[r��	]1J	�;9�
�:ϊ����
�������}d�A�aވ������E�@��A-5�$�ۆ�^!�Q�Z�M�"�oIKkf�'�YXuݕ -ˋ������AD��<��0����OM�����s�gI�!{��V|>�p"z���OJ�+���C0��$�T� ���^�PS:������"JW��8=����;�,�[�A�aW]�S͟������=�SB>�a����7i�����L��16_ðj��p���&�y�� 7���Ts
E�*�)@��H1�OǕ��;�$���f����5(U�Ѫ�!�9��	��B=�:�'�|s��_��eߵA��lRz�E��lJ3�*�i���փ�G���y:O�n�_���<��z�e�r���*wp_�[9�/v�t>�-����X�����MH���""�������^��`!��A&*"���y/;�7��t�!�]˻K|�Lc�6��5����"nB��ٽi&;�T�<�!7�L�Xv/���7^�k*PS��;=hL��(��M�_�Mnد��t8::v�B+١�)�QsQ�}T7�6g<j�@�>��y�E��[���a�]�F��r�	��J&�/����42v���E6��\�����ݟ+dT��<Y�0���X�)Y	
P���������L��}��4�Љ�лV�M@��0�D|�-�oR�]I��u�O���jQ
��Q�6�3�s>ufU�E�E��l�轤r<�f��	�5�>��q��Tq�r�#0����5:�nV�*��H��L�\]KJ���Ru��ۇO��2֞D��s[TU�u���\Hh�UV��������J�id��SG��J;�n�Q�1.�w�퇚 �PR�{7Ll�ʥ�d�q����K�p�оe���0�I9yn�Ny���p��p��p��4��1Vx.�7��܇�t�Zb$5+MvP<{ �� ��|N�`�:ɬp��ڷ@l�?���&�FVP��)d@K|����e0�囊�1��.�b\�����G���yZ�f�Gl5���;c�jS�<'�G$P1��f�����&?��Lys�*%��dbQx���vbUH�JPT�)�ʜ�Q��`j��2�#H\i7��q�����"����U������`�xtD�P���	h�AVp���y�%"8�b�iW�x�ѵ��Q��g����:����&ј��mZ0�XQ�k@vБ����h}g��&A 2�uD�v#�vJ��d��D��C�p̓�	fx1�e��PD_��Q�����|G��h�������a��7�jٔ��Iu��f�ءXe����x���oX'�~4�dγ���)fE��9�V�YQ�3ۖA����-wKLI/��Dc�_�$t��[yD�X�Z@_fP�P�P�u!��s��sE�U�U��0�gR4^B8�q�~��xwI�tw��O`Lk�\��72N��]����;>e�;��Oq}
e�s�zz�6ǒ(tm��n�jp� '�N'y��}"d-����K�������� T�xɞ
2���}$���Աs��W�Bu�X4_q~ �֠bT[��ͤT�m���Cf����Q�cۡ��Xw�ߛ�]s3٣FvO�a&q���Rtٗ(A��F�Ч�k^�ʢ��"J{�ܒ��W
:Ў�K\|X�[ʑ|qPo4"�E�׿��󨒬���5� �[%����3�RL��n��C;.̤����þ'��y�R��t*��b�r���}�f���!V����/}�񱾘j����M^�����vb�Lw�ɻ>�Y�g!��X�c^Lc{n����K~顠Ց����9��o��7p��n�Y�D�&�i	��s��x�W�ԯ�.��Q�$�GZ�������:���:��T_�/�g���N�i09�q׃�
��NG��ML�f/���R�jD�#�,LfP���	�j�[)����y[���Ǩ�XRW����PQ��l!�S�0�e�|n�A� ���'3�X��oM��<k��g�-����ΝY�����ԣ9��T�YU���ȹ�("���	�L'I���aS�_@�ޕץ�5�1��ar����Dy'wr����EpD�9)w�7��]��O&��5�pω�33�
�ʆ�
�Pf�����(�����8mR�~�\t���[����.��<�4���U7y�a�oC�5%�YFw^�p*�\/>TSm"�^KQޔ��q%IӠ����8p�����ӯI�~p��&�ʿ���"P���5�֘�q��C��E�(|�q}����@P
9c���Kf9�<�>��1��ߕ���������S�5�j��7jV�_����Um�t���w�n�cϿ��T0=�s�@�1�އ�!l�x��X��o����`��߸����q0�����n��̯Uhz��ȱZ��e����f����7���"
`C�����ֵV��[�Ө�2�܁'�<�B����n�<H ����B�bk���p_C�X����{���������J9:̬����[���@���� ����?�/7с���Gb�</V�_�/�&��$�����ʑ�	8����T6�U��U�MU<\�7k��s%i�����S�v�#H��ʘ���4F$H��o�r�Cb�*�ú�֧�X(p�`�L��T�c*����U��p�3A�<��T �/d<��o�)�&���ah��664�0���4o�~G�,6���0�$ɢ[�Kt<�j<�¹���Tg��O�ƒ�B�Z�\�پ�,��6-p�������NД@䮒J/S����?0k��kBo*�	b:z����a�3���7��6�-�9�:⫪_�H��M�3<=]������}d\ڒ�U��bh%JNH�0Z��W�1ȁ�J�"a_�y��)�y�e��PF�VU|��[��*���;eG�U=���@�E�.�&s�bM�z����7��r&੖Pԫ�����'��8`ힴ�\�E�8P���2:=�0��P�zW;������{�������>�t>�Kv�h{9���<���4[�r���q�Z�S�-���_k�?/��S���`���
����O��R����'^�d@i	�0��Rk�Pяa�#r#�EƠ#O���hN���i��R�7�3G3�z��E�%�%���J���g�����T TB+z�u��v�}���ͤ��:�k*�/�^֮bē þ���ngEο8x��BB�W�52�"ӹA�ԛ���!@v2݀c�����T�@d��-oD��.��-F��sP,?-G�x��*|*���Gxz,�v��'*�}�ؑ*(H����R�V��i�$J�i�-o9��ͼ�}QH<�+c�-֨E�[�k�p�9�����Ggh8,�`��q��N�m/�8\�"��i�)�v�MA��ӭ3���:�𻭏�n�MN�x�^�	8}&sd�e�;\���;.ǜ|�>��</���rl<5P5��D�o �uP�g��̂q�=��m��z�숙�|����$�p&W ���|���|^/}x�Rl(�#��r�z��j���Rm�sqv槜�O�<� ��I��+�������g�yLlq|\(��3·�׌�?�ɏ'_{ =S:�W�M��ck�b9P�����$����)���%�B��I(���np4�|<�D2�BE+�*�%��ݕ�}gCK�+�SW-�yz1�H�]9��"NI�p�7��u���7�W�4]s�L�ǫ �{
Pd;�n�򘀚1�`�
1��@,���f9zb������Y�k�7YUs=WX��&:Q~��Q�G�;#]�I�*�)��*F�3z�����~	�~�x
�Z��&������m0�k1��מ��?�g��n�ś��FU'Z2P�|3&�J�]�mϹĉ�m�)�A62�����)�4�#��ᄈ��a	�}�E�"/�ػ��eɾ�o��?����x�,��zۺ��GV�$�o������+�,�M��+��|��KJ�������XF��i��0���=㷓@R���u��z5�	5�Ԛ(7���۶[3 w���C�Y4s�{����nG�]��sl+��>�g$@�~Z�� �r�@���u
.Q��#�B�ԕ"�*��Js(���.6���l��Ǒ$yT��`���`h�2�2 ��S�kJ��J�ca�u-� ����\�贈�ym_�r��������u�c������I)���Zw�����]=k��6OW��=�E2����λ��?�b>3wҶ��������ҕ�t�3�r�Ms��A�m��\�Qs�gIe�����
���.�ה�Q�D�YbG�*ݤ�W�e`��V�[n������ʢ����z[J�]������+7urnmJ7ߞy���9�-���_Z�ڎ�>�qg�0�Ҋ�(lh�/���b��}�#�+ ay� ��K,�����/"V��lLe4���{1��B�Y�kh?=+ Ycj���DOh_�ە��K�f�؃8�����RYU:x`���=�?͒�X��X�z����U�XG���:�IR?�������F�CX�(��b��&�5a5��{X�i
��&A��@�GT�l�D:
>�?L��S�w@��� g��gS:�&! _��.!�ȟ���X�Tf^BdJ�Z��R*4 Xqk�^��H.ļ@�œQ�y����ҧ�+d7�)k�n�(�^�8^�٦ P�*����=�ur�X�����z�PD&�^c
ZE"�lҗa�ŧ&�p����	����a �X�]o�_Fĺ�}����y����Vl�+��&Z<����؏5�:=zs<���x1��,9��Cr�(�+�O�:;]��#�Ժ���"8���t��yZ)�GX�o�I��X��ۤ��x�_���0������,V���q�8]�LiwJ[-N�c���G�O�
����}{]��fq�v�汊�����������_��)�j[�qFƵO�V�X�?T֚hz�x>�~}��~�K���f��߁%�?���_�e4ၲ���6~>���W� b����=�޸����;?_���^y���O�>y__Z��k���|;/p~*�")��ڀ�����HR\H�������f�F`5Ĕ��0ҀWMW79��c���u�>���p8p�mj����� ��K����̐�����6%�hr���զw6�\b��Ut\"KY�;��j7UW�.����d����2�텵ȵ�#Ç07�1&�~BW�K�P覤�"��h\D������"��FV���W\@��Q.�-a�ȹ�؛��mѨ�%s��s~��d� (lF�.�3,Q1� �Ƨ	�Y��ȆN�Y���9��H��z�~Ʋ&�(�co��l��~�b�tTR:(�Adċ���~*����xkp���>k2����>y�����s��C���V<��D���<�y����q��j����t|��Nhb�q�Z�>^W� 
�0����k�Ĕ2c�#A��#E�ܽ]Am\��:"�3��w�%���̯@ʂh0��6�1�6�I�+%���\N�'N��.ED�v ���c�}�}ů����,Gz�O+�C�h%�x��J���G֩���/%�չ���v"�e���Q�6$p]-�}\��۔ߊ/�N�K&="�3!=�I�fv\3�U}gd��5hq5�!�������[*�%�s�����~�q�����+q6]1���V����ҙ��(&Es��/�Q�0�jѦejL$�7��AmcR���{�ax�\���d� -GOqOӚ�Ui�0�L��*\�0"��d���zm�tv�U��K���X�o�Y�;Q�Ԡl2� ���ʘ���ǘ'��r���r��2����قbbb	B\	��Ѥi<�̮t�$jqE�� 1q�G���ÿU���aBz�q�����̓�zo���_�Z�h������������N�F3wÅ���t���هV�����z�J���$�D�w��Rlߵ�5�����r�X�/	����I��R`0e�	[���"k���V�1��<�Fc���X�� ��@�|:�� ��T��RAQ�
��.�����<f��*�$~4=��S�GM~��8]�A*����co_����""��vXVRG�o�_'�B���*�i^tz�q��Obј�q�{��}��Nq��x��Z�����mL8oIE�u|�qj��@��@Bk�S�#|���|�41�<�~��6{��Fg�uI��C�C{�9_�6�Ք��|�j/�6J��!K[��:������$c-�G7��[�Ʈ:C�!�S�lA2���E���+���My��e�)~�ͫ�x�`��{e\rl_��$��'�Ҏ�T����.���'���hû����ځ}61{N�B&MUhbpWڞ2��?�Uӫ�5�e�d����1�4�Hu�����i�uM}�s�!����bۛs(cT�KQ�W@�f��P�(�P�Q!0ح6ma9_?��.���V�Ħ�1�'3��=�6f̥���J�X{��zt2�2�#��&��q{'��k�ʡ���a���O��@̢Y�兣����W�9G�7��!_�FQ`��I�T�j�D�ʰZ|w�z���Ջ�l�ݷ����;I�.<1�/��mpˇ����� �cҫzg8�W���(�YEu\1�W)ؚG�D�����yG3�������l���#����A�3"��e�֠ij6S��i�@���W��?������U
ڱ�O	��F��b��m�:cZ,s�uW��X9@I(�
lv��h�PijAY8�����L�S���Oťd!����E���0r�a��G361&�����?wD
	8;���vSb��U�*�6��W���A�-@����] f�J$�%@�F��!��Q�C���P���0��X�QO1@�����U3�;(T������C󭗦a�&��z��� S����^��`@5�W�A����]QF-.��A��@��e�I AI}�'�L�
S�}Q�AV���!A�l<#��S��m�
�I��jC�^���|G���o�N��zm��vð��f�s�q�mk�T�a�ܙz3R�%��H���c�c������|��}a���J����|4�}��X<���ۡ�
q��逻^C���z(kC��z�T>�Y��J�o����m��%�)N��"jr��?V���wT����˸!沏%V��C'����6|.�s�A���z��c��FN�M��r�f[���U��g��#����@߿'�����_����/�ו���<�݊.E�W?��4�0HT�X�u�D��`x��FT�hz�[��q}�[��sz�͖�`��L��XX*�kCmD�&ᣛ���=v���U�0���}�rnb3�$�%\Ͷi�vx66=�P��z�D���"!���(z�q�d6��Q��������*�qWs2���!�#3=q�v��*X�K�ʆ�	(���bn��@t�4�p|@Q�����:L|
�PTц3G����(r�1*)O�U��@/)Ut.ʇ��'�%��0(�&n����t5��+cc�0�K��z� �:^��z�66����^4�d�d��Zq��b�����/����W�s��|���Ð���ı�#���x�,�`/,4�.����A�lc��z��Tja�K�>K����1�0�DIx���f��I-�M��ԸyXG�K��hH#�٬fI�!�ǋ�Cv�~��K[��!�@Z-i�ݔ����m��	'8k�/�<��"�~�6G6Ă��{ ssW٥/�E�v=*�����x��I��4���� 	ٜ�d��N��s�_�N�f�w��G��8yw"ҽ`���T��K���#5^2?�y�6W�V���Ǹ���us�G���X<;"�o	�P�z�މ,0U)�L�}>Id�T�\%s��K���@8�4>�r��P������U�6�A�K�\0�z|#ǡ���_:��㘁)�G�_��U|"�~
�m�g�&���D$m�+\n�|����#�y������Gc���em����H���\��)&���I�2EX<�����^_v�N?�>�]>��v���*��1�$}���K�Zh�='��P�8Y?�R�������w�tl��'O/3A�"c��mQ��(����c���6�+�zj�▎>.>�n)�,��{1�i�fْآ97TTr��jkuTp���چ�=$��n���vgBJ�TR �e��c�Z��.��n��Z霓�^���mm디*:��H��/�)o7s����tb���Q�4cJ���OM����&�	x�,]9�jU6K��!�h�D��1�0Id���a\��A��7�#�G���M�'�&�����5�F�ڟ �@����"��?E�:q.e�
ɖ���b����D�)����´�=5��:�`�dp�b�禽��*%��*�ςr��"g����	QUe{�Fl�����i2�rE2�z�hm1�>1�k���:^��~?�g�����e�M��Pg��&��S�D�Lħ�2�k��0�r�U�� #���+��)Qkp���R���� �`�Z*a�X}�������΀�ފ �6��X��,���]�����L����C4Z�8JH}04�'����D��K`�N�Y(���cUI�� ht�	*�B()=��=.�`�G.\��y�v�]��k^&�̽�I&����U�I::�.�7��P���O������-,k�?J����@�j����&�/��&!}�S�ދ�B��G�o���Q�TI���:�K�G��'��p�� �T4�m��pr9y֖�5����O ����*[�9#�����="ڇ�%�֡+߱b�A�R��%G���:�]QʂP�<�'Tl>g^F53�_��$?{C
�"��D��ē�~nl����P���b��)��q0ntNޝf�l�������Hj��N��"ZX�\9��G@�|B��G2��.�����>O|n��,�'��]�����1a3]�@�mY��4�G��'���M'�[����%����+�{oL��i�|�\m �%#���C��R��2ay"Nrf�wA�i�R�ر����<0���|���� �_�6Q��-ΕC&*-:���!ৣw�>)V����qV�cO��!聓oV����Jad��az��_䒌��6��
"`u��/$�ɥC٣ 4^�[�Kj�sl]��^��'�Z��h�z�9�{�[�W�k�v�A�n��=^v�����;�_�@Q��C���{��"|���f�o���^��ƊE��ک-����c�r�˸p��=Z�1_Gg��<���^�����^j��l�ܱV����w~��棜�ϓ�w
�J;�MR�*0��]�����_ږˠώ�Nڵ>��S[5�~]�6zT��.����W��;��9�,�L���� �����V���Ə�'�����[��2X�J���V�r�Ii~�ǮF�Gg�};�cg�vl,�c{�u���^��Y���Y�8j�n��pN���"�ct� 	�� �'0�K7l	Эc���&��F�KB��۷�3@E���3Ǧ�g���1׎��1��R��rb�f�|#�Ҡ���*{�5��{-�N�0������h�]��y����B"������\r4�gy~����S´B���?f�u5)�:BAYl���k'll�
jD��H�$;mQ*�r���:9y8~��
��<��Cͬ�&�Z���ίi
ޕ�A0�B�1W�aFWW�F�X1��Q���.>a�kn	3���~5&A�pK���`淏��f�GT�y�g���4x�C�a��yg����A'������S�׀����Y{���T`� �䥒SQ_+^=ۘ�_p|��C?|7�� �6��C9{��_���T,Rp1��,cE��&�t�K�0���O%�i@��YH+����L�����$���\��W=�i<����T �Mw���� `�(�E)х�(`y��`䬍�c*߻M:��5�%��z���J�.Xmn�_*Y!�M�:�Cb�&�]�jNiӡۧ���R��!��ЦH�5�0L�V>A��?�z�V^P�T:z���$!�[����O";E�(%AS��͞I�$6J߻9t,㾴|c!�;����fm�s���6�0����|@��9z�)|����tKc���+
�C.�GmbJ���s�����E)$��y��QnS&�?�G��3ځ���M�ɗ��γ���*����3ȣ�qɔZR=��oeFV��O��We�W����f��ײu0`�t5?���ײxˑ����p>�6>\Q_`M �\�F��Cݷ�+�\�t����9�]�]"��p��2wL;m�Qb3�T�i������$�Jl
ڠL�V� =ʰ��vu"Z1
ZDh9���Z@����tY�6� �qE���dRˮ��_們 ����Tom=��K`3�!ء#8�Y�w&�-	sw:�(ꛥ�I����n��wy'΋NU���ʈ_u��Xb�o��k�R�>"�~T�J)��dn�ħ�� D���P��v��Dϖ)-R����c�@�m����M�(8wp8��]��9І?�)+���`T�"}��%�M�Wj[D�'e�����D?�����*�-I\��̍�q�[��H rE�{7�8'w?�/�����#t���<�BgE;W�^WD'L�W���6x�P��W�9,#ɷ,����6S8����!��Y�=�)�#r���N�����,�E2=����%@��8�x6�Z�}I'����\	�Zz(����4�x�7�8視x�6�8Od����ȅ,�.�0��ͤE��B �������R�o�ƒ*�.-�/僪�^�����o<^���O��r4�>�@�(��z+��I��d�O������Q��G��~�6�f�Zvt y����JW=�4��j(+^m��ֳ,U� ��ʭ�����CyjV��/im�';�z!������>�"+�x/�ɯ~���>��s�nY�s��r����2ſ�p�����:���{�5�`r'/B1w�T����ZAOy�� Ѝw��/X>&�e#�H�����3
��o�AW���{�e�ܽ�*��oe�
2�ɘ���g�sq�X^��ǝW*��`\��˺�H���59�(�R�Zٗ��=d��Ԇ&�笄�.�/����=���{��}���$dc�(bβ��v"�G�D��%e������'��O�H�_���s5��)�a{���ר�\��H�?N���`
"C^V�����l��8 oD� ���VX�Zu!?Y�G�7�"z�D��~&�����?f��|�C�ʽN �������4�� �l����i� �P�*\��-��9c��?M�͟���9ni��[���M��tXnqx�����W�Z�<��sX��^�k��yV��kez1ڙ!�t���d��s-�ꡕ�~QB잝u��~{�W�����#�+���i�7?�]9��j��{��y�:�6�w�q/_�n>;���sY���U`cNg7�#2Kf��-dISW :��Ӯ�j1����k��$:�h7�':��~h_�`��n;�%�P=X���d�O���.��������T��n�rqkI��8�zk������"j����|��q{��u}���Jֺ���#��xc��l�R8�$g���f�	k��Y2/��Drm\���{�ƨg��Ue"�ykcӵ��uԕ��U҅��SBLb�t�7@@���.�f��MK�>�Wח��?/���H̺*(2�� �&b�:�ٱ�i(�At	V{Lu�	��\�4#�H�����F�0��2�]T=��'[�������������K�r&ׅj�T�2��5H�X�
%2S���ϣ��*q�J��&!`�ѿ'��m #�O��U
ھ�B]����%�cs�$�k��w>��&cp�B�̱�P��3ar���6A��З�6��͑��������������k�/�;�����s�K�� �<�?���L����52ORSZB��̹a"�ˣ�}��n��*���3.W�8����-ZsR7�U���`��[3K��=Uz ��>��t
�Wa�1�v�Ɩ�O04�Z�L{�?����i���v}�S�������k����R�f��esm���]�*�����q�W{a�h�9{8$�FUa�����W��&?����]�ۧ���L�&�%U�(�,�v�g]�ӭ�>g�B��/�H�\�E����S\Ā�?�� B�ymهk��@�o��bM^���c�\c}r����;^��_��_C60c�n�޴�?��H���:+s�m�b� <�� ���Ȋ�yq5����_��23���a���Ǐkt*`oB��DϤL�h���]Q<Cc����L�^U�h��~�����ߍ�����a�"O1�d}.9(�\ID<�	Q��C�� {��3�9�"�ݘ�a�쬿�Mi����i���˩҃����}����Y�s�ɽ�eO�� �g�,��L"�?=��M���[����K������"PKB�c/C��N�E3��������mq_O����Kv���X5
���vJ���]�sʶBőv�_�|J����x5~�2=�����zhw�XU�ܰ�;�TJ�rX� ���H��|��^���j�$���fr�ja.���4����u�����j�����UM�����iV��]\�]\�x����b��7�2Sp����d輣0�&oɱ�����z�Ы�N��~S��"��8� -�t��Ϯw�g<���m@Y`b��.�/�-@,FȮ�	!4�J;��U�T���Ƌ'/�by���{ڼ�:I��0Z9���R�ԙ=�?� �u�Ac[&u��Es�K�!�71"M"m|�FR#����G�X��F��z ۗ(,���&��-�T���4���\SI�U��WB�Y8ۛ��E5���O�!���v�3�.V64��p�j\Tl[�k��J?���0��o`� �Q�ac� ƞ�-�L�@��.��ն�Ug��!�;�ߥX��T^q��b_�	zn�}����#%U�{ݻp��?�Q�ًͬ����G�u�*���~���� �Χ�*Q��_K�[Uҧ�k�������H��E�h��q�A�W��)��A�gt-1�Qiu� *v���t`��8޾�8+w:_:�1,�7��,_���W1*�V@D��x��֏���״��Fn�<[>���l�����v�a���:Tڛ]oݨ.��M�3o!�T�:��20����%��V	�1 R��
$�@��k��2�ʣ%[��N�8�3�Q�!�"p��S�p��2����͚~���L���Y�%��[�ޯTSֿ���7y�-m��e��F&4:S%�5�gKu�	��0cl6������ f��9�xw����p�ҵ;�8��W��v�����V��1.^�~lX\T���/Od"Q��"5Y��Ud���/�r`�rK�y`��@G�v䵱n?�nXs��� ʲ=�)C�G�\gW����0��Fwv<��[�)V�N����ڔ���S1+������,�H�Ç&�Z�(R0S&?��â�tX����IE��&*�</m�W"8d�ET��ZRA��#�&hWY��l������8]|�?�}Œ�#�ƪ�?���C�%�Y��m�k�秋��o=�O�{���~�{�1��!�ٺf��ۺ����I��A�rR�m��w�P��4An���:w��{�Z����s#�Q�_�绖�X��گg�n��wt�o߳t�?̈́I)?a>J�&�YVTo&X��Y�]k�8^a��ү}�$�ժ�~yn����4m8q^�q_����@8��X＝��}�{�0o��D�r�4���ٟ|����������p��������^�7�`����M�֬��֊ի�^�n��k�]�jӪU��~{úu�o�jo�H�8D2�H����L܅�<6�G_���x<��XxBe45"�Hl-��Y0���� 
���hjq�38C�]�jj@�14�!:�[\����1� ��ё"t�p-)�b�h(���iP���h^r?7�S��g̈�ʎ�ˍ*J�,�I�*N�.˪.�<T��X�W������}��0�0X�ֲ�Zf���Z��� ���Jހ59JK��R �庑���r��n�$W䷄��Dkja4aM�7���J�+������a���p)�~Scj�+|=��h"�p�wYP���Ԡ���.��.�ucjj
��4W͎������15����o�����ɳ�W��?�2~�����Ʃ�#ő��WJ�;%ן��C)�C�����"�#�lM����"�%�����d\���1X:�Ac"�5�d�!"��FAejjX,�2��ChA,�u&ԂiP���i��ٳ���>1@�O�y��[MM�����3|N px��@���(Z��a��b��	f~�7��g��� a5K��0���i��8�:� qW���N*�Ie�B���Z�ʠU5j��C�5+��1@��vW�G�<"��`���{'�|�]�R\�S!niFKhu��܀�"��BKx�oh��_��e���󲄚=}=L�:��A��rӄ�+���t�55��fadL0���L�`�z�lMM�'���p�Ea1.I�ه���K�����<ݛ>y:��X�����cigF�Ύ���8?�v���)@��i+��W�s/O�\�̾8Ƚ8�wi���tѕ��k���<�}Pq�|孋Uw.�{�������
f&rF��N�*9�od���-����������k�g��F[b��h��,�0�����X�EF�e>�ƺ�؟W�ǫV��[_���AM��h��XձD݉$Cc��!^��m�T��K}D���F�AC���O�uBl-��ס�mw���8kw3�4�<̄�4+C{��>���i����yOy�G,�4(���	�����L���S
�
55�tV#kn9�o;��[��h�=��md45� @S5���hj���P�@#3�40P}�;�y�,��}���U6H|�؏��:a C�$�qNĻ ]P/h$�:$�f�$w�#���,����
[|�M��� � ��au��*�2��EH4�5��p(�cg�/��?������P>T3�beU1RP�.8)�U3XY��T٠�f���jd`Z�djt�y�b5)PʠzT���05h�;��7�,8��� 	a9jj��BSӔ�k+AL�5�9k^46t�/Ps�*`ISӹߧ�_g�?��`@����áH��#'kb���:�u� ��ԼSc55U�-���iy!klu�+X�ŧ}�ɇ��>��?��w������/_����s��wn>��Y�~�-����9���*�={]��{"��wo�W�>��R��"Sk!XU���M�դ��u�-g�����Wx���th��U��<}O�k�W_����2T�?�?�Ծ�����B��KWY@����}���'+�E�>UZ:��}�s=�g�@����\�֔oj�36��t'�4���]Q�,�IKF�K��H��*аKC���-���C��b���G���x��HPM�b�4m鈦�H�/ij:�5��z$IM��l�K�憯�u?������w|��̷4�<�9���L[5��6Ke!<O7��(b�����:�8�hsď:���oc
��:#�c��g����S���O���=?vw{�V_��Α)g��Y<i9Ss�Y���"k�:�G��!<�yDA4�C*�	��1��	�5�5��8�PY֠a5�(���9&m�Ma��&���Ț4��L=�$"�+��ZΠY��.i5��4��r��\�):���%���H��e��	����d�yS#_Z� ��Y`j�NIR\��`�5�fN�3�tl/A��FԄ][vnZ�uݚ�6���ޮ��vnڶ�m��y�ֿͫ�,��&����m{v�(vx�vG�Gs����X�&�s�Z��@)�,�N,y�v�76lY�z㊕�W�.b�uo�ܰf��7�����m~��+7�Z�m�����r���I3�F.OL ��H{���ڲf�{k��zw���v��ٵ����Z�ފ7w�^�yg�5;7�ܽc�㦷�gxv[O�������۟������]o��r5����7Vl��k6�~sͺ��׭޴���o���nݖw�ݱc7���(
MD�����AwS��[����5b�X"��yj����H$d�'0zC/8�Z\�����������f�:.���j����Q����yL)FO��S�u@�����i� 59H�ȣ 5��?�O��V0=$TO)�OË2�S�=sb��JҢ�f&T�.�>R�{�8�`Aj롲�iIA�a*?-�[Ɏ�PE!>�5AV��		�Ӭ��A
j����"3�T�-=ZG�ꨀ=o�&�!���*k�<�p��,.ԑ�5ެ<_va N��&[�S_Oй�7WP��PӠ���.}�]����4���(��8Zza��7_>D����W}�`��T��hǕ��k��������j+bMI�T3�0X�������nLMn �$�g�PS�.%��T���P�<��M�15<Vâ2aL�sS3�42�԰�6�jP@hjl�j@A$�U֠�ƺl���P@����f��A��楀���`��y�i�	�H��qɎ>ޢa!��,��䡦� �Y���lL�BSCO�`�z�]Y�>�L}���O+6�9�$��
�\eTh�J�Ai0�Mz��^�i0�L~F� �G�Y�QF�(�'��+������j	I����o��O�9 902'<�(4� T³���\�"���ޖH?��W����C���k�L� W-� �L��s�ǻr��50�&ѓMM�'���N�@L�E�� �&Ƃ�_O���02�3�"���������P~��ܱ�������s�y�S�sSy秭��r!W�r��˻z���T���KcF��J.��^�(�2���́kg Wg^;s����ۗ�ݻZw�F��뇯]�{n�pl�px�t�ԁ��ŝ�u�ZN�v5j�N�O	
v�4���S��~2��z��}��>�ď@����V	.!k`�H�55ա�C���禦>�؜dj�7�Dk���'��7n��ݤe4)��bb� ����q��Xvu�=�����'�N�|촐tY���>6H�hOԼ5�i��J�	ysY0i�h��#2�1��h�GVS���u=
��<�Q��Y�� +@YM�5�� a5�����0g�t����#lg�t�q(�V�9!���PScd���q^.���d�J��ڏ��8:u;8�cqc4�9>�X4'\Rˬa5$��$u���=����v˼�i���5U���P45pէC!�X̫Y��@��`�P���A$N��������݃ϓ�,`IS����e�� �~́C���G����55d�o�5�����й�wL͂�˘��bj��'�Դ>_

��QS���W����r��nj����dԡ���ޣ�}5QK�������5�4U�4�n�AY`d�c���'?��/���~������_|���ٱscmNT%�5f�֧�vf�v��w�Nt�Nu&Ow ��r15c�a�M��!c�c� �k���<�w�v����Jw��Xm��p�p�ݏ����5u���ؠ�[��_�>Xi>Y�ݻ�{�*��wk�������؞}���g[���a��/U8��o�����7F��7g��s�'Rd}%�]��3�1�e��e��eA��!���=%!]�!�����{c�őʲMy��4Z].�
�D�@{Q��Ju���ϳ�������\jҔG��ǐ��H��h��h��TQ}��! �KB��1kMm��&^��f1�v��hs"QV����iLV�X�j:����dB�j��e[��=V�o�1�G�΄/����y��=����n7�=n�����.e�L����1(�Qx�D�&Pg��`d�9���@���r�u���x8p�D��⧝q�[d��i�B�"�֨��4`{G���U�Q*n�D�Y�9�������� ��(w���!�*%���O�� ������|� ���~�g<��Y�����#S���5o(W��d��z�M����ؔA���m�;72�����]B�Vs�����$�0	�L�z먂R)ƕ1����59V�e�����,��j��5"4��S+tB��Ī(�.� 9C����5���	{�ٿ�y���ｽ���׽�v���n|w���VoݶO�Mc�1�{�$�N2ˑ%$bWo�B/q�1F(��j� ��D��dsd����IwS9[�ɛ1��q��0�mN�]��-;ּ�u���o�Z��o�[�v�+֭|s��MTg{�$eQ��V���j]�f��T�f����m��ަ����mǖm��nwض�q�{�7�޸n纍[Wo[�����8lq޹q���h�i�������~��Oo^�{v�rKC����ݍ��lܽ�k�^�n����6�]���7�X�q��-[v�܃���D2�2�O��1�kt��ಘ<�i��v�
�B�X�x��Y��삞`Hc`Le;�z�Gn���a�����A�2�g@O`� ��d�w�,gj�= ��.&f'�CDح�;���L"5LO�22b]q���W�B�߆��F���zZ��~�0#XG�2�� �O`"h�~�EŶh8za�Ah��y����ʳ�B|�ͥ�G��_�xd����[���-G�ӣ�}]B<4��787�Md��9�jV���ch��J���4@�
!XI	�У��h+ZGC�CiHqFz�'х�h��J�'%�̂dx3s-��)���f����oj��O��b�/��-�{�����Dp�*|"E �୴6E^�,;��p VP����UT��S=��YqU����ʼκ�+�}���g���g�����_��_|����閩S�w.��=wjv�e��xe�w~�4�����fx#:� ���G��#
|)Vh��"���̳��} $�&�����A0 f��`���|�L7� &��d	�ȥ��t��Åyj4�F�L%�(x ��'�H�f�Pkuc�u�`aZW�hr	�I�S>(�=n+k@��a����<-����e����p�'����ECi�!b0XgK�H"��'�p�3��ħbT���h@iJ�Hӽx���ɳ�.���,S���D�j��ɞ�dwR�;%ŝ��x�R�eIfE���O#�TJ�j��N��ub�^�2�5�*��������3���k�����p�sqӻ��\B��ZRq�1�& ��-�)��I>ɾA��!�� P�N��	�
MN�����{���Z��J����FI��&�GcB�t�7ѝHp��(Lpg"����y���Z�'y�nA��N�b�y��\)�.��(MVqD��􂺂�֊}}5eC͹���G�'��΍����{�L�峀�S�W��ua��ق�ys�%W��si����{�n��u�����q���.�<������.�_��~v���ީS{'O���8{�ƕ��Wkf�;q�l����}ݕ-�53���b�|���!��A��@uV�"�O���Ϸp�}ž��)�#X�ԟ�7@���@�¬4/s$B~8Zq0J^��n��7Gi���j\Yn�f�Y�lQ�[d�!���o�a�N5ԝG�[��w�2�z9�!���v�(~`�<ҋ?Љ�jO���2�G�G<��,Ƈ�4�m�C�	��@ |H ")��<"С���5���p>ԝ��jn�� 7��#"8�/9b/c�W�D�������%g"�"�0��������M�<ys>�����88��c�
�h@#ണ�)Gjg�� w�Lt&`�3n�@�f2�H�w��K*�E���A6k�M%&�t�K��-��uYDmְ���c��#��CA|D�� [�35�D�ET�#jf� P!�*��v�(k�l5����_[�ˢ�G$O͒@�����f|��Y��5�@YcEל�4��4�hp����^�0lo)2���t��u�{�"��V��a]:���
XL_��yO0��*��ph��ȓ����� d�n���`FaP��Pcjz�Yc55{�Y��l+k�z����k=q�� ZlYlj~��/����ݺ0yq�w����2�dC.���Z15�M������� T����%M�,���_�	Y��,�i �eFH�^So����n<+�]e�}�,���'@�fi��Q��i(2�W>�(��Ӯ���o���I�o�8U��nW� � ��L�P�o���cI��a����E!͹�'2|���N�>�`8�պ/�Hv��$si�k~�.�O���8�+p� %>ƍ]��H�:���\��V�՜�q<�x<CW���<,U�kS�u)bt�S}�k�35�廳@�<Gt<^v"Ae��� ���9g�6M��/�!�溷隗��eo��f�k���\L7Ԛ+<�y:�m	S�`55瞯���W���l_ �4���H�%��8'�����({�ͼ���Ҫ�k�w]�\��;j�u��"�9K$��Kx�|��\����A3
Ø��T�GVYckj;S��h]��>�z�@�N�\"S.�isl�}�Ef���vY����r�Bj��գ�vk�]:^���f�5jY�J�a	�B�\$t�!�_�#q\��8g��545��f	S#pL@V}Z��D+H�j���*��$n�������ּ��5+V�]�ֺ7V�Y�v��w�ٽ۞ɤ��ۘ,G���a���b�����TV��%����J
O4�m�<�s�r���Ee��(��A������v���@�E���Dذ}��-�X�nśo�\�r�ʷ6�y{�����{T����3�j.Eç+�4��)粙D����[6��yû��޶�[wnݶg۶=����޻;6�߾qӶ5[�]�e�;�͎��n�2���O|��������_�����}�\ߧV��ߌu�glڰ�ݍ�C6mܺ~ݖ�k�]�jӆ������9�܃sp�a�l�K�p)��7������p�yMc��Cf3qlL��:��*j�M(��-��������򺦆�l�ഋ鰃�C�ߥf8��q�Jz���eDY�&�$���O��8��h��: \�� �Zz���ckفZ :_5�W��Q��R�Y��Q��H�17>,���랛QU��X}`��qvt�Υ�S�'J3�#|\�]T�&$e�Y�	qSD5�G�\6@��U�|�4���U2�4 ��*�J*��D�Y�ϩ�Ei�qv�;������#���dx�3�9�\ � �ʚ�SeM�5�0jjleMu�ʚE���15��(<_F��b� x�bSS��o���I�U%H��T��e��Uq�\Y���pZ`wuacEngM��ɞ�}��ٿ��������?��G�gFO��h�~��T�Pcթ������CU��@A����K�������|��|9�Bͷ��> �@YS����g������� ~A�� LV.Gg?���~:���aQ�|��I��Q@g1�t�F'�($$+0�L ���h-�������yQIc-��r���0���Y����xScj�450��d��U֐�X2� e�'�(<
O�aD����<��`=/�C��#AM ��\�r�&�B��e�Yi޴3%Ń��A�~�9�>�4e��:�U駑��%nr��B�и(t&��0��Ln:w������%�ܣF?��נ���}5:����x��>S��5Ho�-��P�A#�uu���D��� �<B=�!����n�ޮ>W�����h�5h��@�2�(4Ȃu�?΅��Ɵ75n��	�l��y��XM��I��%{s�ͬHz���@��֕V$n.;�[]3\_3�rx�s������s��.�9re������ �O�5?����f�G������7_����/?lyr����}?��������>�3��î'�z?����fߓ뽏��<��q�b���c�'��O;U5>|dz���L������C��{{kz��;�Zޟ����b��d��aLM�7���Yba-65e�|hj��,p4�#��9���V���4Gi����^��&V��Ѩ�7˩�bR�����6�0L�f������������4��O�����&�c���^�N�Z𱂇h�S�S�#*�)��h`�cS��=M���#p�	���`]��
ՙ���O���3�"wK@Ys�*kf1g�������s�	�1�� ^2愱�Y��8|������d55CX� �����<Ig^In�T���+�%��AvV/�2��L�	ِ���[��#��A�j��u�� ~u�fl}�yi��G�R�z��v������>��Ǘ��F�"f1?���Ga�N���ք5H֑�,ij:�\:J^��X�~�� �Լ��YS���,S�M��~�����ч����r��TgU]eb_c�@s��������c��퉓m��\L�Hc�i��98�h�|�15�������S���xZ��.5��8}$|�h�TCBW��:K�P��[�ō���п|u��_�<��on�{2�3[��j_�mK׵����-Y����Ӽ'y�G����͒XA���������e'!m�9�C߳��
�+X�A��s%�xN����p��Hӑ4�Y���n�3]�gS���G]�7�'Ҥ��OO�-jj�|%�i�Zg0-	춘����%uqR�k��Mɪ�d5�-	��Դ�+;cՃ���(�d�q615�,�>.p��K�.�]״��R�U���w��F�jf����~��@Y]�]��
�ѳD���Pg0�I��d�D�(�]W�o5����?��zjvh������D��{�4Ojj p��GD�8:45O�����$ 45�jPVS���$R���W��Kl��9æ���}b7���D|M;��H]"Z��ѡ`v(YN��ӤaW�j��*1���'|A�![��Ԡ�&C>�T�6�
���Fh't���T������)>HB�U{��ͻ6�ܼjŦ��tܾ��#��B)wq1��租��hn(��=4=U�J���]7�d��G}��^��{���OO��s�n߽�]�nן����{�8�3a�I&4��f*�f���L3� 3�̒�A2��0���C��P&��I6��&Y����E��ds���:ϩs�v5XVu����۝>gnDM���$��*a괴�3�j��*³s5Qˎ
<j�^{e���Ƽ)GʅLn��v0�g �w��.�fг�A���1�^9v��qc���������=~�3�G�1R��,dT�Mc]Ӻ��'�~��W_~��O>��ڵ�M�:�g�hy��5F0
����9*��7�_}u�+���^����ICE�TA(a�Xt����h~1�O��F���j.�lC�/e|=|'�6�ɯ} �00�:��^��=w�/�O��l�;w{��=M��r!)�E��h�A�f�F�%��35da$]A廩�p*�Mg���0&;�d�3n�WӨS\l��Ivh�L��N�i��x�6�mΎqO���M�*�Jl�,n]<g{��#{w�:����i����̄�#-�U�]�_���̈4%���6��N�[�x3g� ��d���x�K��<�N|��p|��p���*-�����T��|ja0q�-�������xS33S˗�,ȷ��5��^�𦆗5���PA3����5�����+`˫~$:t0�>ˋLMW������T[ ��֦J��B��\�\���s��+�mo��z���9gm�j?��ϟ��������W����ز����v�]�>�~������9��iY\>�)i̔trz99bjd�iR�i���#�L�� xS33�6��>-�R��-�#s���p&�A�yj,,�"
R��T�RE���.j%�P��
�T��@��75|X�����=t�%x�gj�,'������Pp�zp��s��O�������{��bj��YY����K �w�w��L%��TO(�:,��dG��L	ƺDݔ�o��7��^Z���O'ySS��e��K���'i�S�����W~�#�n�2�4z��n���6���P[l���-���ZIC���b: 
�H܄"z5����M�J�T�`/�R
9CZ3Ҕ�e� 5�`h�����c�â���6���
�u8���gnlxn�;3ܖb�{��Fx���:����T%���D�<�)Ib
���Lc}u���eZ��]رkE��m�Xw��'�/���zv���6^;������O�߿�������n��{c��ަ㻖ں� ���h<�}qߦE{֯<ݷ�ľ�'{מ9��T_ב݀�'���\?oê��։m�]m3׬�߽nawwǎ�+w�\�{��=�7o[���4g������E��ѓs�ySӐ����NK&}153�pe�L͒,��L^ּ��p�;J\+Kݫ��VM��H֯�U��b���*3�� ��*W������ua�դ�
\�'D��ʃF씍���݉�ݏ�=��r+���GV�#�HK��P��#�� �`����Q(�*U�{��dj^(k�[�P�N�A�j�+v����2�]R�>Ss^�x_���9�I%|B������BuBN�����7)��~��'�z��}.���15>MÛ�>ܫ����� �S�U �$�=k2��Y�;�����p�q��p��p$��fO�i{�q[�qS2�jM�~E��=SǇ��S6�ո�K���7�fX�^ּ�����,���Y|��n��c�O���1��25�8������4>�_����9�yj^S�s1>S�\�S��;��w����WN�ݷ�yŒ����n��S��S��Ss���`w�����[5л"�cP���H}���9�a��|^��?幦�%15��Fn����K�w/Kܳ<�K��%�64�^Wlm�3w��u/N��;뽋����[O��o���}w��ڷ$eǌ��,�5G����^b[��oH��c�7��@��pRd���r�,@-��ѐ�H�[X�(R4��=�P1�U��WD�~ ���F��E���������v>��:��\fa��v�%�\Qg�
��IjtU��J.|�}�����K��ŧl���<�f /kVV� �+����T��4j��Hnԩ��siQ�S���p�nLH���p.�s:"��~^o�H�a�${��5���Jt{�tC��ۧ0������e�������i�sx#��4C;�~^Ӝ@�SuTq�>N��L��x=.�Qv�'%����$��p8.�5g1�<B|_SskHF�C��<�5�Q.C_��E��GyS��+|�e���	�8H��it�l��M�j���@��=�c»-�z;��dֹ���Â6Y��Z�t�h�^�\d�/�-L����i�:^��� �L�N\�eV�D/��zi�I��W$jTa�:�'��H��m�eddLl�����e��u���v����w�{v~�dǓ�7ݻ�}���o�\s�����7�s������l��Ά[7���/:t`��í���?:�oߔ��K�:�&M������p��R��r�F������� a��J��b3��bR.c�aZ4�HE;�qn�ˠ�d��\��q#Ǐ��7&p�_�x�`��c�ƍ�?�Gc�,�S(�T� E�9�{��_|�˟���~r���S�7�6vۜ�c�Q~�_026P9�_��X�#����2n�+c~����3N��0DC�EY"�@C)��4��4^�Z���fd��a˲4ͥ�7�<�7���W�<g�_�ki����L, �` *	���B�����zep8�H4��;15QxI[�.�d#�y�Ln�5�Fgrk���N�P&�N%X�d�.��Ƙ�X�:��D�x�!#��0x,:��^b�k��iwm�t��ڊ�����x�9���J�ȎO�8�c�ң��N=��D��h
��H-��A�z8ƀ��~8I&8��X�L~J�.�+���J#1>M�/��{>��&U;#C�s4>M�35�ʚee�������*����2��*h�C0��������x������I�9MSii���67�8=Kߐa���ꘔ��yj��e=��6�νpdۯ>���Ͽx��_��?����.�����tp�ʓ�zz�gϯ�_>�pay��3W+:K?��LM嘖�LK�����$ 4��C�����������i��N�6�̷�.tLϷN��U$���Df�:��x�d�����V`R	,��$
�R��K���%R����� p���@�5����[_��4�!�Ԁg��{�g����K�~�'�55��yIL�OրC^� r9"xY�K  �L)�J��P���d�a(�1����u�St\Eyo@��3
���R).[M���>���d��7�ǚ#��v�G�����X%��QF�PbA�@	��U�re�<�����A�o������������B`A�
�BL�����!
���	 ���Aĝ
Ʌ�J!b����� ���ԩ.[nlx^L��H���h��gj<��BUƫ��)�����$�$E�UG,YR�rݢ�[Z�6�.\�tZ���ݛ��liٻ�wmZ�}����\d�6�ۗ��iH�R�1�6w��	��bk�]Ei��$kn�3?�U�j͊c�x����hb�t��kQ�^�0�:�03j�*�jVG�M����Ĵ���ʊ�S-��ѺtE��E3�Ϯo(N�Z3%7bJ�÷�iV
;;��4Iܕ5+�������]��]��,����S��-��,����b�ڒ�5���)��N�qS+��*�j�F��4���Pw��V(�7�^-t�L�w���<��Q��"��Y��t���:��i��1�1�>T���}�'L�PYs�[
�K�����-���9�aWW��8��:+W]Pa �ל�e�>%�NC\D9*�r圎*Tg	��x�`���_�j�0�q;A������<�i���{ab�
�+G���^v�`���r�j9紟uYO��G��CnÁco�eW�q{�qs2�]xm�~e��#CǇ��"k|��E���9�7�f���e�y	�ZSß���ǁT2� ����"S�}���9O������15�:&oꜶ�k:S�}��Dw�������Y������wo}��ݛ�_<����پ�aO�Խ=�{�������:���4}/���_15�0�4xS��1y_Sʾ��-��wο�e���.�}���̮��ف��=��OW9S���_���݃�O�-�4��;'y]�}i
ݘ���@CS��N�F�k�QՕ  ��IDATL�k��O$c~<��#_	�j��_1��F�yuD�������mY�Eڴ�I��$.b|i	7lm�tw�z������5w֘:��U��J��R�V�k{��i*�<��gbg���2ӷ��̲�ܺ��㹦fKiXo���hN����iQWR=���g&��˸��x.���v�[��u�K��<�;I���j^�p+��tC��(P�35�ꤷo[x�2���dojx���m�)�t�4oj���:���䪓*�4A����vԠ~7=�S뾞\��I�_ה��}/*
ܓ.R�e������`:a���W�	��LRÛ��
b���+05\X����
_��Ks��O��!
�Gc;��5>Y��B�jh��6b=Vr��^�W���Ŋ�g���b�"k&a�Y\o�[e�4og||�i��R���h�>MS��D�:I�Q�aP$� .&㠐qv����ӽv��m[��uػ�ྖ���5�w�������Yt�܂K��?���Eg�/>w~��ó��qt���G;n]�����V߻z&��=�wg����v4�;e����=�]%-�鳦��R!�U̒~�`9,U*�$$�r;�p�pB�QÑZ,JO%���a�h�Y�D�c���d�����
7:dܘбcCG�56h�hp���%�W���`���jj�|��ӟ��?���{����`q�GTn���'�H�~f��x+~}��ǣ�?z#�����2v��Р�T�)�\��e�7!�0&0������f��Ѩ�|��Ưl�s7`���|����`&T�S�ͻ��y��4?y{��"SIB �8��|0
%�� T�G
����2������D�%��"��0JS�Ή`�O�al��Lq0�N6��&ٙxc�<z��F�՘��6�Q�[O�;��a��ȰH�Q�´Ja�I#CR�BC@j\edq�Ø�WY�Q��^:!)+6,=ږf��0n��@�Z8B�p��Q���WEk�ZY�^�dVe�P.y���qa��HI��4�TFs�6|�&nH�4��`v����x�
P�d`i鷲��E�<CXs%7l�UA�����o0
�U��"S�g�V�Tr�� -5�Z���g駤��E�n�?�����΍m�6t̿t|�o�|�����櫟�{���]���Z}b_Ϻ�������	de,YGLNSON���LjJ*<���N�$�S����5��i �2�\��\��|۴<ˤ,}u��4Q=!Z���156�"
X"R
�r�X&�JD\̋X*�" ���%�_��r�k|�O��|�i�����_��H$>S6p��[��'���7�	���}�����4�P
X.��BH!(�\̹(�X.	�L�r�$�:+B_c*�5�&h'%k��4ހ�)�ڗ�~"�҈�T�.�M�w��vR��$��u1�F2������p�
�KƄ����$�JƋd2y�B��(,�KH�!rWѨ�TIPX��0k�،j��1�	=8�2�
�P
/2/a�H�/��K�������I��Ia�vCV�3?�5hj��q���o}��Ѱ|OYU�@�&2�ɚ�\ǔ��Sr��O+��QQ=��lZuVUAzUaFEAjinbaVLNjdf�;-Nn3G�9���&�KfQ��j�sj%Ta!;�4��]M��!#A�t���-iS�&J�� �H��R�K%�X�%�BA�0C�jVg1Yl�0�-.ʝ�����Ɋ��r�yj�f�gfge�gg�g�p�8M��55�ԋ�4�ӵ|X����废�5Ϻ"߱&߹*��˶��.��A����EO+)�
R܉�0A�l\�p�
��VBrP��4S�nÃ(�����}��U���y�&Q�{8��A'h�{r%�m���bj|�a�5�3�� C�wq����E��q�m��a��9x��9.W�&�/�K��m�㣤���ދ����Ű�Je�\γO&�J�p�4<ϗ5���i�+�>%�"��4�W`{�h/����>�џ1�ڭg��N�Q���x0ܰ?޲;��3ɸ5ɰ)�Н�_=hjZ��˚����+�|,��}ߘ��ʚ��"S�"|7�a��>st���0�ڙ������gjg����3#ڧf���JL���I;�r��S�}���Kw�4�(�f����M�g��y������:wx��������Z;c��i��O�[_�}���j~��Kj?�����%15[�=����q{�'�6��o�:�Vze��K�g��|n��{�|�����q��_���{����p�ս�-�{Ӷϊ�=-~}i�T��!L^m����pKޠǎ�G����������[������#�ƍ
$�ot���Ѐq �`�8$@Ǝ?��QfL$����ۖ;˜�5޲�Q�"��*S{���R�^�i�d�*��%�5�X�,/d|�Y��>����yM���˚R�u ��ƫi�W�6V����{�<���N�<�q!-�jZ􍌄��I��2��L�M�9���|�6]"���e�1��5Ǽ��75�0�4�8_�RSs`�xV�� _�	4���g�N���4'Q�4J�P�� ���N��!?a�=)��[��_O�����m�įK��}��r��\!��Q�w4>S�M�=��Ӿ�O/25�d\�'kTx�0~'/Q��>MGHt����6��M���R���뼲�Ǆ��Q���j����9Z�� Ϯ�*k��FZg��EO��PMÙ���[�$�i�"���kjr�,�2Q�r�B�2�΢�'�Vv� �@]����YӲ~݂����������ŗOλzz��33/��~����f_8?���E�/Ϳؿ�r��Ӈg�i�sm���V<��y���k�'���Q�g��ͅ�zr7�I_�V�aMngK�ʶ��Ƙ���ȂlK\8�"!c1���;)y!��x5�A��D�^�b���M&%�'}=0�MA�[B����F�G��5*�͑!o�<����Ѳ����q��V2�i��9g�_�����g����?����~V;n�R؂!盡����+�ȈъoG�$p�+�G�p�����~o� U
B��!�� �D��J�r�R�L�M��4��Q���`2z7��k�gM;�1�'� �00��'Q`�~�l��6L��S��n���P2)%D�������2ɂ�o��pK�"�h���34�)�F�K�,$ �Lx�X�
c 3*ӫDy�F.`��Bl" �N�6j�M:3C�2	"�0�%0V9�0�.6ܞ�W��^2!53.2�i���Jv�=fک�m���(�(L��Y��'��sP�0R�&���(A�H5C64���b�r���%� �OU3#C狦�M��#��湲fi)C:L� �q4-��
.��7����F����᳼��tT���O���*kK�����Tan�q,.6�/4Ϝ`��nh�O�߰���-����ڱpcۼ��w�ۗ����O������^�va�����Xur_���KZfV7O-�N2�s��&�0�S��75)*��dxj2:5LO" �� y_��iHgSҹP|���ӤLcm�9?ޔ���yj���QbR�J(���e�T 9!2hj�$2Ro�(�2�]�`W�oU�����𦆗5`�� ^�'kx_ÿ8��}/ȟ6��<��P��y����4\.a�[ҥĕ\5nD!����C!�r_xH�)],��d���і�8#oj�EOހ�P�)��O�kR��$�&�cj��''�x����f�����*@�/� (,*'��	�~"��� �%�8%%9�VjԐ�����$��A�`��M�j�����A4��' R�R���ĸJ�@B$P@�d|�d�8ɘ12�1Dh�QzL�C�<S�� ����^�A�/�c����8�4�*��sc��䪴���e���blj+��jX�FmR3��0+0��)Q��H5a�¢\ �ݤ60JR�G\X\v�=�e���.�"�h���tDڭ.3�f1�:#�R	 E�\
~�����������@������C�H��JBq&uV��0Ƒ���hJ�)��toj�kg%S�&����$Pi�9i�����TN�,���L�0;�%��>�ҙe�J3v�k�6;�e�ט��Z�Z�b+���Rԅ	���څ����wR�F�����Ҿ�6�3=3?v���5O��c�x�$����0�X	?P�����r%��35|{��y��a�]�}g��;����M���4SƱ`X{^	����O�����e�^�ho��#�¾����������SSo�\�� ��Լ0��YMá��AD/L��>ѫ�  �B���)���d�YN:L��cN��p�X��x�D�D�TO�~M��+]מ���jj^��iX��o��15��Oּ�׼�Ԁ�s�og�����@�������ڙ��M/k���̈�=��75�:��15;�.��Ӹk}Ӌbj|.�4��P�~�gM��>z��wn�;��x���=KV6����W���X�ć5�6������d~IL`�|_�i��]K�Z�u��:���⦙g7O��k�+~�a�����??��/}u�;���R�ے�ma|��mu��W	5����g�B薎��~����
x]0R86(p\`���`��� a�@4�?`� 4�!���?vܸQ���!,,N3+*"���+t:/G������#��MM���rmK�����i��41��vfY�4���{���E�?��S��������v�PS��*l[y����#�ǳ#��9S�vz�����9)�rӯf$���>�`w\1X�3�����Ҝ`4��9Nr��W�G�P�35��a5/25>A��e =�d�ˀ8�>MÛnuJ�cT?�Ut:���u�I9��iU��֥��Z��YS�0c�/���ON�n�\�؋u�.�������E����c15wy`��m@�0SsG���p/��F\$�sy�����A��I�E���Jv[�Uf�� �Tsu�Y�L� ����d� ��h�Y��4/h||�it���M#�5oj��<�8K+�0(bY��kЬXwل��	�ږ���lܸfVw״-k۳�ʉ��NM�tlҥuNԞ?Y���Ա�cG+�9~`څ���y��ڟ=���/�?�`�O����/�ݖ��'u㪬m݅����\�qur˒̶���g��3Ȥhu|��@�#d*1R;!ub�HB�B�K!�4���'0F��"�d�7E�7%�7�Ao)�ޔ�zS����^��Z�[������HŸV묪�y���'?���_���#�Ok!mi:ZLG�S�G),o�t?f~8���G�~8R<6�����HD��� � T"�$b01�!�0��bS�4Z����m��!/k|��75�ʼPfb`B�O���?��^��g70g��i��"S� Q  ����� �ԈXi�	D��q&�+�f�˲��6"݂%��D#g�bup�V�G�EIQ:�ͪl�ԌJ�*+��������:6�j�w�#ܱnW���4z���NkFbtuI���53'W՗�LH�N�̌w�DX�̬�Q�	'k԰K������*]��II��N������-��pR�S�O�fQ�AEa�b�r���R��R���d�!�� �K*���V�O�,L0���[Y�[勬yWK�����V�!?�:��P�Ӟ�E�����i��
gj*M����Ŧ��֙��Ru���/�h~�̮��7��_�<��Q����Sx��+���v�m_q|o��-��M�VΫ�LM\�NNSOIc2���dN���Y�i�$��kjdM���`r��!�4-�6� �8ٖ��0".jU�Z"�rT*�\I�x��IdB�P*�8K�U6���w��k|�(�s4�z���|�D�
����hp�x\���`�_���M>�$/�����h ��I1H�BD%U)�����"\)� r;ǚ��� �R�`���LL��fJ��{����FT'�UIHu�M�xS3)Ře��Y�]��c��p�
�)�ұ�
?! A��x��P�!J\ a"�����e#�q�J ,�!r �$͌��D�^�i�&"�iXK�z
� HN���DT!$4
R��S���C̨<J�{Le���1<���5dY,S�e��JRW%�eqTq4���%����E+�	I�("�% �"�A�0,Q�D
�@,�W�B�Ra�P�`I�%%9%UŵE��Κ�hzrvB��fs�"��q�Q��a�������Ą���̄�i����H�"4�
�,
����Kq(-���`�28�Fk%��4������������J�H��{Jħ'`CMͼfA
'k�k��>�f�9�lsk��9�i�$�\X�Ya�V�+�*Z�;�.B�N[qA�)�[%�۠
�S��6��K�m�ayצ�o�?���3���4���`O�	�>R@d�{9Ǡ�y0hj U����A{���i�B}��4�6��I0�0�
�_R�\^a��w4�f>�B�ɔ��*��P�΀����ev�����,*�<��=?��AQ_X�w������M�i���*|�
���Q� ��W}J���35a�(ɜ������v�	���|$�� �/޸;��c��Y�ƙ���Լ(��pA�eQ����Ԁ�PYÛ���/45 ���N7��S3�h�����a��?|��vf(��yF�x|jf����lh�����35+gn[3oǺE;{����������15��Cy���飻�{�ԁGw��ٽxMc�����6N>�q�����7��������T�~��پ(v�|��9g��̍ܽ$�`k��΂3�SN��za�ܫ{�<��������׏�~�p���^�����뫮�j8��j�ܸK�6�Fw���7��Q��x���"�~l��-Bš�X q����!A��B���B���!A���T,S) �@��� �����G!Q��
M3K�"��X.��t�sbuY���X�T�-Sj�� ��圠Q�泀%y��\�X�}.Mź�EW��35/55}��Ccj�N�����nN�͜���b�E�_p����o���iS?�9IkNPj�q�=�55Ϙ��޼����*� ����
N��#���QrD
���$�~	�+��H�}J��a��=���Q���'��1�G�{1'0�$��ǘ�uD�<"��jt7���R�~^S���=��ߦM���S�Oe�I)7���s�/#�e����㪗��^�55w �]�@@_�{XLoj@'oj�}�mzY��w�@��(����ݨj�  ���@Q�n5ԣE���f��B�6��z�U�\���1�g9fy�a�O7�'$�Iƿc�IRk�՚����(T�>*�@�N\�J�"o4̀�)Ҋ|�&S#J�H=�8�8��9i�b#æϝ�l������o鞲iu���G���[yr_噃�OL~�܌�f�}iڥsgOW�7���i�Ͻzv����]��[~�ڬK���-?����>�/��Q�gK��6��mZ�־4u�<sY�)7ݝ���v"j��,ңR*�#7.���	j8�PFH<M�R�����d�<t���r�����T����KF�*��c�7�b�hgL��t��;_������g�}��»�Z�$�̵$�!�B�SG�(��RK�H�&�$��8	�`c%�+X���T���P� ���BEJ�L[0�0�&H֧ixS��y,&��l�[m ��j1��z��[�i����1�+�hj��ۋ6��`���loj�^Sá��D�����@D!�$����P"v��X#�55\y�(�d��s桂��P��\�<ςqDა%Ql�M6�F,N��h�H�*�Q�1J7�
נ�: 6Zi�dZX�Gj�����UHհ�ʒQVsRd��nu���֮�:��WXjBlJ|LvZREq����K��Z<g��U5���c2������E���BA5�#´�S�:X�A)m��JH������x�N2��D�e�F8��q�!.�&�r�x0�sT�Qձ �75<\��8�>��HLI�x_���𦆗5������V�˚g� -\�wGMDgm$ 4��7y���[*b�����g�������05���JKs�����Xnj�s-.�,*�͜`�Kb:&�]����ٝ�uol��f��s����ӻ��/��O_��?��w���G������ulW���=;W._�xr}���CT�����>���L�Ґ�q$�<S@{��4�r��a0�fr�zR��>��5�r̳\sJ�*R-��L�
S+l��U�@
�@8P�i)��$ � �U�B��[���W=��*����� � 
P����U����� \��R�-�=p2�{⊻����b0$	�b�\(�	 �P�D*	Wډ+�PpA4*��  ��(XB��$$�T���R>�0��*���h(�@��ic�������fr*�a���T%!��pU<T����u	��$��d�K�̒@�,<�EB�H�\�/��X��*)�
@! %FH)J�0ZN�JJ1Z��H�ת�R����nSX�%<����aa�zB���b(�0�b�0��HDb!J,a%<�-���ctJ��V{,ecE��2�Tk���Wx4���K�	@I����T�k���I:�/���#��p8ɡ�z<H�zиW������+��`�,�s^�	�����\%y\���V�����ϝ8t����#k6�N��b�¢��0���qG:\aV��	wY�3�b#�sըT��Ԩ����қ=Z&F�b !��?V:�5�?Q��c�������Zq~Q�iH�MMf�&Q3����� 3�Y)��T��dz~2Û��������ڲ�+�-q�F7��@���J+�e�;ղN�4]��t ��pHܩ
Z�� ����+N�-��^��H���I�Ȩybм�c���}{_��'�J�^S�5/15�_��ѣ�|GI n+�a��� �"j�=Ts��������B�0}EE\V�T�e��g�p�^�p�F��+9Ss\�:����
���V�n;��%&|���U~�g�DG_2��Q���Ȕ}R`�T�4<'h|�4oj�P�75�J�&�� L�>��O�Ʃ:�i���f9崞r�N�[�E[Ƙ���{�L�M��kS�+����,C���l/���B�L�O����\�w��;��]�a��J���ߧ|55u�� ��qq45��0@{��s\�����7��Чs����+�9��^lj|鄇��7��9�����S"�Þ����|kjV�޶f���Kv�oڽ�eۚ�m\@���jj>~���>� �ɇO>��_~��'��<y�ʕ�޽[��w�ڸb��5��M��0�w���꼅��s��k��ٷ�l_wiߺ�޵%��r��������������u(������l]�mi�Oր8�ۗ��X�}Q,�f�pŞ�l��sQ����[�o��a��{i���u�v,}ؿ��۾����?=������a��o.����Ǜ��q���pGa����%vLKm�2�ٕ��x��M���	R�A�X� 
B"�J�e�#�H<��E 0r��7��AP0G�xi�[���H��$�T�����_R�^^�X�g\��_�oh*2����J�-���b[s���X�X�]^��M͢
���g(��y�aK�����>��\����ck������YQn�MMg��75��Sf�P�ܜ��=!�`v���+Y�7����J~7;�N~�;��W3�O{�O;��s:�q��<�qt����p& �_�U!{!d�
�Ua�vD �����@�� Y�퀰#f�1{�Q���Ѿ_c�Ov��6�OA�u�`v��<�j��#��$�SJ�����7�a�de�n�Ŀ-����u�;����hv���P�%Rs��_�Ly����u���"�{����Eػ���Ӻ{��.��|B�S��A�;���(�Uz�aw�䳀3oy��\���0z
����Xu V���>�G�{)t�l%�����T�&dkh�j�j�^m@V����U�l4����b4Ϥ�cR�0ɧ�d�M�z�Pk�?�7J�L�滙q�^Vd p�����F�Ɗ��P��Ύ�'�TMH�..��2mݾ�IMM�֬��mSն��;W+�t����'�>;�ڹ�W�6\�t�X����O�y�����/�[t����W��|��ֵ��4�8Rٻ�t�v����6���۞����P=�!zj�kM�K��������JCTlB�R� %nF�`�(�2f��%!�Bƽ�cG��������G�BF�#(��o;�Չs4q�2�V�n8����{O����>����G��\�p�ڪ#��m�X�y�^�i(m5���ׯM��3s����eڤ�z�Q�Ч��I�1Y�� �@	36~k�tL�\ '`B�Rj�d(��Y��Jqk�j�^k0��&��n�lF��`��tF�^ϡ��VCRNP�?�C޵	`�&l�����s���<~����s���ۿ���Ⴥ�}�6�(l��`�(U�B	�*�\!ss9�4�b0�3:�(T&(�� X�C�@��E��Hr��LA��4Nf#��\�y,Y�|?<� =Pq )�@�0��z�"�:7��tR)V*���IH��Ub�0y1�
3�23�M�9���ƍ4�� 1��Pʸ�&��ҸݤwX#������XOJ|�'�FBlzr���u��Κ7{ڬ��͜:�abmEINFJVjbjBLL��jа����q5.=���N�Psd�4bg`3�0�#,2B�TF)<Z4��e8�	.</�,�`�� TqQ���R�1�r��4�\e��D��	8/k��q�����/25͋�,KK�>A34�f`�Ӑ���� g8\�M������\������zOg]�c�����U��+��6�mWg�����^io�r�׺yZ����Ͷ��:��<��<-[[�ե���˽���U�7���n�yr_�/?}��_��~������ڽ����gl?�k��ͫ�k�H4x��25I��T]C�~J�nr*;)�?.."	��A�XC
<%���ٜ�TbZ:5-�V��E�p�nҴ��Y������,�*Z#t�"-�iP�Ar	gB��#T"�K���B�P"���А �T(�$�P h�C�\�RJqX�C��R/$
����D%��oJ�AQ�	0�&!��iB��u#2 hx�aİR�&�.Y."`
.(�[��hD�b�gx*ՠ�А���d�R
�T)��J)0b���`r����o�<�J���7(IS��N�`'�3\�'.1V��T%� .�&�L@���D��TC}��,��0�<��*ԉYa)"�"V!g�2 -�"U ��C�R�����T�"�ba���ä�,H:V@��0�;�툉w'�M�&�lf,:\΁E!����0�Ch#�p��	"�
D-��!�j�@#��_'�b����VVi)ri+"u���p�.V]�! �MSK�R�1L��-��U�k������tCQ�&+�L�!5��(臒��T�q�б��J
+%8� { C"8�R*ĐJJ�FM���%B��'$F?|t��_�����W��Ճ��?�ѳ������0��ȸԸ��,Y����
�Q'	�%B��D���4�0
�ŨL�������CƎEǎd�2F��~�jQ���e��Ӓ�I�ȔxZ<6;�����IT�I`g'��u2�����&���~��hwK��9˸<]�,M۔�o�0 ZSM�t��msЭV�̈́���v-ԡV��.\�����+���ݐ`3"܍S�3z������?p��Y�OL�'��h1�
}L���
�=��L�Dsˠd�;"�]�7��_���=B��0ua`\I
����|t6�GIp�F���m~GA=�� �c��jz5<��O��p�܃��"��{C�~[�\V���t�=��r�����k�
��q�X�'8��\�'����>���8'����G��w�"��l�I�W,�I���
.�]퓩�J��3?����5a� B�=�8���>?���h�F{�h:m������SN�i��d��X�Żʼ%Ѹ.Q�"Yמ�o��7e�gq{�^��^��]Y���̳,��R�<˒bòRSc������]��\n�V9��8��Z�h/vt�8W���,w�(ww��@gK�L ;+�+k�W�GVԄwT���.��4VZ�*�UNp+7���Hp�72/���`P�U�������ɋ��2g[e�.�� ���#/kڽy�AcE}8/n:kdw�bp�������?�O�tO�xM���q�ĭ��=۳~n̆y���@���aA�I&o^��eI�k���?��z}k����;�n隳e��k��X׼��m���k;����������jj �׀�C�����������?�����}�35�Z�wL��5m��i{z��ml8�q���o�?�~��}�7��m�c�.��1�����y�=��w-�ݹ ��po��ܶ qw[���Igw7>�����;qg��><��O�<��̇�+����k�?������cŽK&,N�VۤYĸ����xX�*R�E&�I�P�%�D�K��L	����+g�,/p7��x�h�M�{t�di3+׾0϶8׸4�ؘkj)��;Z�Ú�ݍ���"sS���P�,_�4O�8�Y4�,�e�<
�\^��O{p�\��	 ��� ���o)Է�KL�L͚2`��Km�[\{���D�O�\͎���p'+�nvʻ9�ޤ�9ᰁ/�SZ�Q��-̳�o��#J8�@�����#�`l�
ۯ��J��R�d(|,@y4HuH���^�ݭ�o�w8\�=G�bODƝt�68����J�0a8�j��Tw7��'�iݯ N������$!���?�M�]M�W�7��\���
m�FO˰�0�\Ss��C�/�!����k��;��V34��%���4�@���q%���Ñ^o������B���!�k��R��A]ZU�j�#�����6(�S��IFY�QZk�֘�=�7��LJ@�Q�1��z��*�P��ThĀr��MM�V\jG��p�Z�,�h���Df��U׭ھgZK��5k�o�P�u��{7f�?>���i�O͸�?��9W�̺�?���Y��O?zx��ó��s����'�9��ܙ���N��W�c[ᆞ���e[7���Y�gW���U{�N��
�3%i�)�Dt�:¥�u5�+5z`�dfB��@N.����a��N����2D0&�ǯ�1b��W#�o)��l:e���-c��U7j׼3yͭ%[���h��GǮ���/��k?���;�v��h��swެZ{q��f�xz��s�t�ɯZO}����v=I��-qҦ��.W�b{�,S�$"�P��E�!J}����RDSz��`�35VmP��Ik6k�N�������Qo����x��i8���L�]����F�취O|s����`Qp /kHE��Vx,x���g�c�g��s4�N�� �1PQ,T�x hn���l�.��ě�p5����DHKE�\+5�R���4ff	��v�Y����h����8����/) �m�0.�9���y"��Sb�>1����q9�iS�kϟól��y���WW����p�'�e7t,��5N�Ω�:u�C��Ԕ��m0�J#*7�$������qF2Û^'ϭ.��y j�ה���LeUG55)�qH�yM�/}�S����@����f��ӷ��9�3���6���;�5oj��6�'��p��&lU�{uػ����f.��i�M�+����U����容���$�"[X���X��q��EW-i8�w�7��Ù���5'k��_���Ƿ/<�~��N��ػ�kG�ª$sU��*AS���K1LL3LJ��'s�\VfzJ� IdC2>%�4���LI����ӹ�����.��M�2�ɷ/,qOM7��4�,N/s1R��Q�J�]���	�x�:
������&$� � �H%0���0g�@"J �� �J�Ëo�_.Q�0HDa2�T�)C(@�@$$*{ ���K*! W
����P\. BJ%�!	KYD���E����ԀJu����4$��.��L���S314�kj��$�kj��x�6���l��ӕ�3I�̭
5ǫ\�9B���d�Z�Rb	!"n4�	��P�*qZ��r�"�H��˃e� 9�wF��+��kp�Y��S�Ϣz5f =F�zD� T�bJ�Ra��T�(���))��2*�HN�0"@���U,���2?�Z^a+phK��r7S�«#��(�*
����8gjb��XP�a+b����}Y��4�X��M���m2#yE*x��)�2a���%	KB�C���
E�b�@��$"�	L �D�889#���~�����������?��ӳ7/oڿkn��ܺ��46�l�+�-[�i����K
0U(dS(��J�K,���~cǼ�֛���8n�`�Xi�x8(�	e"�P�k�������7Q�NI�4$����)��8bV57Q����Y��55���,cS��1Mג�o�0 ��t���v�eWw��3�a��uh�F��(�0Q&^���@�����
�H���e�5�+F����S�ġbվoTl�|�W�c?��OX��?����!J��DxS3��������<���ac�G�>� _��Lr�I9gj�tUF�0_s�܅4�B�[J�u��m������dN+Г�S�;�s2/
�35qX"���{D�3z퍘�w�b�$܉��~�f;�h+�^��Xy�[�c���{%�n�@���04��kjp>MÙ�:D3G����b=k��u8�:lg���0��H�a�e_�e{��'�Е�kO��[S�ay����3�C]��E4�ei�pG�3L����Ԕ[yG�Xjm*�𦦵��3>ڋm���BGg�����U�U��,uu�8�~E����E@����Rak�q4q�����U\ jK��Z� x�� �Ua]���
wGyX{��kj\��֊��ʈ��(������\��(��#U��U�����w75��w��f�����6Ύ_7��/���ٰ̊ 鹦�_3��SS���nC�oL�ܭ��XӴ��mWw׎�ۼ�3��'�>��	��Ǜ��?x����W����ؼ�}ꦕ�����o�������<�উ�6M<�q��G6���S�i~��y�f��h�ֹ���bw,��Z�qF�����b��L��^b��'�|q{�/�|�Օ����g�֟�0m��̾��k[���6�@ㄮ*g�]4���J��%��ɤ$�ۤB�
2)T���*(��VA�R����`uI|	`��]�-W�BU�@-�2c�E��MP��4��6,��/�35Z��l�E��"��Bkc��g^x�h�0���2�L��eMS��gj�˚B}k�a��YQ�ɚեV��!�+���w�D�/����ˉ��'+�^Vʽ	�wr3��˸����	?j6��O��㸚��=���Y�g�Qr˝������;�����K��0�Gh�-G��zN�3q�G��~5o�W3�}PV�nj�N�=L�c�>}ѝ��`�i�����
��\Ҙn;��%}��������0��-�,ƾ��_���ػ��9��&�p�4��y@�R_�wqn��=\��� �kj����YSsS��L�i9CG� ��Ca>�f����|X�L������X�
��K���(�t�&�j�^���U���zy�^6��y���4^�L���]�T��LM�N:A�H�@�$�@gG:k�ӧVWUVխٺ}�ʕ���ݲaʖ��o]^z�t��W[�}�坫ͷ��ܸ�r�r��K�/�]��v霏���;�\ ��u���م��>�;��>~?m����噝˓�ΩX�\�x�53�Κuz��D�`J` FBj��,ʀq)W�B9h��p0�� �*$@1z�LE��S�r���k뛳���;�z-?��9�������?[��i+�-�|��͟���/���?���?�y｟�>�d֎[�=ת��.�t#ݕ�U��W^.^y�dŕ���e�*��˛�.�=a����vg�L�S�q��F`Z'���j���,K�oj�joj��Ekq�-N�`7`3q�F �cX�ױ5����1�����9^��n�:~�Mx#o�N���l/��05C�6��'�"AHp`��8W�v<"	4�2�]�`���t^4[�.����LQʸ��gt���5\L�7��kj���0��yQLN�&��$��(bŕ�T����J*�+�dDibp���X�Ic7i�֤�j�¹Q�)��!�fC�����hxS� =�2�M�o\��e����e��M��ϩ�����HM���
Ow;�V�ΤSkj�Z�ih��z�ԘQ�s��dzˊ�k
�4Euq���C�,�����qXM<�35�LKc�uO��Y�o���e��y����_X�%��m����2`j�#���G��ή 4VՇ�15mN���V�p�*��q6V��U��W�/���m���jS��E�i��&�Ω9�g���~�_�<}������?�����?��΃�g�>�wv�C��2�j��5���$.�im��&IW����|]��>�L�bR:)	��MLD�щ)��4b�7[ojxY3-K?'߾�8lf��:�)�$��[-7��� #E�F\}%�"�k'��hxA4L��� �z�	bQ�\&R*$(��^�55����xe�5&��!	�ˇ�����^��J!�u4�����Yt�܈��D�Iը�F� �%���Tp%���x�*���������1��LL6T��
]t-s�Bt��(�q鱤BF��*a���`F�-}"�JB��B�� �2H�`��pLB2��3���
�Sq��!Q#KZ���6���H�K���n1(�4W�[��%�J�"R�TP�R�Q��Z��	�����R��{z�Iɳ���hWI�%߮)r��.�Ȏ��^ӔG���X� ��5��,��)IД&�JSy����a�	��A�k���_,���4^���%L�'|m�[o�-PJ��hʤ�⪴�	�����ӿ�����������ݏ{��������8�m[w����}�]8u�څu�7�ϘRT^����H\,
!R���T��;�=���R1!�A���Qo���0�UD1u	�I�x�>��N��gƓsX oj�idj�d�f8Y3hj����8Z3�Y��tCc�z��nuм�i3�mz�U���vZ��v!�Ո�m����N\��T��#L�sϥ{/������U��Y��Y��Q�S���5�1\X�{$��}�D�� �{r��R�]��_�į{�G(�e���p�B ��<����@�
0����勤�Bw`�Xs���nC4������/+�
ꂜ<� ���)ү�8��Ys^�qA�H�B�a�������58��V��^��_K��u�v�f?�3pa5"E�Xɗg���=��^f�j^bjR�a�=�ў0}���~�a>�2��0�X�ƚ�&��%��Լ0�f��'/� ޥO�2L��XVl\^jh,57{i*1-/�h.�� ���)���[�,��bk{����h/wtV�Vք���XY˭��t�T8�m���
�Z����Tao,s,/�7W��n��Qob`ΡT9��S����oXMe� �D�>^lj��5��a�TL�s�	����c�oL����꧍�7-Jټ8u��gٺ,����ll�����~ڶr��5Kw�m��Ӿ��k�ڎ瘚���=e�x#�BS��{��{���̛�/>|�ɣ[o�ݿ��qm˔�+g�m�ӷi���mn8�i��M��mdS��*��E���0^bj��Y�ma,`�ܨ���̉�:7fǂ����WO��̌]=;sKS��c�����������7���ӿ���Ԛ�}M�}M�W7O}�ѥ���*k�#��-+3	���<�4	�C�1�ܩ��`Ģ7i%+W1J�VA�
"\X�3P� 0�!@����`�#��r��B�Z��F&'jfg�d��9�����}�ni�z��eÛ�i<���]�.k
t-�z�����~ZU±zk�-݅��e����'�/f��̊����0+�Qv�{9��nd��G�������e��-�K��s_Xę�>��~JAV����^��I���/ܞ;����?������Ǐ?ݵ�ߛ:>���U�9S�_NGt'�	��J}J��K�~9~FI��؋������~Ac<���Ux?B_D�`�
��I_SsS�B��^������m�� ��_}��sM�Kbjn(�<8�T(oj�#�Q:�B���^�e_�{-&]��VS�U�|� ti���E/�BK���Z��|�N6E'���;S��4�tLͳ�&H�Ez4��dQ\Ԥ����ե��-+W/[��i��ֽ;���t�r����w��z�J׵�m�4��h:q���Ѧ�G��n<rh��K��Yv� ��{m͚UU�V���=Ӷl��u��m�[ΞZp�7g٢���l2����Z��`n`�&\ngT��	g�ҧH-�V�I-�!�N�Ї��Nj�ݴ�f�ɏ:�~����[ީ�|�p�;��7�ֽS�y5��kN���;���'{��_�^���l�gKߩ�\��R~�ռ���{�嬺��~.��\v녂���gJ�Δ��,X�?o�Όݞ�&Ǆi��\sD�5"������Z3��Sj�/�F��xj��Ţ39���q�,+�j4���F�^��r�@��;���hxM���n�:xp�x#>�l��8a�����vƷzԷ�T( ���cG�%?Z%��c�#�35%�li�?kj^SS�����T^3!B�j�c�p�2�d�(
�GC�H�����L�A5Fu�E��xYcֱ��~-CZ�p�-�������q>S�c��sfM��ִ���yUg`��9��%�2���pW��	�n� �@M��f�[��A�2� |d�]C�Y�J�f����Ȟcj"uE-�낹\���fe��gUƒ\��AYӐB�2
��xA3��PY�S�3Lּ�Դ�E��F9��:�0@{-����P����Ym���:ojZ*->Mh��7s��>�ے2ײ
��"��4uU"Q���Q?1?aIC��]��xr�響~��7������;_��W_��٣۷��rd��]���j��;eBX]��6��I6V%�+9}�Vǩ�㘚8�6���c&Ƴ��x�>�& u�h}61��L�+��5Ӳ��r��
�srSҌ�)��h�G�4�b5"Ad�D(�%�t0S�L ���g ��w4������3n�H�x%h���� �D���Q�0T�P��[���5 ^�"'Q)��B��T �TҸ��gmhD
��yA�;.p�+e�$�,Ri"��k&ע
5�dP�#q�����$�>M39S?9S;)C�]bjj��D]y�z�O�B��$jeZ.ĥb\&�>��6(h��RK	FL�"��x(�����2�BpD�`b5.�`2�T��Lp)�h ؂�6�
3��6�UG�q:}��X�X�
D�H��E�LB�d��АA�i��y�H	�d��U�c��,ͦ+�/�v�9�E.uI]�@K���H�2+��~�E�E�dA(�b�c��q��8ui��8Y��${p�6���l�x���U(����C�)$"h
I5�Mё	�9`�L���Ls�&�#\9�էn_��ӧz��O���?��_~u�ѝCo��x�@�����];w�����7/>�s������s��Y0���E�ɩI��Qf�g�BL�+Q�)B!�3V��O�~v��8B4�Wz�I	��	�I�S3-��j������,L�,��
?-�6�y;�i�&�S4�i��cg��5E�<�Z��Z��i��D�ig�6J�A�ZU!+ �:D��lŤ�����,rΈ_1�8�܆",?u[>u�?��>�>7�?3�>ѩ?�0OX�=�xB��Ü�y_��Lu_��'�?P�f��M�W�p��1�yB��'�P��}/k�(0b�G�\bn��^nB� ޿&^S��+*겒��$ ��Y%�35���K0qL(�G��cJ�O"�4~<W';�u!>�R��\���|�h���N��>�pS�������4|������j�q���|�j�MM��t�i<n:e�k�cjV$�oLͰ�ߒ7���4�h����F��"���9M�<S�Vfo/��[[�,���ڥ��rGG���*l�7�ZgUX{��bM��m˫i�1;��%��r;����q�f��h�f��� /�R��w@��O/45������F�%����V�}cj��O<V������l��K'�}��k���nݳ�s�U�Ә�?���#����ɻ7.ھ�qM�mkg��2�75�L9�y��͓|����UL�?��ƋL��E\�'�m��X��}q�%)[$l]��kY��	��=�%���yp��Gg{~���_>;����t�v���K��,�=�ZԿ��HK��:WC�0O�ƴdJ4�͖9�88 L���<8��V�L�BATJR�����o�^Ƨf�D�8�$�%)5Ekh��$u$��!"1�!N4(�(��c_�L��,/4-+�/�� ��ky��/>;3/��I d��d��eP>�ɚ�|ms��OUÛ��e�55�l�J��{NM�\���H�����^Vړ������d^K��w9���~;�ď+I��<�a:�р�w��kj���S�����P_(|@�����8��`:=!�������}O�_xz��ӛן:����{�՛Q� m>�j�d�1{Ҝ�ѧ��)�/B�%�ivZ��T' ��*��=SWI�eLsV�_R�ﲦ�����^S�g�yD3��ޗ��K��2w����=cj��ѫJ��
=!��9�1x���e�=��F�1�:\ƙb@֬d+��.��U�j�B�4�EZ�\�|�V�0hj���|ߘ�R�̗Q�X+�&O���dh�$-����梄��	�S��Z�ۚ;;ۺ׮ܳ��ogہ�s��L��^�ZҲ,w�܌Y�ҦLI���\WY^VZ�,.�����̟�q�u�u���*wY�5?ϐ�媬��T�*���yr'����Sb�#\v=��a>�^l�n��@nZ� ��F�MN�͢si��	%�WOj?T�u�d���o�o����Rj�ռ�w���)Xq���r���m�������GO�>���c?�U��ǵ�.�7Ki�Z~$��tꪋ�+.�5��,<��H���)KOd,;���/qֶ�����ׄ״�ͳŗ�����ڢRu�(�`�4zZ�eԬZ�h5�N�6ju���3Y�fN��8S�2r��i��,6��f3�-^�jPZ��eY��}��n��G��7N��3��#lp���|�l/���#h|��WGO�?~����Ǽ�7R2V��p��L�r=����	��pO�b�!/��)�E�bp0����"�)6£V��TL%%�"8$
�t��KYXe q���jY�Q�]V��b��u��%15��XʤS;�&O�+1֓���+������ȘHw��YV�?o���-kVt��j���gT��d�&:",���f5h�Ө��4��:�ʒf5���a��M�#cM���0�[���>Es����Uͥ����b��8�Ǘ�fh�'��	����"S���.k�j#;�=�uQ��ЛAS��5#E�nE[��Ze�`�
⇏�іJKG�˛X��ryM�^Y�XR�ZX⚙c���T$0��΢$缺�C;V}����᳧�����?���|���޿}���[�m_Ѳj�칕Ӌ��"�2�U�֊dse��<A_�E*�z�S����5e�tuSOWƢU��:�+=@����u{cj�~���<ۜ\ǴLKC��2єh��ԀKp� �b.M/��w`�Sp� �8>�\����F��;� w���D�J����2�J�g�aPŰ�1<j\�E�!�ZR��j\�bҡ��oA�Lƣ�� � �I�H��T�H��.g1����E��2AS	~�	dM231];%��RS�ɚ�S�y�x]Q�aB��\/
#��r?[�P%V�!���8��q�"�2�����Zy0#�'CǢ�T�FAB�N�0	d���nJ�\1cު�-[��]9efGy����%�`K�[S�E��d�I�2Jz�\'��dR�\JIh��0�/P�7F0�U
̚�xwU���m(qk�"ե�diZ��E��QhqZ��򣱼"?�*�bʢ5��$�?,J�N�aÑ�(Ң��e��~:
�dj���M�q�%��ks�Mɟ9-sr}JmU��Iۚ ]m��N��n\����o����?}�����7������W�?��+�/�l�ۺ�����n�y~ձ�����z��'�]8u����'�wo�ܶfeg��u[7lٵm۞��M�̞TWY��S�����P�	�7	��� ��TD1���ɉ_L/kf�R��h���O��fi���5Y��n���Dfy"ے�S��4ck�fi���X�#ޡ��5H;�����+W�B7��m�|��GA4�1zF�^6����0�G��ϣ?�t�"���������I��^���!�P�{!*Q^�<��J������܇8Y��cj|���5�ǘ�!�އh^ր=b�׽F�S����J�O$|Q�.(P�y%zF��V�g��U���/� �XuZ��A'a|�P�=��;�ff����q������^��C�}J�K,05 ��+������\�k{��9D3�X�Q���9c�55��m��dӪT����.h�,�&b�!��E\�P0��.b���R���'� ��*gG�����Rfi.5��Nk��������_Ɨ�x(\��wuՠ�����w��78/��6��"S��� ��S�VM{�d����}cjz���LͦE)��y[��ߘ��ٱz��u�M���iL����� ����_���<�⃻�/ݽ���m���y��.�W?�4���ɾ�O��U15C��P|jf/25ۗ��-��r�,�ݲ n�������4f�k��gy������%ۗd���jz���E��6�΁�<<��G����/�l9��v���3�7Ĵ�Zf%�j�k]��2�]?%����pQ�pP�40�T%i�p���A�R+� RQJ���*.|�4C�̀��-�t�z Zcf�:Ө�Xt�*�C
É�D������,�W/̡�P����<˜4tn:�����Ƨi|�|X�3L�p�i�����U��]���о7�}hBĉ���7���ƿ���ф�'�n�ǜ�ێ�tH.U�!	rT��F�<˰P����Du�[�i �Fř�^%�_����m/��i0KO�x��z���������?�xx篇|0�̜��G��#�>	qLN��3�E�I1~J��a^֜��'$�1tD�E�}�����*�^Q1W�CLojR�ǌ����5<`��(�=\}e�
��55/���&C�(��J�75'P�8���^���^�O�}���Yl�n ݄|!�e�ZF��U�� j�U7k8Y�@������P@�D�|������LMɠ�)�5�34A�H��q�2ͤ.��L/)X0y�ڎ���m�3�Ϯ�ݐS[nM�E�V�eV�M"�:�"�!�O.'��K^
~,
�ah�B��aȫ��21`4��	�Q9�h����R:]dt��`���b�Xl��IQ��1aFcT$�U)��a�2�QŰX�����#u����Z]���ܲ�nŉ�����V]L]�vr����s�=�
��6]�X�_����o|y�ߞ�����~��]�}�����U'�Nh:��ٟ��jᎻ���O辑�q)��\J����S�O��/b�FG�J[U����^8בX�k��0�t�H���h���M�A�6k����i,��45a&NӄY�n��n��p��`��t|(�1�����0G���s4�+�|���������	
	�7��Ƞ1#��G+B�j`A�N�35�1LI����`@�<?�ƛ��KZ��I�RQ�҆Ju���J0������K�d�IK�LM�����դիi��5��$��vX�#��#��4��I������� w��Y�Vuu�^������i���5����iI�q�pfBL�'�ޚ�F��ș�� 3�z�kjp��Q�a���Q�����\j��0�_ U�F҅�d��,���=���*vǢ����E��С��gv��ld��M�������jj��O�a����i��Jsk�����Y��Fs���6���=�i����[�_���R�i�b�B��ˤTMy<]�dˎ6ͬ�9�m��[���돟�������|���;�߷w�ՍZ�L]4�jJaƔ����*S�%	��8CQ���D2y�T��*���"�(���u���Yy4Z�W���$ 4�Ⰹ)�䴁<5ޤ�\|��l��lsC��!�V�f�pQz����**����˺͛IH�((h��?f���ƍzs��7��gj������/�ﳦ�4�ˍ�!�:�[xS��|�q�s�v�'h|s4<Ra"ef�Kѭ��㘚�D�0S3%K�5/35U�oj*b5�.:YGRJ�JL��H�I���!b�@��C�~�h<!`$��8X-	шB��P�Dh�K�J�V�a(B�F�le�$-�=�Y�L�������O�>�ͮcw���7�h.xH�GZҭ�BKT�����g��$����N��"U�2&0P�7.$( 4�o|��X���XwUrTA��8BW��>E��PSS��4�PS�'��؂u���w���A-D� ����ڨdτ����S+�-��jԮꚽms���ug�{ﾻ���էO��ۧ��[�c�����{���?��/���O��w��{�w�����ذ�o��{��?�����<�{��;{n_�}����x��sϜ�=y|���+6�4�h��t��铫�JkJ
�K
j�3s�"��DM�SԊ\Z�L�WONPO��'���=H���N�&f�Rs����R4%�3� ^�4�j�%0���DMG��+I��.s��-�ҮC���䝘�������m�|7��4��b'��Yzـݶ2�]��FX��8�	����s��+����gz�O���={��Wr��#��y$U>��KdޥO����| �_��35���A�d�s!6sS�]� \q�o��|������Λ^�55�eܣ���)���~�߃Դ�k*�V�\��<u�b�UkvB��P!�<�O�w��K^#�rм���Ŧ�)8e���f;���D��H��7޺+ɺ)Ų&��}cj��{�(G� �9<�h8�qs�兾?�s�����Rbm+����8Jܭ�^�\]5.�ttԸ�����S�y��9�$��J~E�P�JR��֦2[s��R�n���r���
n��i����[*���y����h|�z���Ԭ����L����15=� ���@mY��2�٘��75�㘚��������|���/>�{���7��tN߳q�����}�&�X�-�=�Q����ULh<���KL����l^��0/�gN�Z73z��'�i)<������9��,`d35�rp��?~x����������k�ZP`Ꞟ~�L`��+kÂk�A3���r4��I�̔8]u�:]�H�I<AM{�E�#��5(��\�L����⦡�3z���h8eCkX���Z�d\,�Nh�3,Pu�zj�~a>W�mq;?�X��-�{N�<��T0'�e�PS�5`�x0[ojxY�ս�fy��)_�Zdfj��QxS�cW�c��x��\��FB䃔��2�~:!�fl�q�~'��PA�*d�:$��JЃ^��,G(��9,�����AG��`���S�lQ��(���hB��K������?��Ϟ�������_����<|�'RһQfi��^1~TJ��PGC��T|Z �rJN
!nɮ�ybo�����??���r ̰�O|LVs��p�0�\S󒘚�bj��DK�e9Y��Pn$����&�h%_��K�aG�n�B���yZ�L�|�^6I��������15e:Y)�S����S�$B���
�m5����'L�������	�V���`�p�k?��#���7^��OF����������W^��5r�[o�x��o�1b����Z@����#F��9�{��WG���?�Ɉ��J@�h��2Y��Ӳ�KKKS�c:&dF�Q��IE����1,����j�V�V��Z��kqefV.M�ԕ�`Gފ�	�Ư��l?�j=�ԟ�u5��J���q��.9V����#����s��������N=(Zw6��DZǅ�g�z��n����f��+\X���Q',=���X��>ה����vcy��h�5���N�Zb��5:���Q�V3-��2�<_����$ܻ�I�w�.��e4�͖p��m����N��a��
w��V�a5j�gL��fj�:���Bh7�R�k��y��5�/��gjxY�?�o,7�?F4N)�ca�S����.2'��M��	��|oS�5��SS��2�1��(m���cjt� �bb1�T�a��&�eѰ�7�]6��j���%��c���{�]1��ب�X^� ���� 'k��Y֭�ؽf͊��-�/�9uranvfj/wb�"��-�+�w���af#g���^cQ�&7�����Q��F�uT��N��r���g�#��H� ��?��2�1oj 510oj����Lͳ��E��E������Q�i�����D�s�Dk{�����k��jKs�����Xin�5��������Zgs��;��*��7#�
�VE6�D5VE-*�W�]蘙o����HԔ$�2��3krz�uݾz�W_=��?~������>{�o˦u��[/�=yn]�����5��Y1e)�KV�>í�r�3\T���pYad���us��+m�bYCs�p��8�<�,��꒘�)��LJ���Qi��mC��>I;1�T�j΋bRlX��#R���T� � X)UB��O�����~!��Ǎ�3�oԛ�F�1���A0v�'�����B!I"	�d�|�_��yd|	e|�t�
`�!#~�zJ�#� -!hp)� =�!pγ�s��75FB�ù���@�㗘���*��Ma��`C��妦205qW7*F��c5��pQ�R�RK��H���j��"��J$!�q&�֦0��1g�)m�ƚg	/s�O�˘���0�hIX����1s	%�~j��+���£�m9�`��;=ߙ�u�n���wT�ߐUۘS۔]הY�<�|Q|��ȌIaI�G:c�W�����Q�H& ��B�r=��$wN�� \S���fˢ��P�E"�Qh����y���aE�4�m�fF�qN(ڍ�2���)J��]?i��yM�{w,=�����ֳg;.\Xs�ڊ˗[Μ�<����_s��<�x�x{���>������������O�?�޽�/�:{t�ƕs�m^w��G7�߾ �7ϭ�y~�;W��9��ر���۷�w�ێ��u�����V��Z�l�����ϙ�`R]턌�pg�U�m��lTQU�ak�Yna11���f����������}S��%Uג�m�g�㘶8�#N��n��]�R����{RuҊ.\҅�V�BV)���C�@�ݸ���1�a9�����E~�D�ke;���?�}��e��k��k��+��s�����&�#�'�D}�D?��
P����"P#Wq���{^�(|@�a�<� j����ӗ��"�C�yG��R"���%���*ǮȱK
Ⲓ���9�~p]]�K�QgU�T�%uQ�EE�Q� ��;	����z�|V\���y�̟����ny��ܜ+		G��mR�.�j��M?�?��L�PMsh��fj�pb?A��~�Xe���[�<5'#-Gcl��R��m�2��7�fX"a��4���a��gq�W��̳xM�Zf�F�x)o)Dr�y�+*�Վ�z��ɑ�����jWs��[��XVlm,�5�y������e���x�za���@Ep{c���,��,��ܽ�̾���5P4���\mm��6U�^Ac�����\S3D3 h@?�[Z�/��Y9��lXM����S�=�+�=t�Kd��%i�tL��i׺���;��_�?��y�������75�<�����^;ٻ�}C�ލ�o[�W�޿aҁ���=����W���3C�a���l]�ea���Q�F���fFĪ�]S#VL�������pWM_Gm���8<�*^X�yiխ�+�����61����^=w�nZ
1-��A/��6��尋s�r,ӒS�̓���a��:ͤ�$�X���4c�	���W�C,
�0<T��A4:�[� 0h����#k���V�fڠ�)F���J�$X/��WU�ꦤ�[�Y�1���Y�b>hxW9�3>f�� >���w4/Z��$���^�<�Ԭ�����xn�����m閾$��8��X����I���}:!�ݶ�V��*���1r\�w4<>S�����@Ǥ�Q�o���35
r�=��3�]z����������G�����O����ӯ?�˽�_��ye�Խ���zi�S��	Уb⤘<��O���!*^֜!��bp4@zAF\Q1��T�ꢜ�k�!����Bٛs�˻�~zD�j ���< A���<�Լ$��m)<�Ԝ�ѣ:��`��,���{Y|��D(7�����Tl�UYx�_�FWh�N�,�*���|����L�?S�35\�n�P���yjI&#IgUY*ˢ��2�D�7��#�����o��G#F�`Ĉ�xĈ�xk�H��#~��O^�ͱo�	�/ 8*0`d�?؏	���*��Ac�P �<j��^��O~���?9���ヤh�HE���ؤ����SK"�VQ��%	�)�Jc$�uD��JҲ	Z]���:e5������򦘩�'t���t+��F��I��I]s-}����˹�n����z�z�����~��C�����������s��ly;��B��k�o�U��N��[�k�$���.9��p��}���{��k�h�[e��T��K�b���x\��+��j���AQ�ZCi5�AØ��U3`j��oMM��n�DXm�6;oj\�a1�LF�A�Ӫ�	S�5��z-��ƿ�o��k�'��Kcj���)(�?�o\��Q��,x<,����Z�35`������4ω�)��xSS�����l��r�JNH��H&u�X����<q#C�Ռՠfj#h��-�N[d���2�W<�F��y"b�xSN��L[8w����l�^��sUg[GK�҅�
s���SҒ�Sb��.;xe���&��b
����F�Aka�AS�`��Q��ԤX�t;����j�½��d���0�+��+�1����E��)���32433�`ϯ�����P;3�gM8���1b{��kj�i|�L��i���>�mbDsmXcuXg���&��*��"d�*+���`^�c~�k^a��לB��"��\{m��4Օe�Q��o����g���/����{W�ؾy]��֥s&UWLH��N�R4�89*7ΑaLvhmt�����f<�A�98e��'�ٜp��{A�:?�.���\��8_��4�Md��I��I /k&%�k���$m}��$V��&L�e��qq $P
U�� D�35�����4c�|�K	� 	�	CT�PX̙T2��h0Ű�2��ѓJ�|S3LӀs �d�i�N��COȍ���S����+xS��Ϛ��l��,�w45���,;�A�$��!R	���z�0B�҄��r5�RCT�5�Ι��5˓;/&Q��uEӺ���O�X0c ���=%����ɞ�6s��Ȓ%�����fǥϖl��|������V�n�S��W:K�����Nm;8c�Q�����CK�F�LϨՆ�a�p\kCH�
��jaIf��(>,+L.a���Ev�Diʛ��A#�(�35�"�h� �Ɉ$b��c)[�ٵ�y��֟�o=���g�.�?�|�J˕��/�]y{��33Zt��a��y��-;yf�w���/�>�������_?��?{rˍ��V��ѷeŵ����ܻ�}������a���Vؿr_��]�۷,�Գl�����7���ٽjyӒ��V6/�Z4~m�����Xwy��<�P�����Ǳ��t}4���L���<��r �&I�0�]��Y���q�q��-Iۚ�n�e�b��h���t���v�Ѥh�);�\��NR��V	�(B�I�7�;U�>Ly�B�1�q=������f����gU�g�}�4��i��i��n��j����s��s������9M��O�G*�c�P�rK�D�{�PSsW�xW>�;2�=��qa5�@�V��a��}z_ߑ#��ћ2���
��R�m9���|[�_��7��M|K����}���4>Sg��y��M��1���v⟻:����_-^��9s?�����R�@�55��\���4����%���؇}$u�a��%fs����~:e=k?��؛�ؚn�β}ߘ���bjru`.�$̶4ܤ��-_���VY�j��n���(�k� �.,�.�p�M�Z9-~����S�&Ew�F.���ey����[j��ж<߼4O�0���E�� f��ˊ��J-�Jl�K�K]���E6�G-.�/)��VؖUڽ���\�35C5��_dj��x�����񯊩y��|ߘ���y�Wx���;�gLͦ���:�nY1c�����,45+��15�|�����k����O�/��ޣ[߽z�ԡ�=��7tMݷq���{7L��8q����|�������������� }�{���- �������^���W<M$�}Y�sٶ4��iJܹ,a�B��1=�T��S���Ee�ճ��v�Z;c���ya�E�M1e��yr�։�f�קj��Ӳ�tbِL���,�36{��ZK-�%�e����#�g8�-1��HKA�mB�=�f�7�tKIT�qYLI�(����)�A3$OkC���Ԣ�W�a���`�R�S��p(�ťŶ���9Ԣbi97�s1s�С��4 �o�k|����hxq���MMS����c��S�����%�)�uW:yS�]�X_��tr���,[R����.s6�q/-�^B�%��(�w��&8p�T�C��%����cR쬊9(R>�Cb�a	tD
@���{C��E��b�a���U����^�O��ʩ���~G�>gԉ���:q��������O��������?���ˣw?ں��n�ȸmj�~�ܧ��2���<��,�P�C8/B��y)~QN^RP���ŭ��2�rK|/C���p�e�����^����{��!kx�6>fH�]�y"�@\�^� �*��ޘ��
�w��%q[E�P`W��n�Y܏��p����8��@�X��@�e����|�f#���@���Z^�F��H�i�B�u*>��A'��@��(�1�xA3^��\#.V��R�O��:U��'VI1~���1���?|�#^1���7�� �1�cǍ9z�[��|c��o�z��o���W��B,������bQ@H0�K�
�D,�J ~�����W~��o�1j�o�/�����Z�5)9=!!�n�Y��1�ƽ�J�[?A~&D� nZ�%bX"AM�k��>Lc���&}�֜�ɞ�\�۰.~�ނMד�\t����~/}��	k.�y;��Y-�s��M�r���ミ�~�/���d�O;/�t�޻�k�9��6\.�v�r��ҭ�r֜Oj9��@����;��-�7k���+jꚨ����s)[���5{�&��h��Z�N�U�j��5Ԗ���� �"M���ٙ����{uuU��w������		 @pw��2�0�0�����ݳ��w�����b;{���N]��^oUw:!�Uu�{�G&��$���{��Lf���J�E�ݟ�Z5���0jU�^-�($B�X(�p8��bX^k��������t:�kT�p.`�=eq�o�60���
O؞ij�Մ��߂Ш�`BX9<�E�3#�<�S	᫟r�h���Wηq���B'���η� `v�O|T��X�9.6����᫟�ř6q���.E�d@d
3� F��0�(�#��b�Z*�(�Z�B�V����2�\j?�Ɨ���/�V��o-a|�xfQ^v}u����C���۷o�Νۺ׵6���e��$Ă'�Lz𲘦�:@I0�b�X ��P%8a	1�A�.`�EL����	a��W?���T7U�I7B�V^�S�k��+���*�1��L@������8��ۢ�'h���NVK8�ҽ��!��ڮ" w4����Yhg�&�F��E�jW���E�aW�yk���\�]��i�+L�Ֆ�jkO������)�v��zʜ�� WW��-�Ԕ�oH�֥�k�U����DeI�*3Z�kJ�+���F�����_���_~��O���-*/Ȩ,Ȭ��.NIL���M�x�*�(siE6b�p-�M±K�.7V�$��~�����*(FɊ�34�?�.ȱ���3��3�,����&j㑚8n]�m��UAu��&QQ��*vI�\?h�	=�b�PB��a!���a��/d�_�߲��K`�b9 E�&�Q�Ci����p1�C
�ȡ05�G��(d��G¥Ja@ƣ{�|�3�z�������q
��<
��A�����I_�N�t*yIFQ�C^䒖��e~y,Z/�N�&K�S%i�5�`7��R��)HM2�:	�J�V'��c��.N�)�`�S�B����E�C�(.�Χ��#q�h3�M�]1��S[g�?���l��s���7�Mh9�p �|"��l⺳�m��6���5]�s*�騥�7�n~� �=q���>�x�ƃ׫�f�{F�6_��t!��Lv�ɬ��m��'�ۏ�v�hܛX��Ȯ���l	r�S�6��r�I�hU�9��e�M��?/��Ɨ��b5vLր߮|;��l'�*�H�I���ژ8����}g�o<��qw���G�]<�v|�nf���\��K���k������g6ߺ�6w�ef�mf�nh���Ş�/M}��_�����z�����w���χ���<3�ue���L��+}o��{���{�w�~}�+�w޾�5<����cGێ\���G�N�>~��؁���k[6�o�^��VU^��Q��\�䬎3UD��<�6n��Wͭv�k�z���h�Ņ����n����X>`s��am�Qo���#�-��v��]&x�ڮamW�{E�>}7J��!������OsȃsR��B�i�=��g��Y���"�\�3_s�V��U	�W
?���V�~�U�Z���\�s�����.�!��>��gj>cr���&R�Ȁ�ej|]�qS��� �(<Y����������~H�E�����9��h��!�;D�%"�F�N�v$�N�u&�2�1M�\��ku�Gx�#z�)�IC�4/�W�m��*9�:�hP�m�m���������������
KnX�7��A:�"�y!���'i�Yw���1G���,L���	�	0	!�9w��d����A6�M� y�(_0!O��J�M��U{ũ�q�G����ǒ4��O=)��iw�tK��;Qҕ(ڔ*ܐ�48 �9����fa��|Ug�lc���m/��(��(�m-����LW���0zS�sC��#�֒ahH���(��k:��
u��]u�=u����
k���>K�����W�_��]j��Q��k�Gm��Sk���W�6�4y�����۲T�	����,���:{_�g{�����Sa�Zi�*U�V鶗k��*{��[�$�m���Ŋ���޲���*� 
�5 0�{j,��ŏ�k�֙q���/���Gx�����8}����ofj��pSsd}���0 ���Sx���{?��N;�5�Զ���sN���M͹]������[qno��=����O�8�[udG��K����S�������L͙�{�&?���>z���>���|���o�2{i��Ѿ����>45O�Ԍ~oj��L�����-SsnV��p��@�eO�yC��.�Ӑ. g�Z���Ƿ��j�)KPǫ	:�voȱm�Jj)��HPT�+֦�Z3��-[��6�}������5�{*m�U�kKilgQl[��.�V��4�St�x�75!�F92��-���.W�C|�qS�x;=aekp_b6
�|1G �WQ�j�����kM�r]�zc�|SSoc*Ԟ�P������fj �����4[r�>M�;�������z|���)3*�c���T�\�Uvͥ�a�*�i��B�GE�$��0���>;A�����=Nx���<�ԌDP'��$�8�1N�й�4�$󆩂c�9]��1z����.�a�����r��~;��_���ov����֘S�b����G#�sd�235W���H&`����q#��A�n��T�-r���f�o2xO45����{�>���ujpY���>��GL�<`���`�&�����1��5�(_���>��N���\:��<)���Bh���G��!����bz���(�ॅ�J��hղG�#��G��)� 8�- ��XY28a�)Q@�%�?Y�l���[���/<�z�+��/_�d11,�J
����ZB\��|���!𗃰8l���ՊU+�Vc�LV-�^�*2  *"�J��C�#^�)��	\�<p��+�p��L��K��	-�EB�35f�J+֩dv�*ƞ\�Vߗ�r$q���7�\5�L$�Ur�Պ�V�x��؛U�^�?������j�?]��?�����?�_|��'?h:���So�9�����.�Vu����W3vL�t��v�&oN���M\�ٰ����ݡ�\+5%˵.��"��b�X���V��r�P)�e"�T��J X�F*7�d���(*�U���טuj�V�����D|� ]hj��M,�l���`�0�9��4��rq���?�G���0SàP���!�C)a�lb�����U\��x�F�ƴ�S�!�55N�Ѕɚ�5\�F���|�[��8DL-L��Y0�=#��*nj6[�R>_.*��B�Va��5f��b�Z�:�I�������P�'߂&p<�8?�em������{`oߡ}{�����(/;;=<��^� g@���(�*���x� ��a�35"35T�*��:!l��񺇫���h��0�9�^�kj��f���z����`j��X�`���U�],��zovT�{*L����E��E��%ƍe��"`c�\�v�[:�m����gk��1�Z��+�S��Y6~�N4"-�c�L0��%�۵q|�����G��[��PZ����������v�.�¡�[�"�ы�:>G/�E\�v����b4�[�s�!��mP��&��(9IZ8Y��0q��?��-q!U���L� ��	��X��;NR/�����ęFn��i���P8r5=x%9x5)8��k���qM�CW�_�j��aD��	O55.�4���{+�.�2O�S���z������gdj�,2nj
8� ̲�����O��4^��gj
�e�F�K%�)�v���J�$�z��]ծ�5��VCi��n���h��Ӊ��&l<��l��	]��<��/�7x6z6Ł��DV�P^�Xr�Y��#����5���v�|�����}�
�O�G�s�6\H]w.��Lj��擉M'��[���Kn�[�c�m�'j��*K�BoW��n�6ѮN��fF�����͵����u���!S�35�<x��������h�[�z��i��Z����ȁ���K/��UNOU��TOOj�g����MN�ML���k���0:Yv�b��ؖ��>�����/���/��mWgZ�.4�_h�^wm���W��qÍ�uW�7\[7t����cG�9�|�p���G�?���辖������7�7嗥$�'�T�Z*<�r���..��e6����v�5vN���ש�6C�`�����o����{�;���q������e���]�9}���˧�B)غ'f�^Z�j�yyf]"W�5|�Ͻ�g��Y3(s�G�)`�*��Q��W
?�?���QH�R�J.��L���;��k�������������������4ֻ$�}���7M�BSv��}H������~A�� q>��S��D�>M�6K�*U�:S�G�
Cp���j^!3oGn)�I�)2{�]��n�/�����7G`MDІ����|�	�
�8yE�����u���ً���q}חe5���n�lc� b9�	*s�	M38�t����4���G���4��45�075�b	nj�5W����K��~��:5����#�g���+2��3���fs��[f�Vb�Zd�.�u��:���r�홦�t�T�iM�yM��.�R���I�ԥ�jS��xњ4պ<��B˺\mw�����w練�lO��1k�+�dK�5	G��nLٖ;қ3�#{dgNO�fW�}}�jS��-�X���,��,��q�l����S��0�TZz*�]��dM�zk����0MS"�-Qn-V�j~���������#<��n�>ڎ��kj��,45�7%,45���35��9����}z_�������â/>����;@}��g����?���/�{��ݹ���G����o8�zv��25C�J�ず����s�M��h��v����M{��!m�WV';��{���(\W��j��O�I�Ni�S�n�$�J��3��5I�U�[��v�%��M>Ԝr�)��.ng���ܳ�&eg}VOUfkv|�ǒaT%iq�"L)��EF��(\�H`��⑙GLq�UQ�k`D��,D̆%������)LJ�p�8�:n�Sؘ$�H�����I�����'h�DY����� L|�Gp�.ݽ�r��p�75���ޢj\րq��@��G|�.�ʦL�q	r�J<z$4��|�F9�düD8���hm��x"D��$�vǢ裑��H�8�2AfL0�L������T�oB�4�\����������o�����������?����y��'oT5\4{�C�A�d��	�̑��Dx6�u����\&���ע0�G�oF`��u�Հs�:�k�'��WY�kl��:5xR�}D��/�M͇B�{��]����>��6���35�x+�����̏75�0��FE� 
�(t��:ɥ��h�`�i�}��<ćKx���9o���QLoQ��M�Bj�j�ߑ�	q55�"r���+G��,#�(	a��x������.._�|�ʥ/�X��ٲ��B�"�BA�aa!�Q�0"1�L���	a°%::>5���A/,�rE`�2l�:((�F�
��Z�j��ŋW�X>K��~\B�sӲH�/�;E<��-yM�B'�hd���L��[�3w��䎣y�&�^�9t���k5'oW�Z��z��[��n7|i��W{���ͼv����>����?�|�����r�W��N���fm=���d����dl<��5��y1��B��IM{����k�iR�5�t�!V���"5"���R�B��Ƚ����	pSc�H�҇��"�Z�2�Bf�֑��%�I��)$J�P*��� &�I�n���p����p����x���ej�����c�L*�gj�D�3L�W�E��!;J��\j�ҝ� 7$p�W��_�����n��#*pKs��� Z�҃�P.��X2�1y,�d�Q�}����%J�B����z��h2b˝ 6��~_��N��$��$ƺq_S���޼v�������{x���;�������HON �W+�b�D�H�(�H%Xw�[ ;.@$|����
X�I�3(bCŇ�R^�����eYf~���i���\p���L^��>Y�(�5~�_45���}eZoC���c��Ub�P�k��4�h�s��y��\}c��5�ҜmY�i�O7֥ �`�a�˲T��
�T�vq���VCN�.g����dgYNBIN|myfCMAMUnuu~IIFiQfyqVQvjNr\Ajb������NiRJ��F�Ӊ��*9�&8T�h�Щ@mR�$d�L�$���\��Ou�(q*z���m�ع�n^e,�:�����s�$"���im�P+.w��p������H)����"*�?2pux` ��Y�,p�0�[�r |���U�� Rp5,��55�`.1&� �0>-BȈ1	bQΥ�(`�9�GWy3ᙗg��Fi 5����e(��H��ȼ^��:5<&75Z>�.�⫟
���O65X��{S��T&@Uq�r���)u�e1�B�*ݪ��c��es'�d�ɨ\�R�W��챮�gn=�X&z�9��s��S���֓�����3�����dk����O�ZOۚOz�OƮ;��j=���-���>�v��i�Cq���o8���<=�����5���=�j8�h8b_8�\{����Y�m�m�&�h=Y:G���7X<NC�K���fx4؅���c{V��y�4nj��%��Ip)�=��5������\г�too����3'��������''�����*�Gk�'�&��F'�G����<}��'_}y��؞�W�_��>1�6=�45P?~n��@ە��k�Wƚg��-ロ��M��՝8Vs�P������=��i��C}-�65nhn�hl��(�Jɉu�{l�m�CUjW�:$�vA��Wn�+��*��Ϊ������Hk����_��op#=�f����������D{l�>#ܧ���X;e��B�6���G�;�}�������a6m��"/��;bpSȹ�g���)鶀��z �L��
��2��2��e�_I��K~!��/�A����r���/ؼ� �3�R5��O35�(nj>�%>M����GpY�!����N�}LBߥ��a��d�^f��Bͯ�ڗX���»\��\�e&�&�~��pg���4�Sx�%�Eܠ�����$��`�5H|]��	?N�XV��G揟����^Z�'�e_d��s�Ϣ�q2Dfh�T�$�3�d�kx_����Ƈ/P�k�g�p[�~�Kf�9��W��(|&N}$A�/I��fj��z�c�ƇO��4��\eO�a{�uG�s[�}s��#�ВahN7V�*�<�b��Э)�5�ę�cM�}�K��eX��m?NAI׳��h�[Д�^����A��_���Z0؝7����漋������ܙ���ά}�b��skv�����2o���f�3mpe��:U��µ�>�wm¶����j�7X��)g^�"ew�|k�|{�bG�rg�f��|�{��uj������䉦fO�鉲Ƨfቦ�P��p;�Yhj�.8�������j�(��4�#{?��M͙}=��o;��������>���O?|�_��/���_|���o߿;7q��������;P��L͈���uj����ڟ�:5�L��\�-��E��,q[��%��۔޿���1�&3�.e���<�����!	é��%[���q��Ƽ��䮊Ğ��޺�k���M�Y�S��X��2i{mVWEzcfL�۔nR%�n�4Z!�ʄ&1�Bj�%G�RS��"��&������v��)p/�y"p)�`�ِ�ł)$NT7"���F���:�"Z؜ �Hv$�Z=��XfK<�qk�5�R���d�k >5��5��m�R������)�d;"��U�
�5��4������ڳ.�zF�>�"� ��!��#�ǩ�0<.]I/�td��yD�,d�Ȝ"����$�W�PqS3EeaV�śb��t�8�?B\��GĖak��?N�����_~;?��������?�������ߜ8s�r��}�!�	"�C��Y"35Q�+dx��,�5�����MV��̽N�]c ��ej�21Y�Wּa��w`	*yW ������$|�#x���:_����n?np >S�~���rF��ac������ޘ!(t�C?Ţ��,�����R�1��Z�Ko3ڄ�f1�Q�-��+S#�UI�J��G�����؋wN�Q��P�M�Mt�<"��ڟ�li��2<r��jE�� p���^�[�t����!a��(
�@#��+����
YI�ht�ٹ9%eJ�9�DY�x��~+��K���V�G-Y�|E�R��%+�V/�[�t�_HH����{���,&�k�h���:E<���R�Y,Ӌ�Z�A��'�VT���t$�m��Mgnm��u��C7>�=u������< c���}S��}��+7x�A��ф�N����+E����ZIj� ��+ĕK��u��漍1���ҭq����'TmI��)۠M(683��X��&��B�P$�HDr�H)��|�L��
R1nj�R��,Ĭ���5f5�k����\���l\.��f3�ujpM6���=� ������O�<q�=���g�����'*��lSH ��K	��P<Z$�"�v
��J����-4�S�dj�'dj�<H�-�zd���T��-��([	�|�Ke 6`&�r-�b�Z�26�-::��v��n���ؽ�� |�njRbqY���LM�35�wl���ڿg��OiI�.�E���P�s�(	�B /����D� �$%��S�b t*B#	Y4�6��n%7Ig���VI�U�eF�L`zZ��WQo�Ԓ*���25;K}e��r����
��̖"�foa��,]]��*YV���LQW$���U)��$}I�\ J�e)��T[q�� ޘ�R'Y�n=?Z��t�G/�Ov֗f6�T�f�&�f���'��d��&WV�4֬�)�.�[SQ\���2�]N��l�k����N��m��Y�6�ܩ�J�M.0�y:>G��l���'��(�rz��i�U�43��*v`�+=�����֦Heu�XQ�GP�B˜H���qb���!��"�%x�[���%���	]���4��=9(����D�A���L[�i�(�P�<��� �=�c�nj���	aQll5��j�����6i�S�SS�*�jКd�TMe��.��J�V�9V^�Ve84	V�]g�Y=6w�-�ĒVg�mq�l�W��04�0��2���4�7������=�h>#�;�,�C+�ū:�l:�ᢽ����e�g�ɘ��b7���x��½҃7;-'\��7]9O�O{֜qԟ��1T�V��V�jv[j�L����kT��O�֙���M��hc�[�k��h2�e��ɳ�-k�LM���<jj�x�F౉�nuNUv�����u���ӷw��ٙz�Xҹ����r�r
��JFF�FF�F�+�F������\n����0X{���ᡆS'Z/�����4�85\?1�83�ver���K-ӣ-�íí#�M��g�Ԝ<V}�P������ݿ��G��M͛�Z;�K�3��c�ynk�I�o�[e�I�ST�@*�p��Smc��X�X^��5Z��D׻Ѝ.�&7�مtG�[]�^'�����uP���KJ�)�l�EuC�[9�ۙ�i!�)!G����I.��$@�
�����J/Kx7�9m�CzY�zS�} C?R�>WJ��K���&�R$��P�s��g|�w(�[���|����X �OY�X��������W����W~���	�2��Yhj ���Я��G��{D���[L�+,�]�r܏rhY�ѕQgBHCQ�Y�����.3�9:r��\��o�D/��/11Ys�)�Õ��n!�;"�M�r�+���X�f�����-�ߖ��e���R
o)-���YH4J�h#����&V��qM3Ά�4S\�lS3�CpS3%���V1����t��Q���K����<�tѺ�'������Sl�S��R��5t;��{z�c;��I�b�"^��(�)��!�9�|��I�vH 3��aE��n�GD���+�kRUtn�d_�Ů��#�
g��^?�|�hӕ�uwη��烫=�Mt�*�W����ڙ'��AZ^���i�U�)7Uyv6��hL�Z�Ua�,5m���ڮBՖ��B��b����RͶ"ն���^�s������'k O���5-�5��y����?�a	<V��<�ԴF�fa�\���������;���Z�Ssv�V����?��|���8���W�}���������^��xrǱ��guk�ph��25x�'���*
��}vE���M͙-��]Iw�oq��1�u�|ES�jK]�����U)E�F��'����WB� .)P'b)x$�*�rWf��R��[�������I�I�V���&ys��#�V��[�ei�v֦9�c�VU�^��Sz��)��B�"���R�4��M�O��F y�e��}���Ha��IG�4!������`z�*3��#'�Y&�Ɖ�u!-.n����a6�2 �q������d�BY�����9��9���Y��M��P��@�7_��P�����U����e�O9�GU�1��|�u�L<G��c3'$�f�m��R=�/�W��qc2��L�3$�,� �i"k�H�"R�(؉��7�g9�Y�`�"�B'���\͘5�M������?�n�?��_������/�����^�h�Ŝ��(��P�p0}�ȝ#��Q�Kd���O���� �E<45WI�U
�
;�]e�ן��y��yW `K��ʏD���r��<ɻ܇���a��wY|l��g{'L�׼M�I������ ��L
�I� 0#F��s�$�r�C?��O��'���2�)���Z�[�뒲:�4��Y(kj�*)�G�������MM���$�,+����@��+W����H��*��+�b�iV,_I%ӈDrDDTPp���A�W.Y��ŕ���>�88x���c��ʚ��b��"�OW��ɪUKBB^
ZJ�G�C�̀p�ʐp���EK�,znыK^x������@
Zɉ�BL���N��v1�2r�U&6I$z�� ��&�#%�����+�|cJMw��9g��'�vE�R�Iͺ�f��N�T�;s�Mi���D��JDMD�FE��T���O "�+h���:��$�$��N�ZsԮsR�1�HbL��b�LaI5B��/����2�_���,���&� �r���F�ج�Z�2�à��b�L��	EB>��z�2l_q_\�|ojpM��4Sv�����?L����?�1��4x��4��&,48<8 <ȟ��M
CD����Z��Na�β`���lSS��>�gdjpSS#�s)�-��,d�`er`�(��cq�{>x��#�H ��dZ��b��c<	I�����qX7�h��nqZM�(|�ĺ�������8޷;#%qm]���=��ٻ�wkצ������iө�"�q�`����W ��P��aXȃ����g�y4
L#�L�f��K%j�Y&a�]�kdYxY&(��yZ��-��{?5%����{���[l�Uj�]a�Si�Yn�ZbޜoX��oJW�&�K=X7�\�0�%d�����,��������E���4Wa�3?ٞoJtj��ۢL�֧�Z��;[k�z:vt��o�iZ[��PRSW\^��fM庶5m���k��ZZk��b<)qq��h��d3fC�ݚmO�v��z�A�W�52�Rl��uBX�Bj$�S�DL��!RZ������4�t=#��,�f���Unfm,�!^�,nH���	k<h��W���%(���XG�%��R����V.]�dI��� 0	Y�,��/|Ŋ( 1 �H	������������Y�R j>U)�JQҏG��T(M�Pe<��������pS��Q-v�ɰbUf�fj�SE���~����Tİ|���#�w�3��D�%���/0%��Rj�٭֒-��=��=��}����CҪ��� q�m�9]��������|?�ⰲ���kҽi��rR��a�Qc�1[���ީ�w[G?�9�FƮY�j��	ݣ��C��S��s�5gl�'��G�U����>eE��|���C�V+�/P�34�L��hu;	nMj�6=F��e8X�'�[�Sc�ɚL����ϰ�IV���w����i�Y�Z6�&m�Lܳ+�̉ԋ�2�.fd\ȼx>�����GǪ�&�F�*�Ƨ�]��>wu��X��h����ѡ��������N�΍W�m�l�m�<�qej��D��h��H��X��D��X��p��s5gNT?\wt���{����Ի�eKG���k�J����1��$�$)�HqSS����2+��ά�1km,��`����v'�.�6E�8���ׁ{m��F�n5{���KL��'m�F��B[i��䠽����Q�q��}YĿ�@��y���7��We�	���u��"d�!���O��5��?�IqS�+��K������g<�[��}�����36���>��O������Ê¾X�O�,7���E_��_���oo��/��7y�7��ټ㷕?+�� 5��F.�� �r�'��_c
��D�9җ9�W8�;,�t8\3_ef��8�r��c���a�s|�eS�m[���O���,�.���Xw��Q�!"}��g�'X�Q&s��Z�ip;�÷�	�4�0��dj�~�S�fu�i�bܮt�OǪ�{������YxL��t���>S����<EW��3_Ӗ�i�2���e��+�lYV�CLSQ�jN�?#d=t554�D	@���d��DD#B��Rb�������C%��_9�<��v�;�dG�ho�����ty���w~r{�������o_�~�j��@����\y	R!s%#bI��EP�O����TMw}Ү洭��]�-e��E��=�����=��mE�Ś�eX�)��|����~��L����O�<��<��j���9���74��c1G�p���v�w�8����<nj��~f���i�O����O?�������_~���'��>��e�Ȇ��mG���>X<p�4�����o�����=�#{2.�H��#��ƄM��MgM|KIL�M$�т�Q���#EljT�R\mp�F9R�]����$e[k�������MU�%���1m��5���D58u�X�~�Q��&h�1*�K!��P�I�E�N��M��G����[B������xS� ���ʆ�b� J'��$pь2hlb-,���I�*V�KHKU0r�����\kg5��k=���#���#��qe���k|�͙��9��ى/�*TpS�gj|�f_��H���MxL��C��I�hT��Ȱ����I��徟����2��f9�k��ǘ�9
�P֐sT�%&�*Ļ��"�+��]8C�ó\�)�|ܒ��cۯ'��r��������?��������n������.k�P{�RD#d�p(4̜%��Yg*�5G���8Sd,Y�0V�ɚ(��52�
���]b!WX�u�35O[���P��H���|,V}F��#��CTΩ���V?[�>G�-0��#?��Cl��5s���i�`V*�SJ�h�)��"�u�A9Ǧ��9�wF���O���Ԣ~%�Mm�2}�����h�����<"h|<����I�RV���1�4�"2\D[���G�d���� K�,�Z@��y�%��\n�i�6g5���@XI&�s��-���n�悵kS��P�aID֥�����4,2�H!�"��� "yI@�%�_�[��O��{!*Џ�/!�Y��x'�m�U��0S#4I�F��(U�������ʖ��ݕk��T�O(j�'W ���&�*Y.Z"}1P��E~�E��~������[���EK#�`�����9�OV-X�ӕ��\�ӐE/D.z���c��� v0AI��`Ւ�R:$gBR6$��"l�$�:8����5��N����ɾ752�E��2�RbVIqSc��+H,	�B�� ^ZЛ	��W-�L��
l�����25�E��L����(�3LMDHpx�ꈀU���R��K2��qA�]��~��Y&6�3)�C�����<9S�ש)��
=2�Ԙ�1
�"��l���RO35:���t�%ħe�ggg'&�%ƺc]������&!ƕ���:Ź���I5�۶l޷{����z�vm\W]^�����D�*� A�l!����� ���Y	�  �80�̥�Y1�(���Ԕ;������ҍ7~��~�oj�v��wW��VF�,wvZ7d[ҵձ�b�(ۊ��d�j⧘E�I�U�lW�Ek�b���6pIP�[�W��T�����g��6Ź�iI����M-����N�?{�졃��uww�m��o���+kl�lYSݱ�~K{뺆������x�3�f2[F�������%�bv�.�ΡUZU2�j��BT���X,!��'F��br��aT�4--�L/�����hz��^é�Ek��u��R��T���Ѽ:��6VV�ȷ��|5��#��BV�Ė;-[��5��	]�<|�
��ո�!QCB~��y��'����y��� G�2�x�����s�<�f��L!��BL� ��Q�!���D�5/�"�w��aj��OX��A��s�=�r���-v��.q�S���%:lq�xO|�;�ܙ�Ɯݢ�Y��۬*���쑖�K��c�RTU՝4�\�6^P֟�Ԝ (/�7Lzzfݛ������'lm���Ǵ��⺆+O��1�q�����_I�J�c��q��q����5g�u'4Շ����ݲ�^yI�,�U�Z-��W�ҵ�D�ɣ7X�6m�S��Ѧy�.Y�S��D�x\hj����n�;=��܄Ԇ��M	��v��ޟu�l��@��p.`x0g�b��ł��������3-ӗZg.�L�5�O�[s�b��P��smS��#Ϭ�6W76X39�<3�:3�69�66�::�6:�:=h��nU{���SG�Olܷ��oVLx]SӚ�����<�5�(�3K}�Ɨ����j��zo�f�����6���wr78�������nG�,�3�G��S0wI�}"jJ��Fnc��R�v���S��q(s|���L�:�{S����$�7d�+���%d���B�I���ҟ�տ�k�Z�R�oD��ſ�~���kj��F�%��xSs���M����'e�]`�C��#�[�6��2��]�诉]�V���}?_�����߬iy=#�V���<&�_��n@��,������y�-}��}��|U������9N=K��
�n���� ���2�%�����@7�ƨ��9JcN09c,�#�75���P�<��B\���Tި{J&�Q��Բ��gj�Ū�ū�ujq4?�&�H*x��gj�
��
�����ּ�k�Cn�SP�j!%�n􈁫	���92 0bU �?�G��فhh�(r�$r���0
̬K�^{�@�̞җϴ���`z���|xc��w�}�������y�뽻�����nL�ؔP�cT��F%����-b-r�ɵ��ΚĞ�ĮJOw�����Uh�*�wa]��[ԽE��:0�Z���=�	>�Ya�-3�(7.45`�{�ə���xY�DS�7�>�}�'�Ԁ݃�v���+Z�4>��4M�̿7Sslg�񾵧���ݷ��-�l;{�������L�'����}��_|�!6~��W����ݽ>z���=-�7o>��L��������)ؗ{�?�������]�zSF�������n-6�dj�c�:$��jQزE��e�� .9*<`�&A�1�eVgƷT�V�l��kȏ/�7�8e���|�+"h��(�N1�&�r�.)�%��D7�\#6� �����#F���ą�_��߁�����,��B��i��QI��0jX32��ZJ��B�冥���d�Z}m4��EY��d.h|�Y�4|\�l��ZMO��gjv��
0Y��H�_�~d�Ӿt��x�Q����Z��i'�!.{Z&�03��o�J?��~��,��r����ij�(�%*�5��6�:��
o����\�%�p�$
���LG	�	K�w���(fj~�����������q�˟�_{�Ͻ[�:�t_���)��0�h��LF��)\�G8����������u���'*�j.q�+�i��מRQ�}��1�i>��?��?�j>�>*?����ϯxO�X�fA��G��A60��L�������k��Z�e�t�aR�sC|�� ���N+DGU�~%ګ��(�'�9�RB~���<"h|�xM� 759!OD�rb9T#%J�
����X�r�ʥK�._�<   <<2*�E�B*d�*O	�B�P ��Og��
�B�Rk`�ѐ�Rڱ�y�N0�s�J�r2�����Q�%������xq�"�KBB��_�h�O-}����\�|��Rz�r)!��c%�n>k΢�Y|��o��M"�Y"7˴JT������E�����蹀�,_�B���H]�u�s�E/����$s��@��#�����%/�-�x�/�'�V-z�o�O�=�^aѢ@��c�s�/.�z~qؒ�+��WE�X�ҟ�@
%F(t:�fjd�V�ꤨA*4IpS�9��1KE&�<���
�O֘�R�J�U��
1֫[,�DX���||he�OրG:���6`O>����l����k�g����ఠ�a��!�lR�&%��75Vn���k�<�Ԕ��'�LM~4����w�o��"���t���0`&�p���Y\0"0*@��L��Ym�ظ���̜�����8���:,F�N.k\ފ¾:5>S湙i��k��ܾk{O熎���Ue�Yi�)��9f�F" ' ���'� |v ��ri 
�a��I"y4�b��G'i�L� �"�2#x����Lnj|���X����)��p�t�,sm)�ud�צh��l����*X1JN��ա�zA�M��ˌ5�$9�S=��i�y��	��	Y��)��Gj��(?����g}����&ν�ڵ��'FGO�:spg_��������ֵ:�ۛ�j++J�sc�.��j6Z����tY�v��m�D�N�ΦQ��r�L��"�A�L&J"	H9BJ�q"Br�����e�i6j��Rj'UF����rT����𫣹f��Q��Թ�Z��.^S�hʏ1�uR�f���!�V����._�t)��#>MC	��zx(D���<RJ	��D�13R�q�r�Pp�J�#*��I�F�#�
@�b�F���O�G�#CHj>]�be����1�n�\
a���!���(d�_�4����.E���K7nj�F�fE���-r!yA�M�j��ۭN���I�'����5���6i�Q�fe�nu�m�!u�!M�a]�	���K�EM�E�	m�yG�Dܖ+��Wc:g�v^r�?gl>nm?mh:��?�e���[ͣ�O~�0p?w���S�}�i�f:GR6N$�w�Z֞��QT�V�V쐕n����k�	�jO�ޙ�7��٬����\�$�2�%͈�D��H���25X�Ɨ�qr�hj\���Oe~Һ�䭝��v�=�5p.{l�`r�pj�hb�h|�t|�||�rt�zt�qj��򕖩�5C��f.��}m��l��h��Ů[��.MU_�p�r��p��P��h��D��D��X��H��H��x��t��,�qr�~�B���k�o;{������-[�7�_Ӽ���4� ٓb��YUVy�UVb/�S��!X��Yk�b�h�iw���z;�����=V����e���=N���'��Rw�ɻ�Q;X�̰m�������a�����F�F��T�@*~G"x[�]�{Y̽%���_��pޓ�_�e�2��`1�A���R�;��wb�oE�_D�D��fj����ej�&S���I�A����Bp}�]1~�i���{���H�}+ޠ��׹�	��&���M�.���3�'/�_����~�������.�_z�-��\��3���◘���M�p� ���T�I��a2�Ӹ�kX� ��*�Y�?�u<"�f؊K��
,�c	&(֥���dA�L��>�d?[���43<��L� ��ퟰR5R�\���y4g�5ǒ4R�o�f]
�q: ����4�e`͡pS��@�Uh�X��$�5/�"I�l@IH��,"�Ō��F�Q"#�u�@�FR)���@3�H��,�a���r�_�������|���3���o�hv���7];���oLm}�F�[����wk��v_����J�ԑR�oVJHb4���Z�(l1&k�rښl[wMJOuBW���ı������ʚ<��5�W<nj�5x��gj�.���)�����ˠ�hj�8q)��j|�����6��ο4>�NO����k�����L�M��;����GL�g���{o���w_�:|xW�Ѿ��#�;FN�>-S3�$Ssq/�i�WL �晞����c�
�����K�T�ȰC�fXG�C��CW�"�W�-���@4�B)���I��՗f�f�g��1:�%��(�쐲 V��'�p53��%�Dl�V��(1T���H/��
8j��D�>"��w%�.��&&�����.��0��/�a:�E�����?]61��R@��lfG)+�����
�>�^M^㦮���j|��5��yD�����}_�f��lMW�oՓ-ݚ#۞���W��W�*P�.��-��j�u��y��Lűtͩ8�	�ࠐ�maH�c5~]��aN�GyY�弓���y]����T�i�f"����<�5�u.|E_�nK�7��k0fjfI �b>���?�������Ͽ�����������?�i��o����?<�nYӴ"z�&���'"�c��9<K����3Nbbm���i����@]�v��+�\���X��
���>�Լ
a]���ނ�o�$�2�>����5�x5��2��L�|�W����}��}qS�+Rs�����\���.05�\�8����s��y3�%��N�� �������������.�Dd�Sr�Q�`��S�`_���eP+�U��8e���A��S�O���L^d���&`��$-9L�����^��o�K���GQ��H(P���V�VmB�3�0��6��9��#�}}�ƍ�[�ʶ��toiػg�����^=z�j׹��{v��T#7�ddX��>L*'��a�ȏ�XN�ј+"���n���_X�r�OCV�HX*&�:�X	l�3m�����2�U�7���*SK ~���.���/Z�㧫a}��-Z��OC�.�,�c V�#�#1�ݱ	�F����Cၼ��2���~/,X�,�/.	��O��.{���`�tIȢE+������ �OX��W�$�(��#)�� z)�(�%�Rm�)��"�U&��fJ�F	���&�Ф�Ubl�
35z�H#��$R�X"�B	����[z0�ވ.P|���da��Y�>Ml��M`��� ��`�_�Q�KӨL*�A!��$��7M �h��z%1؟C
��d��� s@��he8$�Na���id��MMa�þQeM��w@��!���-͍���$n%V�QXD
�D�2XX����L�C\���$*��l�yb�RRӳ������t8,f�Ao�� 6��n6�D;�ܮ�����@JB|blL���v�c]�Ue�۶t�tnnj��,-)��KONJKJL��ב�0��㰽?K��_��ఱ����ǠAT2�D��d!���1b4h�M7	�L�L/˄��<+7��.�|oj��b���.q�J���h���k�4&���%�)R@k��-]ў������o��n���?05=���%־J�jώrWW��5�P��ɵ���p�����e�q��.�(5ژc�Ir��e&f$��e��$y�I���8wb�+)ޝ��RS]���iǖu�wu]�x��wn�]�2~�������#{{wt�����ѳ���������4'7%>�㊱[�3��sźm���0�z�M�3���L+k�"�H(�`��I(� �FJ�:��Q�t�Ԙ�Vz��\b#�;ȕNz��Y��u4���(��*���J'R�X�a�I�f9UV)GĈ�D��WE�\��z��.]�&~�HA r0§�c���Pzx D���y� �$���abf��!�D��!��K,�1��S�P�'�������`u��
���Lri�.,�E�J�K�M1�r��
�2FP'�M��'I֤�֦J���ɂ�$~m"�&��� ��X9��ԃ��϶�S-�D�*�n��\kJ�6�N��,�ޤ*��U��U��3�7֝0֞��9�j�]7��iLM�;g��V�~��ײw]�<~'n�Y}�^�} s��=S]s�9������J]��1��7H���n�k��l:e�?���WW�i*z5e���vmz�.���e�N�X�f��b��̲x�2ũ�pJ�`�KP�����X!�_ej��|'֥�aEao�����;3�]�����f�v��[5t>��ٜс©���񲙉��٩���5����j�Ǜ�g�GG�^}���x�_�e�����݁o�����ڑ��S�'�4ό�]�Zwyfå���S�&6NMn��j��0�6;����s��N6�9��챍�mط��{]s[}��Ҝ�8{�ZP�Дؔ�6i�UTf���
��WZ��V���`�4�xMv�Վb8�v��i��X��f�'7����
5���#�쁉}����]���Ġ��)�uW.~O��Ġ�H��@�x��)�����[|�m�ye��g�'F���c1��n����*����{e�o��_�?G�����0o�������i�L	35d���75�  \4��M�;�3T�&]r�ĿiF ��1�u}�s������O]�����[�s���s5�3��\b�gh�
�
�A`P�����F�����l$�Wy%�����=�о����kƸ9����6�Ά1�8�i:2N�&(��b�F��}�	�3�	&0��a��BM����`�I�f��55,�"�3q�a�8� J&����i�3&ŔC=��\�מL�J��L��>-S���%�#Eؑ.^(h��^��Q���Y��9��<MW����Ғco+�_���r*�!�F)a.�D	�����%���B"��4v�@�X�:b�r�J44P 
]� &gi��[K��T�z������/�zm����+�Zޚ����������}߽w�W�ݘ�ڻ-��=#/]/�� �p-����]_�ĕ�q�M���u���;�<��N�w��䪻sT=yʭ��-��"�vo��aj�C�Ya�Ui�U�|�6��X��Z1����B�lj���8�Fnsiw������Y���\��L�H�����U{bw#nj�����`�������0A�}������w^��ׯO�;ڿ������6^<�2z�m�d��Ɇ�u��k'��`��CUc�+�����؛>�'mpw��������]���IOd��9�5�'k�9�{�;�lSsj��tg��m��;3Gv��)��_��q�<j��O1	r$D�s�lp}�"a��s
70�z�ۨ�
�Z��X��S"hA+���A~P�j�"��)r��%�C��(��s���rUȢH�X5G.�ΦSX42�A!�HQ`��@*�Fa��L2�A"�jT-2|�0)%
"1��B�4��1��שy���<b��}ͺk���Cuf�;s$]���\YO��7_��@�3_՛�ؙ�ܕ��[��W�;Pb8Xj<Vb9��>���BG����V������%����aA��iw�k2�%��*$���f�X���(2V-8�&��4�6Ka\��}\eB� �>rM�\��QtF�Y�i*o��a�Ӥ���3
�-��05�>xo�O����?��������z���>��A�z�)�������J�b%�I�)"}�Ș!��\"��t8i&�<E�Bb\��o2�7ټ�8�m0�00G�A�@���Q�����MDr�/{W�|_��X��T��k?i>�?��>k?j>�?CU���r���D+������
��2��^���|�͞a1�X�i��xC4�y
���c��Լ�U�$��
n��ץ�+R���{a�@�ȠJ8����K�k�{�v9�Y�\'�7�h���A���	�����^�`��P��b/�/��#KE���(��$�R3]@�@N��gDHT ���o1f*mzS�ǝ���\_ڵ�d����6�;�u|���\��k{�^�57�}fz�����ɮ��mW��}��o�z������������i�gݺ�����ކ�gz��wl�f��3��"�t��"l�bb�2.%X��uR�YY�\���	m(j��zQp�+lU��痼����/�-�|����Z�4p��AˣBV��^}~Ѫ���Д����Y^Z�P_ۖ��\�$$$���귒�%�{��lY���+/�{��eK���[�jeȊ�aK^|n��E��/Y�b��_|q	�|+�-����R� �w*����\r4NŏU�N1'Z�s����!�Yʵ��5I��3f���� LJ�A.�Ʌ�Q'�hR�F.Qz[w�.Ą8��bӘ,*��'��m!ޖv _A�ǀx0�q�,xe����>Ĥ�d6�Ģ�d�I�
'G��#"��Q!!��&"($"(,*�$�E�C#H�!�� po�
Aɑz��&�I&4���[X��	`7$�|;#�N+p��NFQ4�`	\��m��)�f�8�������hq�K�a���P��r�<�C!2)���Ax\����|�X,���j�No4�`�T�R�L�u�����l�Z��+991%%)6��p:�wtB�'=9� '�������������07'+-���2!��,�� �T��o�4�t�*E3h:��	�F¾Nj¢HQ�V̍V!�a�E�f�g�\3\`�晙fF��	(��0Y�]MV��V�x��*�W��%�DkS$��Ҧ4�9]ޒ�h�R�g�;r4�r���4[�f���9�l�|{�eg�}W�cG�m[�魴� ��'l-3u��ǧipz��X��*[o�sGmlOULk��2Q�j�%q:�S���<��o�(<&]�Y��0��m�μ���Ԣ̔씸ܴ����I�0k�e]uIAn�����}�oݼr��o]�zefl|prj��#{�w�޳c�ޝ��z�:74�W偟KJB���Mv��ewD��N�� ��a2Yt:-�
�<D
��t:�DD�p�!��k�(�����y�
���Fb��\j%Y�E6�7�D/����r�,��E�I��Lmk��*A��&�8A���s�C�ȰH�����$b����ȕK��+ �Е԰U����(fT D�s��aZ �B��|V@̍x"���<"@�����C��	%Aib�*�Q B����H;\
E��d��f��c��t�0φ�:��XqC��)MӜ�iJW7�)�w�>IT�(�MDk��x^U(sAe.�8�W����.E�K�y�)���
Mn��p��|��ᐱ崹匩����������b���䮩��ٴ��ض�;gc��7�x��ob�����'��|����!wG��}oή�k�^]?vw����ޫ?}�e��-�?�84U�j��ټ�É�'���[kvY*�;*{�]�����5�)%vW��mԘ�J�[�L4)�l�L�2�&ɳ

l�Zb�q��b!> �7��'7��M�q,l�����-�%�P�Z^��Q�u]�ޭ�#��Μ�<_8>\>;Y}e��ڥ��s`R}y���솗�\��85]34�82>���<���?�p��p��7��G�F�Z�z4c.�t޼�u�ڦ�7^��u�ʖ��7\�03�nb�}�B����s��O]�`�c���mj��hh�/�Ȋ͎֤�X��*)�Hʬ�r���"�2��H��7�֘���ɂ4[��b㯵s[��F���2��5p���O�2w�0�d���/d0�i��Q}Q����e��TK?�����qX�+�o(į�/I�[�M�uf��2_�����5�_�u�3~o��^����w�o��_ſ�j�ox����	q�bC_�8���O����,�ԼGc�Kg>��ޡ0���t�$�;�y���=�]�!M�z�-�����&zPi�}���/�?�����4��?���_.�|}��u-o�%�!�{� M��$�&]x�&��LF���SAG���_�+�ϟ��c�~�s�������]�4�3���_6L�̰s,�0�}!�6D匱�Q<F�Ӽ,�5���|�Lr�)�?��O!���qo��aB`��iLt�0�"ӨpN(��R\ө�[�W]��8�H��L��H�~W�b[��;Y�%I�9Q�)A�9^�1A�!I�)�$�=�ߖ��9 ?��>E��&nK�105�>ݘ��9M�)E�>Eܑ,iO�w�k�e�;rl�E	[
�bE<R��D�����ÃVG��C��=*�	�z�1	Djx1(8�ߟ�
��5�HΊEVV`�뭜�]��ؖ�O�y�D�K�_����@��Ӎw.��{��۷��������[��m)ݲ&�8ɤ����@z�ʐ�/���V/�{n-|UN�mCC����������m=%��<UG2oK���\��X�]��)gg��2��rp�����+�	� �x��^��-�p_��35{k��u�}����k��ֽk�@_�iw�L�5�4;����{�vĀw4�p���$��Z�x���,t7�p�3�i���}%���� gvW���]uz�S{�O����_z_���[��=wp��25g��9{��q55�y?�]�������������׮O�;ѿ�Ծ��#���h=�8~b������5�G�����O�(���О4���e�#����|�O�,�G��Nϙ��ӝ���n�ٙ;���`kbm��"Q�j��R��C����� $���,���(�(9��h��$��|�#8Σ�����`VDL�S��4"@@%�Q� ��4�P��Z� ̒s����(�ia�[\�0�$:�@%F⻏á��T�_�e��'l2�CC�Bb����rLH�G�lS������M�`s��3[֕#ߒ���Sn+P�(� v�c��kw��������E�)�}n�>︎7j���6?HO�8/���ws���˾�����vM���H�q�WX�+��9M��d�)��{�ϻ��] �2��$;�L�s�n V_Ժ��������>���/��O���������������ߜ<�NU��2L����*�w�_�B�(�2w4�����:�}��!|�M.k|�7���x�7P��<(�*?�?�h?�� ��������`	�CX�,~�+|���i�[�M��{�͙e2��	}�ŞaB��*m ����a�`L�_R�_�I_�7��e1oT�>�g��r��F<l����C�^�U��(a4�hk��)�^ƨ�a��5R�Z�dS(=45�b����5MM���/�&�#�p��G0r	Jv��G3�Ѽ✖-�w�<�w����3��N�}��so���εwo|���o�~��[��o�u��{���u�Ʀ�W�/��{����w�Ov�����_�r�f��L��X��x��d��L�š�m;����u�T�����C�H��Ġ p�"���2B��R����6>#x�;�������#�!BP�ߋ˼�f�O�[���.]�j�b��?Y�8,dy���~?Y�OV
ɞ����DO�VigR��VD�S�d^h}�*��
����e�B�,�_�t��e~K�/[�l���A!������@��U��~�K�-ۋ����u.'�T���6K�N����ep�NP��J�K�r+�h�!�Z����J�f)�(�%�Y���BdTr�^&�I�&�z���I4�B,�	Q!�� �ǁ���as0_�bR�,&�ψ�� l�r� >?	�>.��<�X 0�\6�C'�i�� G�L)"����D�B#ɡQ��rP9(���"fj�M�t�0�&�s��$޲�LM���35�.�)rs~05N��	�8٥ ��C��<�V�kj���$� ¢p�QlJ$�N�Y4��Ƀ!�njT*�Z�`�F*���Q&����Z��f�x<			qqqN�����ޛ�xOLfjZan^iaQq~A^VvVZz��c��D(_iK'S�9��z�|_+�gj����g��d	���h%?� J7Kӌ�=7��-0��"3��B/�ҽ���55�B\�F+�H�����@C�dm��1Eޔ� 4�)[�Um���,mG��gj��txv�>S�۟nj�|�o�����İ��"����ww��5�V��N1�	Fa�Vl��� [ժh��m�'ZM�Ѷ4�3'1�0-)?-13�����k3���Q'o�-��Im\[{���W�޾q���ks���������տ�o���{���ܹ�����0'/7;51	�S�X�0�w�q�ޠU�d��𽦆�#�x�(p�!�E�8�ߛv���k����j��Rl&�Xi^YC+��K@��	(w���!IМ.mLW�`�(-�����^AXIXN�{���Ej�rF�JF�*f�?#r53ʟI\�"pH�������a�j������`��?����0SC�H\��A��'b�I��*>Q'���4�N��l�2�&F�&QՔ�nN�4���RUk��X��Da]��6�_�V��ձH�.q!�"5�l�8�-O�hcb,щqљ�5��N[�NӚ}��G�k�Z;��;�9֝�^7�^7���m�k�P�3�g������gzG��3���4��/���?���}��W�_�ܴ���Dˉ�����W�}郶S�k���Lh����O�p }�!@ƺÀ���s�,X �fKz����5��O���q��cL�x�:լʶkr�|���"(�
Jl��|/k��`�v����05YN8��I�r�VN\��`��yFuF�����u��6�;R9p�tt�rz���lݵK�ګs5Wf[_��py�������K��]��������w���|2?������5?���[��֍�6\����G�y��G�~�v�˷7_������+��_����˻o�l��������#�����<���{����ꂒ����)f:�i�-"@�YTeU���Fa�I�`4��MfA�m�����V+�j�q6Z�یp��wPRpʡ>1c���+�v��{�(�(���r�:�&�,A?1h��[_YLo�ů*E�d�u1|C �D8w��\�k\�!��Z����&=nj�����7"ɯu�`��kfj _0ٟ29�0�x��=���w(��d�=2���,�G����!���z;y��^#¯j�#:�]}��=������_���������^����3����NF�M�y�%�Ɖ�i|�ƿA\���:�|8�HPX���1�`����١>1?ya~��wmͯ��\�ϑ��D��e��H�As��g���8�;I�L�!�$��]�{M��M�$�e�/VF ���.��8)�!:���3���DzE)�jP_��܆�8éݡ$��x9fjeej��^S#�Z�&	�m	|0����{-̺Tq&k��i�u������)�d��4,��>Yڑ,kKV���ZҌMֶ�京x�b��� ���!�c)����`pUC�MT+* Nǔ�0bH !p59x5'"XL�P3#�K���W���9��`p����Ϸ�=�t�\�����W�5����O����_?�ya���k��J˒�:.�����L

Y������/�)�E�I���T�Q��R���Fg���̴�H��@��P�S��R��.��fk����M���lp��,�6�ֽ���:Ǿz����k\�������z��M�8��D��i|j��S25O35��4<nj���yD��8}h�B����� L�.ݟ���'�_�6u�ā���m���x�e�x���#'�G�Ռ��@ᙚ��t{u?�ҍ5����ao�_��˚G��,�5�͏�Ԝ��L͹�R�g��?�.�%Gݔk(���5<L��X0h��|)��D�r��Ц�Z�Q&�p<��K%�.1�D
�D �F $1�"aS��f���(y,9��Q.���0�Ka&��j(�0",
���35,R���e�0����;%�q�5qO65�q�G�A�v��45��l�MM_��� c�W� ���S�b���³єC}'��NZ�٩2Rd�����Fb�m��Tq����o��L��R�d�X񩦆ǽ�pgQx�MC���8�=ə�����<���N��?MMϿ�`��?�������b��~1��/�_��ǎ�+.(F(��{�_#s�R8���-��i�f&�<I��M�BY�38��y�
�@%o����@�>�j?���K�<��|�� �������&�e�&�u�ʼ����9I��QȣT��>NgS�t�K�!12,�N�x7��r�
�r�-	N�2���A	<���c&ňE}ެ8n�2Hv��N9�YD��jE�)�V��x��)�ʚ�'kJ����j��Rb�(2��F�d���q�,�����m��:59|d|�o�잩�#w��|��#o���;�����ҍ�/��q�N�ݻ}����׶�����W7\����݃�櫯.��g`�ij�j`�����5�����Ճ�%g��o�M����ޚ�ґ\Z��:��#�?��pj�j! aGH�����0�(��G<BԆ�,|�"B%§EV-]�䧋�.�[�߲��V�-}q�����/	�{>p�s��WDAt�Ffq;RD����'��G�H\:�Bd�
���$,Y�xY����~+V�X���/.]�lժՁa�AQ����+�V��/[�r���K/Y�t����)�e0�(�E+��УD�TH�����c��8ϭ��r�.e[�L��a��b�N�ԋ�1� ��(��[�X/�J2�V*RI�J�@*B$B���EfA:�Cc�h�3� ���� ����'���qk���jL`6 L�n�\&b��4�I'ER	?�Bh�BSA
�$����AX�����|v�N�n�g8$9Ѣ�h��O��w@yV���H��;����xX�`��Lfj�lpG�צF�CM2��KE�T��U8t2�I��.75�D��$R�X"[X�[����9"�H���F��&r�\,��Jm5�b]��Ĥ��Դ����8��S�E(�Mg��9�N� F�t&�Τ/�t*��A��d&)�Kw�L���P!	Fa�7S���昰uOyFZ�������6�����������Z'0�e�o��a�D���l-3�9�_�L`�=�S3>��m�&p�����[c�^��V��t7�XJ�)F4� p��9_'F��Y)w�4.�&�jLrZSݎ�O^jBVrlJ�3�mK��uj�V%6he�-�eey�����o�y����+Wggf'F�w�m߳w�����ۿk��uU�e�9�Ԕ��h��lqZmX��75`�v-#���	*s�΀�D�H@ɑ"j��C��ߛN���k$�25�Vr��������,��S�j�Fp���h�5��J���
��(�K~ϳ#VX`�`9�`�¥�r)��&��(�j �$`�! )�Dd\�3��D ^W�{�?���25b�S#C�K8�
8R���S�N��6��������w���RL�$�����Sǫ���b��3����|7?ύ���&.��s�3�c��j7Ŭ�n�5����t.a�����Ѵ�C)�.$���[s�T���U�7�n9��µ[_�õ�~sh���׿<y�Am縉����Z�:�����Mi�)X�_��H\�&w�:@|ݖ�������l���v�n��53�9k\���b�+�l�X�6���6��L�t�6۩�s��m�|��Њ[y^S����256�������l��AqV(�#2YxZ�Е]�Z�vwWۑ��S����'Z��vܸ�����wn��s�~�J��X��t��x�+[.]���o�埿����������?����/�~�s|����}wn���w�����7^�;77���;�3~�wb�wlh������}���8vx�ޝ[��w�T�����L��؆�i��Ɨ�1�L�	]cF�����m�"fv����������S���DT0�P�"�0�����j\H�$�Ц��a����+��3��M��9zC½*d_C�7��0���������J���F��uZ,S���V&��T��j~.~��A1Y�%��e͗,��� pS�.�x���e���#.��Bk��]:�	[��}�$x��^%A��cf���?�v���0����˿���������_<�Uy����kb�W>A�'"8�)X��2�;K����A�xh���sX�Ϗ������7��ϟx���ʹ�;Vg߲�"�cT.� ��P�1&2�FG�8�3����)�åO5��A�3��� & �����I4)�Ak��esf�D8��M�U����x�z�jG�lk��;Q���4���3L�eͺTq�W�<�Ԥ�x�fS2��ٜ*Y�,mKV���ZR�ͩ��tKs^B�]-gdl�Q�����.W2��A���zLb$��!F���L
�J� E��C�%��Ң4�(a�r%ay�	�{���P��c=�k�x�����7�7�>�8��j�p�룛?{����]xkf�؁��=u}m�%�V5�
�kݐՌ��Ѐ��� ���/zq�"!D�+Ji��\W�؞o��B��
��MO�xK���HX�k|���삃�����f�Z�B;�����=0��m�G��B4>w4����������>�*>�W
8�W�s���gj�������:5O���΢���������|��'��>���[/]�:{�P��=�g��n<���:5�+F�)9�˚����r1Y��uj~�5��_����5��9�js��-��{��w�l�>�1��ܶ�<�<YgȹT1�M��`��Bl%���+6���C��V��<a΅Ð�8!&��� 0��(!�$��d]�c��`.�D�DS����1�dl��LYhj��6��&������
��X՚x���1��8��y\����橙�=��B��ݞ|-`w��?Gӟ�<+;����c�w�o��=HO|��r?3孴仱��&�5��@~�\��X��t,�2I���L�2��9XM�dAcT��5Κ$����L���^C��F������r�?7��?��#8}:���8�����3t�0���\&x��|oj0�bjf#)>Ss�ºA��b`�i���4��Wa���-Tz�[���xM��r�2����OQ�ǈ�35os�X��ʺNa\%�/����9M��Q�#$�0�4B��R�T� �5*@G��AoHM��R�
���=��D0Ǉƅ�1g@���G5��ZTg,�c�^��G�m����j�FL��3�U������)?�5EB��25Y"B���("Ǌh1r(�,/K�4��m۵uߩcG�����z�D����ӣ����\��<7�1=�21�81�<5�:3�:;����Ks��`�y�Ճt��N�M��l��P��3E��V�9�.&��M��Wv�h�᣹�7%�UYc�0�㰹42�nH�A.���4��nA�.>-��P�U�إb�Tj�8$r�UK�[�xŊ%�V���Y��򈀥+_Y�\���V->(x%12�	 FAt*�F����pfH# ��:���\�����|U����W�X�t��ߊU���#�#W���[�l�e���/�[�ly��Đ �J�sF���$�j4A����(4h���Vr�5B�I�ԣ-��r�"� ��R�A�`�F��ID�d�kt2�~��/�!O�B(njXT[΃k���� �������'�;!���	�kxl*̢����x�	��j�15��0b@)0�R"�(;^/�r�r���.I�[T�/��-45�h�7��{�OW�F�c�94.���jh$�A��4p:�8,��|<;#b-�a
y{l�X,�wc2�xU o}�Tإ��T*<�a�E(_)���p����v��
x��aRd!<",(840($(�H$�S
�D"��
��J� Ea`��0:!|���@�N�����T���r�P���k�����<^�75��n^�.>Ǐ免�qp��joʦ̴�Ҋ=�&��ƽ��ݜ���T?� p�)j�L�Ȥ�[�*�Qo3����1��I��i��)q�1�Zj�)�H&��-�ۛ�k��l��{��k���LN���MNL�������շ}o����ٻs㦎��҂����Դ8��3g4��#���]0�]�ѤWk��/A<��!���(1\@S�"-(%F��+S���YH�V*�#���ͩ�@�r�,�U�kɐ�/��1�  ��IDAT���%�$Z.A�!ș��̠%p�jn�?�A�1S��� �Qj�"`�
�a )�DQ3��?75R䡩Ø�CD��	^V�1C�(儩��f	5N�-��˝��4��|�����I��75���R�ă��<�<�8�#K�bn�5:1����̯���9��\}1���7���:��}!��b����΁���֟�g��T����Ԅ�u�Cק��x�����;9���-���c2K�RF��7t�o>P�q�6����eH�+��e���p^��%�ѵ1�%�g�Y[&ߒ�7$HM�*s���֪mz�Ѣ����T�1ˡϋ��Gk
�B��ȂY�@�BS�}�ɷAE6�����ɲs�m�$�@��&2�h�K��m�<�ӹ�G�M�o�4������o��|{�ݗ �o������߹�޽s�=�ʫ��._������O�zMͽ��~����7�{���33�^=x����[��x��Gﾼcvr������]���m9sj��Cm�w��nkڼ�uV���2�$#&ۣˋ֔z4%�5^M#�6�kM�z�`BMH��Դ���5FV�����0���F����[y���!�D�{`�~�|�C:@Z}S'�*)��X���߹����aԾ!�,C���+�U�q��xf�
��D8�x�+%�i��ҩ�Q�N���Z����R��$2_��;��-�~���9�/Y�/���O蜏����w���<�r|�����Y(h|�K�}Ȓ~�U�C��g��"��hl��o����3l��?���?����0��'�ݞ������'���:���d�x8��w�.�NC�H�K�0�v�@9|�B�M��������1?1�i]���5_��=A%�'���7�@&��7SOС��f�śb{��M�O�`���i� ��6x�f���2/R��sD�Y�Lp:�4�&��B<iP���������J{�]��0>��,�5�9��RDm)��TQ[*V��[fِ�lL�{��H֥�;RUmiږ4}K��1�^��`���4� 2KE��p�%/�F����4%2�N$��D�L䒣8�H�H�`�e�L6!�O!�$-�����A�J�`O��}���v����W�w�>�z�P�؞��=��G�o��3�={b���ʾ��-���V=��F���A!�W�"B8trx�ߋ�-Nͧ7$n���R�؞chM�t�({�[rĝ����B�����75x��`A�R���L�i���pSs�%�ٲ<�D��i�t���̣<%S�4Ssrw��=M��9{`��]����O���� fj�������/����w_�qu�̹cێ�n>��|�H���k���>R5r�j�p�CSs�r�)�fx?��i��^PQاf����9�wr��LW܅�)g���mM?�9cGC��Jwe�.ΈJ�UOX �H� ��`�aH%@�b!�|L��	M
~ǂ�߲D�@y2W�r��0\Ѐ	nm�4��EQ��V��	a �h�x��V?="h|,45�����tR�B�H�"j��GM�"%.Eu�\m��p�zh���d�B_�?��<bj�rՀ=Y����x��X�H��Z��դ�Rbog$����zj�+1�[f�u��Hy�/��ai�iͧi&�Ȁ�ej.sؗ ��3�a�3���pc(�9ID���T�y��횦?�����������w��������ө��T�^6���(�T$�2�J��R8�(�ggj梨��D���ܤC�\e�����.W��[��'��צ��2(����S��cD�O����I����(nj���W(ej�H�!
i�J�чh�a�=*B�%��s&�M����}���^�J|UO�أb�E�R
���a�jȪ>gӜ�����۵H��Q��"J��^�`>�ԔK�I�W�I~�5O����H�rZ��+�ǫ�\�~MaJ{C��3'�\8wx������������S�.O���o��j�4�~e����KsMss3ӕ�c�#��3^����{���c����S��Ce#�`,�x�h�b��P��=��{�N�(���v�3?ߚ�$R(�ڹa��()LV�h*1U#��P���q!�
`�L�˭R�D	^���KV.^�r��*��U~�K�\E���\�4l�A�eKBV�E�Z忊ɦ��$�Z�����|q9q�i�J��U��+�_\^��-[��oUP@`XH1,��B&/[�j��~�V�X��j%1$�K!�94��V
��Rp_�����%��D����k`�
��s�2����iZ>M'`j�L�C_�Ŕ������O�[e��J�J��E<��+D�(̀9T�E�0)<6e1�l&@�a	!6@��Hx�'"Caz1�%A�`"p`v�A�>(ʦ�xd���zT8�"!<�J
�
�B��aĠ`��PC���|J�Q�J0����l�4�-)���܂"�ש)t�j�G��#�����HytD�҉lJ$�B�j�x�,&��f�0�z70a�!�M�ѨT*�B!��>LH$�H������ #8��a������z�����
.|*2^t9*,<,(8xu �}I N ���פ�� rT8Fd(�h�D1I��"�i����� ������I����{�W��L����+0�k�@��Epw� qq�9��$�l;~~�Wu�޳	��ܻ�Ͻ���zVU7�3m��;��]���Շ���i�������25K��K���pB֬�χl��E4��81
l��nDe3���	��!S�|�lvG�@��),�.�9ؠ��	�����r؅�OѢ�������������ƺ��2��춙h����ߵl�foܰz��g_}���KgO�<r��={�߻�֮z�Q��5�?��C�/�?e���I�N����X]^!�Ѭ����P����U�	��UKl��O���p�kM�_P3�E���k���׈���VlO���{����,�p�l���Q�ِK�2hU��jA���[R�������|�̔�Lh	S��!��[�|�{�Yx�z�ܸ3��8��:��'��	��d��h��`O�hj��1��T��l_9�S�w��K�����2wUY�����������u��y��y��e��Y)���J��h�$"Yx$�"�F���U�)��wϙ��]{k��/���C�l��h6�p�2��M�Jʺ�*z�S�1��77�5F�����*Mʐ'e���ӏ�"�J2ME��	d֐��5Y6��c��B��P]�����^��9�#�B����-������ש!��B����+"���`go)����0QUb�ۼk���o����]����[���m���=�c��;g �@_�?�c��;f<�}��]v?�ȑ����]�k���O�X���W������7{�滿��ɷ��w������>�rÑ���x��_��qc���+�n£�4Μ>�%��.��t��%��/�`����3��N��008���R�\l��{*���?�!MswSC�d3���@���b��Z�6ى�&d-���+�!R��Z��7"�a�D�J��W�,�~|)��8��u�ʜ7�Y�4e8GAW�:������m�/�֯��_�m�:�w���ڿ����|EP_��/ⱚ������B�w�Ȼ:�]xG/�Bݑwa�@�{������y�H������o��v�����o��?n�˿����7?~���s7������q�������;��/�Q�)5qL�� U��@�ȔϨU���<��͓�o^>}�M�üy�2c�IκK���5z�@E��}��M��a�F �b�#$+Ԧ�4�p�5�yaJ�Ĩ}0}�sj�v�zK��ɜ�M9�� K����}qS�L�{C���2��
ӲJ��*��cj�V1��F�����N ^r�8��6��=��?�%4��hfK��"�X�.�s>���a�<?G��)�j�
����iH�V�k�����x�;�
�Z;�uc�<�c��CS�,˻�W�ν�u晍=1n��s�WN+��[�ey׳�O8�e��e������&Rd�M:T���䁓���*u������|O�ȤB;6�\�д�ƕ�i��m���`�yY�ci�;ʚ�삃��L`�"��Yф��&h<9���,S���������l[9(����Ϭ��u����=�~�XQxǆG���5�Ǚ��Vm�����L͍w�|��7@��?���O����7��9}h��g{���<1sדs��4��M��<9i黎�7M8�閩9�y¾��~ڻ��om���Q� j�n�o�~��@����w<P���u;��<��a۲�u���+_���<,oG�Tè� ��ߘ��mς-h{�Ɛ� ��Zp#j0�:�� ����A�r	��0��D����� �M���Y�3qSiu���Z��0�Մ9��Ω��J׌j���;����E��6��65w��<����
�j:�	S�����ֹ�ʹ��{���zm��2��M��4V�T_�beٕh��w���Z�h�
5��4?QQX�'�b�0������O�M���x�t�3��p��'L�ˎ�o�x�����ӛ�~u�_޼|��)S�m[��.~P�����*�=�
��	S�	S#N�J ���Fl�G��R5��M�����~��]L͍aEj��:�����)=Ç��}Z�>�v�AwF��I��I���<�����f��������{#�{����O��Fl��`&@��f_ĳ;�{6��Th{��.� �9�$V� 5�,��	S#���5��[��Ϩ�[��ۮo�jM�r^W�a��cv��)k7�{dú�?��U���о��n���{�;����E�.�ta��ssϞ�y�Ԕ�&=<t�h�>v��s/��u���/O:v�{��]/<׶s{�ӛ�<�����g6ׯ]����5,)�8�������4�#�s(��k��k�<���j�.�#���8��j�٭Q��P���2F����H��2&'ml��9i����HF�&+ې_�I�$J�Ԑ9=א��ɒ��HF>,��FI�F+��ȓ�ʒF$��N�75��O��1:slj^Z�4;[�����Q	����������<L�_Dn�~s��X�f�WD���s���K����E�����F,h�7x��<���r���q���!.NP6�6a=o��q�h;O�Y����hLO�:�Ac"q+C�	܃��6��h8y
 `�ʢ1Ӱ��)�A(1��/O�\/��fj ��Uv�2+K��e���dyF�<ģ5SK��^lzK�}%\o	�S�wǰ�b�4�@v7�ˉ��L�W�j)�	� 1���@����"W�T�aQ����*��5l�P�$��ݞ���x�v�nj�LM^Vv^N�T*�H�2�L.���5J�Z�P�
�yJI�Z�mP��` �6���5L�>�у���� �����25K��K�\	��q2�X�&����	���Ԉۄ��o�`�����xE����uF�ո[#暠1�`CfZ8_[�`���b>OUQ���������a��������"�y���s0��;g����vlz��-����]�|����G��}~���[�yr��5O�~���\����L�1y괉�fN�hi����LEI��M��m��X��zX�@�r\!�TH���h@�x!�
5auWHsGY�P�]q؎/Ŧְ���s:�K&�.W�]n-w�m��Q-�}��P���hM��%���,�g��|R�Ki�h]>k�p�t� \uGnS3��ij��J魔�B�25L#<.�4�R��yvD���.L`4�6���c��x0^ޖ���������1O���3#�aէ����zⱚ�rs[�����P�o�+mnm�nnU62�R%��]��7u$k��I��l<)IJ���ܓ��m�7]E�����v��+G�\�v���n�:�LL��,��f@[������M�
6e�,/Ӑ���ς�Ӕ��#�r��d%ݗ�t_jҽ�q2�Fdޗ����ʓhr-�C-,��kC��"WG�����Ud�	��a�/�i�����@�g\��R�EDg��j�d]�\Q�(�8¥��Ά�9S�=��o���[�ͫ�5�b��Є�q��>_O���%��i���WV[be���i���w�����n~��ν����w̝�,-/��yt붳o����+W�u���c��%CQ5A�i3YX����
#ޢh�����|.KC���6h�,�U�͉4M\��� ;-��0���� 37H�2�azn [�R���F�т�c+)�
D�����㊕�r-����B��F�B�7U�_�D~
~[X��p�=���L�f�S��,i�B���5}�#?4��Z�_ZM_[̿��~os|o����$���O�
'�D�/`�3��?2`�kS�^�Լ�' ��� �B��ށ���-`�-�aMG��{�gl�#���n{��?���w���������_޼��_:q�����c�uo��:������z�d��[��j���{T�r�������[���3�m��/fN}�����ǜW7�����~|TG����
5��Q� �I��CM#_��h|����M���Ip %�F,X�]�~:_�);}F��Kb�M��eo����hj*5>Pn\Za������6Y3���g~XP� �2�D�Sg�Wg�S����Z�T�_j�:��ފ��g�j�N	ò�H��|k]`�H���i�3hPH�CZ
ұ���"N��6?�iHv�[?����|q���&�~t`�܆�}�9��]�����ll�'�]:��̮œ:���m��,) wK�÷��l�BB�:�4k�=Iyc�BF���C�j����Z�b�����F�5b�FԀ�}�*Q��L��i�͌��F�5��M��M��5�I�.���� �=�����Ȗ��mY9Y45�mX�ܦ������o[���25�	�[7��`j�:5���G7���_}��k�O
�f�ʍ��ؼj���<�a��'�����M��>9���C��9�y��T޷�m�����X;5	Ys��I��RQ��ҭKcO-*ڹ�b�c�Ϯ�ݾ�n���M��D�չES#�I��Bd0X�s���;x4�F n�4�6�<h�,�B���i;L!�lc>Gu$�T-�;A;�E����A���h+O�4Aa�(���iPo�PB�v�ujkx�ѡz�DQ�����h�o����i5�)e��Rݏ�@%d͜
�LSs�L��n`U�ge���8�:\k�\��OչvT��Uy�T^�-�^S�rM��/7T]���^Sy���J0t��>˘OB�I��,�����u�N��	����}:d�R05g�%ڳ�`�C����O�<~�������o�r���_?�����'d����d�Q~B�	�F��R#�T��O�����)�pF����5w�5��M�8�M�.,�drݰx>�z�=��-�F|�9���>m����Ʒ�M�LB��s�C��a��d8b��O�q� �0Q����,��H���/�moz�7�������}ֳ6� ���fz��x�o;T�9T8P�SY������[l�f�i�V(Uc�M4��fj�[uB�&.k�,���1� ?��i6k*E1�����J�k�1���5�Z���߾��=/<vp�����?�g��ݳ��{���3'�==���i'�O9vt��〩�����s��^:�����_����^�8xp/`����{_���lߞ�ZW������X� <�?6�n��͜��Ÿ�Aw���F����&��
�P��}��"f&f�D�VD����52#ct�{3Gݛ5ft��Q�{GJ�-������ḰsdT��7�^-���J�Aآ:Ɨ�3*0׈��,4)U�4V�4Z�4FrO���TI��̤Q������?&� 9U:6E��R0vLf�،�䌴����EN.��3��4�Au��\��=T�����unP�!� 4��d�/uQK<\�|����܌N�ظ�`��Md�Ɔ���By-��D8M��G-<b�`�I�D�fX(�Jc"6�#N�p�؏����C]F< 4���W`k�a`eP��VBr�^Z���S��(��9� Uv�"3S%���<N/�%���M�=�w���eL_)�[J���������fjT���J�SJ�:;
�Z.Ѩ�B�%�/j� �_��Q~05�L��_��&��~���8����p�F+j�DZ��{��/�ɥ�<���cS�g��y�^ɡ�";Y�c낼hjZ�X�`j���L͒.��N��X�f��jn�5����G'>>1H4�W�I����z�B0{B���G��=4�r~O�P��#f��J�\���\�nڭ�5�t�5%��Օ]M��-�M�U%Q��L���
�}��L�5{��c�{~�{������x�+/^8r������޲���mظ����-^�`��Y���6}R{[K}uMy�PYZ&���x�@�G��@�:�L�-�\B*%��B�ev�·��o��n��w��]!�pY&�5��2TNL�ag4Xf�z���?�d^_tB�����tC%�K�ݤ�,���ܒ5�lJ��5�V>\�An� +��*��	�y;)�-h�ߏ���)������Z	5xDa�pTn��P���iu�UU�I_��b��f���\i�^k�Iq1�y��a��h�Q�M��'UC��rt����z+�޸��*O�w]��$p���婠ѹʤt��<ͨ\�}���T� �G$�'I�7�ޱ�Q)��4�}��Q������~��>�r���;vO�;�S ��f���C�z�:�ApRS�銌��%�MJ��to�=#��u�贑���Y�\U�=)��V!yo�}9����f0&�[[��������*�{����0�	�����3Bm��(�B�ظ"b|�'̍"DY�a�������[\��
+�ц�@E����V\��q�G�+�&���:mR�Q��R�T3�������}'N��z�O?{��O_8|d��E��rI��%3/�0{vqC��F%���Uy��ԌܑcҒ��t���_?''O&-PIsT�)�$�Qc6��E��iء�@<PCO	�ӂԌ 5+H��sC��X�����ǃ�z��In4"O���P�
D� *ȚG0�*T�V=iv�U�=�w����ߗ��$�����C�_�y�o��/Z�3|�ԝ!t�	�Uz�F�a�F�c���g�q�6��%��3Z��Ϳጿb8Q�|EP_���8�O���!ES�1����}
xOO�o `�B���������כ�*���W�qx�U���7��M<S��7�򗛿����������;n>��˶���1�rTǜ�q�AO2^���]�����<�s�/��k��u�}�t���'�q���X���C��i�<�����^��=�i���qMv�F g �e���¤�c��8g`����'f?����v*��d�-��y���4�#��,���=�l�ڟ*s���?X�/+㗔�K*�	S���r7S3����&!kSS���1��fQ�i^�uN���&T�z����搥!d/���N�oa��<c�9��� (� ��3Q���N��nM��P���YI\Xb��C,R��lHO��ɥY9����MϮ�޶���i��z
�w������w��3�M��;�z�������K�V'��B4��'�4J��:�<79sT��`T�E7T�]2[�^��Y�n�pM#�~�M8���Ԭ�Y?+:\��&h�G~VE������y扙;��{~�҄�ٺ��ej��fg�nj>z������~����|��/>|�҉S��۾j��7?6uד�Lͮ�C{6�����<a�]V�޷� ���k��6A�@t4�5ͳ�K�toYݼ�p�򊽏7<�`͎e��h޼�eaѸ:we�1"rYN
蕊�|*l,�2�v��:�hx�f��x,&��"nC.{mIQmqP���-����ڡ���"E�[t����e	;��Eی��?�@�Eg�A��b���t �Ѡ�?��=f�2��B@~-2�eVD�(<��6���L�(k���oj����Vv
����ݽ���d�k[�ko��Te�Ś����U��j^��~���j����s�1�'�DE�D��n��-�!�Y;�cG�x�F�V��H�g�E�q@E�1�7t��+o>����gn�z��9s�U�:� Գz� �ӳ�Uĭ@�
;���*MsP��iSsZ�fj��'Lh'L�[FǻF��f�qM�������u7S���Ĺ7p�L05��� �q�<I���3yC��A>L�'(�(Ib��Fr�?� L�y��U����C���P�H����>����Y�.���h��,|�*z�.�9l[����9&�t^7ը�h�N0j~�� �F45���Դ�T��"�Dy��8��r�`����.}���ٰ��m�<�����m[���%��,;ud�飋ΞXx�Լ�'�95���Y�N�8qlƉ#3O�u��ܳ'�^�����7~|c�W��?�s�3��n:�g���vn�ؾ�䑥5��ٴ���e��ݡΖpS5��V�Ԙ���{X$ȣ��cj,\d��-�"��U�����>��ޤ줤��FI�#O�O�4Z�4V�4F%4�5#2�1�Y��Y#-%�S�zfÍy�S��� O��zO��%�꒲��"SI��2���TK�+�(#[���=:k�̔1�c3�S3��9�B���6L�R�L_㦪ݨ�i ���G6��F/]�$N��(�!��1���^J�u��!.B�IBMM�C(�*V�Yi���IQ��Ih��u��%��F���7�z8�gf`�'a`�ɡ!��@<f�!!�kT����'L�-Y�����P�d
�0Y�Q'0&�s�EL[��1}����+#{K�;���r<ag�󿐩?6��P�ܠ,��T��4_��(�bLF42B��N"�H�RY|~�p,�h���L\�r��@��G�N�-����:|�V'jY~A~v�hj��c��/r�D� W ?[�������r�R5���*=l���9�LM�W����,�t�������M�<<.$^n����(M"\�	�X��\��G�>6���U�zK&6��kT6�8�B+��a!9kج>�9��TF�*�:���Z:[k*ˊ�,<���P�[X�8iܼ���]�����?��ɧ������xY\����������@͜�3�M�4i��ɓ����j���%��MM,�P7@,3�;�F��a)�@��Ti���,njRU"��5L��ր���-��F�5�X`J����`�
�Ǘb�*��5��6����n���O��)���p[11�B��O����
I��<V�K)���E�� � ;���j�S R,q ����13�ʬP��q	Sޜ�=9��!���-��M��MMu��T�=Lw��Ufi�YK���Ԃ��董��yϨԑ��B02��1�#�%��JF���Y06E��&O���4Z��}�����/������x�'Y�w�52C^���M�v6�N���JD��{_Z�謔Qi�陹那�L�JK�JN���5jl��Ԝ1)�#G�$%�u�}��\��D�^k]��Rhk�X:('<%#�pS#�uꋐ�!t0��/$&��#}EDW�3�2�KCU�����wP&
oO�1��'V �9z}�V��Վ�J���J��3�7��06<3#3s$s-yd՚=�>q�ᕫZ;�?�������n���qB�ծ��ZX#��eKS�f��/垤1�$��'i�=I����ތQ��N�r���1h����4��h�yOS�� =#@�Ps���$)��!rY�x0D����r��UC��d"}�=�*� �Ͱz�A�N�v��������/e7���=�}0���s��]����9�!�I�i\{	�_š�(��%?d�O�K���������I05��L�a�_Q��qM�N~C�25_��/�s�� Ț4���V057t���Q���u��(s�=��	�y5�������\�����z���_|s�����˿����{����=�o�^�Ys�)����1g!Ӌ��
d:��.�K�;W�=K�9=���S�|9i�7��}2��	��{��_^p�O��S$P��ii��ڀ�qMsGSs���FL�$L��=�%,�����v(4;����zq�gU:�N�v�j�^��<o����)�l�YW�YWĸ�������nP�Ωc��Ҁ�q���k��m�l�j��m�QS���t�%�.dp������m�L4m7[�N�p ���f��aB_�փ�#��)�(�����]d�
7S�$��!<�ѣ鍠�{B�+��Y8�-8��hV������^}m�l,6��N�mj�*��,�1�(�V":5�B�ʞ88��j)���Ef�>���U=�ٻ�?��'��Ƿ���cM�05b��8��������&b�G~�*�?3S������'���<r�L�m�&�3�W'ILӀ�w�������O�}흗Ο?����+�Y7����wn��k�̽OO߻e���'�j���9�q��M�uj�jnթJ��mEa�X�F�G#����Ih�Ԉ�&�m�f۲q��l[V����͎ʅ���l_ѴuE�����&o���Sj
V��2�����)1R��a���,�a2ٍF���l ��p�bAmIQKuIWcUgCeSeq]ia}YQsUlkb��"_Y�Sr�a���0�Y��	����@ZH��;3�����(�8ᐎ4h���K�>���?f�\i�YMͮ�g���h��4 И^�'@��fx��n��#	_��ո��"h�.���.�#�N��L͓��-;�u���Q版�\I�ry��ʗ��5�\���^^v�(�7t����.S�?����G��m�q-tR���0p��q!_$�Ku#�a�� ���{���G,�t����p���V�nh<+9�<˛�@��a�B(lvTC�R�Y��T '��Q%8����'�᳟DG��⩙��4��Ej^�M�B�o�����w̮�L�w��wy�;��m��c}���MY�!-o�p�U���/��\\��,��٢S� ���P��8N�Gi� ��7{��^y�L7��-<��}��]�m�nD��B���]�h�y<8R<�Xqu�m��z2�z��M���ɜf��nG&��d�ȐE�����q�S���p�>N��+���������>��âj6k�iy�V����-e�'���Y0�C+[���U[�^�k�#�w>���Ug�.;v`ɉC��8��Ա�ϝ\z����|�2h/�|n�ՋK/�]t�$hl�载��fީ�3��r`�ԃ{f����nmۼ�w˺�5u�~�a�\O���:T_i:Y3�qO�M�ʌ(��Ki�.������j|��G�~�Ѵ�6�S��Ji�A��T02E���ױ��*����<ؗ�səj��L�������9�����G_횿��vБ���e��y���In,�A��*��&Y��C��5KAgH�1Y���)����H�u_���sҳ9��B������Wx�
7Y��*�p���"�^�^ F��6�Ԇ�1L�	
q� ��1j�LqH�C�, ��	[ɰ�
لm��)t������I��r�� q�k&>%-�ɠ� �;��A�f�KS�࿻x��"6
1azZ���r ,/��0W��iiz�<3]���4H���a3\�g��LS��(�Ji���0!PS���s��j�0���1��T_�0Z�)&O��Ё6���P&X���a:c��RGs���ǆ턃CiD�W�k�9��in�,?G%+�I$�.�R@A�pP*���$.	q���'
���n�1?�<^^(��h�*Y~�$7O��//���˕2�`y1S~*���������2��$�,�1^�"��X��w�[<���;��	��zA�D�0ҋQ��#'���٩�Blaf�mv�C45	Y#N9��-��m�E���;K�\b���Pf8�k��FP0��b��G�����P�t���	���Mj4��r]d!��k�]x's�(�����e�HUIImyyme 
�m���v;}o[G�M�/^����}�͗���7}�����Ξ;y���c���k璥�̝1o��I��O�1y���]��u5��%�"eű�Ҳ��jQ�DÅ������A�7��� +5�R˥�4�T��`Y���0~�!�ɧn�b������NdjƗbC���*jZ?��8�ñt�����L,���ꈱm���.w@^Jj���ĉ�������^j� $��Q�2��@���;	����;�TnJ	��*��Q��H����;p��l��I(� ���V�/1?�	0�B�.j��,�
;R�!�BL{��3�/�&Up��g<�l0M��g53���̴:zj-5��TM�U`ݕDo%�[I��S�e�ۃ�,���Sh�3�\M~�,;#73k̘䤤#G%�;2��cG�L;6'5� 5Y�<&4r2�٩��%�dp�����������ٛo��q��>oX���2�&N�2yf_�x#oS�2�:5%+7G������Z������9�Yٙ��yi�9�cӓ�SG�5v��Rt��C�ƈ�)jo�X�"��"����)�{���V1E���d�@:����1A�t��W�ZJ\徠�d��(�f�%���c>#��ψQI��H=�������������������1c�[V�6<������>�j�ԙsb�U���L*=�ќRѼ�+�+4z��g��d��L������V�������16-c��Q�fߗ�HNra�ƀ�=���/�4�'�5Arj����g�9Abv ��G���Eajy�{8®
�k�̆x�f�[�*�e�a�a����|�"�i��0
}|Y��M��OE�	�����1�s,���[v��=Mk�ҺӸ���N�35~��>�/y�k������7Y�[�co75_�ԯp��X<V������������E��"�i����zA�|�0�,���6��'8��0~F�>��`v�mn�����]���]�K8�g��t���_��ßo�������ˏn��꿝?�����_�����׋�vH᳄�,d�����-d��e@���D�G�9����i�坆��͘����x���?t����Q�r�Q�-@{8b���A�R5�0���pSs�ᅂ5q}#,��$ʚ��� {�n="&k�u�4�j�6�j;��n�wx��E�M1���G��+*�?�(����Ì'��ܑ�U�P'�
�SMέ���YX�/n4?��^��ReiR5N��Y�U�	��2���SB>�l��-��� ��h��0\X�҃q�8�2�F�i�,YI��R!#Y�t�y�=}��R���(�&T٧7�gwD�6�m]eƶb���n)1wTz:kB-����g�m4e�_�1��`02�PE�,,��륲���QA��=�Oo�,�/��,�/�-鲋�&ag�F��<�C���=�{	e�ظ ��fj6�-�0�x���mӠ6Ή=�C]aq>�O�l�W�iA��E	S m���F�<P�Բ���e�3�l{�mۣ��tm�{�Ja�nq����=�r��;��}׵��&k6�~�5��^�ؖu��F�Ԁ�g���/>��W�y���������ֵ���>�a�hj�?=��SSn��ḾM�k?�_gj���"P;��fv�wb����s2ZL'�Kr���hcq\45�����h�rغ�ք����U�pSeqgC%�����<�X��LM,��xmA��nb-��aILL֠qS#΄�z=n0��F��
�&`=�Ss��M�\nC��do�4��8��^���L)V���;�����w25��f��V���@�O����m���x��l,x���Z}���ʫ�Wk+�U�`jޫ&�e�;a��Q�+��M��9��`�=g@N@�|B �f?���9׋��H�h�]Zj'�m��;x�6��������Y�a�
9��Oh�jj '��q,rR	�fgD~\�&����C4?mj��lo���M΄�5͛��i�MobF�(�
D�i�D�����M��s�P����{̂�9hs��.�G~ϗa�g�'!����E+�S�l��=r���NUF.�Լ<��ɀesԹ�NA�0�,34ӎ���hj�:5b���z�A�����yqoՠY=(�m�I��+�(Y)��:��7/�68wr��U�lڼ~�3�7�|z��6ڳ��ލ�o�rv�sO\>������ʅ'�^Y}��o��鍗6�vm��W��>��;>|g�����>7����-'l�<��g�>�m�s[Z�f霆�s��M+�����ֺ�����Ԉ�M�ڌ���K�|���i�����s�`~�����0[P�<;J��TP�uQ�z	Y����=�=w���S~a֪�+���x���>^w���o}{�o�]�t�񷧭;ؼ`c�C�V�\[1mM��'�&�����a�ڡ�U�6ώ���Orw�ʓ*Œstr%.��ҥY)y�\�V"�5j7CF�|��+w3Un�+��Z7��A�<���k���օ���aL�)6"���Ձ�D����!?X8ȣa���)t�ENr�����w45A�/4 0HD�T�F���p�P�Ԁ�rr���,��:R�$4
D!��s�ES��ʒgd�MM�"+E��K2���W��BtY�J��2�'Fv��1��Mh�Ԉ��M��ޒ[V▩���%�"LW�9nj�~<cv�`�N���d��%9Ҽl�4�Ǧ�@"����ⱚ��f@�׀� k4Z'8��M��$#0�z}&�'�R%��/��M�L"�Y�����5*��MU���V����[�&�	��-�	�_L�K�����J>���-VsGS#fj~�� Gă���yl|���j��/Z�^>�tq�`jC\���1?Ox8�N�v����^K\��|%����Xmyy}u �Y�F����Hk{��;u��[o������w�����x��ׯ]�|���v�\����&N�4n��)�'�M�04PW[][YU+�3��*#�0x�@C���=N���4��0�Ҡ���2�^*�%y�Zb�E��Kv�`�F���6��+,L��#	M�����*��M��f~V�e~�kɸТ�������&�P����\�Ccm�Y1��Ƭ/0C�����Ҫ,J�ɨ�Aہ+�OeC�`ڠ!�Ɗ��x3�aG1��p4	�_�U��	�I1�m����n(���`�i�E\O�i��<T�O�2��$x��ߜf��F�zAӈ�fF;��V�}UTo%�WA z���2���k
QQ���C�LyVF^jZ��1#�9vt��c cG����NO�OO������yNJ����,N����?|��'�~��{<���J��	���7qJGO?ř}�\�����'IK��OM�����槥�ed�f�dg�ee�e��&�%�;f�}icFbZU��^�5�[�����=j�p�E�P0����7�ޒ�QaJ�P� �/�K��Q�+�����0�V�l�D6��'h$+'|�e$g��ö�c�56i�褱ɣ2��MO�'-��1������9�)I��`��h�(�`M:� [��X�^@�B���k6 $h$�M�fKei���y�������Ԝ������Q��ܛ���Fd-sg�4��P���짦��i>b������9~|���C����̣afU�^����<��ԮD�²��L�0$}L'Y�����=#��ߔ����}8�`�/n����;]��Sx�ƞ%o75o3�{�Gf�2i2��7��5��d�g��{��-c�5���d����N����B�/ �S-���T�}�G?�b7��-~CG|�'?4P� ���aĔ�G(�)aLh�/h؂]p��P��xKz��E�c�[�}��_|%dj���n��?�����ϋ������Ι�j���P��<�)�tJ�]4�u�e-{QM�V�Ge��
�L]�-W��w���������j���q�����S$/֣9f�������x����mj�$`?B ek �iu;ڝ8��H���b�fU��bj 3��Y���j��Y�h^��Z��Ze���N�Ă��V�Q���IXHs��7�x������aMF��¸�B�0$%��20b%7Cٌ�>[K�����36A�_f�R_8��xJs�@�����Vbi�p�cC��Xꭊx
�'ǘ@��h�(􃩁DY��I"Oq��r74�ι�7��'x��ה[uj��[	�a�F�����C}?���D�f��m�F�4��yjA���zO����8��Ʌ�O�_�eIu"8��5������S#h����Ih�[���;o~��;�x�����/?~��w_�p��]�z��-kf=�i��k����b����WTm_ѰuEۢ�Ќ�Pg���I0�R��W(%���p��k�q�x����a��n��rG��H��������������:�\S�R[Z_�)WD�eE^@i��8�,�9���f��8q_
֩o4? h|l0�S1	�q���Ԡ����Z3�]XW!7���TO)VO��DDS3�L/���k�fj�vbW�%��fnI�yY�uE��x��45O��v�{_�p�/v��N��K�/֖]�+�\_)��k��5�u����q��NP1M���5M��܊�@�v^+L�:�B������mz��y�r^F�'4�>�M�� Ӭ��7�+���v�u���AvD��b�5�)��P�&��5r���0��g���mT�Ԁ��~c�fj^�mo�o��o[\o��oos��X�k��*�^C�W�5X�%�	��!�"�]���_?Ԉ��0������Gv�P�#r�E^q?�Q��2��4�� h�f#��]�<��q'B�seE��J�v4�2�빲���R3:�N�T���,:�S�,S�3j~�4�A�:��i3)xe))-嵝1�܁�%S{gu/[<{��o^�u��=g�:l��#�/�x��K�_����s�/�Zu��c'�<z��#G.����][�߳����~��so����k[^�8﹧�mY7�����/�S{���ų�iy`A͜)U3&�N�P;q�~BoyK��g�9��!Ә�V���xp���x8m���<�(?Ÿ1ކ���#���31�)霺��fo8>w�����L]st�S��<={�[/.�~y��K�}w��/=���g��y���Nm:�h�+�k��=1a����NZwv�'>طlw=�i��xe����E��)�H��WI2�jU�R��40��h��cd
�l�I�{�
^�ES�腛<pK�[�懈M��h��^�څW�0�c��>Ȃ!��Ok V�!ThA�6�Ў9p@�۱���L�	x� 4ăZ��w(������q���#�	Z(�0g
�CѰ���(q�*���fis�5�Y��LEz�,#M��"���I�$FH2*�Ds�k+�+��r���*�;����; t@����=P���hD+��
�����W��/%uj�J��eΖ��*�:H�V���ϔ�fd�[/ȕJ��]$�
2��pD�(�9P�/J#\DM��P	N^6���K��%����[�&
õJ�$7/?;G����HB]����	�Ѩ-s�?�� �BB-[�NMw�0#�/�Do�j��d͏e'/h�/h�.l���&�I(��d8�� 	e���z��+�./_r�@��C�-�c>rP���Md�+E:y��lu��t�R�L�A���i�h6Ec�eU�5�s�a��.�{���>��?z�7_�{�>�vݪ��&65�zz;�ڛ �M���/�Ѐ;�:].��pv���p��i������q�\���<�:/WW�Ck�.B[h��=D[��*fS�׵����Ft4b���bx\	*dj*���&ff?��<��2��>��9�ݽ��hA_ьV_��5B��J�!f�8��R;P�Q�C+��a�
���M(=�ʅ+l�P�7�rm����U ��҅�܄�Cj�w�
7)K�"�/+�8�� /�	�ISd����r7R���xc�l�M�9(]�P����J��j��j�Z�Fk|ғ0�iN�yV�qv�qx���zjj-1��\��Ӄud_5�W�������`7���"+�(��	e�<35{lr�蔔Q�ic�ǎ3vtrژ�̔��TIv�,3Y��T�IF$��F45��ݍ�?y�����S�Є��\�`����{�PCG�p�.O�����W������Z�����"����ܜ��0*%}����M�_p"+ڛ˃�1WK��Zl�(6wG��(�%�O�����Q�)F��ձqQtb� L�b`;���X����	l_�家�@Y��u)�H��r�S�d�w�{�sψ�I��&%�����_0&'oTV�؜��|i�T�/U��TIcS��{22Gd�䪵2�Fu$�Q C>[�L�)P��� c�3�S�RsES�567}TV�茌1�̼�����#r�L���,=!�7���Ĥ��� 1ŏ�5�� 17$jf{��� �@�|,@=�!�8��&dcX��WA�G�G`٣��H���`�Z�� w[A�	������Gx��q��j���g4��i�u��<O��P곴��8�)�Sz�HG}bda6��b���*N}����G��� k~��e�~C1�!��,���`~�1��1����pS��PO~џ��g�a���0�_��_P�W� ������!��Y�30��ԅx�Jc�̓�n~����|'�~�������|�՛���M��1�ja�5_ls�ꘁ;���i�sj�������O�����P�+���%�W}�#}'OR�)�=��B�1�-��^���hj�3¼���Ԁ�x\ov�f���ny�ƞ�P;㳟6[V������8�������Y�ͮ"��P�ki��,�L��V��ߴZwg�T�&#f�M�x��+���M��g9��i�(��M��#A1S봐V��t4�	�NQEvK��R�7Fl�Q�����C�+�9��W&5D��z�����o���+�|E�T��]F��6�#�!DM�c Ea� (�GJ�&���l?'멶/W���hI8��M!a�Ԉ�&���25��Y73"��D��Ǧ&�{G�@�Ӌ�.F��,���-S��455�x���|��'���>|��_�t���=[j�쭫g=���'S�WS�sy��׊��sj�*��i*�<��L��Ѩ��|*@�H��0���[ˁ��轅|�h�S�Ԗv6Uu5Ww4V�7T ���ʋ*���Hi��8p<N��b�h
�1H'�r��;A���L;��!9� k��Gj���ցt�١;��^��V��-S�"�|��k~�Ԉ�aЋy1V���.��G�Ys7S���+��]�����#EΓQߙ����إ��KuWk+�W�_�Ů#�xC/Y]/2���05��I��:X�5�s슞 �G�38u���͗,�kV�U�~�^6�g5�Q�_�?�ƞS�{T�A5|D��ȓu�@���5�I-~Z��&k9.�&dM�Ԉ\0�b��"D���cj�49�2��M��&c}��������2D�d�^�\�� Qӈ�����m�S��"�}4���w�~>��/۹�����_���/٨��v/�f��v���\Y����k��/���m�8�ۈY�z*��e�f��D]���[�&΀�㬆�~�d4�ӣnɚ^��âi6k*Ye	���,��5{bϚ��v��x���g�t��c�W?�y�sOMX��o����3k�O,��_���h�5��K��0� W ���v�ʨ��*���o/��S5e�~�Į�g�M�P>�U��V;�U���- $�z�r�Z45X�U.T�4V��P���O�N�dFl�<�C��,޾b���?���W�zo�o.��ւ�_�����g�N���Ц�}�O��;5�}�Ow>q������םz��i;_����I[^���j���<޸hoݼ��=r�{�k�=K��U�[R>��i������Fy�0���C�f���;�27%N}�t�k��F�-M� ��i�f%L�rB��b��N_��C�6Hi ~ZduAN_d��W
�X��Z�l&��$|�MMȂ��0�+@�",A�b�6 ?&b#��t(>g
�7�^wP��sz�V �|}^�.7G����Ȑ���2R�����1��1�4�K�&C�o��ʌ�ƾr���B�Q=�6M�(Is����*��
N(H�C��q%��W����b����S�j-qUMEN�B��^)L}�ː�d$;C��3�����|�\)j��s��J�Z��:��p_�Uk�L��SiĀ��3�^�Idj�R�R�����ΏZ�r�0���	7��]�O��5]!]w�.D{#xOT�H
`(�j�j�V��'kf7:nɚf��f�hj�X�hj$���c ���5��p�m<:.�`�8W��/������J'6��L�v�3�6�Z�%uZ��I �:p
&Q�� AzA���<���
��m]���|�ȱ�/��t�ܩ�ǎ�8�k��+W=2w��ں�@�����H4��B*�l]p��'< �W�[�}��Q=�S�*I�D��+�����2:�����r7�\�tF��0�0��!C�]d��iD@[\�{b>�
�ZG������Mk�g������u���t�'�[�G���h*��\lG
�z�t�����Y��w�2pl�p�Q�i6d�Q��P�	���$ +$��Sƕ��C)Es	M<\�ׄ�ڰQ]l����2��Ƈ4���"�#����=%lo��-�����
nb�yJ�mF�mF�yf����:緉��g7������L���ՑSk�ɵ��nb3���@��1�0����6��Z6"�V������::-#93=9%-nm@;;5?7]����N�g%�
��y���F��������o�{��˯n��lY]����Z����;;�׵u@S���4c�r��
F��f��奤���f��d�'LMfj��{��$%i
2�F�&��.l)q��1[g��Sl�2Qr��/����K�E@oư���@��RFO�&��G��rSG�����Q�)���T*E���1#SG�H1:utj���QY9#sr�H$�
F���/H-�fH��2e�\���5V�����1��Q%��3nuO��dꂥ�u��ɩBh5ʌN��L��O͕fH�3
���2Fgg���J����=jL����I�������k��AzB�������d>ՇM�b¤� 17����s=�?�,�?�%V;�Vt=�'�k�*��Q��1T��P?�Vj
6(%O����+8�3�>�C����Ov�9ӷ�;�����K��.��Ӥ�*;�ȯS��xJ�%l���j��������6ǟ,�?��h��3wkԯi�W�[��Ɂ-���K��L}	����O��':�#-��6�i���n��0DY�7&�pS���C�)j� f�E�kyB_ii�y���/���ﾻ���v�����7߾~�¡�ڱ��i3��J_�D��Tճ�T�`�WR���
?����+����m_���������u�7_��gH�$F��'E�	�cS#h�=F�'�xy�d�O���g�%�Nr�S��0E`�=�����l��W�L�XS#V��[M�ղ�L��}Sj��E�
�a�^��F�Ҍ�,bc)+�9ǚ�Mo�O��!QC�H��Y���`lh�	+E��Ơ��8�
W��
�� V�Fbf�!`�.�u�yA'���QWh��1/S�a�v�a�LB�	����M���A��uRT�+S��|���ĺ�����+�UiDDk�7�ɚG���Q�1P#�q��4O/�xjA���J��O��'��S��.�W}e��m����Φ��׮�x��s�_��ئ�3����������Ԕl[����25�o}���e�L��9P6�VR_�(��6p�|$p��h�}(�Р�D�<�8�12��NG��(��jb��5��=�]m����P^_]\U.� e�~p�X�/Z�/
�|.��g�G�kDM#��~��iP��&z�8��!�j�N\�%4����jhP����ZfN2��0=>*��55?F�vA� k���h�%L�n�f]���ߎF���1�"��"ϩb����5%��y��򕲲W�J�F^ux��s()֩MBӈ�F�5�3:�\���}��N�f�U��"�_20��qF��T`�5�q�9��`�L���S  p䤎eM��0qZ���c�~�Ԉ��X�&Lh��+(}7S�*o}�h{�d�m���W(�ˤ�L_��ku�@^���ZpE�
0�O���$v��ejR�F45`��p�5\�P�����?��?�Z_��I���S�ƓAׅ��զ��]M�z[�6�o�8q��[�I�|��eC�[��ej ��8��V�&�i�S�n3)�l�:����T��	M%˦�?�h�c+�_�|��gϝ��YmY��A�C��C���B)8\J��T����uVZe�*c`)��|B�	)@Cc&Q��:��~We�_WZ��Q�Z�.�8��`E�[@4� ���A�@
��!j�q"*���yX(��&��h�v7������r�'?����O��>Q�lOӪ�-�o}�x��G:ܾ����W�m�ֿ�J����O��9ݶ�l��W O^��|��闺6�Թ�Z��KM�_ly�B�#�:97���އO����}�߱��<��8��}z��5RX�Z���i�xIki[���,qbe.�ܩ�t��<�F���chu����i���~��O6��e�*,P��Pl�"�>�hC�F$�j�LP�9�.�"��k�v�ဠXP�x��g��]p�``�1D-BI�b+�aw�؆مr6�����$���P�i�!?O�����T���3S%i��F�2G��t3*djJ]h[�����[��V�=eXW���X���X�������{���3 q�'0��/��K��co�����V�	��n�B0�B����^���������cSW&*��i���W��F��X���ԔǪ��K��E���f72,��+���($Ra�n���fj<���%v�څ�9�x�ڼ�.�@g0.k
�"L\�I�Ԉ�F�V3��̨��X��n��o��o��8V����$���C�A1q�#|��=�q����CK�������L�d�@rZ+%42T)�2X� �a���x��2I~A^^^nn�L!/�Jd*%k2z~���M�6iێ-G��ۿk�6nZ;e�PcSm0���'`��9�m�%)Ԡׂ{��Z� �թԨi z� �0��J�� W������#��T�f���AjC&�̉7��"��oA�A][H�Ux�����菗��P��ņI��*i2�ldͬf���F��6`r�qB3XMw��M�P]�h(�5�̅��!^`n���ȃ�l�X����J/�=�c� �z	�f��!��;����| ��R⥤"�n����*4i�V}��:�]W��PCi��%TO9�_͏�6N�7O�3M��'��S�����-�9�6��,Di�9D�ZY�b��.�!�����)uشvR3���D*�qU�P�qR��=�5�M�v��5��܌�i)c22Rs2S2�Ǧ����L��J��d(s2TYi��Y~�6/Ks_R
G[?������o�����8s��ƭ�Kj�4(�c'��{�����@��* %'/�@::%�V��4�N��L�������f?�ef���H*�ڂ��k�:zjB`��Z�h+�u�L=�\|~"~���w�NPx��A{J�b ��o��TIM�5N�6�����2s[���6�X��$i����8�cSs�3�Rr����|�=9yIi�I�IY�Iٹ�f�ޛ��'3g�Z�����9$��Sh��T�o�{����KWo
U7)>�@ܓ�~�����,InF~VJ^�؜��̱�)��N�w�t�H��hƘB\������ =! h����&���>0#���s��4ǭ��1,
�˃��n|�]g��Һu�z5�Xe�=���Ĕ	S�I%}*?oW���.�g���_��?q��$��|k7�������3��$!;
坂
��w9R45�X-����������G���V�͎?���c5 ��|K��R�_�7(�Ba >3�	S���@3_��/	�s��a��?�֯�~EY~A��m��-�Oa��0�az��O�[��7����կn���7���S�ɍ���K��ɽ��}�/��|1\v�[�9Ku�Oh��:�����$/��J\�r��s0s�6]3;.�Ɨm�k�On����\�9���	;�	N�9e@�NSs�7��F�5w15"����`j��F�0��3�/�Y1S#���*�K*����+������*bv%>���[g�Sg���X�n	A'�K,�����F@�p�x��l5�LF�[)� c>0���3n�)
`H�^J���,��O�vw1����p�U4)}��K
y���W{M��C�<T��(t�>�P5�H�Y�@����N �C�M
�a�A��k�:y�^����-��&5Lo,�Χ����5k�㢩IȚT�&�iDS�av�(eD/3��l����vf8?����Ԉ�&�f?��ʕ�x�w?���G�o]=kדs�����nj♚[�f��ꅓ�Ե7��kb���� �"%0|6DA#:�B�[a��P��zl�"OCM���~|`�����A�5�����PEIP�5%E�X$��g��C��D�/��cM�㢦��F���fd�i�'�s�J?.+�T�n�/�ͮ���pB�L�9��ӝ�F��Q�똅��f��6q�65k[=���U��s,�+t/򜫈���	�������++߈U�ST�;��q���"��ݭ��pM���5���y%8��k�:5Q�N�&�3�?#�O��O�C'��	-y��5(��1tL�2��P��
�&.k�i挒8� ���
���Φ�L��X��8
������x��
�p�:�]����� \��/j0��ZpI�\֣�����C�;�9D�{Yq���2B�Y���m�e��O~קn�n�+��ۍ������T��bu�]�o��~u\�κ�a�c�5�J�!���|7S3����3h��x4��1�e��35�Fe�M_o�W�MA�̞�U�fl|����L}`Ѥq�uEaA���i���2� W�����U�k�2�J�i�$���+�K�JMhu�3&���Z�v��XX�(�d�BC�b�ڍ.;8Y��F ܐ'�JM�V�@�|R'5�6D�B�a�v�:79��d*2��&��:����*�8�x��Ǐ�=|�}�ٚէZ��ڼ�R��K�+��?v�m����ޜ��@�����/ׯ�h�p�e��-/�oy�u�+͛^�_s����KO/<Qz���%'��wU��[6}[�к��G�m����u
K;b�F�+�<V��5��v���d��9�rT��W��u]�n���-Ț� �{��O�{�Ve�*,X�GyC�3�BV'`4 �� ʚ��9���(rR�R�5	YsgScE���g��B��hMc#�6&d�}F�͢.��N�!UrL.�%���g����K�W�>��[IȨ�9�25\�W�wǠ�}O�!�iDS#j��05`8P���1}1�/��A��Dw11��(e�KM}��*oG��6l)��
��Ԉ�IA�hjDM�jҨ�*�hj���|�	Sc�_ �a�_���D1� ��B45��e��K��S��r��~��a!��҇yC��v��.��ehqkۼ�N����	��Hw!�U$�T�/&��O	S3���\�O���&k_�d��dM�1V#ʚ?�5?�4w75�G�U񅢖����/�-�P�m�A^�kpy.*�3�W|W�����50�_�����$;?O�QS�Ӕ�akl��8�����N�߰���	t-\n���B�� �� �ܹ8le�b�I��h����v�pP���r�d9�L�";Q�[Pu�$�:?�RH��ma�-(Ț�M�Jh h'�
F��+���8	hF=7����l�Z��l5�n��l7tZ�������JK�w\C l�K��~�ئ�% f�G��B�*�+�6b��(�������T��Ln�r�H��s��R�eV��6p�P����A���o��������*�{*��j~��4Tg��`��h����b��l��b�����6˼v�����U�5�測�f5�	S3���BMn����q�ظj||55Tk�����Z��bg� u�4+5'59/=� =5KH֌�LO��NW�f�s24Y�ڌTu~�!/[�=���ï���Ͽ����}����W�l���!h�b}��s�M�����Hj�J����+�������$��OK�MI�NMւ���ro���V���[W��%fo�Yۋ����(+������V�a@�4z��_������2_�O�L��*zx>kM�l_�Ufn.��U�[�"�	E5b12��Q��LO��4&=)=')=;)9-)3;)'/�@z�D~_���<�|��"�h�Xc<�bGФ\�(|�J��{��ϝ����}�s;JkPg S	����ҌԜ�cFg��/����#�Fd�N���JM6����S�0u��k����ԐL�a��(`��ꁧ{3=�l�0ǭ���"��ǝ���5�%�kQ�ZH�$_�Wb�դ�1H�J]�Y%�*���^B�o}��ֿ�m�a�����G��g���f��H�BjϢ�S��8&9��:�˽���a�Y�3����[���6�삦��實���j5�ԧ��7$�+\�5_�x���D��#?�S��Ϡ;���(��h��	��̟��/ ��3��>k9Gr�7��|a��/��������_n~����ֿ]8��v���뾙*dj�x���V��SZ�����ᮨh�%5y^����i�8�1�y��&�%�=�S��͝B�s$s�DN�9	�����q����$g>�܊������b5'��#FV05�L͖�Y���X�{q�(�����fF9:�
�S�fU`3��Y�ԬjnF�iz�s\���ǆx��ИQk,��Fa.��Z���as�Mv�h�X+ nj�4��$N� 0�$𸯉��i��I�B�f7�	�9��&Ti�b*E�2�*Ƞ�0�}&�����	=��~�0�A0�dh���M#�g+����u�43)o*wO�.��⿿ǛX�;AB��.k ��LMB�75�y���-�*E;��M����Y�� ��25�U���{�鵏ݡ���/]��ͫ�\:��3��tږ5�v=5���L���DES�}E���ٴ�屹M��߷xfO{c��2��;�
rA��1%(��M`�cB�8�!8����h��-ŅX_W��	�S�z�;{[�nGKucmIuy�hjJ������$�&��"�a��ZT�ٶ�$v���0�v��Q��X��>'��W�Ԡ�<1M��&E� �NM"D��҈��+
�+=��F<n �WG.�g�o2.k����fs�w��9v+t���b}�ƚWjߪ�y��潒��}�7����˔�\�)zD��/U�fjDNi��
�>�0P��h���=z�NXf���pN�H��
��J8�Ѡg40��' :��i�:���4�S:�?�"�)�sr����L�(k@{x�llj.#B͚;����e� �U/"�e�gu.���ZpE�.i`rA�\0�`�<����D��ļ���A���a��A{M�38h�Op�Ey�e����+��c��}'��;EꞃԻY��|.�����Ƀ_Ι���IW�wl�W؈Nj
&�
O�5?�� &��	VH�J�e�Idj:,����S���Ůy��͙�l���Bs�M`����{rr�͗���3!B��;&#/%+?#_��PJ�Z5�ȇ7RFe�Ҝ��9 fC����<�"Gk��ncs� D���L!MMO������HI��6J����da�|^/T}s�z�wc:/	yi$��a�TdrD,�Bkq�Q��4��i��%��>r����kϗ�9[��b��[�_kX}��3e���]}�qõ���۶�V��j��+�k/��:W��r���|�~�ku�^�^�J�C��٧��rLx���g�>4~}��'c�Vz�[g�[#�:���a��~c2����MD�+�#�N�ܩ�ej��V���|�0Y#��V?���"\w��Yȵ��� S�"jD�-1C�F}���Z�~�Q�!�@�Y�B�N4�$��T�E
�Ɓ�m��	Z���F��d m 8�O��b� ,�k�J��T ��1��R5!4�a+Yhc #�e����0��s:%�V�r	�����Rd�����$I��-�4h�;���l[)�S��Vҽ�xo)�[������O�iDDS�_%L��-%z��Y°��`˸�2s�#nj�u�����P�;�~nj���J�F�ւ#�������L8[	�t�Љ#)�]*
���w{J���M8}��
��V'���;����R�u1"����Y05�N���˚0�Y�v
u�1"�i�ʘ�f��MͬF�&�f�(k���M�k�˚;���V��[����=�A������K���&�yC��U.,�2Hs��ي�LYV��@*ϗ�W� O"�>�����Qkt9����t��X*j�W<��ࡽ.�ٸimsK���r�m����Uj���z�Z�S��R!D���h In�B"/�J&��R*S���`֤ʂ\yNfANzn^fn~f�,3���^2!1V�ś�T[!�V�������ш�v�EbQaaT)>���Q�ͪ4��~f#7���D��s�,�;�s�����m�:m�[�Ӻ"s� ӻ��|=���rsw������kCxu ������Zք����,� �.2��<��0o�Q
?#�"���f(s���KԅX�δ��{�<u������V��VG��6��6�v��v˼�.����6˜V��v��v�[���r4s[,�Z#`N;����H	���Z�Nn@'5���u�P1���P��X��y�J��n�	G52Uv�$-M��*IO�NM�H���������Rgg�23��i��<$/�wD�yn|��o���o~���o|r����_hm�H�ȇ�ҹs͙���w<Ip2�Z!���H�UFznF����R�SR�Ǝ�56{䘌�cҒ�S3�S�z_�׈4Ĝuac[LX�����Rlj�r]�;B�FP�щ�f����
���)�߄��)�B(����*���\Wlj��4{�F,�QhLZ֨���1I#��R2�*4�0���R�Ea��N�ӥu�`��G�%2�G*�szt�R\���]�]LY���z�ݣ��w���;7����	��ME%.���x��hP�����l��v��ˁӓ�̱aD������-S�G'�M�05S���.�L�n�G?ǭ]�3,	c�R��:�`j����`jVÊ'`�JL��^i��VK�Q+��ˏ*u�����?����t�t{��b����f�5���5Ty��ĤG�}��Ú����-
�A���W&�-���?Xo�~����������ha��oH�78����w��`j~��_Bd�`�_M�g�9�
�7@��I��/	h|�r��ǐ���B�/a��S�a������K%U߭�x��o~���_�������k��p|��v=��O�����.c�ܑ'3���	sA�]V�WT�j沆��&N��8�CO�+$w�6^@�30~�O��I�̙�k��������Ԝ4ZDS���wEMs��ESs��O���<������;<���Y\��ej���3���
�U��(C����K=��8���[b�p�nJeF�&Lo�a3�����H�mfp��۝`���V����jh��WqJ,r(p���-e	�H1��Q|�Q��$ɪ�{��I��{��TN%�Aj��@r�t�;���zW�S z���:�Z�A���ȭ@F �(N�jp��e��ib����9�-4��u�U\�IT6��I4DS��5��L��h�ƺ����h�^X�����UQ��`�f�U����V�~��ŏ޼���#��<���[W�ڽ����[�f����ٿ�o���w25{���;�W�W�.߾��m������Dv<�|�d�e�.��v����˚7,���Ĭ�K&u5W��>�L� 0��Q�ĩ��I�p �Fo�A8����h��P]:��:u������{��u��m�nkh�-�)�V���J#�Xa V��C��̱�Ai5au�;�8G�&��M���f����,!>���&פ�t����Ƣ�	���2�`P1QM�i���gU@�Eif�O�t���̫��ʪc��.��`j�\�Z��}��xv�8�F���
]g+�.Ԕ\i���T�zS���uoW׼_Q�V��M��e��
o�@��K��R��@.�A��9�6 N�Wt�%��9���i{���:��W�9&5�SbW��U=+̄�Qg������PJ8y`�I����Sz���>�%�ia���SN|���_5�	���\8��W�N��D�?�5��	����P�w��(�oi�����4���%*rA���z�<����3��$25"Gh�����}&l��oA����<r���w��	���:>��n��W��iB�S��EG\�s%�o��|�`�o\���y�MX�7.a�m�B5�T�2C��l�I'r��M�m�f������Dn����XTNC�QY�T0���sAw�ܮ���"pVct�Ҵ��I:E:
�tyz}Ah	B�c3�8��^K��0�ш�l��m��,~�@�:R��e)���8�q�yP�R&'�IMMN;r�Ȥ��dI�XU^*���r'��:?.���0D��#fg����¾�X��P��e�z?Z�dw�c'C�+Zu��ѳU�/׭�Z����WZ�|�{�;};�m���M/ul}�sۛ�O^�{�zӖWk7]�>r�t���׫V^-y�|dщ��c���;����{���ђ�kcV�Z�j&��
�n{���w[<V�h�/G�y��,�P�mp�]_��׻ͷ25Z�fj�|pg��.b�c��RK_�����U�7��z7Y��ʬP̤d�I����4 Ў�kh��,uS`sQ;�	Ղ�f����Q�F
���L��Pl�c60�D��ۈX��8a3�C�E� l"���6�"���(h���C�9�L�4�>D�nC�!#��Z"B��rv PF�R3���3�_���{�]W!T�W���S}%�X�A�5���J�r^45՞�rO}�����h��+��e~&s�g�K����B�"�S�Ԩ������������I$p�F�Me� (�b�eY�I���]�V���mQ0�u��郧p�(k���'+
��MM6�	��Sd��R��j;!T��*7Y���H�[�qY����:z!Sƺ�p�`	=�����e�_c5�ֹ������j ï.q~�hD��������L�L���9��]A�:/G��)����B�%� /'7'+���#Z3�$2�ؔd�F-djl��ꪇY~�����N?q�䩣k׭jko��y��͈b�E��v�j�P�F��(�Bug1�_�+aj���s���2y9��̼�����l��I3ҵ�ٔ� dĊ�h��h
Q�ET{��65b��5ܴ*fr=���V�̨�f5񳚍S��Y-��`N�ea�s�}^�cf��`l��g�?4�aŴ��S�3��&5�z+-%\[1�\D��
�������?�.h�F������.��A�ۉ2;\ᄫ=X}�j.�څ(���������j���Ќ��잒y}�}��}~��^ϼn��.׼.��N��^עn�N��vA��`j,�4���������'�����I����Zr��_�V�}�e����KZ�&7G��&MI)�L����>6339?+M������e�	��b�yȈ��x������w���_���><s���mϷ�v�GS�` 2uʜ�78��R�\���QJ���LYz�,-U��"M[0fL�Q�#G���<vtrVZꨤ��Ia+�Z���,�Qss�(���E4���a�E�jK�;a��a��8����r|IN�b�����
���i/3�D؆
wKc����R=�Wa��2���&������������q��������'5.X���C��n��	Oo����w>7e˶i[wT.�����n8{��W�����;������>���k7�Z��}p|uSGy]KIe}(\l����@0%����X��A��d:]�8/9��y��d�- ��z�K;ͭ����q���A+B�az��hDֳ�5�f�Z�(�P����ի���ꂝ*�^��F�>�����7���{��iw���GQ�����$?��?I��������/ ��	�
����4�ߘͿ����b����/�����7��3��澧�ߒ�o�78������|�J� >��C�0�%��3�@�� ����A���#�(jv��-_ Ə��Ǹ����s��7�/�y�囯�v�Ïn~��^>�����i�����7C������CO���R'��y}IM_Q�/���B�=�S*�����Z�
J�H��i�K��Μ��ˬ�6A8c �[�a�L� F'��4�r3�R��+��cw�G�F4�IR��9���<��'�fc̺��:�Ԉܲ6U��j�U��J0���?�THӔ��J�����lZ93��*�vFL%Ԏ���ʄA���D�������hf93ř ��a���K��������'YK<{�@��c!R��tM�(}�hT�n�I��y&���H���l��Jiy\M䰺@��@%��a[2�e����0�I��qt0�V�U�*RrS������)��ۜ���ڶ�ӱ�˹���@�P�&�Y��<��<��MMɚ�w�Ԉ�F䎦&ag~����U�㙚�������`jV	�f�C�WMxf��?*S�u�*Q��25�@؂�'7����7�y���C�wl~p������ܦY�o��{���OMڻyh��!1S#����l�߿�ٷ�k���m{׷�Y׼{mӮ5�/��{���V��ZygS��C�wd��
�gWT�vG�{�ݶ8�y^�����+*�=T��g�۱�e���Nxtn��撊��J�ʼl�B���@���_@'8q����=�c����:����ٹ��f�&N�����ok�oh���+-�-)���TE�C��h�(p٬E���ׁ-�"��4e�X h�$�2�F��l�������X;O����ԛ`��X�}���II%'i�H:�ʁ�x���T��T��R��V��^��Yi�]ͩ��V�	M�cS#&h��L(A�4S�n���f]�n{���p���6;��6�c��U.�Ԭ�����llunnrl�wn��?[�x�ض7b?W�X�R_z�����Wk*^�.����h�+��U���r��N��Q=|H�;e@�����9:�4�R�Oʅ� n�ZDX�I/Lv=a O���z����s����O�#:�ޯG��:☚8�c�Ȱ��Z�D	b�R�� ��#J�Q�pL�9���j��t'��S}bԥau��VT6����:���d_���J� .��=r� �om�9�6�V���3r� ��s� �����a 
���8z$�>7�����<��D�R�l�Q3y�C_� m@���ޱ�p:�r;?��?v�>�خ���2�V�vE��(�p��O�ι�d֧/|m��Ō~���9&�t�v�E?�SsG_�@,X3�b�h�'���fC�f��V�8�z���2)zl�ZR���wT�)� *��$��$C�hV���uN�!%�, trL#G�
D�"=Oaf||h��0�H����X����f�ye	`fq��q�h#	#5�"2�6W�� �bIA�$/S��!�NQ�$�����f��p��P��"�h��ɨ��e���t��K�j�����|�����V�<[s�t����*�_���r��k�뮵o~���W��^�X�k㵞�_���j���{�}���wny�s���������骅�Jg�l]r�n���qk#=�F;*lY꫙�.���|enG�c�,g����gB��R�0}�ց�;�F�䀚\�&��٭m�� �>=��o����DW)�cJ�q��rK[�k
�u~�҅�م�nE�L�,LYg-�����@̅;�b�c ����h���"+Rd��~
��[Xד�70R� �y(؆h8�����ي����1��Q�챸4|UYu�U�Z$�Wi�Pi_F�/�&�
��xU�4��IH��u��fb���J삃��Jf���3.��S_�_a,7TX�U9�ո��x�*=�ހ�1�A���͐f�奥�eJs�d�Y�TQ Ԏ�i�z�O�R*��F��2�X�4ą��	�����8��d4Y�����@��tF"����X,��f�x�a������g�B~Q�T2�R*Q��K����Y��<�\�kTFL0!e��C�x�F?�@�|�� ��׵���>}{��B�#x/���uj�˚)U���E��"5����d��Fζy���m���E�n��n��n�gjDY��@ ��q����^�}�������/zhB���"a�S!�e4�4]����͖�d��%39U�Κ�-��H�r��
���:@��Hr)H�Y�%��G[q���O^�v���l}����8V��{�F�@�A�P�"N[S(����+��}e���j�r����*�D������������)�ʐge�y�V�g�
�HV��F?����F��=���:�j@WH�05b[45bх.5�-MM����1��٩���f�`z3?����b��a��e�����-��?P�d\D`������PTO0�;<�#0��?��5TmWek�ۢ��B�[l[#Ǝ�����W�No�����]f�-5��x�2w1�_j�Pew5��7��3�+$>���������e�������y��q/�v-�t��@cA�0��:��&e��pՂ`a�И�&�~�m��L�&  U��j����Y�(����:�B��*qoF����9�2s��f��O%�LQK���ъ��N�ߓ��q�n������o����x�ة�KW<(��T������� DX�zF�!��XZ�vT�,))�{s�$KG��KJJK���%I��r����)II���JlK�]��ۣN���EX@G��Edg�*�zc�X0GlO(g ��n}������R�#F��5���YV�9H�f#����x�?6i|��ՋU-[Z��C��u�����8<���g�.:{t�����^Y��K�_{��7�x��7|���W^\v����/m|�-o������\{��˛_|i�ًY�c�#�l}詭��lX���Y����4���Jp����a\[mƻƁ '��aCnd��l7Lt&��<�~�n������q]��>��o�m7�Ak�g�{��y��133�Q�,[f�cffY,Yf��Bv�n������;G�(����+��>�9s5�]I�w>Pg�7�s���z�f+~�!;a��wIX[���(m����J���ғ7Ғv�S�2��i�*���.��\������j�O��j�/�_(���+\�uF�8�4����I���V�>�U���yW��D��������E�ߊ%�߉$��E�b�D� ?�	�DĿ�O���a�p%Z���M4�|�|�~�ÿ� ������|���1��'|ȟ�}A>�O�#��-��5�������~��k�<�1���K�/����_�X�Ӎ���~(�}��.*"�G��7�m&v�*�EC `r�ʻN%��G�� &YAtK<�#��Ec�+�hX| ��gx�����_a	.��k� *Jp� �ˇ%�k�L�UT��(,�`�K���HrE,%�J�($�)��;d��ls����Z��'(Y�t�+�"@�_�û3e�2� hj�l�_��ç�}(d��?��#�
 ����{�Π�6]�c��b�?a�q&gs�|.ػ��"�\E��F%���2	��P$Y\	�0%*��R�T�KdD��K�\����<r�4���M��Rr����еB�R@�#t����a��$=�M#��l�ˠ
X,�G�+ ���}������a��qZ�pv����3f[D���m�*��+M�ˍKK���t`�]Sk�2D5Mo��Xv!��k��-���m����ɦ��V����mO�4����m�M�V0�9/}�b?�y"P�׀�c�R{�L�����C�����Ƭ�t��ܳ"��'r�7�`o������J�l 4ͱ�UG7�FM�iojؿ�a߆���:m�t���;{��\{t׺�;7<kL��1ej����Go��������W��ػ��օG�/8�k��g�����z�Ŗ�4M��\�]{iO���Հ���M͚���{#�q�'�DN��d���
��n��U��+�V�O����;���얹;�74�y|z9�+�NK����>�bv<b����,hjDT!�ӽ-�um��%�u��e�M�5�E�E�9��p�7������n�v�4[t*5���^ � $��Ha_pY���(dr�Ɇ�F��iR�L��bz	�FY
U�#+��
N���j��A	9[�Z��UX�nV����e��m@�Ԅ����=�J��yO+
�݅
hjzK���T����	��L��D��H�7Os0K{4�9�מ�ЌF��#�[��{���3���"�WB�W<��F�u�zL.�E<�U{�# Bi(�c��#����Qk�L�0���=��2�� C0��`��	2Ac_�s��0�E���|���[r5Mx�*�$	'R�t�8!���Y�tl��+S�O�_�hP�DM}��a����i`]a ���@tCMC �$_x�#�d�cL0�P�Ğ����T��3��B��Ao�O�j��h�k8zM$�"�.+E�բ�j�
�P�^RHޒ������'&��V�+*���C4�I��zv���]�Y�Fwכ+羶��W!X#l2H���bF��֮`�ɿ⿔5Jv���&�CY}�AE�Wӊ��RiZ��=��M*���X)��F��8 NI�RR���I���*�IW���P�\�*��J&V��29.S��*�Z#��R�R�T�����O ����q��NH%�dpXN�?��Y/��<O��'y���ᤙ�MH���� L�!E�U
�X��5:m��[Vи�|�����ll�o�캝������]��n��7�{�ѷV_���҇��[r���N��v���#w��)�:R�e�t�p����˹��d/8�ܟӹ/ܰ�S�&�pUFa�'�3s�����(t��&�ͤ6�C���$"�͐ 9��Ds�h�����5�|=3�@�32�ML��MQ�.���>"y�. /'�i�϶"� l�ͤ􂩌$%0��� ��� �N���=Z��q v)�!��r�)�T<���WB�%sl��hE�%V".
n�U��XJEBM�H�������ϱ� L�Iؓ��jV�[Z�5�-AY�o� �^A�m����� &�4�h�baG��-"j	a�
���E��01O���Ƌ�o �����Au]H�14���A]�OoW
��KJ�%�N�5#�I3f��%��I%%�()d�I�ur�l�A�>�Ԁ�0��d�����q\"�@S���222�v{��B����Ԥ��RR�SgǓ�Xi�N�	���k����L�0όZ�fn��Sja���*�r��H��v�Dg����j������Φf����֦�}�05՚�*Mo��#�ջ��|K*�M9�\��,f����3(�qiqsfΎ{~F��ĥ&ΙJ{Dr��:��H)|6����4��{�ݟ�qs���ޛ�L�p�t�yj"��� �F���AMC�V=���>���dMrRBb����3Rf�L�5�4k'9ID'Y�|��������̈́�)��M�R�3���,�%o�����:d��E��dA�zQ� &K*�K�6��B(�:������jǚf��ѿ����ֳ�ҵ�̾��^���k+�2��ܯ�
i����SS�����Y��;���ƶck��%S�Q�ek���͋�l�����ip�ti�eIxj]��Zn}�ye��0,/?<:(h�)@��b5�PB���K0�fi�
�.(���O�y�ҎiG��=[Ҟ-j�"�Vs��(U����6��b	��a��Ri/����7��������=��璞'�ı�^�������{rB�0>�Pe��}�7���o������~�ǡ�;WF'w:^R�$�ۤ:����T�b`:�PK���Dϧ�����̿y�����{s����8�{�{����=���<���w���mʲ(�<�b��8�j���ƍ ��=�����|06$������:��}����>q���D�*#]e0I�F��e0�Ë��7��ܶ��Ћ�g�w\�0wh���;+^�������Y���Uo��y�Ϊ7�uݻ�y����_Y���/�����%wn/�q��ΝM�>��്w�m�q{�ͻ�o��4:vpbr����W��ru�s����۳o�ھ�������`Fa�5�,/4I*��
#
MM��תᴪX�v���`bW�&f��V��uih+u�&��Mqƪ8��b��Bz�����������������t��z��:JI{���G��R>�jZ-��V���Q+~��}(Bp��L�$�>Φ��ȣl�->�%��:��P�����^���W2�oĒ�I��K �Ä��
�A��c1S ����)��	��K �?�a�����0��\�'�c.�tS3�i���ėL�>~�I'���&�/|�o�Ã/><~���m����pۦw,�we��ll<�y�ľ�����2Q����ܠp'��:��'������&ް�Alȧ��!�Ww4��)�� LM?��a��� "B%�B�F�"�&
�B�T|y���4�%��DzE*�$�\VJ�)��*�-v�"��nu�ץ���$�����W�E^�;jj�G��5!�h�[����(`���
�z����
��x�O��SU�ej�6M�d��\1�x<�7UHp�}�h�O%WJE ����"!x�A������B%��͞M�3˕j!�KT(*�T2+%�.�q3H3���4���?m���,�Q
���dK*`�yt�CGX>�ġ��4�J�ӣ����>��.�IKM�IIx^�IU����T����ܾ�ܼ��F�X���x�$jj�T���/:�>�\�6ڷ;&k�lj�U�@S�nj�-	<��S��ڿ:����Ckr��;�[ph]�#SSstS���MG7���|xc���O15�5���L͇���{�|��+o��z�����v.9�k���s��l;���ԋMg�4���p~wÅ]Qv��Ϛ��0��k����M��+'zC��FN���������9�Wr`y���w-���\��v(E*!e1��!����6Rp5x35l6��b#l��ŵ댥9�5�e�E��%倆��Hv�/N���>�+�氛-��H �q�u*5cSJePӨ�
�RF�LF�R�P(�&[�Vj5*�Z�WɢB�Qa,%��T����i�iV���d)y*R��Rm�է�[�L�i���L�?�4+
�.��Ԭ.QCS��L���`C�nc�>fj�.��]%����򵇲u��ړ�9�n h�o��oG<�2�Լ<�e��v޳Yn�74�	�|HHԊ��L��=Da�P���B£$� �6@�_��hl�;�����O�uD��G8IGn0��ʹ�]���3�K��x�H~3Mr�LTG���A
�(�Ft��#k�D}��Fj�:PcjF�q&�1S��h�i���o��<�h	&X�q&�c ve�����h�A&��}�Á�f��B�*���~�%��� ���"�_%���.jD�T��
�TI��Doʤ��u?5���������@�8��|��>���̋|�=�uK^_���wz�n��6���Z�\$�CDn�u(Y튯h�Ң$hV�r�`T��Ӫ��y�
N�5�F5�AC��ҫT�:�Z���R��ٮ��l������������l��CW��*C-`k1� �F���>�����_$L.Ĥ`��8X�j
�Ab�s0�L!'�IIj*�Ig��T;�DM!SR�R���f�z>~�s�9����$�S���BScA)1S�V�Mb�F�6�C������fٞ��V��[w.w�բ]cᵗ�6o)�2Z��z׋wh��{n/�sc����;��v6��o�10�ŉ�{o��zǶ�ƾK5+��v�lXy2�qK�j����W�4P��_�ԛ��lv��l�t�ҬW2�^,7��v�W�l�5�LM4�扦���+uLU���}����
����#+t��x�]�c� -ϯ��5|5�j�#0�~#/�k �j�K�u�86	`�����oWq�*�_�S���a�UD�o��P�J�C&0c\�~Z�,������>�^Q�t��;b�W��~YcH����4y�M^B�|S� �3�m"+J�i �aa��4�zZ�'dMm@R�V��Au}H�
hK�:�U
�|j"=1.m�̘�I��LJ �I4��	C0〵����nj`�X��z�`u�E*�J*��d2�D&�����z����6�훦��b=��a��y4
8�Z<p"[$Yf,߂Z�Ϗ��������,	+�Xu:
M�VM�5maYG�b*�)��\�w���.k`45�ڀ�BS��F���֘�ݏLSc�0�91S�8+.~Ƭh(�Rr9% MҜY�c�Τ�P[�a��,&�mظ��K7n�{����#�G�������J�<���[ ��������,Gh4��N�>��W�݁-ا�29-%9>!~V��D�!kf0��qZ�Y�sJ��$?�(ȷ���=�Ly���� Ҕ)l��ZsDm�☦��&VCL�iW�`VQ�Ԭ��v�:���k�o�o� �Z�k����+������B{C��.� hʳt���Uxڋ�s�3�ԅ���W��h�Z\\P�YV�]Z�^\f_Tj��
�j��ڌ�Z��FϚf���t�O/�2w��z�+kM�]i���hb��k���������e�jVe`~�d~��+O�̕-�sD��xK6ޜ-�,17ڂv�?	���/$�����П��ĨC����%~�o���y�s	M`O�iI#��/�X�ୟ����������7޻|��}[M�|����^�Ү�ȕ�3qK3EPC���	�s��d�n6IB��$�X�dr�))L���s��K���e%��h��nc�M]��=����G�8�i`�`���Kr�xȅ�e.���P��\��e�ڊ-���l;�������_q��һ7݇L.~��◮/~y|��7�n]o�u���͎[7;oMν99�����ɥ��W߽��޽�7W���_3:�vpp������\������g�n:v�o߾6��]�h^����y�EAG�C]m�V�F����o�q���5Фc�YzZ��^��6h�]*j���݈�J�9�'u��R�V�����WГ���t������$%��\�����^�>a�i��q�ڭ4�~�Q�\)�P���cܢ�n�(7��	}�C��n��Q�kB�۸�3���t����Q�+��A&��L��R���ߊ�_c�/Q����䛦 M�g,��L~��|�%��#���|ĉ����k>��DJG�[�6{�������D7Q�%�e���p����Y4�+�n�rW�|�'�I卧2oP�/q�W���l쉦l�'���4`�·�5�K��Ԁ�=���!��A]���*!�����d��L�L�,�H��45Gu�A��E�lk�t}�������Y��L�� S3p2]���DMMg:����L���
�$��a}�KR�<2N�IR�`
ylʗ���02P٨咘�L75r&�E,����d��ե3�r�B��0�����8iI���� �=�M��I~A@�-e���cd�]+1*p��H�
�/B���cR9tb��ө|&��AT��
�F<�AcP�RfҒfHx$��vny.ɳ���Gm��˚��5�S��� �]�3�Ĺ��{W��fZ�s�/��Z@���%G7V<S�_����������~���?��͗߼7>q���C��Zv|������zjO�=�gw7}�i�L͚��5���4ͷ��S}٧�d���>�6����Sk��,;�����U�&�W�B�@@�og�}0�2�A�������!,����Ә�,��F�+��J+jK��r��rs�L�?��c0Û��U��_�_���p��z�Q�����m&��h2���^��Z�R��:�ڨ՘�*�FiTʌ
�Q��p�'��k��O�#d���R�d)�ʴ"=��B�sӢ�fJ�<��yLӬ���'R���YM}ZSFh��2=`c)�4������9�����_�g�Y&�[ጻ�K� ��H�Հ��"���r�d���LHe�B|!j�1�b�c4.X  cd��4�52��5H���L�1�h�/�K�2�8"�_:��rķ8�,�,E�I��hr$9� 8'�:��,}���M_O#JՌ�`��ɚ(DٚA*0Dc�	FD���h�n�}��K ���㏙�.X��1F��汧�C��0X1S3�� ȈE"�PAL�\p�sY�8:���k��d�i�{Q����d�����/-�/��ϭ��l�WT���)���R~=;���O�/}cE�ˋ?\��H��ǩޠ��"i�bJ��ԥ�<��iQ�Z�%}aj��z=������r�d7yV:eN@@��ĉIIRZ��I%ދ`Q���4��%��2)&W�e
�X!���\�#l	K,`�,���(�Ġ �h�J*8o�I����=sN\
�O�œ��dZR)>1aNQ�?��<7e�����,(�.��FHu�Y��� �
�E"Չ�V�;,�j\V;SQצ��;K{���6�ح��W���s��m������>8|�݃g�|���o��1���|���T��Zѹ5�vm~�����@�r[�C�i4y��������ެN�p�����T��!�Ң�5"�VVk�M75S15�h@�ejʜ��dV���ĵDw$EE@Y�W�z��ҢtI�KZ��D�h؀�B@H��tXP+ꐰY� A� 0"~��o@>=��8��i1lV4��������c�ƭ"�����j>��A��q�V1׈����GӒ1�$u�:Cƈ7cԠ�_h��AES@F����FҘ�k <�4��ĤL{�x���
�/k`�HS������DXM}HW�V�5�m�,4��
�$���f��NL��DJ ��L\��$R�L"�(B�pV'�H�01SV"p�~�:��f�Ţ��֗E��錙�J�a(J�3��L�ўfj(�i�MiN"=9�CJ��F�7�"Vi�/�
��"��L��R�Uf�U8�r'^��j�h��k�����td*b���15P�|�X||
v�`︶F��ZK�������K+ӛr�yN�U�B�����9�Sg�%ΊK�='5��!�$RR����8'iNT�̙EJN 9*�j��	��7�y��w�N<x��������s���L�����8����b�l'�=��>�L&�_�$k�k`&TZjrJB\R��ԸY�(�6s&3!���p�S����&��2ej�̄�y����aj�4�y�J�&�� b�fY�yy�ey�mE����u�U�����������:ow�o~yFg��9�ڐc�%f�g,�	,��qyc��������������-�k���?����Ӑ���nj����5�tSeMl�MY�YV�,�Ѐ\�V���/��q��ɻr���2"5,�15����"sc�5ӥ�IB>�Lb̚Ez~&%�,L$�ITYS��Π�g1͉H��Q���#�b���a���{���?�����������d�����n9�pǉ�.7������_���p�.P�j��2��D�2*Z[��4
�C����,�� �K��:���Q��Ybj��F\�à������҃�yEyn<��\�]�tk��3ۻ畯Y�rx�3��O�r~�P�е�ѡ�����!@��@�صƱ����G�4�k�omin�_p}|��ز�+oLvO�u��\>0���՞sgW=����S�V<���e۶�_�ji��y����V��m6e�MVk5XPhjZ��%s����:*�ZK�WS�T�U�#v�"��P�ҋ�ʸ�0����#-�%-I�ݝ<kM��)s�Q�/SR�i���KD��S156���_��?������ �dQn�<B�\�3��y���"KD�����d������J՟��S(�(��^"�.���Q"�&FL� ~&��+���@�����: l�M���C������.k�����\�,�GL�{t�;t�t�U&���Dǹةd���I��m�r
[�8�Bo�7(܉4�M*��e��yZLL���f�Λ`��.�F&45�l45�L`�ɿƌ6�~djx؀@4����R 45S	P�����8�i���4�U���\zQ!>��N��G���d�[��#[����jjb5�xL�Ĉ9���|�<��+���b�9Yn�<�paH�8S������GT����M�M�=�OMLr�`� �\��D!�����Υ8*
��T�bt�D����gq�,`u�@S#�pC�g��D������|���<�B�P��Mʠ��6���U�0�$J	&FyP�5ajX���/!k�TX�Rf2SgKx$���iW�d���ԬzTu��!T��|�� ��:5{�j��D����J�<�*"��p_��y��
�-:���ئ������4��~�����[�'&��8sdӑ�ˎ�Yrb�<hj�ObjN���\�eͷ;���Q�㪬3�.l�:��b���[��l.���p�dz���q?�`o6O����tM�N<�Do3.�)�v�9��)�έ-��)�(�ʙNQN^i~aEQIcm]UYyANn$�gx<.��fwX�^w:x�x��i�YF�N���Z-�s:�Qo1h-z�E+7k$�H'ᩅthj4�QHu˘�
z��\���)U6�w���ihj��F�] �.�M�>Ej��Y_��Ta$�FE�e�����E�}�����Y�S!Å���4䷌�7C�w¾{�"��(U�}��x%������v�h��VOJd���MeF;a���t�(�s�̸Jf@S3�BF��q>>!�	$�|U��J��@6ȓ�%�L�0]q�&?C��+�3�g��KL��d��ЉD��4ݭ4�d*v�!�A�R�)��(��25�a*�+��`�1�ш"�B�FL>��o�0V}�"��3�?�
?cW�EP��&LP��QdH�c�!����cQQ�_Bx�5	֯�\T�G1�A.��|�C�+�ߒ˾0~n���3��=�\���]�Eg�A����>_��ݞyo-o��w��<m�Q��.P0[$�.�C��P�!mQZU��H�n�|E#��V%�@ō��դa5j�:F��V,N)��e���A��Ļ��*��Qr2JM��d��f��2���s�JqD��J1��s�r�V!Ы1�^�(�zo���ɮ*�G���'� r�ۮ�TJD�����|R
�)	ii3��͚5#!�r�,Z���YbZ��G2c4F���萲�baj�R�Db+\z{N���yI��M-�����;w�%{.�=:���{N������'�;�,���9M�R�Kʱ�Yӌ��"���R�]+���!�\�.�Z8L³�1�V���DT�L�&K��h��juP�p(�*�pq9W�Q���B��eH�� �dk���i9��'��b7VK���˪��
�P�%2�J3�%�y6�k��l�me�L�0�
@" lFB&AȄ�v->���`�%L��n3�2"wɡd9������V��Jf��;�z�<��P�ӕ|���pm"�c��,��)c$Kh�"J��6P��r��>���ꢇ�J�/��Á��1M��ʚ龦9�D��GM��.��O�XLM��x��w[�Le�$��̆�&eVB��dr"�Cg!�
"Y].�E(Xc`A���Ԕ�������$hj��`�۝N��dR���ȀG����'�!pQ$	�B��U:�o75��Դ�����iq	`[�LK�15�4�.ϵ�mX�?BEf&45�6"���!�e���H���{���@Y���G�0
ҕ�x֘ha 0�f:`˸�����{�j����*-�S���s�l2���HK�I�wd6Q�wNBZRb,�L��!��f��+���g3$��`�m2j�o��ҍ�w�_}pgtl���Cy�Y^�[,�Q��e�(
p;�������&���)�΀yl��1e�d҉��)	DB��53�qBJ�A�v��a��x���Zi�!��%��i`��W��O�dQ�vI���,�4�XVe����,.�,��-�r��vw�d VT�/���*u�ٛ���ن�cK����5�ҳ�6��ƿ���%u�����y}]���sֵF�6�����S�]���4��8W�ٗU��T��XQ5�i���@M�YSB�8}S� VTj��Dk+��FM}�["hSHP=ಔ�ن�t�C/�(�<.���N���OF��$}���%��K|,k��be��#�M����Y�wׯ;�����o�j���|������-9rm�����r��OO����Co,<0T��TU���u'*���9ܾ�|[ߩ��͚@�Ԟ,mͫ갸�2��QJP�B��rݺ<��0CY�.~������4 ��҃��l�0��eN�̕�+����]Բk������|z���yc��#�-���7&ZoN��o�i�j�ԏ_��>T71\7:X3|�n��et�cbd����룋'F�M�u_Y>:��ڕ�����/��_Y}����g�Ν�>rxپ��ܾp͚��66�4���eJl�b���*m�K��H��פ%�M6��D/�o��J��Z�!7�)�T���.#~�&��P�ҋ��&S�%L͢��˒gBSs��|��v�N~��T&�7���V��d���1��A��Jُ%�8������g���&45/���{"�/4�?Y-�������F�g�����S��U&���5��3N�&|""�k��%�)�	�1[  &\�hj>a=��L�5�p�%?cH���>�ߧߥ�oS�7�=���w-�~9�6JC�sD�4��3A�ߦ}HoP�7���L��$s�S��@Yv��)YC����=�4C� �{�ɇ���t0��4,��`2�0.��&��L�U\xT���4�ԜS�N(ѣ*���g��J�m���|_�������jo��D��M�����w�9mNV����d�����E��\k]��/�ȩ�̸�H3^ �"����hj�(�Q0*$8x
F��%���16�Kb�RX)d�P�1�g�ɜn2�4j�\jR�zU�E�}V�Ϭv�.�$� �0+3�*�MN�z������N)��PL�E8L�� X,>�EdaO�"�,i��ؤ98;Ū�����g55+������w���l�r휗��������EjSӗ{���5G6�>25��15��|���>��/>~��w���uSsd������3�������S}��M�ўБUA�t;�pO�po��59VE�=8ғw2�i�4ֶ�t�d����:�J�U�*"���`WD����x%�������|&[�b:�ʪ7F|���Қ����06T�4��AZ���k�J�B>�Ù�ty��`t��Y�pv8 Wl&�Yo0��&�l�-f��lr�v��aЂ_E�^i��Z!K��4��XD�������fv���Դ�XߡNt4�k�i,��'P������Ra�\n��"�D��X��P�7_35����p�:rE�|w#~����Ր�5��Uo���鮗lֻz��rR"��x�hT��@�Q:��5P�����1�p����O��	�j\�CՃ�U��2S~�����_E���aS���䥌��3j&0�x�p��>�8�$�H�ﲔ7��Q��+Y3�׌P�#�(�3NeM����7�q�]0�(�)�u���t�kb����Ca@)3���.�dEj��=AS�����5QD�A	~E����{�)iI'�)�B���Ncj>5~dP���0�TvR.�䲼�^��u�>Y�佞yo.j�Z�����"[.c-�p�ŤN-�YMM�j�Դ���넩iԲ��r�@L)�3�e쀀l�&j�	RZ*?-�2gfʬ�H	3�.���\�+�T����Jl��&���,+tU��k��Z��uV/_�ܻ�}ݚξ5ٍ�R��&��
�l�9�7��M��I\~2�1;!q���gEMM�,nj�����S�B�g�F�tJyv1��XbK�k�'���kɢ�K�n^޻g�ڽ�V�Z�bgg����y��J�>Ӏ;�l��c�#6u�\�$���D3��08Ga��4��KI�^|��KJ�����_Ҝ���/)��d������|J���&&��*K�ckD<��"`�0�$6N�J�-�o��x��d����� ������/��I*���h+|������K�ݲ"���!+�K�m�<�8�"ʵ�l( ӊD�6�6��A�Q�\rV�c��2���]̷ ^�R� ��x4����
 �vQ<���q�&a���iy�Z^�!"ۀ�f��B����> �����A����f?��K�LOz�:�5�CMӑ%@_�4¦� 
�4�ƀ�> �v}�ZLM,�)`��(΢pҒ����9��$
��!�B&W�J�D*����t:9Z�F^�C{�Ԁ������ȰZ����XL����z�.�|�E�r�9��4SCNI�nj ��dFr��O�*��U��P��%Ev�Ȇ���b�&&45A�-s``�v!�.>�5�v��״%���^� 0֘��&�jy���?^���5굕��0�s�Y�<��.�`�$Z�̴�3�g�J��'%&G�r�iR��HI�p�4�P���t*�F!���A��u��޻~���K/��?q�paQn8��1>��Z���p������Zp�F�T*�2vw�K��j5p��(��A�RӒ��	�hw*ҬȲx!%E��\2~�	/���ɷ�
,�+�;��@S3�H�3���%*0�	!h�K*��JK+M�%���5DԒ
+45�5�+k=��,���Y[
�����#��-�Ŏ�Rג���j���t0�����֜�����,�<�������sGqVԀ����Dk'-t41b�f�����RB�<M����ј�G�&jj��mYb��Oi�kXUPVT�dh}v��f�&�̤0��M��+{���l�9P�w>͹�W�6Tl+\�n�hՖ�������p��;['?�q�Ý�?Z��j���'o������w���0���o���Yu4��@��+�N��=����vf�m�T,�Y��u���Fk���t8mFp094���m�[�l����D��dLӀ���Ud]H�;q�[�r�����쎞U�z���k=w��̑��Ks�F�FG���Z�O4]o�o�i��V7�h�jn���46�61�59�����cK&�W�[}kb��Ȓ�+K/����^Y}�lυ3=�O.���;�lݶ`�%+W47���T�2
L�b-^c�4X��f���{�F5�Iɀ��N�(�P*��-�IEY����r��ħl��6�i�O�ن16!��<"�iYڜ�)���g�IK8EK�&Է����?����TN�����X��'�¦ޤ��`�c15�bM�+<���/5�?�m��6�Co�O��?t�?��R�~'�Z,��H�K\�OB�/Q�&J �@b�����'�)����s�"k������Y�.<]�|��ƒ��.�1U����}D�ާ�ާ��e�ޠ�PE���/1ķ���,�����I�e��XB�enӉ�i�'���曦�c�w^��0xטS5�,�W8$AM3���8!k������fj�ER����dJ�����S2�Q���R�_/|�&ޑ.���"5D@M�	�汀�':�N��活ح&45��./>�/oJ��Q'B���a�͠ωc���X��1S�ps��\!�˧1Y)Tr\"-!E�CӍ��O$=#��dy�33ܙg�ו�s��]�^[�i�ua��oץ�n��c�y�F@���2�MZ�Z&�`.��\6�a!l������s�� u�w,��8�x��`�q�B��Ҍ�S�MS�bj`4�c-��/��yVS�E�ɬ|������D4�^_�(��7���MT�y�G�}���?������˓�N�:5Gw/>�w�������:��T_&�5�M�ᕁ�&��]WphM�%�-�[�V7z:��]�M�R�� c|&@�T���E��"�΂s�[�s�������#��q�"�F��V[Q^~EIis}CGK��ή]s;[�Zk�jjK

s"��O��	�g���?�e�� hj�f�Yo0���l�v��as�-n��mѹ���McQa���E�� ��6K-�*�΅6y�V��5�m��Z|D@�w05������,��,&�>�Oрhj6T�T�	*Y�5*k6G�l*Ro)Ro/��������ҝ�f lٯG�oez�d�oG|��	z_	y_x^�g<�e<��r�59P7e��dT ���'8�+O��e��a&E9����q�8fj�������Sy�g�W�ozj�*_�q���,���;~9w�k��+L[�~�a�O���I�z���P���25�޼12�{W X�0��N���Nha��1��~p0� :|h�ʥb�29`�]#�W��rA3( �^�f@H�B�D��Q Q�GG�k�,�?����(�٤��T��`Ros9�+�?1?7�aL�-)6 ^�KO�E��Ʒګ�ܸ�'�~�3�vC��܌K9�,ҕJ�R-�OjQ�:U�N��MM@��p��_��Y�k����H�bhұt����(��	JԼB5�)��Yi��ٴ���2!W)�Tr�ޠN��s���^�a����o۰xK��m��ٶ��'�t�8�����ӧ�Ν�t�Ҏk���O޹������w����_��Իа�G��3� ��!T�HlVBjbR�����Y�8�05�i�	Ycs\2d���%��!��L[zeNiMAUYveEA}i^]�_p�h9Jq<������P���{���z��J��S0�8D�eє9�(l�)�m�g��D�.��Ih҄*2F�~
�9
u6����&�)I|r����g��q��I��^YD���,3ʝ25
~D����򴄦�ӱ�fj��V3=��'��k�����>�l�����ڠ�&�"z�x��Ey���-/uɊ�B�$�!�s �vA�ͱ!�V�,31
Bz^@����r�SBw�iV�!�;Կ���.�e(�^ӧ�O��Ѻ9|���Qr2l���S	�j̉�J�_��2!E.1��Ä�������ك���	Y�451M3��tfK��y���ꃄ��Ja��*
�lJ�R(�R�Ƈ����g&ό'%���T�)�dR1�~�B"�4! V��%Z��ƀ�� ��z���}>��n�j�0�	�����t����F�P(����f��!�I�&%�yT����r��|���!�15Fz��Yf�T؉ݕN�̉�:��1S�b9P�R51Mә-�n15�� �h �J4P�|�Ԭ�TVU�WV�{���K��zp�u(�����H�$͘�����!���J����8fBq�4�F�Á����XW[ѷn��;��w�N^>q�piYaNn|�1U�T�D"����������\(k��N"�@G&����f^�hJ�Y45|��Dr�Rܬh��T�t��1�,�O��"�Ycj#hK6ޑ/�W��_�cW�<�shjW蠩!&В����VZ�W;�k]K+m˪�р��LͲ���BK�#ڊ��Ŷ�{g�cQ�wAUƼ
wW���k}+��=����`4��L��>}e�V�YYg﮵-�1A�U�V��G��bJ�<M�@S3%k�ihj�����0�)Z�f*�in�֩i��bjj���<����������C����y��.e�JkǶHω����/^�;�R�ٷ�wߨ>� o�Xա��;�2�_�<�Z��e���5��]�z���G;O��8u�����g_Yr�÷��]v/�|�����է�zNU����=�;K��;��Y��q���^���
z-�63]U���gȞ5�&Z�f����V���R��@�v����r��TY��ջ(�gQ�ޭ�����W�L��`��P��H��p�(A��@�H�����+������C-C�ׇ;&G��Yxkl��U�&�o���3������'������w}x���+Ξ\v�آ#۶mm߼q��M�֮\����XW�[�9��fy�UVg��L�z�^�nP� �jz��Q��Ti��J���HE_���7K��U�-��^	{���	���)���+�	�I��������I�4�&�-�M�_����i�����̿ѩ�TH�Ey/�(���I	֩�f?M�w!k���gP����x�������d~h4>4��U�I)��\���7bɯp�/���G�C��p�%W�3�'�\�'<��\��O�(�k8�c��)�)S�Ө����B�?��>fH?fʾ����ФoP����WH�{$�6��&ң`�o���SC쐧e?�-1�4�8����f��`p�1�W��6��c�0""dML���nP�bjM55�r45�$�9o���[����ܒ�j���%z��,���B�鵄c�N��h���hs���nsr[]�V7^ad)�^�8m'a+1�O��L��I0F�����p昀�����!Ә�TJB2-)U�C�&kn X��U	��fW���d�s�yaoq��(����>{��ɰx�:�I�����0���V)��(�z�|B	!\8�
x���_!* �55�C�g��ԉh�!sK���c��4O55ߚ��s�й���bj�����QE�9� ��+~B����hj>����?��ǟ|��{o�����O�_wpۢ��ٻ�̾y�W��N�ˉ��[���[L͞�్E�7�l[�i�/��u�<Ұ��3�(C̢�H)\:��b�R�ܨ���.��MR��L=���уÅ�GP��7h�9�̲�⎖�]s�.\�x�0�����"�`f0Ơ�����173���LB>�x����d��f��n��-��i�p:<N[�Úa5eX��ѡkP��K"?	�N97�,����\�f��=$�caA����}���������4��X@45}D@͆
��j˖*��JB�L75U�U�
Ի���r��3�'Æ�A�@�c4��̈��[aﭠ祰����j���5�nj�7��b�(����1��o�- d<K �jV&�	_�È"5�r�b�+�9��(K{I�5�oz���˵�~�������t����+��y�y�e9� ���3������f*��(aC�Sxd�%�$�7I�ܠs����f���qF����WDM�41)3ʜ�>�Ԍ�y�<���1S;=]A�fOW�hj����$`L)cgP��0�v�O?ɣ�cQΧ&�Ө�E��t���[MZ�wb�I.�$'�+.�;����y����k�8t!츜��i�@SS���I����fj��O45�R)�R�.S�̐���u�d���M��ʲ-�ן<u�ԙ�/��>r���&^��;&�}}䇯]}�+o�2��[�_|8��W>����?:��G^}������;x��֡�-�.]�;waՉS��oذ��{UQׂ¶μ��PE���G�
�EcPӒ�P��8i	"z��ϰ`l;������DM��%��bqXo�4Zr�.�T#��tT���d�8�mL���9L	�� 	ͤ��e6	�#�q	UJ@�`��H		��<�lw"۞�2%�Tqt�L����h"%C,��2�J�Ӓ��Du6%���n�9�9)X*I�dX��J�A�w75Su������1Kٜ�4ei3�Mm����+��ʊ�#_#)p�y䑬De� ۊ��ܰ��q�n�����"�Ksʿ&b���t�W�ƯaCS���Q_C�`�F�h�Eȵb�6��|����9�nʈ&&n~u:�%am!��si~P5�-"j�wfK�rd`sp����;_��iJ�'�*`����1b Ԅ�e~Cġ��p	�MM���P�(���D81.Rȥ
9ѧ��>	��P�D+(���'� 5����;hj�R)8烹��
�J��|�)45�����&��KSCJLN�K�25	��� !�2ץ*pʠ�)2q
����t"�Na�+�#UNA��W�"ޟ���U�y��|ט��fY�扦�=�J���\��L��L��ƾ�.}A��.��w)�J45)3_H|aFr\<5%�����xJ�=#1n&��?J�R*����U]m�-���5���w���yktd�*��]<q�pyEqAa��R��h4�;���SPPPZZ^SSWZZ���3�L�h�!q��5D��|��b��tR
=%	�J\;)��j�\�c��8��v��R�Ycj�Ä���NJ��45�"45��fQ�~��Y\nYRa]V�\^�Z^�^V�ZZ�\\��(�t�ػʜs�]�*� 0OV{ �j��k}K��C�M�����yO1S��ƾ���5+j̀�:`y�qE�ׂh�(k��ʚoԀ\\m�MMT����h��+��o���X}Xܘ����r=�L�573��ST]�ޱrۺ�:Nݯ�7Q���Н��7���=���璘,:p?�������?*|�zӹ����V���ፗ��7���u���cw�O�k=�2�����'�7�g�9_�w�3wO��Í�/����,�o˯�5�#yN����~�&3]U��x�9�&�i��Chj����T���k滭B�S�Zk��[V�����ަӇ�O�vy�����띓�7nE��q�z׍q��c��񡎉�y�G��Yt�p4Ko�-�5���k�L��;���ۛ�����tst��@���=�t�86��E�v�޻o�Ν�W�jm��+�n���f���f��1SӨ��LM��Z���i�m*�Rc���,�hמ7�N�н"�6��eD�t��$'�%'n!'���c���[����2鿩TS15V�C�������4�
8/1������i��u.}�K�3��L�}.�M��*�]·��Z--��f�C��?t�S)~/��V*�m��745P�<fj 1S�3�s.�3��\��/��P��Q"ĆK0��|��?g�>g�?��>�������S��C���C�G�&Y�j��M��5���k��.�|�o� ѱ�QQ�	QTx��e��6T`���
5_75c"�1S�/�5��_:P�����ʸ��ܝ:�6+��-^���`@��/|����hjb5O�4�X4͔�iup�����Ҍ�(96I�6�OB1�HqT�J#���@S#B�b� �#<!��p��$��J�ђR)$1I7ۊ2��
���ޒ���Ң����P^�[��(�.�gz %���PF�m��4v��i�9�z�Io�kt*9��W"F���PlE���A1�������!�3��נ�b����񬦦�R�̀��V��bjb�f�b?��O�YM�<��+�O����S���?�"5_|���>��g�蝗'��pb����K�����|���s�;�h����¾f(k.�n��������� �wV��Q8���`G!���|hj��9�5��Ƭ3��tqs�/8��S�BL}��N��/;ڛubS��]�G�
{[lK*�`���7�s����7!eѹL��㰈�+�
��Ȃ�1�2pk���B%�
��`d��_`2��PYIiEYyeyEyiYQAa^NnNV6 ?;'/+;��l��+'�Y������x�A�5juSyO��'Sc�Yvk����#�ҼP$�bU�`�l��e�$5���"Z�V�E�^IWDՕ)k 0��3��1ڃ��(s���LT3�	�X4��yw���X�[�XS�Y[��4��2n�6m��l��v�;j�;jl;�,�+�ۢ�fC�jS�z[�fw�v_��P��HP{ҫ�4���C>�h�q=�~#칕黓��x)ş~/�y�i�c1�2���tw4��
��l�G�Q��N���D��8�7��q���l��r�_y� f:�֜㛮h#�V�����9}�G'~zx�ˣc??0�//��`��P�I��t"E|<	9��] ��\�8G�OF��pH����K	"��Ic���7���4�ƺNb�d`�4/������ �	 v6�z"t��=�⌰���Q.?V<xz��*�@;sU�^���5�h\�UH��3��:�2�iGXi'(���m.�ML�#��C��'�{&��y��>�	NȄ�2�o4�}����ߞW{�<s$�{.`�k���p�$iM��6�;��(�|��h9:N�AP�bW������ţ�?pK���?|`Ͼ{=p�s�.��v�h�����]=�����k�\�6ti���#�6�\���3puյ+����W	�/�_t���C[_�Ӱm[���������[��l�����@I�#��`ad�Iz�H���j̈́2�b�[�s�\���Ĉ�Dh�T�a_�J��8��b&��3y?���8���LOf���V���&#y4��.*a���2���)�e)k��j��<UX�,�Nbg��C�,+=��Hd��$�.��J�IR�x%�y�|F"�:�F�MbƑXs��qɜ9IXj���_�O�HXɏ�9�ZN����gr�= }ML�<��T�D��҇�����1Kѐ�����B��LuS�.��!��i���J��ȍ�#��MW 88�|�0�̏�ӯf�1�������V�]
�SNX�h�CF��ӼZ�_�x`��8 0	��?�m���2!�L#|ڰ� �4�,ȱ �V�c��[�R�|y�aucX�R6e�!YSPL������� �"
� ���	D�D�QQx�NM[��9SӖgj˳4e�r����2�!lW�4"	��JIH�=3e��q)�R�Rh)4.�#�`�'��J���Q0`%�Q0�hqY0�UI���t:=45r���!��v;����0+
�Ԁ��2��JJ��C��L�HdRrJZB���6�J�uj�J~�.�q*���0��?NEf"����*�r`��X�jR��e��>�9 n���
@g,*G1/� F�@Y�����|�7���dU�~u���T��B����Sc[��YV�cj2���Ka$�N��BҌ�I��$��'̞5g��q3�K�=����c��vV��|����y�9������;z�g���k��ܝ�}g�����.vv��Xp�z���������)**���)//�D"`�W*����X,F����6�'B�͠�)�I0��NM�iiF�����y�]�k�晙z������*
��tN��MMsx�Ew[��X<l����\��+ B�LE�L��D�Li�*;�SC�=Ee��
Gk�����^b�,�u���V8 �ݐ�5�K�˛+[ë��kZ�k�}�=��ӻk˪��-����FG��bjbR�MG��@A�4����DK��������(`"��!u7FкV�������,of0PXP�ں�y���Mg�w���9�:�2�q=��Nh�m@p׭���{n�]r�~�����^o��f���v��\)�5\��z�����n��Q�g�x�`κK��ӡ�'rzN�:��}�p���E;#-=饭��}z ��H���2�9�B��i��"*k��z�T~b���"ѮOSuj`dxY�˳�r�x$]�
�&��7�7�.X��n˚�ۚ��{��kW�u���������U������U��[q�ƒ��+���?������7ּt���w'zn��x��<X=>�핛��/x�~�x�Е�#�F7]����UG�,۳{ɖ��ׯ�Z0�������!�_�n��(k��Z���$�5>����V��ޮ�.S1��cV�9���?���w
i��ze-��KO�N��:���3�Q�n�6�_�؟���T��C��]T�8m�j6�B%�D��!`M���%��OMa�'�B�]�ο55�qY�H�r�fg����&ӿk5��T�A!�V!��L�;��7"�/Q!�W�k\ �F�o�O�O�/����|�O�"���|���	�O��P6\�3��3����C��}��=��G��whDԻl���7(�d���-��G�
O�2Wt���c	a���tx
淢�k&�0ʆ·�O�Q*�O�g� �15��ar��56
����P:&RLHT�b%��D	�~��&�9P�
Q�摩!>��dW0q�H: W)Ճ*�5��DzV��P�u�&�f�p�C��.��4M��|ep�l͒ >]���t���6���OۢjZ�f���lw�������).2"Vk�����Vb+9�G��e9AM#�֣�\ ����(O3��0HZ*%5>���,��+?3����7�U5�V�f�F|y����̢L_q��$; &9Aw0����9`֩��N%�j���J$B��`(�}`<� �����4�������JJ|��B�R��
��X�WTU�{�L�7E�+tQ4 prco���JY]mX[g^�`���eͦ�6745ۻ�c^����r�u���k~���=�Ț�B�T�Ȁ b��q�L��kbF�
5��ݑ��}=���3��!����+=��plK��9��pxK�M���=�m45Gw�9�c����Ss��-G_��M���zh��;6�߾�O>x�hj��ⓟ|�λn���w��֝}헏�9������/�k�����o��5D��_o��m�f��Oo-=��hSg��*�Rku�ԍ��p�G4���y:Q�ʚ�L�<���x|�/ �	�j��a��,V�ݑ�rg���N����IN$3?;'73+�DA0/���G<.��h���b��b0�O��|��p�0'�03���F�F����4��O�"�U��S�CS37K�D[��6?�3���b�f^���F��d͊|��BI�Ԩ֔�hjv58�ij �՛�5ۋ�{�t���tGC��>�ŀ�(*<��܌xoG|w��w������;n����t�h����VknH���h���2���5�p�����J��u� p�� f �i�aM���o���������|�������n��ߜ����3�W�s�]y�J�ű��
�R�Kd�U2z!��J�_N�^I��L��4��?I ���`}��D���\#��<� �9�`ASCh�o55�Q>J#����+8�A�dB��K����0�q�ua�ю�I'�)���m��L��F���}�va�ЋR���O7��T����ί{��j�84��q�o�g��V���iUӞfj�X�Р�Ey����R�T��$l���Ik2�g�ݵ{۶=;vس�đ�O�;r׹�[ϟ�z���+g����vn���ށ=�z�./��l�*`�+���\����Ņg��=q���Ѷ����mܱ�f��U�勖崴+�ܹ���I8\��M��4���3LB�M�1�"~�I�.\��̅	�\���11X&2ӘJ��2$�����x�i��4 ���%!yd�OF(�"^ΔU�5LE5UZA��a�)��^(��Kd��9TCUG�PP=E���*�dK��!ф��d^�7�ę�̙��%��X'�L35Y�#SÄ��15D�/^�C�� ^�G$��(��<m[�!��%�Дe�k�B�J^��R��ȍ�;��6~�ɱ"B�dyY&~T��#F�_��hX ���P3�J�O�	xA#2���-�L� ˄�Z1p"-p��|;�g:E�NR����,]T�V�D�^ycHْ�i�R7G�MaysH���(��������G��zS3�`LM�_\痴��3umy��\sc�35!�ҪI�tfr|��M5�ʡ�Q."DPhj$DZ��Wk�5`.J�ݸc��e��tk4�͖}��n�J>��0�|*�F"���԰RS�שɵ���|3/O�x��S�)s`�Na��YLM�j^�L���&�9Ȫr}o�zU���8V�{�mk�˫=Y�|�2C�*xTfr�~��&iN���8�I%�M�J&6h�`�kԪ�B��¼��S��ݻr�у���v_�0yc��͑S��^�0w^{Aa�Z���;�B(��������������ζ����'zT�F�N�50���t
55���@��cj`����eV<���51
,�b��@YSn��d�MD��5S��T�L������ ��Դ�Z�Lm���KG�ʚy�΅5��45=���L��j۲*��J"�雦fE�nE�T(M��@bc�*�e�D=�o��350�i^�z^�rn��3Wܖ�7�����6�,�+K���HF�Ԕ55-���W�{,o�����ۇ3��6����_n��6�6��q=w�d��E{'[.�Y{�~����}5Gﴜy����Go�(�9T�k�l�@ɦ�e[���i;x#k��Ђ}�ΝYsw,ؖ۱�[�j	�#9�H$���9>K�G������'��0���	���+�O����%	��y������]{6uڳ����k�z'F�޸�������ֿ�`�+�m~����^����o��������scͭ�}��k'G{�W]�v�ƅO�?�я����[�;o�-;w|�s+��=���ឃ�z��۳oî��.X��:����8�#���1�9�-vY�L,UӠg6j��r�
%c�;iQ\0)��%���{'��,���{�i�)ɫg��{~W���4�-�!���cT(�����C��K� %$����X�I�:º���������k���o�Ƈ^�_l�?���i��R��R���wJB��^*���b��p ��+������#_��/�O��|Atz�>�@Y���/�@ ��Ǉ( o1$�d?��f+^�K^��_���`�_�>�Ԁ9���A�BnRy������M��9S+
� �A�p�3Ő@4�Ԍ�r�Ew���d��L�U\rM,�nj�He礢c���	�n�6ٱ�.le�u�M���ү��򞦛�6;뛦&
���ms#��Z;^�G��$�K��+1���Ƨ1%(*��� Lt�^ e$fj�T:��d�(L2U�&K���}�lX]VTS^\V�]�,�	�ddz#ނ�'/�x�>��i1X�^mҪ�*�S)5jhj�������Ũ�6�K�p�4=��:�����O�r(+B��B��2��
˒R#X�����XL�W���cj�zS�ipߒ ��W���4O�YL`��G��'�����k
��<25���15�45�v,����ξ���?-��1A���-�vm>�sӔ���������ї_|���o}���K'w�?�u�Ʈs������Ø�鍺c��4S�gyƹ�%�W�^^Uk���+2����FID+�(%���H8���\5�N'"��n��\'�e��������W��\./�^o�Z�6��r���{�ޠ?��s����d����?��X�Z�V�ҫ5`b�h�������鰅����܊��¬@�c��u^�:ӭ��F��C�N9Q�a���cmA^{�cj �AzW�MLw���s40�)�k�ī���K�kʔk+��Ԭ�6m�1CS���6��쬶�d��2�2ݎ2��b��álݑ��_{�g��3^�Y�����{"�AȚ���u;����z]w=�{.�=��%����|O���Tð�>:�A�1��ԌF5�.r����7Q�*j����$�����_�����?O|��<��?~������ϯ��_G���}oun��]�y�&wΠN枥	/�$W����
���t� ]8D�2�!2o�̻NL�"�¿�~S��$�љ�k��fsG��f�Ǐ	����r�]�W$«RpM.���t�a���=-��#�1�-u�M����H*�D��T���f�􋐳b�a�M�jm��4���������,�E�q�UܣbtIS���M*�3�bä��\�q����-f�D�)P	�8+߮�,��j9~h��]�6�ٱi/�{v`��#[�[�H��k/�X}����'�_9�������];������_��������]�0���y�ͽp������  ��IDAT�3';No?q������Z�n=p�jM_uOo�����u���KЧ4酸@$�I6��aM��+��e�W���tL��.�of3T�)�4�%��Hc���>7LE�����,c>E�K�r�dѰ�$�%�g)�تB���"�Ig%3Ix���R��$�-�m����1��4�:U�H�)��.�0p��
Ӹ�8
?�̏O��N�ΎǓ��L���h@�)95+K���2s�\�SMM�*
�� 
 ����4eɚ�Ѻ�0��DPh�*0w�[�u������>"��k��*?^���EA�G��v��.,r`�N��v��@l�쀎ư�1����� �N��%*t�c8�%Ni�[Z�!��*�}�j��!r����*��& �)���Z���Q�e�;r��9��lu[��%,nc��4��AAs�(��4ĩu��y�aa�TS�:50��5�35-y�R�>hUXT��K����Ys����C����h�mMXb��&f��=�8��U,1`q#�CS`�X,��0aV8���>�$���0�R�<j��S�U�oA��<�Tj����)�q�l<@�] ����yL�Ę.hb�*ׯ�֬,���Ү����9��|+j����|�ܣ*�4V�p_`E�9	��D����x%展R�A���z�<�k�Io7������7����22z��͑3g��_��d�¢\����q��ܗ�����������⬬,�ʃ$
��ƣw��n��e&Dy,&���DJ�'�ǁ/��0[���02�h�U�k�rL��)�h�VJ��L�5�N&�T����Ԥs���t�KaU(h�����a5�jj:�Mm�ƖB=����Qj�[a[P�\X�#�,�K_���n	�j�i��i��6e�4��t�+�J�3����� �t?����1�����rz1S��D�H���(��������lUiPU4�ӳá���ƹ�m��Kw�>V��|����mC9[�6E���[��^����V�W�喓���~����{�jN��^��f�h�����矼3����C�[/�m8S��\��-ۮV��*^��t�5+vW.X�Y����2}��x��^s��P������Ԕz��$3C�(�!Saq����migKߊ�Mk��oj{qg����G��=�~�t����{�lݙ�vC��5ykזn\_�us���%�7m\W�nMa_o�ꕑ�KB��-?s�����\?�����4n_��h�[<�a�ꦞ���UuKW�,\Z3wAM{g}K{g{���EuU�
���6��[LM��V��7*�R�J%�E��Yq�(�h��V	I��P�f>����CM^�� M͞ĸK����� �T��A&��R���05645?WJ�p_fQ&HIC�����1u�� �ri7�]��*&xS�_��L%��A�'��ߍ��k��U�A-��J�;��wJ�����A�_
�_��_10��O䗨�y�_�Ā�sE_rpB�p�j������@>��G$�r�B�{��}\�>��ɑ�ŕ��S��U�Β�Ɣ��R<�<���	L�����cj�bjx�l����bC<|�
����@S3����̷��~�����\|D+�k�v��mVl�[�ƺ=�RF4x�|���^��]n�xj��b�f?AS��`���T��|��J`�����8�$X�曉N`e�� ��pY��d!��$N�6�m�㲇|�Y�¼�¼p~NP��	u�3}�P���4�m&�Ig3jM:5X��*�ˤ�@�P(dR1�
�"�"�P��G����2i,j
-i-�Z������X:K�L+*�`�tw���������ꊙ�X��_oj�����t��cjnn;�e����9�s푝}Gv�֘���9�c#�	�������_?wt��c[�oYpfߊ#��/Z�S�כ�����%�wT�]{�����,�@SC2~�N�~j%FO��">�IK�Qɰ �5��0y�#�i��
���`0X����t����n,//���03�������
����a7[�F�A�U�*�\��B�B�U��E��6v���y�2Cّܠ/����8�C�%!wȦ6�-B�IX^�̊5���AyW��+�w�AnG��0�B��0ga&oq�4G35P���41��yP�X[�U���h@��:B� v7�v58w��&fj �+�[��;�/���菄u����^�%���k��f<�>� \�;'}�[~��u���qŚv��5��I�t\(EDl|�#���\l�G8��|�� ��I'P��>�R�Ib��ʛ�p��ξ���_>|�����߼��߾��^���F��r��+-k�؋N �=	�=3Ǔyg����"K|����N&�Φr/�q�&2FY�A�`���!���&��55P��8�l�(�?���O35.��$^����a�lD��)%�U9�r`L�1��r�Ab���y(?1�0>���5���xg��C�vf�!9�z�����������!��i�E�ZA���Q��:5O35�>���%d��+S�j����Ez,c�9�+�6��X�m��m��l9�����t����6\8���UO��tjɥ����{�T��SWNv\9�q�L��s��Kg�.�i9w����SǪ���"���޺C�k���;�zzJ�W,\����oT�;�2u��*�DJU	�Z�55|����2�/A����'�31h�f�g'��S�	TG<5=�H�d� yiX^�(7M�CgR��,D�X� S�g)}L��.w���$�:[`��s�I���-EhJh��8�tK4��!�J�P��II���a$�����3�4,�*�C�N�ϊ�54�C���hj�*f��	MM,�鉦�]��&�a�.��P�4DD-9��<U����s�L����\�'rT�9
@S��1KQ�Յe�!iCDU�W�	j�� aX*���mEB �"�w�E���)�Ҙkn�1�P�m���W5U^u�_[�6��M�Ɩls[��-�4���Yhn��7f)�#D��J�r5�EG��3KݕKЙ�j�R�eJ["88�6���A�1(h
!���<������[dM[�B��n��CX��5[�Ѷ�[rL�Kmͱ@S���JLĦ2��ΚMM��Dhj�4��MDhFel��j����e�2p�sp����1S�r���#������f3|����,s�!�F£��|�I�J�-x�-���
;������+����cjV<����M�U�z�Ew���R�Wk][�X����5��]J�S#N�==uv\�Ԥ&΁%��8
v�f��QH�4)E�����B�����>948t��݉+W�_�[����D�V�ly��p���s��C�PF��0�e�Cp�n��{�P(��%D���DN��6{V������9*.�%�g�Eyfa��MM��^b�@�5O65A!�|����=����i�'�e�3���s[���@ה�c{�i^�}a�M͢Z����&��o���)cuc:45ݵ��樬y��YQ�뎚��U&Ȫj3���'��WʦB7��Ā�j������E�y������y�<��pS�ujJ���0�Q��]UY�ں��ce���E�Wm<װs��ű���U{&+vO��[�^��Z���q���g,>�ƒ��������_�d��G+.��yxb�������?<���#ˏM�:us��[���/?4ܽd��K-�GV�_����;\���������p�s<�"��ȫ��.��S�k�d���ʰW��Pg夷tT�X��}�����kV-�X��d�Ҽ�K�-�,\�l�2T7Jr�����f�l�����t:i6�b!��$�)E��W�g����V�׸nu릾@s� �@}���0U)�����#��������.�##���uiffMV�1�o�;�݆��քU�5&n�n��4+�QSS��ԩ���N)y��M���.�W���j�0aj�x�5�������U�3�Ž�/%�*�8�����E�/%��I$���C��O�v��y��|�I� %��G�	m�G�����|�]��@��%B���OD�����4��`��Q�$d�F���'C;3�Ԁ�I`��ሠ����-|�F�q��s����"��} T@ޅ�*�[\�[|�[<՛\���l���[L�V�T�50� ��@�h0�	l��}2� ֗��hɂ���FP	45c�:5#��MML�<���F"�nj�����#z�3�ˊo��\xo��i���(kb�fz��������6;���|��iupZ��f�����S�L�d���3f=�JL঑�,�v/420vL��c��@S���2Y�h_�����u*�A�vZM�t�ŗ��]�;�s��m�k�e�9�6�x�ͨ��>ip�Tq4��}���L"��\�HPT*ĥ��maL��L������S�58��鮲�j��^�j�g�����fS�3�i�25�d�_oj��vf��5����'�?Sspsۡ��l_x|�c�V�:5Gvlx֘�C�6CS3U��ޅ�&����[���g?:y`���[�\rlϒ�;;���?��yL�yJ�����ٍ�Wv�����lY�'�Q���VI�JX��P�שǸ-U@O%~I��n5*k�[�`�vNp����]���w���
l���[d��#�HNNN~~~QAaan^v8�x�V�A��*U:�Z!���Qj� & �[��6��(Uc1��ƀۚ�s����J�ʳ3<���xi&��Uq��J+�1o��"xg��VW��f΍2?�Y�Ňvfq��r�V^U$���@_j֖��*�}U��ԧh@45���]�Ν��]��j�T�UvU��9��;��iNy���~�u$��O�2�xL|�u���q���%d�+7Ѵ��|�6%k�(�7e�I�b��
��tR ��`wP�.���.�.�$���}d�q��vђ��~8�ѿ������/?��/����>�՝����+�<<z�~�u�]}8	=��=��9��<��=��:N�I��M:��:G���6̑�S�S9���r��N�@���1�П@?���b�9C\�0�?�'�	CS�M͠R2�S��Z�5�\?���"�#B�1�y�O;Ǣ�hw���5�[�_�5o����������2g;�t֡ʴ_Y��+n�P�z5`:`�(�se)͊�E�3��yu&^���d���z �E/h��tX�]�	r]�5K�m^׻aS��/n:zx��Ck�_{��g���Yy��˧�\9���鮫�ڮ�l�?�t���ⱦ����՟;R{�@��+�.zqkў-��=[�^�V�{K���������pg����[W�(sfg\N�A�Q˵R���3ƍ���L�20N:΋�Ur�!��Hc��r�)�`2?+�I�2�D�$Q E�M�Sp{��H��5)
Y�"IU�2E�D� ����T�&�x*M��s�l�7����e��"�P%R�TL�I��E�L�dV�`�qB��Fv ,"�L�	*�!%#�afj�:zL�|��@M3=�	�����>$���H}ǒ�lY{��#Oݙ�����-0��3Oߞ�m�Q���
���BUg���X?�J����<mK� s�������2���-.t�`��+�����bgOKNwc沺��� `a�\l�57e�Y��KG����1��1�Թ��5���Qhh�Q5f��5O�Q�iϚr���,Y{�pK�aS����7�-�5S�B� �MMg��td����O����MicH֒�n��[r�Դd��sm%^��$5)P�M�'Y6�M���gs�<���E!�C���>���"8�+�J���L8���8σ)
��.fdd�:5�߳��i)".�$�xM��E�eƠ�??���M����O��<&hb<�h �Ԭ*W��Ү�����L�� ]�3���#'Q����O�䦤&	8L�LlԪ�{\�C�T5-9�� /������Ko���������'������֨Ѩ
"�	���l�z��4��:�\����%�z���Q��dP�)��	q)�g&�x�7��'g��bNĈ��,hj�l�"��L����p0��ł֦��n�[sD1S�j O�5�hj����%ƖB]S�����U�E���5N��j L�ԧ/k��h��4y���	KCS����<b*�&�izj,�k�1�S�l�|M�aE��[X�+<-�F1�PE����M�����R�Sq��8?�����kYsWoq{_Ἥ���V��]�f�Ŋ��K�_n�=h�5ְs�a�@�֫�.�n�P��Lن�N�n=[��L��ӝ�/u�p����][Nvn<�x���{..�|�}����[��n���Pڲ��nanYk$�*3�0�ED�]��tK��V�3f�ܪ�t�KLM����²���6'۞W�+*�U��F�݀�4��"�%�E�BE�J}�D5C����7$�ߦ��65���H	�(�g�9B,��Qt��<���T�x���K�ͷ�ej��I3��9$zB
#.�:#.�3��������?���P&G��1�O.�׈ˍ�j��Ό�LM��cj����^��)%����m��z�U���=m3����ܝ�<q��9/l��y��<�c�"oa�G8���7"џ��?����n���TH��`�1J��{?�p�,���x�I�o��bȻ�>�W���?�1�dP�A� �Q���R���7��WB��
 �A`|�L!k�_35��hj���?�~�H~*��S|��>��	� �wy�r�o�~�S��S��U��Q��u��U��i�f���q�·��!�K7�?������!>"�"���d��O��\C�������* r�B5�T]S(��*�a�x��a�7;�>7�:�(�$�/�HgL75DJ�Sz?�Z�0���ƌɚ��!dMV��+
��8����ċ�>c��	�T���F8L�e��.h��	�l&�r�L���:�J�V) F�F�Uj5r�Ni2��f���Щ%.��e�:M�Ae֩LZ%X� j�L� p��A�T(�j��x/G6�P�aR���"L� D�'ؐp�49�4����l*^E�#fjVV�WTZWT�?���fj6���k��S�@M�iV��J�<��pL͡-퇶�;�c��+���=����{?=-�
�k DE���!���������{��o���Ȟ�G�߳���'v��?����h��9���4Ssz}�������Օ�E����UŮ�s3�3�6�t7T��"z*3e=5.-5l[��ld�����=�'>��
ֵ��l���
�6���v�j�4MQQeyE~v����/�A�8���H)��DbL������~���F!���J	n�k�\��o(�.
8�R���J��:%�V��U�xM^�3�ue��!^{���tEX��Ej����<fj���)������T�W�^W�[We�5j̛�[�	M��䆦fW�c��� 45;��K{������#�)����p-`	�&"��a�5�~��Lx���I��v����r��'�A�����f{�d~�`|I���1ܐ�n�u7E�;��.&����P�]!~G(d/��St�!����V��?n|8�ſ�����~���߿���<��w�>����ߟ�|�����w��<����`ג�gfQN��Ӑ!���1*տdp�n��a��2Ep>�y%�;L���8C8�D��L�4���7��
�o15��p�V�ƍ�	�fD�RI�b�%�wJ�:& 4�	�uZ@���AS�^�O�QH_#C|��j'#y'e��s@-�#c�Sp/X��`�z�*^���W���R�%���t�z3�h�7��F^��ߦGZ�5�B�6z-�Fy�Ϲi�����o۽}힝k��9��w,?���'z/�Y|���˄�����*�h����BPu�P�À����N�/=��h߶�=���n���8:��ܘ�ymV�*��y��y��VWu����]Zj��Ի�Z�Q�Wi��c|3Ƴ��/�%�����8f?YX,3�e&1��gۛ�%!�A(&J|I���+Ua#)���R�4r�V�2(xf�0`n��g�Ҡ�0!�:�C�2I�Z<M�$I�Ibn���r��$!�*D�0>8$&���a\�0.���Μ#IL00�N���L��V�"j�����~��)w�-;:���/�H�h}�mCic͙��lY[��-Gٞ�"��t��M[��5��#Ej@W�v^�qa�eI�sY�{A�m^�en�u^�mA�c~����֞o��,�%�2�,}Y]heSVOK������iχ�j�^T��,v����r�`�ȷw�畸��U����(Է�iZr���|EG��=S���#LD��DkʴE�ְ�9�6���L}B[3	����t�ȞHg��-dӖ)m�Ț#����%K��4g�!]K6�?�{�^�� C0&���2󅘩I��LI���L���py\6�G��<��,1��0�	�����ɤP(�~��c�V��`k|#��*
�RSD�Q��Ћ�&QĈ晑B����)�r���$(��`�����m���c���zJ录ڵ5�����'8���c�)��r|Bj|" �)l��J�IG44���|6������+%-~�`LwX.脦���޸sw��ͱs�O-]�����t���A�
5�P���n
�T*|���l*�O�~�y�������N�9#���gq��H�)V��!�A���kb٘�6F��05P�LO�����h�'hj�h[֔�iϓtȠ�����MYC���djڊ�Ez0�*�̯�/�qBY35��҆���+\��]+��S�&��􍘚)S��z�N�51S�[g�.k�\Se��=hj���,*V.(R/(��
s�9b�'�!"�	+���␥$�W��SUY�޾��s��M�n<1㉹����v��O�[��u��n�N�,f::��������8��c'�C'333����nۅn���n��M���~o��������\�ѱ��X��[�<3i�Ɏէ&�<U5�@��}��;
�m��X�ڴ8�z��r���W[�!�h���M^6y����g��Z��L�u����"�;O���-ibm��]dK��ϪKɩOϭ�ί.)����OKH�MN*�H��L*O�'�
=�"����sLͳcjjҕyI�-ʱ6�疖g�L�hJ8�C�r��LJ$�J��QF�QG��F��cD`��1#G�C0��;.`4��px眾K�L�nMMR���HQTJ@������ƍx.hԈ����Ə
<6  $ �6v�<:�ͣ�)��V���1Scj�u�Z�VAi��p�2#�ۥ=�43���4�Ao����K���7*tv��eQ�ۨ����}Eߗa�+B��d�F�?65o����k�Ez���t�G?�'�A�D�d��Լ��~���a�}g�|o��ۢ�ʠ|m�~���K���\�7�2��<*��/���G���ȚOx��ل�!v��>㿓(��� ��V���D��X�H�O�&[�*S�
C�_�W�*���
�[��%���Y��3�0��bs����P\�[+�O|�ODӜG�Ą����,���;!�C��y��9�PN�4��@YsH��j��u�V;e�n٢xٜ$b��i�g���945��j ~S��`O����<��yhjZ�F;��&(�s�"��"��
ϊ��Ƒ�l�����P�75~qu�")1@Sc5[�v��h��F�ƕ
�c2Ä ��/sMZܢŭ:�U�2i�F��_ �JA����JP(�`D��0�LBD�H1�L!���P���cj��cY��=:�&��_�4��9��1�
|�:�؟oj��y�_S㏦�o��ύ����6�r����v̂�f���?���c�����K���m��[��F����'�������7��{`G��M}�Vt�Z7�����[15��w4[g�@�nj����>۽n�}y���ѹ�#{���+'T�U,i���֐���S�Qc��!��(���`�4|�2O,���p�<�P DDb	
�.r��z��2�2s�r�
��J��*++�s���No�%V�
���q8_ ���D!�@�������oդ��x��Q�A)u��NCQ�7ŮV	�Jn,@��4
b�1��b��+hKCS31�Օ����L�A$��u�=�R�?7���9%���JPB_o�/W/��-��/�1.��Ij|5�Ԭnt�k�4z����,�4�W�VU�J��
��S4[�U{��ŞҜ�3����2���T��ׅD�y���v�k��u��:�'z_L�����r��t�hw�d��hq���okl��滸�Lq��5�-DrU(>�F�d���,�^<�͊9߭�<t����d�/�����~���z�w?��g+\+�܋�v�G��3��K1����<����n^����h�[C�_j'��J;#�Q{c��I�S�Y���5L⋂���9��>Ps^���H�@Gs\Fp��'T�s�e�pZ�<��CE��N!���p�"��|�)6��P������^��T|U�>Ρ���v���B�jy����-�VI����s)���έ�\5c��:QOi�ĵi�O55m����DM�UXo6X������Մ���jAS��ȩ/�H�_ط~���kV�^��oӺ�k'�韲q͜�;��?���)G�t��zlOӱ�u�vV�YytGő��{7U��X�wc՞e;
���Y�8c����K��,.X��p`Iު�K����z�:�:\�M��jGy���Ė�i�v+��*����)Gqq���&�Jy�^�T�������98|3��%��)�pnz$�*H�K�R$�tIs�����f��Y�򜴆��������Ңi�e3�+z�*gW�M-˞T�:1�S�h*q��LX���2�(]+��
."�qv����P$�$Ih�8$R��D[X�x���Rpn����f@S�e�e�ij`@͏�>��.EԐ.l��`ך#���A_#k:��yzB��;�u�Ś�"P�L*5L�0Ϩv̬uuW�gT�fT���=3k���V��*!�gڋ]��R�8�>}΄�y�P��m���E��K�*�v�:\���<GG����1��9��5��6���Ub�(ҷj m��)۳�]Y��L�#kϔ �2P�,��LIK�i��i�B'fK`��p��yL�C�58!k�ĺ�leK��%��d�%�MMK���Dfą(�Ĉ"�z�԰i,����q >[(��|�Ưi@_ ��p�&�Z��oj���V+��C.hj�^o����tj51?J ��l���ܘ)�j�s�h�Y�75E6n�������I\�A��15���ps4�QxV�bN�n^-1�|�Q�T�J1ˌR��If��Т���xd49&	�t
���z�ͤ�*�RD Z�\(i�%..*�E#�M����+WϞ<u�ߺw���kN�>6A_yy��n/�P(�~M�T�Db�R	.+�� ��F����w�O�(��L��u1�!������i!��H=Ɗ�R��� ���Ԕ��EVJ��򤬩p2a�ʷK7�T{8���?��-_�^�����e�������Ui�T��hj&W;A	na5���z4?�h|h@�]����gU��45���̮1?fg����7<,��gjԏL�|06ea�i�UY��4'9;=� ������qjN�Ą�&SR��U,���"{�V�Hk�S'ȓ$�����ϡ+R(X�(��9�* J�G-���VL��Ȫ���v|,ol8s|4+,�AQ9*W�Q�U�v���N[B�#��5�:e�)�Y��)�B���c,�7�<S�옚�,Ma�<3+̶��&'&[�쨀������??"`Ĩ���vf���1�ύ9>,*42&"26<:.�����(�+�ɍbp"h�P%`����֩S����z��b��
�GtR8=:�66z�����>�3r\@@p@@T@ /p�..4������hj&++,����S�I���A�O%�*�i˸��L"IMoLجp���dP/�����Q��2���/��/eү���ϔ���U1�&�M�E>���\D����Q�=����M��T��H�;\�7��[�<ȷ6�?��/���t�tߪU���_a2 �]��J�����_P��?
��P������#�5�D �-"��D�9����Ia��T�;T����H�_�>���͖��S���_e�0�׸*�+,�}��Y���>SZ`�U���0.����FtN 9'�.��K�E)�Y��I��<�ԜUj �M�N��"_㔭tɖyd~05ӳ�Ӳ050U45�¨t�l5���	5cgA���m�D�_ja��4�8�^��Wh:
�
d����cEL����������|�7���K�A�w�����j�jT*%&�2)"A��+2(Q[�!:�)1�7h:�Q`j\~D�c`< ��X��+T���˵�T%�)1�-�ԀΈ�!��`�b)�� ���qUe��3+�}���5ξ��M�õN�x(k�=����M���@M��Gvf8�嘚��+'�X3}���]���Z�h���;��ܘ�M����Լ��k�w�x����o>x��7���O6��;�}پ�s7/o߳n245�6M<�i�c15jT���ٿ2w�/���;�i��&C�jjv�K�6+~Go�����ӓ���?����҉�n�V;�4��*�ʄ��\��ˎb�FR���,�F"��*���9|.aj8?,6�=���x`�0#*0�����SSTT�q�5
%�2j\J>�â�� ]�oH��P���`�F�`�����ϓ!���P�1�h���TK��X%��⒥�0-�!�HB�s���5��@;�ES�]Y|�i �3��rD3��3�S�75sK���T~YM͂
ajj�uO0�������m!L�V�
������-�4.�4�,7�.5�4�R��;SR�'2\��/�\�I���x1#�Baj�'��y�<��.�5����A�~���������}��}���6�w���j�m\}S&��ʈ����I��(W�������'��f�ж�CW>�Ǳ�����?o|�����v����0t��:���*�m������d�9:z���ֹ>�m�~�¯:z�������f�I�� ��;�~0�}�. LMx��(��jj�GSsZ 8#�K���j���i|��Oi�L��v�e���Nq'�>�v�;�]{��{H�=�c�f1o	E���ƿ�����M?L'm��n�� �u"�:	k�X��6)��M��&۽ե��aM��;t_Fᇦ汀�v�@���h��b&�i�(�-[MH�m��*a��T�4�f$-��ۿ|�E��V�ݲq������O�40�ȞE���=�����;'��xxG��mU��n�8��l׆�]�wo�ܹ�tpu��e٫�/���?��b^Ί��+d-����'i���is55Z�����kV�>ޭwX&=�ش�D/�e�S�ƫ�^	?I&J�
A�+Cq�W*�	����F�1<m��Iפp,�t�-N��5�X.�$3�RY��QW�7���cʺ�wM��g���S��:�����/8 �1g�ԙ;�'m�kZQT6'#{rBr��S�P�vU�̅Fm�F�(لL-7e��xa$~8�+����L<xbIra����䤩��d��z����4�����da}aj`�
0���M|�<1W�[��,�:
t��ڶ<MW����B(�J��ˌS+�=u��5�޺�Y�	��Q�Z��*��@�i�����ަ��ƴ��}�@Tf�d�oϛז�]��U��,vu9�m��kg�uR�}r�͗4�2�� ���X~{G��#�̒:21����g���%b��LqK�PC,}���%���,S3)W��#Y�������i�PN�ַ���5-9�	���Du�Ib�CS�35q1�a��*���x�/p��3���
���k�� Sw��h�Z��<����0�yj@#�z�^���8~<xX�s1�_Sc�����$Ä@SSj�X8?ޥ[\�V{$�혚�����y�qN���L�W�'�v���6e���T��(�HYv\����K���1`�l3�V�@�:�.�ʠ���Xf���$�����O�����p����/�^�dQuue|�\>�ʃ�` �^o�\V:�.�`,!𭧆�گi��;���4&"<&,�H{D��bPZ�e&�� �@�~*v�˝�b�SL੦�)iˑ=ij`��5P?�Դ��;�,]��U�)�Ω5.��:ϴZ7��FP�Q��n �	�,�56���==�5~����r�Lߞ�0��IS�?��<� �S3��Y�h��,�*+KUUd;K��=i��%5��)Ez[&�F�A,����Þ���f�aBX�#)ϓF�>OD�FF��$���uE�0c�w1�%	���܈��G��Gz~Dt@@��υF�O������ct��f��)��k�K_�5T���<r�i�= ��	SӘ��Ԁ�ϊ��L���������z�M.Eѱ���0n���G�GP���a�ƅ�7.�I�!r@�#��1 jX,-����GǍ��x~T^YENa��h�"���%3�a��1�qq!���؈q�ac#��D��
	DF;�>z$/p�""�ŊΑ1Ku����,���}��E��YǪS�j��F9i����&;�d<o>i����*�[$�!c���I�Dώ	��<*b�vQ,���L�G�����K��J���8���_���Ub���7%��l�eZ�y�"�z�O;ǧ^EyW��kb�-1�%��M��])�+	�).��N��6�r|o3}m��Ө�Ƭ2��j�V���c�/eҿK�g ��P�g���@���VB>a���P���s��Or�_���)͟��@t��?�>DL�!�Ŗ7�|�\�}����U��u��U�"E�*G�W����ˑ�aKo�$���M��
�s�̻E�f"�Y�����4?��\D�$�K245g��s(O"2hj���LqJ��@�%��s*�Y��JuB�:��Vu��^��Wx��^lI� 	����������jhj[ �TS�S3���z+���-3r�L"7JE�c��A�#d0������� 0T$�]�T"�c(.��J�S�
�ݑ��J�F�ab;��8t�P�F�|*PH�B����hUr)x("�F:)*�J�B�%aj�Z.Ua�S�q"�0*C�"��g3x�8JD ��5J+�]�)zhj�Թ�j]�ҧ:�Z�j�3��-�����3 �l ?�3���15�27���ؗ��������I�VN߱�g�@߮u~���xL��ٴj���K�,߶n ��W_z�A����~���o���wOذ{���g�_6a��)�6��Y߼g}����Z_wx]ݑ���k�!����)߿�|���U�{W�_���?oߊ����{�g�]�u`Y�%���ih��
�3?��;�A`L͓@M��g���M�13c{7Q���ٷ���򊣫�/k�6�~`fmwmn����dJ&����8
�Bg�� ���q�l&���� ������I��8<���@�#!�T�H�Y���$R!_ ���Re��xN��5Z@"�Ǥ3�4:�xpl����~�A2�[%q̦ƭ*�Y.�!<9�"�E��ByQA���H�s��QNaD����E;��]��I®tޤ�i��]Y�IټI��I��i�(`z���H6��)������˕ P��4�kt�kK��p˧��vSX���׬ir�re���ֶ�ڲ���_eZ]mY[eY[fY��_��Y��ؘ�ݞnܗi?��:��=�>'�r~�������Ƌ���^�E������~���w��9]�|�� !�7��{���ݲ[oYm7��k���"���4�Bu��=<�v���>�Ӗ�����<:��ߏ��ݥ��<��g��}{�ա��wW��D��E���#�q��0d+��5oh����C����i��9�wm��͞X�֠�}�ST�Y:�<] ��s,�6�IN�8O�$�y�I�1�Q6�1�8�u��>)��rO�yGQ�	﨔8&�r\��P�Ok�Mʫ6�%��ZrPJ�{�-d��v�Y����<�	>�,�w�Ƹ/�?��~c�������.09�y��,�jz�
Z�*v�>e%���O^���ؕ�Ṡ��[�L�i*j�"����s�?�f$h5r[�l#0��m�� �EO����"�h��Z��hDj��R=Ҕdɵ(JS�k�&�OX�h����-]ܷyӜm['�Yվr����{�l��g�i����+k6��ܲ�b���5�� U��6�Tm][=��d���U�sW.e��堽bê�����/��>����bk�1U�Z*J����LSz�--Y�jM:�
�T�餈U!q�0�q˥^��en\�K1�P*����S�aB�4!�U���UU�?}����Ó��������/�9���S�?���3�����/�l�;m�I믵�����eٙ�e�ۗ����Düõ}����\~~ƺ�U�v�vn�kX�Q6;)w�3���0�s�����#)�H���R#�I�ZeB�IR��t�L=?KO���o����GSS���~�M�6�I�č�hs��%��4�9򉹸�k ��Ug���X��'�v%�)�z��j�ӰO*5L)�L��AfԸ{洤����jL�՜�7!mvkFoK�̦�I�.���|cs�aB����4��6���V�#(P�)�sO�5��x�I&d��Y�[3�����*��u ��x��lYW�lr�|r gN̔M���l�1k�T��j���r�u��<^�7c�G�S#1��00�	�������(L"UG � |�o9�������T*�ZJ0����&�?`bb���X,P�C.��O���஄���~
��Q�!��|>�͎%�őI� l�5d�4�
�F"S�c�t-��!���r!È��1\��c�[��v^���0��QLM�T�5a]<R� %�1IҜ"�khj � �Ưf�ǂ�f��`6Y𰽕�yu�3+����n,�*s)
.�C'�莋�a�(��E�|�T�S(4rbP,�qYL:�M���.�"��`Е��^�x�ڵ+�n�x���ܹ�,hjjW������EpAE"˷�:<8�<5�I�Rp/��� �k
�,0V����	��
	!GGpi��X'^�M7{��[�E6N��Yl�75~YS1l�/�6�W���M�w������Y�w7`j�aZ� M��j'A�ۇ�]M�R�*�w��:J���)U���nȴdz��]����)���M3���|�k�)��T����4��<�� p֟dv� �����5X�7��� @��5P3ʴ��t�
�i��)Exg��-�xŪ���ƪ,Sn��</��0�j��i��X��и�1a�}�eT������$?� �cF��EFG��Ȃ�X��!䀠���"ENi����u6��*@�Xz��1c�G�0fԈ�Q#�#G�F�
5z��Q�F>?�a�P^�I��P�;E.E�GQ斕�%�r���+��J��=�:��&I\���R$u)��T�>UJ� �"����gJ*�U)�m�w�Q���c��FG���8.$$,:����ǅD�G��	�F��!�XQ�q`���T>K��1x����ǅ�<7��`Z���4z���Ee���F��Ƈ�	8�6~<7h�8t�::���LR�e�J��Jǯ����f�E�nV�5"��"�Zс�-3�v{�'���.�Q�b�J���W�8���,�<J�¸�E��[Hq�E���m�� �^(�R�YmCބ!���:�Wzݿ��/��q�%>�:�t�{�K:�%���]B����b�����@�y�+�F.����F��V��N��A��Q?d1�[��F�|���[���R~��e�oR���P	�b�g�7����W!�g��<�s��l�﹒?�/D�?�5A��� ����
��HlH]oa	�(���3.IR���[��2��9�W��둂w8�T�KђWH�W隗��,�6Cz���g�PE/Q/��(�;4��"�{�Ż�]�>�W|\�
�x�9�G.K�K��(%8/#8�J �%'qB*;*��{r����X�����	vǎ��cZ�!#~�(�g��Z��n"7͜$Y_��/�/q�F��2��
C��I�f� ��$])�$Q[�`��iqs�]l@�����9���Lp0������+3sr4l7J��ܘ`zd03.�C�@S��ب�+%�L�p�X!C��P��19�+�J%zpЃ�a �>`���SQ&�N�Q `�*��b���F�\.Ѩq�F�`�)F�1�2�}�<&F��]\��ĸρ���@�"��"�R"�1�R.١��X�\��l��}���*;�{+-���)�ϫ� �W�| }��Z�Z��(��Y6ؖ�v}�O���L�s�|ͪ���]�U� T3�� `#��fR��db+�SaL͓������l�I�ԛ�yV��Y[��a98'g��\P����=��� >Y��qn��y�[�..\T�ci��;���-oغ��eY���S����kͼ=kK��,�1�t׺�P�l[K �d���ly���p`daj o��2\����%L͛�Oذw��fn\6a��I�6���в}Ӂ�P��9��zߺL��fξ��{��|S3�qA��1G�>;cWo������Y;ff옕�g~����K�-��4�x餼�bo�	wH�F�XBf�#�Xѱ��d�ĲId0Pp�<.��g�l��gP9T*��esx,6��p�,!�'!*�B��� p�s'�=C�~05:�
�O�<&45O�N#�8����)�"�^&1�])7c��9t15ZΏ�E�C�Sčq
�����ig�rr6%��Ο�����@Mӕ���L/��(�BS5�3P� ��YP�_\kZVg��4�Ԁre� o�U[�UWT�WW[�TY�-k
���+�T��5;3���G��'s��\*J�V�r>�u>�~%�q5�~�a�j3�u9^��?p{�9<�\�{ބ{	�����=�k.�5���v�f�n�]�[/�L�KJ�i��(j:"��������7��w�Wk��}��֟:��Ѝ�>|���5.XD7�Ǩ6F(v�*Q�i�6~T�})����u����-=_v-��a�o�_vg��;�X;¨�c9gi�3�8�i2��qG�Ӝb�N1'Y?p�M 5�1.�8�uL�>!��	GsXF �Q�rR��RK���W��kv�%��R|@�ߍpw�d�^� �u�K�'u�ͻ�ܓ���-X���Kl�a}��O��a���5<�Zs����$�oؓjY�Q���]Jj��6���5455M��05��	D:�$k3c�y�E�lF�h���Ȫ����,�5��fZW��sf/�7���ݻ���;{��ik��l�4k���훛�7��[�_���jc������7,�X�_�fy�@Ն� P7+֭�\�
�%�Yп(kќ�y��}3�&���j��%��"sq�1;ݘ�dIM2��:�A��A��KD��(�XUr�Ra�q�\n�0P��
���&�hU	���m}Z��Xz�w�՞�o�8�6`���&�z�u�����U+/�o{�m��	��5m�]��F�ꫠ���|�Ӏ�ŧJ�(�s�p����g��/W�?Y�w�l�΢�Mٍ���-)���)Y��\)�-D�F�0�	C�
q�
I�	3t<�Qw��[l��545P���35
b�Q��`)P��?��G�%�멀9޴rb�����U��{o�wNKRO�Tf�$���Κ��Ӝ<�!aZ�����Zlj)44��Z
t��]���営B��m[�zb�
�B����$�N�/O45]yJ�5� <Ɣ<դllr6%W��5��[}�@M��&d���'�k��$<Q+�ɹ
���ȇ�&2"66�B���,��y"��qxй�6Sw�GFfZ�����lnj@;Ɓ�8�Y��@	�jM�(����(DX�SM)4D.�1�W/I�Ȳ,(45�6A���cS��9QPV:�iT�UP�(pHpw�����]lq��݂'��ⶸ;���.��%H� ��_�>܇���y���>��5}���	���XT����I �=��%��N%�?pd�>�������m"3�/�=�&;v�F\� Q�sS��B?�������]s'cbg��-�֡���!EONN�����=~�����v>��!��b�����n���r&��I� ^�@Q"��N�ŀ��=�#";AK�fY�-s����X�̐W|�	6U�*��\m�c,l��۩L-�dw/]0t!�+����<�e�S���t��4{u�d=	����@�
���Xɕ뢷�B�߹G�}X�W�:��?�KXyz�Ґ��3�d�1���`�Fi)_�dHq2F�B�/�����u&��%�H`\=�8'~SM޼Pb�F�I�l�U���G#(3���/DD(���wu蓺���/-nR���&��1��#����j�#�If��dfѬn��4��T���������%�jG6,���Rc�p: n�,H6�Xܴ�GK�crR���A �^����ct�K݇f<գ���!�m�}���+�a)P��n�m�[x���(��[&�@���b�A�/�N&4�#�~��j'88�w��{d�X��/���'�#!� �����+Pm���2�ScFqɨ���s�`������R�u�3�H�XO�bX�{��+:`�� �w*�.@�������@�����qnɩ�ˌ�L�j0ZKQ�(��C��|.�̵G�Sm�o:�}=t��@�PT��C�Շ�^��x�gJ���bW�^iEޏ"e��>�r�H��mn�j���z�1�5�`���(��1tϦ�|����_',�B�1bw�lZ�lnf�$VS�v������8��|��6�\}�.��-_�wx�işh�����U��$]�u�J��y	��t��>��s�Q�z�p�R
nO
&�;�\�r����w~ӥ�z����HK����ݷ�_xtf����>)�7���z�Q��_��X��A	�ь��\P�c£2�'>�v�T��<����+x�T�K�p��֗��*��ELx78W�IN@��1$f/�wl.3i4���@����q�Eӈ�^:Ʋ$G�2�!�N�9 f鎼��0�cf��	Tx��Yn��`�UH~���{��H<���ґ`���_qҖ�YQcip�l�wK��%�B
�?�1J3S'}`�N�#��]@�S�\�@�A�3!��ƚ�6	���eLs�4|�T.Uu
�!�
p��4H7���$QL3�������f
�e4b4�\��3������8�j����7��Jn�Q)�d�������M��m�D+�R_��~�o<����V�&��R�M��L ����s���|f�#�X��ݧ'��� J9��9z[�Q)���-G��@��E��Ŏ�a��oʃ0�+. �
� %�s(����l���
+}X���.x����֎~{ϸ�]Ƶ�*��[�Xpة8�[��V��v[�c�/3fMDF[��p�����(����EZ\{��������!g)��[r-��$��͖�����j}�$A7(;�3��~�4Ӌ1�;q#�o] ����4�8n��ƣO���wZf�@�s^v�Wa#8,�b��s�3�FQ��ˡ�J"N�v��$}g��H����<4��*�+�S�P�E������5v�����YCu!�Y��۰��$�D��I!^�Brh��u���2��������=��5����@4���b�.�ħ�H��̸���ӑ����̘�E:y]>�ѨRK<�7�q�寿���<t�.6<|΅�<�/VohW}�ڳ��2���?�����uV5�_��d�7�|�'��O�\��ð�rur_�F8z�Wg�W�وL���:C�S�f�����'W�v�Q���"�	�{���	m0�w���_{��T�5�k��Gᔹ^;_9Z+�kc��`�ׄ11�(��OJ���(�����9&t?�T�}7�I�Z���O�.T���UC����E�c�f��z��_��u
.�����bC&�{5*�?��?d���Z��p���`���>8PU0�V$�V [m������ rR�.�
$mݱ����Ob�>z��d�>�'@�?Ǆ�eV�Ey��Uu
Jvα����G����|�*������K&[�5��GB�J��V���$�E��'���d\dm~�*��ngQ��쟲������[R�:ﳺ0P���W���`�_p�wK
ʀn�O��c�HKe煔�,l2��hQ�a�!� �P�b��c�<����Ա˩b�LL:W�;�0�w�b8�b�lx��>~�����20�/��f������r���~<�ϮE�c�I7:1_ٮ�~�=��X6�ͬe�|ҩ��$b=��S��R��4�q�b�'P��Qkr�t]*�ONђ�*�/��C�!	�REW2�f�G��V61;v��5��U���)�jGZǣUvYAt�d��Ӆf�A�is�͠��,�����b�'����SfJ�:��),�� �e3얗A�:6G}缢�9U��8�����Jʻ/>����O����ﳉx��}�bv�0�y�����"F[z�0g�s0=ϧы��M�6�Cu1��B��U$23�zXDQT
u伊���yD�If�+=���C�w��N��g�����sn]?}':�\�.�C����4�����͎"����e��\��߇*2�K���M�j�M�	>�J��VKd���U&��t1�#qpy����8�}��Xu�,!��-^̱�$���� AV���P(k������T<P��ק���-5��t�� �i�{�˶���UUbN�}�,چ>g���U�m��Е=GԮ)�0�z	?�S�-t�[Ir�WD��\���do�G�'�p��%^m��G���o�B}/ly����,e��r{�z�����i$o�l�AEB/	n�Y�1�3�;�2��bz\��4��ŕ��"1�qn+�4��q��D����'�7�������YM)8ښU��6C�x���@W4AN��4��X~ӛ�٘o��S%]?r9���X���.a9[�D���-PX�A�eM뷻�h`q�)R_V��&*SZ@ݭ���-�L���J+���m�J�����{�NJJ��L|��@Am�*�c����U��ίuލ"���U{�H�;�/�	p[��SJe���<b�1�+}f��mb�Չ+5ݶ|�
G#!p6����3ّ�����DA�HD����l�k�Ur��)�%�Y6~G��4a$��	�0��j4�.:��D0�N�{�lFc&5�Z:QX��ʍ����I��6issj�`0���Q���Q�SUGC�H�6��_DԱ����bW���<ƨ���O#)�!i���iW�*K�sgT�>I0���؃������U�׏���d��H,�5v^�,����^�G9�Rn�EZ|�\dĜ$��Oշ'n�������2k�������j^ik_t;-��tnik�c�G�Ň��"��'��E5.m��]����8�k��*��^|:��oX7�j���b|e���ETG�,�����p���="�@����W��s��� ܷ]�_X��!%���ZvO����N�WZ������^MWR�A��ä��ե<F�b�$��'F�ɿf~�����v�u�������d��1=�[z7�̮8���rl!�yu��-���<��!{2���9��?��U��p�5��+R)yY�.��������W�r����|-����"����ΩJ�)���gdt�^Թ����R���Y/�.UbLM:����|�<,N�OX�_dbF��C%1���O]�fgf""#GGG������������o�1���!G��"%�TvkBZ%��?K �E��5�+�}�թ4w�C�̸��"�q݈.&���<|h�Z�e��#F�Ɋ��2����v��*��f3Ȧw	�_�x���x::��`.��
��{�i�ܦ��P$�ARi�fC���E#�4�������`f��vBH����!�����ׯ\�v�����P���山�Hӯ��֣�T<;hb;��K��q�� CȐ�ѬD�/��%�6?Q �� w�b��9q<̄׀3�Y��$�4�.L�a5z�-@ֱZe�I�ʀ��ʽN[Q5g���ƿd�:a���
�яU{��)�sĘ�tP�L��5V�Y�v�o��X/����@�s��ĸ-K'�3rړ����ѣ�Q� J���i	,i	����a�0[������;F�����/�C����Sd�E�MCk\9�i��]����BcrS�E
zhJ������ ��:�A�va�q�h}���z�D8գ�����~VB��V�ń,�զQ�믱�`�Nk�-&��^�;މ�^;�k͢���Y^i�/��b�^�.�'��m% z�x�X��s�Ɵ��_-���u�'#@��U]��xG��]��ű�ĉY:Ff7�3�_������n�:�lDi ��Q+��K����Y��S�;N7�����qA����-�I��8�O�O���b�Z�\p��p�U��"��]��T#Lѣ`��Z_�O�ۢr�c���$�9F6��w�1����2�.�j�՟dB�A�{���t���w��Y����~���?�ֺؚ�9�ͬd�4��鯟�Qp�f�ncg+��:�+\��DD�~	��/ȃ�4��U�[�Cq�k��n[���6��'Y��w?��[��`n.��k���Y�HtVZM������V��Z�����+��_VZ�uG�q�*o�΂D�����;��?�Y��D�(L2g�כ�������Z��R2,&���
�q�R|�.y���NE�٦�>qOZ \YW��,X��ҋ�OI��\l�^��#���6l?4��wc��ckט�V��_���:�eTI�b�z';ߖ�g[������3���`=��+r�|L,i̓�j��TplE�|*v��sp��w�����v����I�#�ױ��RgwI	9S���_kiIn�(���߰�H�t�� �wE�Ꝙ��FϤ���[���y}��z*P�[(�Y�b�[zd�����q1Ѿ�S�\iÓ� ��b�nb9�UGz���Kf�@���i��Ly0x�d�&��H1�10�Iy��u|8��2ܟ�� I;��2N��g�ع}�
)04�
���}�͗4��,��푢��1�6-��W���G���1�>����'�]H���G�ʛ���ꗝu."ۦa�,=I �������7q�e� �wy�w�
yj�S�X�0�G�ð4��DX���z��w˥]A>�lc���4(�͟W�(%p�F�����c/�?h1:gK��_���}xHc�X�k��L�Hj>���&	^�#[���e\?�J��~|������ �UU�O�I�r��;k��܉�>�4��v[ksKNNޜ	X48W�*��f��$��]/��(Q��߉B�Ȉ�!\�;N@$!6 ����]�=6�˞wc�y#hr��q}M|v���B��r놧(j��L65�f�K,Rk�7)���%p�"Y=v�f4v;�6Y�:S�9֤춟��ty���b�r��~T�k�]��f�Ѡ�`��tKd&;KF��n�Ց�锿�Oc4�=���iys�F3M"��T��[R��l�HGE��_8�E�?�)��Kا~�u �l������	F'^���&N����w�dB�Q(�H!Ha�1?�~ �$�=nhⴆD$ �`	�n���#��g�ʬ�eA��	���菳W��>=e�F�$@�r�rd�m>�C�%_��������0��l1�����Z���z�����k�(�*;�tB���k?��ɂY��S�����}.���6^��n��g�L	�uC��ճ��(s����9-�mF��z�{qj\1��S��p��HpH��!�!!����E�$\nC
�O�}Z��Me�����D��6�v�	?���̓)jv��F�����T�W>��e�~Q�����gv��wB��\:%��"��l��r	����S���I|���/ߣ���	��Iu��MĴ��|!P��q�vu�(���>�N�F��}�-�LZڈ^q�:pQ1��V`������m�6�9�C4��mET�!��l)�|S���W�o榃�x�S�1@�e����� �b��_,�m\�v�lX0Z��~�����
��v@��&�pџw{�m��^�w����=ؾD�.����Ξ�?8��lsq�ލ�=�����98s��o7򫐾c8CK��������9�x�Yq�QßB��G��C�;< ǧ4E�HJޭ_G�0�1RM�?�$O����fo�p�00Kd��S' �©.#k9�ff���*�㓲��민d���xMs>����h�����p�="h��D�ҺA�}{�EEEɩ���c��.��ؘ����rNm555�_�&t��u��(q�,���J�$@��I�P�A�^�$ݠy��� A��I�l�vO�@=ΰ"��^���<#]��R�Ym�mی�Y���4��0��e�a���,&���|�18�|]XA\e��%��� Z���)��qֆ�}yΏ���R�W���8�����)��ʇN6��{0���X!�(��%�4���d�I�A8%�����V���mF��:C[0V����w�Z%9D�SJ��S؟@d.�8a�� ]E�Jb�+�>DÈ�
�D2�BP�#h@�b��J�������p/v%��T@��Io��"`Ǟ�W܏zH��H�����؍�3*C_�9��U� �C4��(@B8FA����W��B�^eXSy��r�G4J�<��U&Tf�1a��I�G��7�\�5���b�ַt74�lH�c�	C��(Pn ����ƫe���>W~������nf[jf���w�)sܿ�Y�S�}`T=ܡ��S����~^Y��Ho�Np(���>�κc���ߋXV"���p���4�7x�JI��.��r5\�6r)�u�N��H��s�Ms�8+�Ry�����qϋi4�nˏ�b3�v/Wo���bH��1�EJ�{��edbc��-U��{�����!���
R���5�n1�A�a�3%�L\�;b�����r���r�/Xc�_����7st]ɨD��h�@��1Lq;�W
��I��z,������Ƕ����H�B���	�����6]0��VE�u�_?��oU[�W��sX�j�)��`&ׅ�~"u*�5/��UG� 1��,ֈ���,���.����cl�Cg�WT�A|��u��1�9^L:�4��5�º�8FOh���ת��C��a&�7c�ذ�����K
�A��ö�;����_�g3�)n��Me]�'�wU'���f�+�_H��젭>;s_�ȋc�n��J*gF�v�K�M��~��e�<'���\L��\�yB�e}����iYzi' '��q�-&m�~E�iy�,�$m���θl�pI*K2w�h����o���������xw�姝�����{g�J��$-�����|���b}Mwbt�����g ��&R�xB<[��z%� x$���$�S���k[�eTV��[�:�����z$)�"|�W��M]�<���|������P��wP�j����DXLj��.qk��z"64���BJ<�r���Gލ�$��7e{O��B�*�>��%T���Wi<<��E���R1��|���o5��vL�����Z�N���x�C+y*[ɼ�j�5��Ne!`dVĦ�F6��]��="�VU��ϿuK(�!�@��a���<ٰ�`\l
�}7'^��X:n� �T�>�^�~�A���0�#{��zͿ� ]-l\\���R`���{��oW����#�ܗ�.�>���*�?A��0;y.C��c��(d>DҢ`��+���q��1hg݈�[	�����# ��t@ �l���p%],���^��E\qԄ@�/�ӵDK!����e���F�;URNзH�,�e�����GCjk��| Lցwnq��w�EO�G���;���竭���Uz�e���$�:��I�G����2j֐ϨU(-�S�'H��Nd�A>�S���<9��c���d�؊����sD�6�w<���4h1j����͕�_%�.�J�%�����0�	�&�
�ȟ3�c9D/� 85����R�V��J�R�
à�eiZA*���	AC͚{��v%6y�rj��CJANB$b���;�4E�yZ���EG'#��!#'  $����Tk1'O�C�+�9�Qvd���	Kf��l�����D/J�� ��=A:�@�{"��X����|���f�K��]Nf�>1d�e���@j	E"��)�!�o����+<:&��٘o&vre�7��1;(&K����iG��ӽ�9T��RJ�ɐ�D�o���w����x��Db�1	$���)����)Rf��K,#;�}7��^�Tr��e���ߌ�|vk��ʯ��JA��]�\n�v��,��6f�{�|rx�0r��wRbRBb|<AK����h��K.33�X�(R�H�Fn��;T�׷��H�x��zr��?m�O
�,k�[w�t�R��a��:��]��#G�R8%���6L5�d��1��,��p��[��U r��P����y���3���з��_�E��U�C��I��+����=���OƐ�
m��v��i�̧�k��q��Y�����4`3^�"����U��忒Y�7�#�v�[���v��#���i�H��
=˄�u��H�K��^�؟��^е�>ȼ$t=�Q�K��vkO���wxC*u�N��<<�E�2����1?�2U��ѩtˢ��\��G�`�����uD���ٿ8FҵL��|`G�_�3�S��QtԒ�d��$�����d@q�5�)�7��F�i�SC��5Η��jV(�0�p����p���#�2�y�v����.�ʑ���s�tZ&aa_SU�3��	r���;?���� iqR�pi��0Y�Z,}�
q~�溺��Z��x����������Ƕ
��~K~	#8|8<~�`�e,b���h�"<r�zAמ)j<wl?��1��̧1�������/��e.�$7 �Ϳ�jg�@t�D�7)M�SR�����{�L��GoV4}�[�7�7����~�7e���n�W�����-&`
	z����ϻ< }+z����U�N7呉~��s�F��U�Xc�r�4�D�#n6��u�.�t��\�::;!�0|9Sp:�P�8V1J$���}l���0�5�ڕsf�V����]�8ᵮU�6ʧ\v�{ {�4�+Ahw^m�+_l���/31�5�����ͱEL盨a�r	d��0-��Cb!(�S`�^��#7���h�0�N��&�UƓA��*���C2�T��H������j���=-�2�#�Ұ��?#)��Q�v�.z���ߥ���?�<U�<�^n+�����>-A�r���XpU抌�~��yח��^��*��JS�x�6����{Rˮ��-WUZ��t'�A�Q�Q�@�N�h�q�U�u�����繂Oo:��|�]��/��*.����=χ� �
�Ջ�[�T�r�Q����/\�)���Q���_�d�s�T��W>��͖��e=]�x���z����H.8�u��<u?�P֐�5ئ�/���<�!�\��� `04s�/�8vfJ�,��t&�f��l�L�q�&����X�2��x������ .�%dR�i3��?X��>�3w^|�]��a)�m���O�ːøj��\ ɟ����J%��B���8u���fU�l�[b�_��p�a�UbC���u��ɜN��q��M�8��ux�(V���.Y��T�5�_C���w��kW�ָ��U�c8|q3w���l��u0�|�:��5�+�k2k�X�7�^G�+	Ny)&8]p�P@�$�wMU9��uľb����1��4�΢8"����V��\��,]��x��� �
i]�s��)�����5�3;�̤NE���G��q_���ex�;�V�%Կ�0BI�����S����j�Yeq &�Q�s�vz	�{`H�'���p9<3�i[\m�]�;���=]ۿ�m\mt^�e�"��5�	j
bm�E�yV.Tͧ�0g�kq����n��(���o�&�1��qxA�_�מ�єF@�ڛ���[H&g����J��3OD�$����? ]����ܔ/('H��n=V��,��Ͷ�%q=۰��#"�#�OL��ZzB�ĨlsK����s4>ۙ(�Ei:�L�Y���1!��\�f
`0�9@�{ËT�{߉"2����!?�K�ƽ"�%A���S,r 3�%�P����i=:6TPp����Dp��M��Nm���S���G��tX�!U>�c�I]YE>H�b"��N���>�mKf\����)�Uۀ�qZWb�L+��+����"��Кyz��5�s?������s�h��h��9��q�ʓq�|��hp�6�T��p¥��B�藭/��3��=���׾Xk�xyz�]����D�BGF��'
��Ef�Zh���1�3���b��u${��n@��U��e��D��+�dr�����m����8���%=['���"�A�`�[�Jrr�-�ѩ����W����.�+<q���f�.�s��͌>�ظ).��� 
wh�Ŗ1O�T�7k���X��%��,�ۑ��D~��F.*fT�b�����=��K�u������J�'�����2=�ԏ��h�����R�������s� :f
*R��������!��w���1����O���PJ`|���,��ԭ�b��N`�i|�'=%{��ʅ� {�A�ܝ���0cMPXuo\V�W���N����N����ltQ�d˩��D�R+�pP��KAk-�WY���e��Vc��M�[F��=6��3Ğč�=]�:t4�=����z��z7����w�ܜ%�o5�a��L���dV4�ɴd2�.��qVU�4
��O�h&A�V�ě����5�0	���&��y�Ji\��F���*V����̃5����o#�Z*Bw[��������E�lqϊ��(i�t'o��I�sl���� �h����"�y���ź��?SU�@(؇���8�D�Ge�xJ�n�\�)�M��E��X�oY��p�Ks�MǛ����I��=uƱJ�Q�<�sX�s!��Ɗ]�H%�T�)�K_1��K_��~t�W���l�@��"o7p�,{�B���p4��^��y~Rr��kOև/��>N��*��q��	b�G=3*�����M<� ��'W�V�\�dRN?|q�Yϋt��׷��:ġF4���U�g��7��2����j����L��/3�-9����}�9�gg���ߛ$�̦%����S�y�%@�&8kF8�����a��)8���)�뙔�H0d8 (#cv���g�^q�*��<V��VZ�(�S��!�n%O2��d�����y�Cn;>�ӛ�?��ʠ����i.��������IN
yee��_�6l�߉��3�j0���+x�S�]_�Q�
ѽ��s�Nܼ��BQzL?��r�����DM-��Z'^Ϗ���D4g+���W{�T�Q��r�]��/F1�˵&�*C$��M���,~C���ōo��~'�Fߴ���l_���S��9:J=w�a��4��mw1����386F.j,:����w������) ~�5���2��"��P�{4F��TD�9P+J��o��d`ޫ�%k
'��~�ܓ�f.��W���:��)�%��(%=,�V�)c�������M���&	Gp=���ֈ�idım��q�8� �*���{K�qҟ1�TR�6��jN�{Q��$=�9߹ ��y�м��L��<!|y6���C"�Y�K�xs�ڊb��w���Sc��?z~@�ؚ�ٔ�ۤ%���^ᠢ'�?Br�ۭ��]�k^x�������Β�Ɋig;ߕ��y�]�~b����{�N�5Öq۳��L�@��YGSjǊ��@_D�I����Bt�[v��2)Z�ۣ�w�n�UԀ��Okn��%{���gW+�Fut�� �eđ9�#L`i3HL�@�g��iOv[Qa�{�և܅v){�¨���,,!e.�c�-ڎ[��;�S��w��mJ�R�-o8O~B���S�[�Р�`if������c�UK�x7��#ڜ͐�_��8�A�}�Hs�q�� ��!.��$�h��ѕ�%��/ QhY��sd���,��K�v�
�9.]�l8�Rq��7?QZ�{���9O�Tkr$6���ͧ����r3c�ԙɂ�D���v�6r�5�b�@	Np/fZ�j�Q�7LՅ;j�j� ��������`������z��|
��6M(������ve�ZvkI��l�rpy�9�j���k|p;�����A7���R��ظ�r���5���0~A����&1��*JJ0�Ӟ���m������ j�B����ycijۑ}�p������ai-������U��jt�-���v�L�j���M�}b���G�d �s�����%��BiE.��q�P$C}CEG�����H��o�VB�����3���=ru<����o^"�˫�1&�<ꍟ�T'���\�,���NE�����B�Y1¦�9��c��o��%���n�f�g�f�p��:�j����.��>�aQG{��R�I�Ɯ�.������8Ι�No��j��/��s������]7:s�[��Vy+G��'�-�{�N�f?��1����PNk�ϵ屴qi.�8�<0�,eM�&h�f8�7n�,:g�黂�1�w���?6%ń�0BƼң �7�q��ك�g�@wɪ2.)�����{z[�N[T����@iOi�t`��.�QM��Jt�^(K9O՚���o�otY&&�\�-��NJb"�}P�1
�)'Q�2QU``���;~nbW^2�����}3-��d��G��'�:HDc䙁�?�m�{B������izA�?J��V�����U�i��ʉ�e<����#o*")���w�i�@_�ܬ)%��ZͬE="O{�y�&Mw7��A$I��a�0��X:�ߋ�N���"��ς^��N0�>��p��V/J���w����1���l��n�:JH�|v��M[:������t'������!M,{�1��DU���"�ļ��S^k4d��M�c6_�_+qz]M��6��n4����FE�9�QD\L�4�\(+#��*a3pbu0m�6�f�Y%|p�ޗP}�$1���E�]>�C�h�c+���Sw�VA��,bX4F8)��96	!��i�����}B:ݎ)�>��'?�{�یک�������)?��NP�^sPV-�7�����
�ﯶ$�zbщ��\]��Jj%hd�Gs;#
�����ud�y���PSv%ڗ�7YA�r'��!
�|Cz3{�6D@I0B �+��c�ZЗ�f*f i�ɼC��=��{v*�c	kc=ea6��S�,e<��ݕ\T��~i��5GD�h*����s��T'9���ɷ��~����r3�s�vG��+3%�����tm#AǓ����l�_s{J�����V<�������s��X��:ڒ6�;]*oG�Q�2l��N11:��_����c^Z"0�\�����n��8v�s5�of��QD۽!�*�K
��G������i��=ڴ3���*�#
{��^�x0JM�;��8��rj7��(��զ�)�q�]S�}R�=�'[>b�V�,�T����H��ޓob4.��w��w�םva���=FՕ�^ �f�C�- J��\��\ED��>	��j|�I�.z񉾲5�f���o:���=D�~쳕���Q����;쭯��1;.��X:)�n�)�Ʌ�/8>���N?�������a��菴{fQM?R�	�{�y���]�M<���Uk�O�J/�)�����f@�ep}��8���2�	�'����,q��]���VV�f���ϗ������{�4�Z���ټ���Pʝ\P�;[�Q�A�L%���a1I��e���ԬQ�ɗ�Mp��q3>�z�K_FE����/�`������ͭ�����(//olt�	A�������mWPTtn���q��dgA�T����6�%Z�k�!����Z��T�f���wP ?������)�F=��c��,v{��� .�W���x9��b��R�������$��� ���r�Wo��W������z����a�;3Fl�rgۇ�o���l������tbS%�������E������:D��S�$����8,{��S���3��3�|��>�PTo�]���8�$N�����4)J�q��p���T<%�6�����E#8.��Ц����ʊ���Md�����)�I�/�gF C��N��L�Q�<EE��mZ���t��aG\���j�O��3�n�M����I�wc,��N�cl�T�I�H��Qۮ����ߙ�晷�̎1&< ���!����bl�MU���;W^���4���0��N����L[�}��"���
���ߘǾ��aB���4u'���E�H��s�Ƌ��/^�3F�)ݗ���f����?�뷙s�L�����_Ҵ\4��X�)z�5Wf!�^�Ge����m������Q�շ�L��Ƴ�g�L{)\GP���/C�_.`��~+�a�3�7���́MA��,�'Hm�x
޴Z���ȢSL8�1Ԃ����y��c���.�p�����DdM(��&j���:50�IQ��$u�е��
v�i�ǖN���&��B�i=��X3����_1�\�ڇ.3�z���6'	��=���t(���O��dIvy��=����2�v&	��%�s�b�5r_���{B}N�%2L��d�ʗg�nJ���E���Ps��l�JE�;�i_�=�����"X��e<Ι��q;3+�~�r����Ҩ�X�Wy�L}La;��[�9�z&��я����Q�UL +&�G�"WMd�����Fq�꼵��0{Y%[A�<�b-�����u�+:zc+ ٫	�/�׿L�E'Szdsuu��Y�P�ۢH���X��LŜ�!1��V�A*3�	[��� ,X�ׂM ��Р'H	5����%��X��|j��Pכ�d���	�tt���OB}@a�Ua����
�$�c�o��I��ƗEe�w�!�^З�Z��F��K1^�����s�xr�7�$Rٌ�ƕ/z���ֳL!ۆZ�h/Y����^����d��]F���k@�,3O��2��^N�N�p�95��$^�7YM؃24�N�A�ܒ���]~ �`�����<�4��d� w������R ǜ;���\Þ�~������#��[�<c@�0�;�;����!�p/D��D$ء9w�bџ_��=E������rC�����F,� �
���"��J���nG� �if���y���K���G�h�$�M %�[�I0�C
r���^��Mj�\ �}�����+\ᯢ����U�=T�k�1��gi �l��V% 5N_��'� ����q,�l���"�LF,Ѝ_����X�-V���u=S��]e���쭤�����:5`�(��&�5��e��2&�SUjv�hLB��0z^f�$2r��Ytg�|x�o����R��_��UT֊H�� �sc�`�<X` AϢ��7{ �謷���-<?+�?�� B`V�e�8����h�Xj�p�VM�phvG��^�٬�_��c=�W�ʃ#�hD$`
�st�?��|�^�T�������?DED��HO"�G��ϭG�:aQS�G��������` ���>���۽U�����L��@�l
B>�O��S-���T;�bPID�W���;�36_�ލ�B�h4�U	,�A�T��Zk�S?AM�]q�Ȗ�D�� �!(�.��8^��B�,\cZ�"���V6\�e8�y�\��-�#V�?��׺;[�����UF&�}��hs0	j����ʃK��r�8�7K.�7���a���q|�/���m���������������7Z��f>�{��s\tz}=�*����i�y���PJi ���i����'�9p���t?|_UfF�K6>\�/��ha��ʞ�;mVh�c+�г�"t�ktvE�7�����Y@�8�'�`��S�np���Z �*Z0��&�s��k���_�������@d�_+o��{<�eZ�Yj�iZ��ojn �{��r�[Jɛ2��b�[�#\��Q����V���/u��u�o����~��C�����	0_p�"�5�!��CӐ�1�5�]���/��=W�G���2�ʤ�=U����U����5��o ���Ƈ�O��e��/ږ~3a񻦢��+1�<�kJ�����x���(���gY�%��Sr����!ׄ�+( �.���B��>�!�e�C.�Ŀ�Ԝ��'1�\q@���Ử�N��x��d��4��������ԧ���٪���i�p;��v/�-^��ֺ�2;�c&*�v�$a�%\\ĕ�a��,��˒��*��t��v�&�	�e�T*�V+��MMM=8rssKKK���@%--t�&��l&\��av��.� e�?���k`��V�CSc1��f�Y��^��لNҩ��h$���&�9鿺K��cj�#��Lq�S�5�����-���5�|뵗��������>x���ڴ���%��l_;y���=&�h>����Ɔ�ꏬ��齟v-��ݟ�������˲v/�ص�P3?LͶ���٩���R ����! r	�$K����g�7���Ύ�%m���m^ƶ���l�_�sI횙�=M�
Ui��Du�G���x52.�""9O e	Q�H������X0P������/؈���fb�o	:��C�L�`|��Ǘp�(��0Y"SHg�F\(R�Q�T��� ��K�v�ܩ�:��FL�B .�P+��d,;�6In��)�#����v��<+�>Yؙ�u+gJ�f{
�3�����D�S��U��150�J�E���&P��%��M�e���-��	vL�pM��-V�B;8�X ��ɵ�ѳ�1~Gc�ަ�SJϴ��J�_�ٛ�ܕl��5lq��:��gޛ\����W�־9���Κ�/חݯ,���y1�{�j>�Q���R�BuH�:�ԞӘ.i̗T���s��ė��/ZS��o/�'P�1TuT�y-���Sެ��^s�3��}֯K'��Pz]�:N���#t�Q��Wv��^��ϑ�g��3�9��]t�)<��f�N1�'��t�1��s���b��Y�x��� ���'h|�昈s�G�'1�i\|V)9��W���N�dP� @�V
��e�}R�n1k����Cd�ws���}�Q�TrU�_�堼��NK�G�A�ox7��M�$2��`@�Z/�ꤻl��F�b�I<Oϟe��0q�؝FV���>AS�ev�D �k�mB@�C��Dh�Ci��m`�i���S�s�s淔��2�nnOa��8-!�kNu��mJ�Qf҈�*�J��BKi9U�S(��q:_�dc:J0�4P�1q�h�(.�EEH|%G�Q��,R��&&s�\�Z�j�2�7����bқMF��j'��jTj��"b0=H�B%*�`�JN|�4�0�ۑS]ٽ�j��¹{2f�O�9��u�1�k�E�˩�.�-;���lʒ3��^u9sqW�b"� *�=w������Sv��6k;���2Lީ��fj4O�hnYcnXf�Y`��c)�u�L�d�Ƨ�rl�T��m�[�Z�Y��k^�<ل���&$�,ʷ"E����pX�hj %~�SP�Uz��	��D�I�6YX��@Y�75-Y2P��H�YfxL��yL���f"CM�L����\n�Ra�a5�Z��LL�ב5�32�!����~��VV��jӤ�YxK.�l3e���l�nʐ4�� ��)Sܜ��� 0�LJ���S�5p�Mw�V~�oԓ�����)����B+�<5�J��KL����B][��)SY�(M��6_!��1lR)*<&"��������w�=25��x��]PP���	Fc���%%%UUU�111�`0��=���	N��vxh����>Ѡ��#:/�g��B���.���O>S�ۥ���p3V%�85�t+�k����~������*������iHDa4\�41Cў�"	�h:��9J���IS_�'.b�3<=����n_ ׌r0�6��8��{��m���
�<� 2"T�͉��Gǐ"��â�橑߲���[��r}K��q$�FEE���EGG�� ���۷_�|��իW�\�{��3g���v���r�\�R��M�"��ϕ�K�ľ�V�(\8p�9���\2�����Ԅ�@S䏩�����H�UX� �
��+}��)w0����é�rA	eMC��9�xk�wx_���]L$��Œ��RSʴ���д���/)�mF�uZ�uj�;����+	Y�S����8} �O�my_��w�545��z����FB��Yg7��6�e�/XfA�}a�[��'np��!|�ﷀ'�~i�vF�Q橙Za�R�X��u秺�fpQ#C�Ə0~D@���Q#>$  hĘȀ�B��X����b��iʂ��嫷��������Ke�D�5���),R�C��
�z�D�)"H����1b���G�x����G?7*pĘ�Ϗ	�;N�b&���IΒ[q��$I[���xd������tץY���4i��T�.E�4r��4$?�SS�"��֔��3���mN��jW������G�N]��}���v�?{r��Sݗ�O�zi�k/�ܿ�v�L��3�/��޳e�}�?z�o���o��dh蝯�:���{���q���+ל:����ݷo �޽�.��~���G��<�������6�ݻr˖ūW-\�d���kj�2��=�4^@ICh?SS��Ø�%	���Ȉ�OV��r�߬��U�Wb�
�
�sY,�z2i0:�8�zO |G.�S|�H?�����|o��de����k�4��b��^gx_�xY,��e]fR�1�WDl��骐}Mȼ%bߗp_��o�wp�]\�B��J��F�;���:���7ӿ��o��o-��L�o���5��!\�aHg$bgT�!��{L�-&�|'ǿ�}�l� 8�[��K���b�o٢�X¿�T����9��u[��mC�{�������Ͽ0���^���������WKw��c��E�?vV�,��g�E!�(=C]�:�|V����ֻ��;r����/R�c�y�s<�%� �%@w�-DzS$�&_��S��TyU���'$�r��Zu���c�����ڍ��$U�bY�bq*� �����4�yY*�5`V���59*@o��'[ѝ)��.��.LN�LJE;���$Q{�p��y70��}S�&�hi�G�h�c�Tׅ1r�K��01����A�b>G�db!�Scj��A}��΀`���A�п������h��b1�H�ɬ3[�6��ᴸ=v����;�\ Pq���^�Uo��L&�^�4��N+aj@�Ǣ�d|�B,B�L	��DX2ɤ�5��iI�u-hJ ���Գ+Ms�-�k��5fF�"_9��5͂z��ۢF��&ǒf��V����-������e45�':�khjS0�1<g�p6�L�@S�̳���<5�W�XZ�����5+�;V4��.�ޱj�{�.ڱf�����Y5�SMͳ��f��cj�z�e�����g���;/�֝�[�ݵb��	��:v��Z7�������i ϊ���+�5�$������17�瘚�m=>zS{�Όl��l��l�M����/e�\"Zg����/*�_���pIg&I��벌���c�ۘj�y�����b!�͈"b�)�1ԸX ]�6�F��às�>�%d��T
B�A��ɔs8
O%��B=��R3��
�R�P�@iS�=��K	���v�E.�Э�D��A�Y�dƚ��jV�N�b!^^{.>�D�[��)�w 3���J��r%����=��g �� �k�U\0��g���6�	M͖���]�I�S��y��ط��&�xt�]��Ŷd��b����{�e�u7�jN��}oOo~{r��m�/֖�,Ⱥ��i=l0�jw��{��ø���tAg���\����ݷu�-����uC㹢v��[���������߶v�nҴ�L��t���_1�v篊[^�/�(�������C<�8=�]�ϓ�gI�
���!8�i�I&!kN0X ��y����4�9�S\��Ԝ�qL@�9�@��9�F�k$���h�sf%����
�4{%�G����E��a���sY������%\8/�����{��B�l2Wq(k��"�:��eo���e���m.�:�|�	!6~�s�9��1<�4��tY�O����oj:\�����.���陖ŵ��z۶̞4���,ѝj�9U�E.4b\���D踐�	)2��+��(M*c $���:D�Ju"��b����x� g`�ł�0.�F��EG����9:*,*2<2"<<:Vߎ�L�-`�A��!(�42T�ɔ*����[�y��3R;��;��̝�͓wY���Ny�v�>��;?�X���O�,:��� �$�;���$�g.����jѺ�en��_H�w�1}��s��s��}�a�K�V[�[�jGC��v����^��.��L�r%ٽ9f{���1�F�ᡩ�ɶ�L��e�[�Q�/05u)�'M��үi���R�������3ÙYm%v}�0�)\�4��:���]���75�r �-)Sk=�e��bSS��&CMMs���oj``�����?��QM�H����0�nj�˚i0yJ�nZ�rz����Ej�V�f�����������-��.�	X�U�T
�|
e���"�����X2�M����4�L�͡��2T�d�`0��O����****//���C4�^M�������`��� ~�\.�� �A�ej�d
45䨘�Ј��0�Ԅ;tj���X���9$��'�Y15��cj��ϊ�����<&h�<�h ��Z���]�[��.wL���`jh1��hjbã��12M�(�R�D��B.��d�(T
�^���興���X�1�Meee;v�z�����Ay�֭3gδ��gdd��a����75J�R"��M�p���].�vV_h�>��Ձ����SC����I3�9�:�_bjZ��֬�Ag������ZEhj��hj�Ed��N��@S3���]�Y��������V�C"�5��0���Uj�����i��Z�������75แ���:ۼ�������}M��dÖY5��[O�if���ܷ �T9�D�U��\�l��/�r�8�&.ds���b��ᬠ�1�q�ƒF����%<	�0D�E-���x�>�j��kS�S*��:����T��)��,��;��O�Q&�E�vDc��ǋcs\a�86dD���c���$�Q=ZEQ��4�^�D�~*��,S#!4��LMI��<S[��KO�:]
�IZ\��~ߖ[�NY��{�����>wr��S/_�zq��k�/5�?�~�l��S�;75ܵ��W�#bj�~?4���w�~����w6_:�������vݺ~��]P�_����ٍ�Om9sbӱ�k��Z�k������lY�n풕�K�,�=m��Β��&S�˒��$�g��4�ujJ�"�SA�15�M�N�|�J6 GWbH�T�R"Z��e37Pȃ�Q'(��B�;��#\�;��OJ�ߴ���C����!w�_5ƿ��_茟�����"�;\�u���_�t�\GطP�})�%��u9!k�U �ЏT�_k$��H>�H�j���f��i��a��d�J����H3��N?����F�����gj�W����N���B�O��+\�1�9_�g�����9�eS�GmCKw�<���W����=t��?����]�Y�����f���V��4�J���x��e�}���%o��־w�Jho���x��"�Ty_C7%45���;"���\�##kDW��\FПkj΢�YTyR"?��G��CZ�~�f��X��9Q�>E�:Uݟ�\��\��X������Y�*hjfd`S3Y��zyO�# �yx�vV렱�-�s�+��B�$]/LԊ�u�N���P�#�!<�ķ���IL��42D"CA�й���LF�	��w�n�d2�t���Da���tY=^G|�+!ѝ�䁲���]n�=��j0�T��O:��l�����CcH�<�<��F̊U���ˬƤY����k������̀�kj���iVu$�LJ��fx@�����g��l[\�}I���u���XѴ���hj�|���^{��W^�?x����W������w�<�o�ʅ���nYټ}MӁ��oj�yj|u\W��15������'4����[��gi��65�w�M{R� �v�qf�n�M�֛4ؓ8ؓ e͖n�/�&~ko���;�힗�g~���y;���92в{i͊�9����BKK�����\�X��X�����5J��#�	�4>�
��(\*�ͿU��ϕ	x ������R�9� A̘Ċ��J�o�_�[�����-$��N2�MX�Q��K�Z�G#t��n�"�ۤ4��j��P�U�a�1*z@�.�%�YI��ήP�*�{�%��t ���ҙ�XO���B=�Ѻ'����%�f�M�?���ձr�sU�ku��4��4�{�'X��5���f����z��Z�`�wS�mC�qm�v�W�έ���lr�7:[���Y�S�I7&������ɟ.�������u��=����nf_HO<�>�rlð�2|/�>�5��YϨL�p�E����vQn>/3���H�e�����#��0q���.^�͚�_�����6�}=���#�4��K�"���yx�c��{��=CaCNS�g�ܳt�i:�����b)�_�<<�[�rxg|���}R�Ƀ��c"�#>Ms��
��9�$6�>�F�i%'�Y��C{ަ>m�A�!�h���G��-a�BY;��mB�V.y'����:��౏	�~Ss�Nc���>1o��=(dn0��+8�|�jc@�Z'�nR!�M�]N��b�E�H/�����IV���i"�~z� �*���4�� M���%nwI����!�h�ڑ	vqw�y^y���3+�RN�V0�j]J��" =B̈��%�X��	)rG�
���9\��)�S�zT�K�|�J �z+nv�A	n�Q:GDa���:��`R 4̆|�1!A����������s���H���JL�PjUF�ʑ�*j)�9�ѹ2i�:����ۼ3���I�"m��9GR��X|"{��������g �&��[����Yr*}Y��3v:&o�vn�v�[-��l-P��*f�J�����y���2�7���0Z�tF�Vg�i�F�ڦUx�x�	O5�����B;���Lp�\�*���F�ti�����:0���'�VCȚ
3A�.�"�j��35s�2�'U9�ˬ-:hj2儦��2�~S�P��X��M����j���X�ዩ@G���km��F�L/�N/Ru�������zלZ��RSw91k�Tl�,6t雳T�I�,�̩�D4��3���(�/O��fȣ�O`��75ğel,�N�0�LOO�랊��JJJ@%55�8�nj����]�p8� P1ǳM��M9"L�&iQ�['�r(
݊��؁9�����YU�9���r[[��2�0�Lb���{?ń{us�4_���:�J)����d1��
�KTT��Ĉ�d,,,ܱc����oݺu�w�>}z�̙���V��Ԁ����:mCM#��U�^��p���a��
��DF����jl��T��SSda�ܘ�L�-��,R��0x��M�c���45SJA�>��9�6~NCҜ����Y�	=���}	h�4���Nhj:K,���r���z;M�_�@˳bj�������c���p���PCX!���=�����i����
G[E|Y��m�q1�oc�i����!�Q���q̀`�s�1h��ηd+��Ⱥ�1�u��o���˿�����/��r��o]E����KK�,���<�mvZ�{~�"� s��=�2W�Мh��Gmn��kM��ۓ�tQH�ŊE
�Q(�� �V��,K������L8�&�059.AQ�"/]�����e&��uF����;�͟�a��c]85�ԑ�3G�.�k�|��̱��Ξh�xz�c�[���\�ʃ_}<��o}���g�9�½ugO�ٹm��=�=��k�o��~��Λ�6_:?p���'�?����U�w�ܽ�p뢁�s�.�?��9��gN�Q_Q�`)6a�$KB��15�,ʽ&��|�
��2�r�h*\%����(���Ǩ��"��8��B�������j��t�omޡ��!w�?��?��Sˣ~%�^!�y�[\�6�,�r�C=�g\E87Q�]�����"&xI���B�U��k��ſR�~%�Z)��Y��������W��-�y�cXg �A)5��D�������J�J��J��B�5���u�o4��I�?�d��귔��i�W��s����C���~��}��ȗ˷��o����:��#w�G��wd��sQ�p����������J����|3�I�b�����K�33�,&K�d�[�Af�1�c�'q椓�t�4sw:ѿO���a&}�~��Z��k׮�\���9���7z�6����MV�U�Kl�8�m�%2�.�q�J�E#>jj�ԧ�d:�
�u�C�Q����x{?-1��8�3�)��F<o�N[%c�H���%<��u��x�ܼ��Ǜ8��5��%x���tP��f���򈩁eM�����(�V���b�E*�E� �h�7�D:	��h��0ķ��i
�E�өKip��{n��3�L�Ã:���L.�hF��j3�f�P��j�h����Uo0(�j1T�F)�*er��M�P*�NEE#�.E�N��Ӳ�o�4(�5Sך���+�RQ��ۼ���W� �J�0^GeBUB9M����rJF0�Cl��75O��񚚹�|��L,��'�8��[Z��y���^��q��O?��/~�Ϋ�>z��٣�k�F:G��ȝ�=9^|z����<���yRL���Ԝ�=���c��+I��-��!�a�#k`󟘚V�l�0���oe�e��8Q��!�|��X{ĉ��]�G;�OJ]�;;�3��Ud�MS�ǫ���j2�U��4w~�#���I�
&IB'
i$�!b����S":Yʢ)y,��P��j.�&�����Hy^�.�"xԮJ�C%t�צ`[�t��
.Ō���9h�q4�j�������w����`�1� p!Ց�ݛ#oM�7'1���1��Ok�nJᷤ@���i�t'��(P��4�9�2�ǹ|�)�X����Y���D�~"^3)?��
���)�t�,�1��m�.���嬰{{2��,��@�Կ�Q�nKٛ{�^-ͺ��t+9�ZL���S
�	��8_tZ 9/��e	���+t��l�,8��#pϑxgH��D�i2o���yi�ơ#��:�������c������	7��%<���/�T�,��H � ��!YC|�jj���@�����Q�48�*k�Un��[������Pm�U6�kj���e	sMι�^Չ/��.�iN0q�����cX�i��%2��y�ǽ�㬳�,�ii���$�ƈ��ĐaR�l�!|P?�S�GX�)}^�=�Q0���N!�Y��BEj S#�<t4
b��4�J ��r�B����0���2=�YC�Zr��R��V;D�q�(.V��o|������d"|t�/���r	!2JD�(�$)��%����
F�D��h4���	�\>��ƁQ"c&�ݩQ�y�QK�"��c1!x4��A��D�C���|w��������;��'0�l_ј4O��|&���f�1ʜX�Z?�8�4�4��@��O���	�8�u>�{)�w5��: L�{�#�-�y¡ x���O;[OZkg��� K휩f�X=&��c��a]^�.k�6�][+s��ybK��/�GJ�.�b�P�	�R>_-�o25���b��\���#?�^΄jJ��`Ɗ8 �S&Չb���R���n�`/�(�*8��5��4%lj�2�PXM���ع���55�����}y��0V��b�۩Y���0 65��y(k�4�h�G5Me,$��Ԕ� x}�CM�(mL5%���PMɒ}���E��s}2��.U��$B��0B�a�F�&UHFP����ٽ}��P�n��
ש��HpEa8�	6���P�Z
���f��펏�O��!��
����:��j�:��w6{���ݞۓLMH@ � ��@�%���yf�o����N@S�c��#AKyJ����Ԁ��4E}��9Mݚ�oHі������"���~� ?�����ؾ�$�e\�B$s�tppPh��s0���:ph����422rvv�ƍ���|����rOOOVV\!D��3ljX,8(���R��\.�5��kj��Ap`P���ߎ]���� 0�ݹ#�o	 �a�B�SF�P��5�����
à |R���<��a!���B\\Y��ؓ��MMS��-��Y��,ݛ�hͶ6g�3���l3L��TMe��<A�HTV%����o%:m���(�%yMMk��I15^5�����f_؛�n�T��W���iN�4���2$��XAy��$Ŕ��k�B&������=���+})� �%
��9����JsAGl㨳��Z�W������Y�ɛ}����w�v��z���_�7|�գ�?Xy�z�dr㡨��m WI�)�L����϶������o���$��c�qF>7ެIs��D��{������cMM���2P�Z��ʵ8��hcamn��Ѽ��#Ý�g���Ν,Y=_���܋k)Kg�.�d�-�/.�K��;:3q���7�y����뿾��?�����_yixm�yzb�±�7�?�ɇ/ݙ�y�37�\>;�x���ى���N��k>��~okMmu[c�������4E��Pr�R��I15�Lc�M�c�0H}4�0�4J�Akj��q�����(~�5����֘7����/
�Ϲ���18ЙoQi�I��x�M<f᷌�_�]!�o�qwY��ِ���½�&��'�'�} ���'��ƿ���� |.`�Z#��I�g��O:�_u�o��o4��rC��d�25P��;�.����� �`S�!�o�T�~IeN�'4�&��S8Xc�Y�UK�Ɓ鍃�=_�~U����=��>�~ķ����ǋ^f���m@fgfc�����)��М���y'}�����o��W��[��0,kn�!nz�Ea nR!n�r�����f��\�q༧3R�)���Q:k�O:�GB��a�~��[����xxRLMk�ͣi �т�H^c8��ͮu'k��Pb&<	PA(7���zB���ka���NI�����$L2�%@��D��jHx�STx��a��8�Cgv��}��������G����	�,�ɍ�J��Fn2���3�
p8-�.�6#������&��l�h�:�V��*2��E�P� ༦������)��5�(��NT�_ߙkhπJ�<�NMg��P�55���͡4p���J;`��6Xi�+�,�¦f��8Te~���"b�S����xr������Ys�r`M3s0w�@��?��l�QS�������3�+������/;�;՟�0V�0�wj,��h��Ð���?�d>)��x_̉�XH��Ǟ�X��x�VA�e������VY�d�m��6�L�e��5P��:�t�}��1�z�9�xk�B{􉎘�6�|G���c������1��ºJ�%�������<wU�+?Μ�TF���*�����PUl
�k�,R�C���M�����,�X�2� ��I��K%U�r�f�
X���N��m�ӭR�YL6	�F�"��85�OE�U�wJp�rC����?�g�-��LYW��=GҜ�iL�7Ē���q��:$nR8-)��4!`���l�4�-�4C�F�p�i����\��g��2Tf,5�¥j��s�G��㩺�d�x�j�%;bO�e369��:k����ZE'\��󍂘W���������w�V��Z�Vc�{�T�=(�}P�{-:f�b?�Ҟ�(Od�X�St�9�p�%>C`�@SO���c8�$�{��Vt�>*�{#������;tM��ҞG0N�bN�"�c1�%,f�ZF!`V� �2	 �U�&Y�)vf���j��8��4K$,�hVh T9�S<��"��)�\HӬ��kBƲ��"c�)��4��ZѺ�wNH[`�3q�4�,	��� 3d�4>h��>K#����%6�y>djV��sL�	a��#"������~b�\�A|P1d���g$̣*޼V0,���1�|d�	���ˤ�J���JI�VA��ڣi��T8��BK��25FF��V��±6Pd��Zl`��R�!����#k�(��6!&DJI(���S1R:N�"*�$����R�,H�ȹd�,�L<�K��)B1C"c�$L��.W�L�T���v�N��bp(�`��A�cB��@2��"��AP��A�!�C�}��v���$#0\2���
�r�ک�%:��Sj�"+��U�a�G��'ݍ3�M���3��٘��ѝg��'�_J�]��,��Q�c�΂�䃫)�� Фw%�a.�qટ��LY+�lUӎ�)[�a{Ѡ-�ג�f��U��$�t�>^j���"DJ'_j扴|����x\�����r�S���j�����M�7�	�4e1<0���fSS� ���`Sk��z,^S�KW����((�&��Z��lj��1�V�i�H���&�F�e�k\�-�汚�جi���x�i�ep�<�;��($nN�a5���)���\���*�qMQV'+Jc$�.^��g��E4���۹m׶�v���B#qx,��#Q h����`(v���:�D;|��w������[ZZZRRRll,��æ\�����z��j���S����>�=`�6|�.�_��9�NM��~���Ԁ���te}
8�ʖtMC��2N�n�˩
���������|��v���؅�b�r�P-�˅b&��Gcp,2�1�q�Ш"�������֭[7o޼p�������Hyy98r����65��H�R0��฀�
.���S(��l6�F�Zש�`� �����	 ?<�;����&���T�A@t�HJ�?fj
\4���$S�Y�(������&IQ�(��i�27�X�x5�>Ӹ'�$R/W��	
OX��!Jt�� ����xI`��В���uj�s���~&djr� ��T4gJ[2� ��T&JJEI�K�U�s��hJ��bDb��dK/�J��n.�3���J��msq�F��L^�?v��ح�c7���ݻ�jә��n�\|}������������z`�^����W�G�����N��k��6��\�����d�� e��L�S.M��SC5�VI���=��S��`��yNI�&�,K�<,ɞ[��4�U|��lt�~a����G��Η=){}%s}9��������Eg�dLMT.?�ƃ�76>��_?�����o�������L:{z��7_��3�^Zx����^9~����b��?�v���������C͇z;�zk�47�4W�Gī)j^���($�15
ތ�}D@�R�ؔ�L�!y�A9B�AO��>|�L�bjx����?�K~#Q�Mk�jLί5�(���~�������z��x�F�G"��c�C|υ�,!�ֱ�7���Ļl�K̫,��!�]�m�6�u:��m&�S�W:�ס�H�۾a3muz�Z�!�-��M �+��W�g�φp6�!C(��6$ү��?�_��R�WB�x�_��o+�w���L٫*��
��_����?���!��I��
M�Xd{��������z)���?�:N��䲍���������d��$��}���E4��zC��A]Eæ�&��
�6��O15��"�u��=��O)%'t�Y�l�.sJG\ҁ0ѡpсp�����I��-��%h�Z����u�`Y�%�f����b3	��5gj�j5�zR��^��JbT4!cS(��542lj�D�7��ﳟ(�\N��g�D&�������}�	S���2�H�WYmFW�����6��b5��:�̰��s�U��X-z�N�QH�|�L%�0D���PPjY����/2z`��U����|��i�P>�NM�G���O^Ms���xS�I}��`M�==�Ԍ���A��{�����L��jfd�̞=����<����������W���&�L���-��:Rpj4׫i�F�O��9����q����a5'z��f;��aG;��;ܛe�S}�c��:�n@����I��C��3��ن��F�|S���c-��[��։�l�{�;���������i�﯋�_�Qٔ�H��ŨS]��6Ѧ�1��5�P�!� �r�]ʆ'.%<�T�"�"�p���
`�J�CU �s��b�����T2
�MF�J(1�"$�$�e@5�"� 2�3Q���js��#_ٚ%jJf�Ǔ�c�-	��Z[2k��xp{��-Cܞ��ǓW�<���`Ms��2Zf���k�_3\b(1¦f��t��t$�8�i�L7l65�6�U6c�͘ųZ=c�-�)������o)������{��_�Qo㧽M��6}���ž�/;[�.-})%�����6�޲"�.	K<�Ov��>���"�OS8�X�<��@✧k�0�w�2?�o����w��{������:A�H[����c�C��H�2
qr��E.ar�\��o}�wՂ�Ėh��8�%<�"��B�Úf�JX���U& �xj�\��/��B���Y�s��u%�,e�摏1�G����R��44 ܝ%"O�p�)�e
i�DX��/sX���|��r�N:J�M�P#��|�AB �!�OB�б�|ʌ�5��Ψ��b�~!�����!`SS)�T�qP(�G�@h(�*-65�H�T�F�T�
#��ĄM��5%Zj��h�ns�\L��#�-l3�GE'*�9/��`�L��E���rID����M1�\
V���x>�
�pH ��g�i��\֨(�V+	��������Cбh&�"��d"T9��F������@���A>;v�������("�@"�hQ&wVh���>wqox�@L�Xb�LJ籌�����zOg���8��uh-��B����ţ�J�\��K`1��jJ�����1�'b��S:N%�I㜻f�V6j*����+�D��,�sgu:�L�eG��m�H��IL\��˕r9B�;S�&Q��15�_V��������O��B��|wףif���^�G=	O�\�25�iP9a��p-�E皡R5�a���W����T`ߓe�Jו$Ȳܜt;5�Ad:�١�JzrA/;�I��M^3x�Uq<���4����iZ�U0���}Ms��%Yڒ,iL�:@5&�;���,�ej�䍩*�_�M�)u]��2AQ!�7�l2����caS��gwl����D!�4�����q�
	���ސH$�؃M>��;�΄�����,�-555..l��n\��5�T
����}���� |��w��}v��<��m�a�3�~J6�.�E��1*J�����w������$yS��!E[����� ���h��=`�_��](�@� ��52�R,�0�D,��yM�[J�R�BAdd����իW�ܹs�޽+W�������755�C ��v����Ԁ	|�_[��J�2�d���R���78jh4���`pP�ٽ}lj��o����x�/����	v	��� �������L�M��� lj�O@T�	65�f?5g�[sm-y��\+`��i�2զ�+�T�q��	+�5�j�k��h�d<`Y�����'�U�w[r��9�'��x��Ox�9^S�yk��9KӒ	�OC(Qc:xs�{R����+Hvf'�'D��;B-�Xpj�o���:]п^>v�f���3Z��;t�gu��T-�Y��~��#G.E��<�B�܍�7�N�*��Vq���[���w3o�b��_|�����Y�;|�x|�z�r��eG/5��Y6�QsȞ�_�7>��jK��#�r�M���k��d���3��)15��q[�N+�d�JuLK����b��Ğ#�G�+f��O/>s�d}����+�]-�q=}�pq�rq�t�x��s��S���o����ӏϾ����]� �@~���������s��[~p�ĝ[������9=���t��Puo���##G��t�t�5�՗��G$���*n���,�|�:5j�I%N���y�~�����0�2JƏ"��}w�	�M"���~������+��\�a��ܰ�m�S��(��J$�G�	����6��*��Ԝ	�u&`�b��B�M:�6{��y������������������`���3q��(?�J6�)1�Q��v�����k��+���W|���q4�!�4"��X!��M �3O�P��X��D���l��09�������)_�ޕY>�9��?S�>�8~$s�Hd}�*{�(��&��"ɽ����
��ME��57Z��\��W�5�t~&�|�$��f�Ő_�aobP��^H����E:��?#�i��<�����
g���1��#�첑PɠK�	�f🚚�1��!lj�9u�	��Z���L.�P`Rn&W��f�e&��YZr���oūiz&Zť�X.��"�" J}"�)d<�B�P��°��T��|� �x0�8�fsL��G�
8�H$"�R�ӫ,V�3��v�Ý��Q�n@dTXD���J���tMF�QC,�Yt"���BT,��a����o2z`��'A
�Q*Y�]`��+�r�]Yj��,�9��3v}�i��X����1�O�C����{z?x�`��75O������L�f¦f�`�􁜉ނ�������(���?}絛�vm~��챃C����*g�K�N)<q$��쓇�N�<�4'�!M�$S�0i���31��9q����f�://k`S�dY��k��k�dM�Փ�i
�ntyZwG�7|��������d�e��1��k�<��`�遼���Ѷ����C	��э���i��XMA�5;Ғ���(����&\#p��a*�K�Up `�R�!T,�05{3`�r: LB�L���T2!M���T��b���H�X�Xa���*�N�9#�/B�΋`T�
[����~K*�1�Z�oK��'�:����,Qg�do��=S�/G��a��y�<lj �V�!�W�<%j���_l(1����Ǌ����d�	65Gܐ��r*fCUGC�'�c���3���Z��ɉh���7���=P����O�[?���H�����P�/z~���aE������s^KL�튺��]R.�Tgh��<Sx�ş'Rgp��d��?k
!Y�^�)��h/�Nh�q�b��\E��}��|���c/#V��!�b���B�,$n�!�a_��@.� �B��\B `k�(�j��+ć5�T����$��(�l�E>B�\� %��EM�]�sVd�e)뜐v�C<J��j65��1�5d�i2n�F^�����U�
�}UȻ�眧�OщsT�8	9D:�؏����$�07)���ٳ
΄�5 "�𰩁Zt�0U
l�[�$���Fi��������J�I���M��@+דPX���6�s�lT��,ک��yL*XE'+h$9��҈rYɢ��4-��`R���F g;����3��D�|>��&��x&��T
CCM���11�����p��	
�E&�)D�OBRP*Ià�و���hTp2�_��ݻv�����͗�!��"�Do��;���iu�%=q�}�5�i-����<U��t�t������ٽ��gӺN�v�#�g�?�{p�`%��hT�tX����ph�Hj۱�����ö�KA�)�.�G��i�;��?<�+<�ݕTg�*5���lirS��)R��$&�@����,>��R�z���9ӥ�G��Sw���>�5pm��8�fS���� ^So����lj���*YQ�$�N�Ҡ�s<�6�0i)r6�Yk�M����h!���f?��qRkj
7u��yT���I|��Ԑ�nNS�����[_#kJ�$K���DQK*$w�ċj�%���X\��m��צj��	6�M��2�\6��w�s;�}fǶ�������a�$��!�����oAP�������>�h4FDD$''gee��䤦���Ā�=���5p���K���(����yf���簁;X8_NRQ&���S��O����Դd���.
�iHQ�$�3��MIG2��� ?������}�o �19j�\%��Xl2�������4p��@�$����x�ĉk׮ݻw��߾u�֕+W����Q �`׮]��p�\����H$s��?�Ep��J%8Xp���x<p��!�~�BaS�s`��m~��#|p!>\2R�Ãk�p65	*�����?) �3R��0�����+k����ͦ�:Q^� �\E�,s[��5��}�fYS���HT��J���`�$@���z������ �G[s5���'��t���	�����J�����F�/fz4��N͞Qm��,QY���Ord%�3���J��J���R<�B������j8�N�ٷ�ϼYr�A��{)3/&�܍��:z=�ȍ��k΃�����8t:��8�.�=��������k?��N婛�s�sƗ��G��D�ϙ�Pt�j��zJ�\L�@La�+��dI��b�P��g6'�	Y���`d}OSC��"�cLMR(;�LspM6._A6Dh���sdi�iz���`��������ⵥ�k�+o�Pz�z�/�\X/[Yn�p��Թ�3�G��෿y�׿|�Ox�����'���2{��3���\:����_�w��˯��t���^�z���K�VN����8:�>3�ov������d����ʒ�����L�*U�OWqRd�����9��R��	1sX@���qh�,��:J�	:�{�)���[l�G\��ї��e�[�FX�=b��armT�C ��+��+|��}�D��A����:���S~��P~�Ȩ�4�T�]&�%�6�5.��������x�#�)�|(c��Y�U�}#%z#5v#9f���pZ7̆���j%}-x�h�"�G�=�F�_�W�+���J��+7�֍ȸ��̍�����iq"ֿǔ�M=@s�ŋ���?&�?��>��>��?��>$��#Iޠ�o��[�^��̆?���Uz��%?w���y@V�	���$��b�`1��yG�F"65w�JE�%�<�w^ :'�UJO���F��Ez�&r��]�0�0A��(�?������Q��M�oT]8�5����lu4�Rb�dM���]���@M�-�B#)]��0P
��t�%���V1�ɡ������	 2	A�`_C�@�Q��&0zcj�iL�78�,�'s��%��
�Z#��&O��W�DǄ`k�2�T:�L��E\>���A��X<���t3	H1�@F��=�b#l|_p�Ӛ��M;|S[���д/[��VyP �{�}9*����x�>m�(\a�-R,���`#3�m�͓L͑:�c�"h�|/S󔘚ɮd���Ț95��皚ɡ����|���^���+���8;�;�����c���G
=�&a4���S�٧�� �Ssf0~��Y��X�
�������8��ms{-��i�ϴ�aS3�6��o��k� �6�{���>�1�6Zk����7��)j�9�Hk�đ��Ց���4Cy�� ֜�M���L�?Z/�1�͒X�8J'Ws�*�[ɋP"��-?\��j&T�t* ���p`Yk���1 �t���(N	`���`+'��	��vj(��bT��.�����I[��5�Ӝe?�%3�S��鼮,(ѩ+[ڙ%��f�����H�P��p�i��v��˚��Ԕ������(���2^b�,�N䛧r,Si���h�x�r6Rs,�x2�|&�x*T}�&=jO�#���{*�v�&띞����t�����χ;~|��G��~2��eO�g-M���xϞ�*�df�
��b���4�9�&gI Y⋏��x�I2w��Yf�938����u���F���.1���W�I7�I7x���o65K��L�"
�0�&�r>(�\`�� oz�f�Q�5,���.��	�:��L�-QpPm:q�AZcA%iֹ4�� .�ـKR�*O���ȸ�b���y�G[`��pG��92z����`�����=K�BiVi��\Ɐy�����q:a��9LF������~�z��3q"ڌ�=)g���D�.�������=2��Z��L��<�7��ZG�MP���T��&Flm�����j����G<+����Q~JL���r�*:Y�52:I�$��T%��0���G��`�+V�`PK-����h�2�`G,�ۜ���8g�U�WDE���G������t0H'�<�4p��PId&�����h<�C#q!A� �n��;�vn��{f'E��D��a��ɏJ�L,hK(�H*�I��n�k=��6��r8�i$��pr�PT�~GF�)�A�F_kH�7�69�;�K��9��2]�w>�r0*�ۑ�jOi	��r���ev����:[\�+~�;�*,���g���,IZs��.U;�R#��f��y�ǥ3��M�F�p)��jZ�����<O���Ԁ	�恝�G�{�G��xp���QU&�+eUɊ�tm]��� 65Q]����b��c�KÛC�m{2%	��haQ� �JN�S3C��a��0 �E������5��x>���f<���-S��M��;SS�6Aؘ$���E���Ğ������i��u�]�T�d��yvǳ�ln��_@` �S�����aS�F����-�s�b�L&���T*��������������Igp��Tf��f��b�$R:���������B%��nj��;w�<��y�YB����C�7A�J�ѓ5�Gbj S��͘��L���4$�R�{�4ߙT !(�aL�n��]>H� �c�T���Pć���?<3�cj�D6��ř3gnܸq����?��޽{/��¥K�z{{ǣ�F"��C����1
�^S���
x&����=��@15�������P��?`j����O
�h@ݝ<�O��M,k�O�p0����H�$�PD��>]ߐal̄�t�8`Y5�{Y���IQ���	��$�wB}��1Kݒ��cא�/�%G�XӴe���j;�u�ȗǘ��"�c�>a�jпҞ�i�R�dH������Sm��q�d�L�%Ą&%�W�4t�Oi���{6�g9m�r��ͬɛ�#W��V��/���N8z7|��q'^��{�2��2{+i����K��O���,�9��O������/��_/=~�p�r��z���䁅ԑs��I{�TL��̾�����}��R�3ˠ�2k�.�-�jM��bMpi�`�Y�F��	�41���,3�B˶B���t�P��cjX��d�iF���Pa����Vi�XӞ��#���Uh;=?�¥�W�*�N�^����k�^j�v�zu�au�������O���vc�W���ƫ_~��/~v��/��ʩ��ϝx�ʙ�7N�p����꽗�]=~��;׏]�8{q�蕵W.�-/LM��v74�g�%�G�
b�r��t�0]�I���$�L)KDȅdB��A159��|(�&�]��S����Z�Y��VpT�����<� ��ϡ�hC� "p�g� �牄7X�9��$_rĿ�i�h���GĆ=|#4z������K�������9�WȤk�&�tண��9�����KĐ�����E�%6�U�u�m�]�}	�!�=9�s��v�­�������P(�n�ڠ��Z���OR�_%�oD���4�4͆T�G�O\���\��P(7���c#)u��}��c���/q9?Ѻ?��?fh�`�>ċ�Gs?#L��}F����}M�yϿ@y��yG�@�-�mM�Gڸ/�	��C_���A]���@�D!���cj^��_brm�w�J�.S������,3 ���X�3�RV"<���J��b�cVɠ]��r��	���=.��t�B]�;�8�a��p`o k�ǚ�����lI��lg6�15`����1�Vj�����e��E.q�Ko�L1��?���F�1��H!`ID,��#�!_C���T8�	ܨ�:5P=aO-aʷ72�L"���8�@�����Nbs�|[,�KeB�T ���*�Z#��\!�Ʌ2O"��Ƣ�$�@�aqP�M
	`Bd,���xN�G�ρ���l�^�.0v��[��J,�9Z�\uO@�e_�îO�S���^_�5���|Łb�@�v1CU��r���'v��"h�l4^����h�����lj���L�Ϙ���h����܉�[*
wA�f��S�˚�����}�Λ`|���?��~�·n߼p��D�DߞɁ�١�c�KO�-8>�wb$��p��P6��`Ƃ�Tͣ�fa �D�ɾ�Q���P�15p\����	�<��N�fA3���r w������D�e��:�d�l�O7�N4�a&SMN X̶�M�� S�a��&�D�k��=�>Z��q�U:U8�*��5au`��P�*JԤ��I^�S�`�kv���憫�n%ϭ�)��(���hxn'L�v)�6� ��n��lb*����
n��i�lr��
���L��d��h�L�]N�_��a��;h{3�홒���t!DЖ������t'8�	�`�����fs9a��-{CE:�p�~�� 8\j�����ź�Rhe��4^l�(4M噧rM3Y��L�q&I?�����E��\�	�|�"�4ˆռi��JV��Z��n����s�?��{�P�k�u�t�x���ޖw�j�i������ڗ
2V���bM�e��y����x�ɚ�N��4�2C|��;��C�Β9�d�4���� �"I��+(�U�*�p��_Š��[��-^��t�*X�"�x�X'b���G��z��[�Z;�ϳq��2���'�	)�"�1pQB�,c^Q�a.+X���Jᚌ�,f���N��'��p�����gɄE~O,I���E�<�~�Ø!a�I�a�����I �A
� )�1��h
֨�9 ����rr��(�4�p
��B�.W��4�r-�BG�2������L�0��JO�Б�@�Q:z"+ ��f �� .PM@*	##�4
��ecQ<*�C'2�D��)��j�D%�8r��hQ��X!��$J��N�:YxRTnU�����n���	cp�Z�J���q(�c��A���ɌF%3(d:���x�@��vo۵{�o��?��|���;�}l�U���[\v[xxxrLBNNQ}RFEXL�5,��Lј��0��L	����Hp��9Z����)$9�� �2V�D�(>-@c�8���c0$R��JY,�T���2I�Vi�F�QzU�A�֩\:�]����F�D+�˄����J� ���0׭a�i�n)B��Uc�5h@�H�a��8@��b$���ifR���i��+r@���R�fx5�e�j�2^���@�+���� 0;:�O�`�W���M����<}K��1K[���IUU%+ʓ�����Xqe��:C�'��V�V�R�U�]�6��"�� �>�vG9���Q���JOu�Ӝ��(fN$#�E��f9��at�ŗDq�.�S��Z�}�U	"8:�.Yܐ,�]=�)U֜&�e�Z3�`��"�S%��1�>Iu�򴅪�����$�뒔�ɐ�K5����F�ABcw����g��v�޹�����?�Ġ�Dpa�F�k#�B �n�H$�k���ÁK1����t���QQQ��O.���`�0X���p�b��`t�� �]�T1��!G��� ?�Z������@70�����4����~���}v;���F�ga�d�I@	�Т�=YGK�L>EC��.���J�FR���m����5�NVQ(��ŁeMy� �5Q��h܁����U����!�8�� P���Y��hNS7���ѩ�Wf;��j���faA~(?���l�U�ݵ�T"I)�i�*>��C���Pp5��`���D�H LMM=v�ؽ{��{｟���o�����ʥK�:;;����R)�W�B�P�P�<��E",k������n�[�V�^��d2�G#p��+	��^���c���m~;�#���d�A@t��qzz���W&Y�����&ˌϳ�=�o-*��4�$K7U�;=A�.U��oT&=�"ITϯH�T�@���W�*�ӵ�ή���Bwk��%�ޞ
 ��,[U��0\\!)��J��e���O}�Lu}�"C��L5�5Kh�LD{6�T��8vf�����l汦|��L%TN8]֒&lN�6%��XuIܺYE�&;���I�M�+ɯ�*�N�Z��<�1y�B����#c�\��z>r�R����髑��!���O^u�]���=r9�o�up)n�B��ukou���i�A��+{N�*���9t*i�\l�xL�D�����ɸ�c����҃�u#	e�<m�ޖh�F9�a�6K�Me�E��(�汦&�� �.&�� �;!kw��s��E=�NͱQ�y!�H���9ť���	��ҢĖ��m�C�5#]����ON����~q���}� ��K�]8?tii�����ջ����~��o�ޗ_�}睫/�t�ҥ�ӧ�O��|���������/�\y~�����'�������9zbh�Ⱦ}=�{;��+�*ʪ2���mYVU����`���rZ���+%�HH�b|��%D�QYܐnP� ]#Dױ=RʸQ0���q��9gu�gF��2���>{J-�1jv���oǑ`�y?�$�],�K��?�_�44ھvGnD�mDD}��to؜��"�|"�/�<�3^dS.���A'�}O#|��!������Y�k�K�=�%6�>w��y�D} ��)d�%�~���Ȥ����{��/�ί�	1a���0�7�Ư,��k���	��A^�3 (�	��oD�od��岯�ʯu��T_��P
Uv�FK�F��F��ƞ�N,�@������1[�M�!Q���1��)��	��1��C��<�u$�n �N�.�q���!���z�){�̻����$�Bbo!ѷP��x�m<T��6�S���Z��h����kD�5<�*�t�@�L$_�P��闘�sd��=K%���N�(�9�3\��vJ%8�7��M�i���E8`��Z��=n�>7���:��O�N���ڣ�m���vK8���l
g�Es�Q@K$��j�dՆ��"�=nZ��R� �Zq�fL� s@�_n' ��; &ТWn�����&l�	_d���	Y:R��^*����fF�tR���$aȘ`*A���`D�/�!0<��@z��18O���9�Dc0(L�Ƅ`�<E�z s��Nbd  L�"�J�3H����D��aPYT�'#Q�K�	)!!&*��&1ƥ�eXI�1�y{��-]ޑ������k��4��y��3Gޙ#�ʕ�����
@o��@�n�������O<�4W[Fk�[��f`��(O25Sm��� �.XO8huikw��GLt�Lv�O�K��N�{?A15����*�>X:u�vn���ᮓGz���7;�ɚ���H/`�p�G�@̎����'�	�3�����^�35��೏���÷?}���G SS=������c�PL��Ѽ�ð���=>����tAIO��Ԅ�0�h��L6����F+,n�+03mS�&S�l
o;\:Ti�pW��	��8P�Z�*O�fF�S]ܴ0A���c�knr1rN���r 	��eN�Q�*�c_@4�	 0�	�v>�ƣX�d��R�D�0!�%�Fˈbl�08B�D��h�1��E{�to��#C��G�Y��q4��y��b-�fS3R�п<������i��`�H�qPd/0�����Ӏl�L�y:�4�b�J�M���Z����#FٌU=��L�e����[�_�/}�Z�A_�Ǉ��n���O�z?��|��Ӂ��5������w۫�W�\��bf����Wc�]�U�e�p�/\e�X����tK\�0�i�eG\� k�{թYE�W��ǲE�x�L6��Y���kD�*�NF��Q+$�2�DF�P�kt�
r4�<���, ��(kb꺄vAJ\�1.+X�4s]�Z��W$�%�,�v�I^�O�P	�3����`M�J$��)KT�"�v�I;ŦMѣDT?1���C�&v����*r��?"�Q0��~9퀂�)%��q�\��ت&7��PX�R0�F�f�L��4߱�D�52�i�z��Z�)d����B©Z�6b���0��:&MN&�8�.�S�L��;�P�*
��#�K�v�!�����������^�����n����I�m�.�j�\=s��dew��e%�Y
�^i�3x@ �C`B�AA��&v�;����~������s��6	��%
��I,:��`��VWDh�Ak�K�l��J��<�H܍!�(�h = �B��X���y<�O��B^��pih6���ѐl:�FJ �|�D�PdL5@LS)2Y
&�R̓��B!G$`
xt���\"�ij�(f8L��.��B��O15�����6�����W����fO��(�Uk��9Gߐ��M�T�(+��eI��Dyn��|*3��������ʘ���=�jS��z��Z����%���0 +��+Ȏd
�yy1�75'���_<�¦�4�Mu��r�I�������LK:��gj�]��X��{\ ���C����I��duS��!͔�VFEf)�M
��o�;~�k׎�^S�Cb�h ��y�Ԁ	ط��d��W�����p�\���0��7�l:���RD>�#K�FSd�j��Tj.���h�І�����WL���aS���6\�,��Bz���dūi)Zj�
j���Ԁ1�@�4��5�MM�����xdP�����<�iV�{�t��iH�C1\)20iJU5�hjU�q��P1lj�� |���K��nO��n/��r���a� �$��L�]���[�������/>x���/�x�7��ׯ]���Ғ����%�HB�P.�K$��S�s���mߙ3N��-:E�|�ǚ�"����f��I�U'	��yИ$�J��LJ�����d)�4Y(OUT�i���-�ٚ�؛��lj�#�%Q��Ei�P��L�@�u�Np���,mC��9�-[E��@x*�<�H��M��<������~��5Uؚ�mNb6&1��5ɢ�yz�>>����\X�]ߛ�o.����q*��r��Z���kh%�ȅ�ѵ�#�a����	��ň�K1�עG�F^���2~=��ݚ����i8�jݙ��Ǯ�L��>�?t�p�L��bD�z0�v�U�o�i�,�	ͬ'	m*s��f�9��H�.ڦ��I�-�T+C��40YFF���m�r� �b<!oPԛ�^��LM���15,����(�VZ���f�%h�:Z����%9�K��80�;trtr���峓��,����ȅž�SǧkG������T&�$V��O]<w��ڱ��NL�8~dnv`t���e`�pg������Ʀ���g����s22�bb�#3���2s3��R㓳�R�;:�:�:+����Ì�~���.���h�������,	>S��cr�>2��,��x��CB2
&M�y=�uN�A-����HpX"��c�5A��|�;�3��%4�e*��l�ْ/E�_�Mr�����:"��а�k����N�R�g"��b�}�&��N�,b���'~����%�*��yID}EH~�GxS@y�����@�xG�O%�X��¬_hV�  ��IDAT�����P��̿��5���_��q��
5�ٮ��I�;��/2	T`X$����H���d�I��R|�S�Q���Q��m��m�m��8��3�Q�����ϴ���">�>b(? ?"r?!�?#�>%�?!���<�,�]�M$	E~�&��G�N���!�Bbo"07��[(�,dj �4X�@��)8�i��wo��7=m��)WI�x�N��b.RI���,
��=ç�2ψY�d���A0o�XE�6ል�g���8�a��pAW8 �:��q����(>�c�F�2�55�z�CSSN�OMM��\�l25�ͦ�؄�MM���k�F�+��qv�I)�щ$t�O W�� p�~ؐ���Nxp 7,�ţp4 L�X�@� a�|3!� $*����������Ԁ'�uG��	�`<> �	�cBh	� !��R�O$p	(.HD
а�6֭%�EnZ}oo��=C֚&or�c��Ulq4=J�S=�5�I�f�'cz�Lo�to�́B ljf�[��t.��;6�o~�sf�sv�k���V����lj&��٬i ��7��������|��[��{��K�7������a����#�'G��<��0�{b(��p�?������}cj�E0�l�{�`����UMM�k�%t���j��ht��d�H��cu�Q#�I���4�Y�y:7J�!Is
��(��d�+����%e�J�N�qQ�r��pɨ^�09<d,|������G�HN�U"R� �`�p	6R�q�B�x�n�����'���3K�Y�l��h�D'�A㥿D3P�����bj6k��k�Jt��9Rb<Rl-0����-�ֹ<��<�\�u:�4�����-$:�݆�hD'����t��J��E�ZU��U����\�`_�;����`�󣡶�u9���ᎏ�Z>�k��P����X�Yk����f�}��a0\Q��x�5��<�}
O=M������us�L]'R���5n�^
A�
<6��-0���,�aV�!+`��\!!ש�Uf����aV��u&~�CXᓖD�e1eEB]���d�u9悂yQɺ�b���I���'�9.�4��@'��Nzx����H��'p���@'��F�!|�!|�~|`r4�(�=���!*����G%��rƐ��'�����R|��Ъ&��Mr��Xg��Xh�f*��Dl�6[��� u���@�ԑ�F݉<D=P��%C�a��� .:���0�x�&�	-v�=�j	�:�\��1)%�E��u]����fF&OLM.��ih>T���jp��h������}g�j��L��iѢ��`��A#y�@:я�	$`Pd�B%�(x<q׎�AP��]�������s�;|�|�	!��ʌ
�Yc��v�Cʖp�<2��	$� �/��FQ�(2�� �C���	,)�/�	���*��\"�G("6��@�i& LX.���"��~$�.�@�"�,J���T4��&RQ8
�#����E0�HN91LMtk���kj(p�'8�	v4^6�0�S�`GS� ��N���i�<�?[s50`ޒ�k���g���������D9 /ZT���ɶ48�V�v��6���u4etUĶ�JUI6Z���d���1�$@N;+��� �����!Ú��uO���T��P{���,k�Ҥ��a5�����%Jj�(�OT�9UےfhL7gE������!æ&�g���������!�H�"�P��A��!H��@��:
�m
�ի�j�F��ju:�J�;(��c�L�L$���1�Q�p��a�h�\x�In
������S� �>m�j��5�P���@9�h��"��X;NE�W��Fݏ�ԤH"� ���:Y���M�ð�(��NMUv4�{�7@�� Sk��4��t��e�H�=kR�Ɋ=	�Xy~�4V�V3��.���e~���ٱs�s���C��\,�����p$x��A�-+ .�SSSs���۷o߻w��?����K�nܸQUU��r�X,8|�@*��D�'����)8�^S�?xU��T��}|w�5�߮���?)�&U�ҝ�{��x?&�O
�kҤ5�B/�)"@���)K��$I�%�ɲ�Tu[���8�^�j��(r�Is��!�R��)����*��%1r �*U���lCS��9�Ԓk��ֶ���s4P�S��+_�W���i�ڥ�H����X�����j<��!mI㷤r[�YM��$nE"??F�����ǧ�����vg��%v���^�=��t��ı��#����G/�Ǯ��_��x>j���磎\��=r5v�z��I�7�'n���->�J���j�ܯ;�j��{��oU�^-[�8��{,u�lZ�|\ӑ������������N�)Fi3v��m3D;4qy�S�b~/S��d�~gjyv*ljrlp�H��S�L�Z������#�)��������Բ���촚���tsZ�<�E5(4��nTp�J�M%qhN�Ф҆Y��N���ń�c��pGCW���������L�pt�B%�r��M��4[]V��d����DE'�B�"\�c�^��&+Y�Rr���##�J!M�1&[U�)�K��r.���l��Y�츑wV�_4��t��*�D0��`3[��ӑ�C"�^l� ݻc�q�H���	��G�S��6���Q߄Gl�ܐ�q��f2�F��R!�T.zC@��$\&cV��El�)��q���؀*�
w��yQL�'��*"�%c�%"����/a|��~�W|jTn��ئ��M�3���V�o���:������4���g��/&՟ү�P͚������� V���V�I%��Z��E��訯��6jnt�otMnT��!�����/��ru�1��R������y_�9?$2>#�?��?��>!��o�ȯ�^@�Mf�N��Ò�𰩁j����;Xʋ8H��!@���v�[��xM��6�y�L]%S�Pi��,��r�E׽��Ep,�.)<����&ѼE4cM�E#vA�����q?45gj8-�,���*X�<)��cM��	)X�l�4b��X�$� �2;�̆-�`*�ef,lj2��t9��ȱs#4���0�F)`�q!���H���`2�A��<E�c��7�#k�	������&��`%���ypP@Hp ��Š����������� �T*�JB�	Hec�0L<�E�sI8>�GP�.5%��Kw�3Ø����4Ig��-]ڒ*nϐ=E�t競�����"5�����oM����Ψɮ��}	ߚ���������ʚ�%��{f�Z�w�8�5?�9;�wf�5�����>8�S��[�~�����ŧ}��?z�廗Ol65���3�p��SG
N�柄e�p��H��YS��}cj�+���E��_x����j�ÏԆ���QcM1�iC��]�����$ea�<�-J�rbt�h-�5*�[�tI��SL��\2b���V�`�"մp%���< L�dD���b���X5=\�w�1RL���D��D��p��	.j�fk��J}��CE����*X���30�.\�<
��-��f��.5l�2^�+���
ˑr3��55��)Ճ�c�&8�f,253ֹB������\�l�e2�0�hXH	=c�*F�q�lH�뗲'tҗJ�߬/{���~s�����կ�������5�52��wz���m����㞆�۪~qh�/{Z�)ιq'�u�f��T��e+<�9:�$�~�B_���Y��L���N���+x�}�<r.8x�^�?�%�,㑐��h�Ѭ�Q��:�&��&�s�k|Һ����v &����	uYD;/`��A��$�t�F8N�/P�O15����LY��ט�e�,�z�B�!a�1A���؀\@!p?)x?�KC�"���!6~D@��Fd�9퐔�!���p�R|��آ"5�I*b�
��ٙG�"h���X{�L@��^a��hJ|��
psvZA
�lCl�W��N
��25:�=̑��TXSV�TS�X]�^�ob������'��/>�~���[�_����K����2ta���|�����5�����,�+�H��L�n����:ؙ��Vxh�0����:M-�h�<��)SX,<���`}��پ�ٝ>�!�]A!��_��;���������+5�tV�ɮ2�*[""q�x����y 	���p�4���Ր�R��rl����
5&���W�XR9]P0�R���e��t�!�sEͤ��
3�J�'`w ���������H,�`��C���@Zp0,!!tl�SB�P��0�(�����8�꼅�L������xM�û	|������v��jZs5myڽ��BCG�	��;18�	 �fUi��TMS�����V�]��S��ۘz�3�@�Ѿ������}U1��D+ �@|�5R�����ͤ#6��ύ���p3���HFa���� x^�c���i�F���l�4-�
X�<jj���y(k<�8�S�O�6i]k��)Ò���ʬrlj|�����۟��ْ���t0
�@�HoL��Ԁ�&�T*����B8(����|.�N����MgHB���p�tz�B#��HTH@`����dj���Ȏ]>۠� ��<�b�2@�$9��h?^ÍSQ��'�Ԥ��fY���lI���s�"�^S;��d�fM�ij���M��%��y��xEy���-{hj��X_��_0���	��	��#xӸL�T(���eRiT"	�@�u�ʢ��"x����ܹs��y���߿���+W�:�N�.�i4�@ �D����XSc6�aS��ǃC�lм��o�ο35S��Ǧ�я�XS�Xk�fs��S�FS�*TCH=�F\�$)K�'J��%I��deK���Ƚ�4����06��kR�����(iq� &%1��DMU��:J��z�g�s��9��\}G��3_��@�]h�)2�o��A����-��8^Y��)�����=�K[��i��dNS2��*�JR#4����Ԕ�ª�ʽ�uC)��c��'�_I?r3e�f���თ"�.G�>3z;z-�𵄑k	��'=�4x=e�F�����7s�oN�)��S1{�h�J�����Z��i��jt=��xr�xJ�hLՁ8@EoBپ��ބ�z�!Rot[L�0�%Ҫ�����$�8��O��I���$#=�Ȍ5���X�"�)3Z�J_�asUL��E�0���9$�Na��,2�G�\	���c8$��M�rq|:�ϠIy41Ǧd��̎�L���+MZ*�IbP��`:�@�@���}�Ǘ�D�}w�B�H?%���B���IbB���-%AyO�LM��#��0%"\	Y��f#�x��1��M�h�,$K:�)�lR��P���~c�����9�~���`_U�й�Q�2�?��g�$@E�l�Gm�"6�"6�a1�m��D�|_�}�K�N#\��H�3Ȁc�;���:G���]��^���I/	Hoʘo�i�s�o���dU��4��|iQ�Ģ��U���WV����ܦo"�߸�߄�6h64��岯�⯄����",�Z,�e͟e��KER��h��"*��i���{�7�������)�W*���4�����Q������a�㘟؟����w0��C/b^ǐ_Ð^B�� ��C0���۰�A��b(/zd���"�5/�7<xK�\���hL�o7�v�D�D�\�R/�ik,��z�C;�g��`M���ӉN���,�9�x�&s�����PA���>E����cj���pfs�k`G��<���15^S��M�
%W8�^Y&���NJ��Zꠔ;�Т�\�	_b&�ӟ���"&���:f�I�n�r�*��A$��"�v��&�o"��5D,�ECn��d���� ((��}}}�y���|(<�r��]p08��gAP�@Dp��;A��A �HX����S� ��1K�b8����b*�($F8�ҢDUi����dg:��i��Tqg�r��@��'_�x
�[́b࿅�yJLTN�;}�'kz����������{l�cn�cf�}z��)�fz�� ������!hq��@����4~�������|��/>�w���㇪f��+f�����SϽ+^G󨦁���/������f�Dc(`�)0��o��h��j�o��ڗ6ޕ9؜�Y�n�5W�h�$�v��+�n9)LF�"�CH�pa2�[�Wb"TX0��QNI�C� ��H5.ZK�3�L�x#���r
3�4+;���r�
���I\/[p�r��v�.|�9v�-n��5^�8Rc�0��i`_�X�l�D��1[*7���˓bj&�l�Ͳp��x��0Zn+�e��RSs$O?Uh�-��:�8��9�m���4˩�����S�Y�a¢T���)��Jz�{J?�i����~S���%w�o�ܪ�{�����W;*�������ކ��V��R��C�?�iy�(�F��fT��}M�\W�W���l�����b-�+l�y*i�JZ"�IP��<!`�
�H�e"b��P�@�NT�*�B�\`Aj��t�G�P ���2��l�2����W��&�/�)�B�9�4�r����<%�p�L^�R�R�L�9�$�4K����C����n�7>���C{hj��a>	
���e���/#�	�mb\��(�7(�r\�_��W��>����L��@Q6^e���D-ѓ�4�:E�	��h�R�.!џOE��t�YUXS��ko���������+g��-�.��\_���t����W��ܼ�����~�O?���S/ݞz���+k�˧�/�+=3Ww�lۍ��;��޼�tu���٪s�JO�Ԝ�=p�|�cM�cuG��{�Z����"RR�zS(�ә��o۹���'0��l��o�w�ێ��|q~(6��`�4\��+U2

W�g�qt)�� 2�d���5�9v��ᛙ��:�H�6Je�V�#TF�Lo(�l��%ճe�LI��,)���"�Hd�A$N0��~8�/@���@�k|���!�]�����)�~tp媥!"l���"D+�q��S7~*�`�͛WЀ	,h��滻���fM��Դ��:���J�ݥ��|Cs��ԧ�T؏5�[ۊ���4$��&hJ��eM,;6���H���ʱ΂�洺k���F'Z�)z���J{²yA��0�_�;y_6�nӻ��:�膧SxC�c4\�f��ns��P֤H=�
��IVx��4ͩ��t}[��9Ӛ���I-
���_}���߮�۞{\c���+*�B
���Cz����#�D#�HpWN��[}���*��'I��aP�"?�fO������p�Y�&�PD'S`Sv��v�|���jv��n߹���ފ¾�>�c%�O� :��� AˋW��ħ��<��xe�wa5�z?U�
�'��|��w�����dEM�65q:���a���(?��0��v���dRi�-��`��,�{b�|6��F����wyy��_~���|���_�tiqq1''�d2Q(|���)�F�ՂG7�����~�����uj�.���cj���yJL�w�w��;MU���He	��$�'��cj��	��$Ec���(��,f_i4��<��8�%7�<^S)�s���%R@Y�zO�aO��6� ~- �(��Жё��*0t��zK�J-O1�%���}�`��Hd���d)[3emB�Ԥr�R8��<�4A��K�s&''f��6�W�i�s����\J껒2r=~�* a�ZʑR�nf��Ιx�h�岙W��^�3��r�^��K%cwJ��*��g�Ŧ����v�F����������s����+�GV��M�.h̭=�W�]Pљ�Yi���-n��e���u�6E�M�h�$�<Ej�15�đb�����&V�Ek���j	I���Ex:I��H<G`��O.�Hl�š3�d����S���D\������VD҃H������ks�N,LU6U%�ȍ
�F�g�D,���0��K$��0H�_�����8_=$���a�	��b�wH	�).W��c�d�">��R���q1]
����r�(_�+֌�U��Z=��S���/��~13�fk�k�%'��I&c]$~��{��y���\���Ѿ�ڈ�߈��&��Q߄�����f��V�����~�N<�9��h��S8�e
r�t����D����3H���oJ�����5���?���0�̮��65��i��2~e݈ulD�7"�PC(�ià�F��j�x��<�C�Q`�+��b�$�?j���G�2<��伍ܪ��ʍ����ԍЄ���?�KJ����)��*��dS��}���G� K}KyK~K~�{�{	�}��Ac_��^�^B� _C�������%P��7���u"��|��P|�z�D�@$��H����¤-�i����Y댌sV�;���	OZ$G�b(��&u���P���55p�`8��J�_45M��=nlj p��J'	�5[4��$��RJN(��܎��b+-efl��Xl�d�ɩ*b�#'F*�1fY�Uj�k�,	�ڍ�݆���=�7*���"�q�0��!h$�k�	��� 5p����Ags??�E x4�oA��C�! ������E1H2�	�@����|b�YLI	�����2M{�uu���|m}��-]ڞ!kI�&=�Z����c(���f��9X��oaj�S�15��=����}(k&{���¦ ��?=��kj�8������������?�ⳏ޾����ݹx�ؑ��������F�燋����d?}���-�65�V���� �/�jj�Ț�F7`�10�5�;ّ2�;��Ƅ}e��lSi�,��	�� .1*`��S��#"��h5:V��I���h0�n��h$�Z��Nf^8� R���F����U��=)P�����|#�F�)6T��7E��?ޕp�#~��=�6Q�eM��5[��������k�J�^5�����<��<^e���B�[ YSh�7LZg
 ��<�l�0��8�z.;�zY�9���#f��1�l֢Yp��g'��\�������j�z����披��+� /��>��dd�G�ouռ�T�qw��m5�
�_H���u3�}�j��׮�e��T�*-��X�E�<��H#/���t�*��F#��I �+��X�e�JX�`a;X�c�8�
w�K��'_R/�hW����%�l���x�o�i��g��S,�Ii�����St�i�I�f�F]�� ��ԓT�<	7�C�{M�>��>|�>RP75���8@Gp����Q9cDF�P�I=RP�,'4�j�F-��D����<����C��Ra�*-�2��H����D:F����B�]) �'���֎�N.9�0��<uqm��K��ܘ�q����ы+�׎�/�\��t��o���G���/?�կo����_}y�՗;�^�<���b��B������%ϖ_Y,�|�h�T�����f2�OԜ?���l����ɺ��ꡁ�Ύ�ZGb����9�|�r�_�����P�T��������AD?Ibi<C���0T9��@��h�K���B�[h3� 'G)��*u	c���1������93Gf�+����hb-U$ñ�!�?�S��H�,�.@PyH����HA8�����y���N��ݴ�;yA�5��P>FI�U���ijhy.ƣ� vk���o��"Pk�zO����O����bSO�����Qdm�5��O���Bہ����ԉC%G��jJ�mL�ߐ�ߖ5�Wy����p�Ѿ����ю��"W����bjb�p5:ƀώ��F	R��4'�(
�s�����k���x+n���	�)^ƫi`S��2Upua�״dl�5P�ޘ���15͙��pU�Il�2X�������m��k;S��B�`�ؐ"]�}T�a�X2�sl6l��}>�I$0�8\2� ��,�����Ĥ�������,��:�P~��߹}�SL�<�f7�����̳�ߚ����=IM~JL�c�����߇���.*���'��9
�5[\�ӁM8��e?%��$(+b�y.I�����8�`RH\�weT��`���]�0�b� ��\&��'���+\vGvz���.ܿ��w����_�up�ĉ�����D"�p8&����`M�GM��d�h4�Q�ԀCn�H��]P@�np�<����w��>��{e?=%��?�k�'ݓ�F(��:YR�.�
��)��deq��[S��φLMOy���8@oe|WITKnhi�� B��憉����HYM�ʐ*
m)��䙛r���H�diޘ��(��4ˬJM0�%�;ƻ��s�����"k���YJ�3i���Aa5ͩ��!�5R��)L0gĹRb3�����ڎ��=���`�F�����{���7�z���M'�j;�vǩw����й�G�~xx������_x�5��ޙ��f^:p���o�/��p���s�w�ܰ�TM�=��ڎ��ޙ������U��+*iJM.�r�E�\QVk�͘dצX��fa���l�/S��q('��K�pb���P+$��B��W��������g��������R�/�����'!X$���P�� ��Dt C�f�8h:�ـm-�m���/\�;9��ݚU����:&ď�f�0��F�� *���C�h_vw83$��J�dK�Y"\��������yR|�U.'P%\D��P�A���'"�i�lQ���݉������5��IĿ:>�q����������9�~�F���Bc���}"��Fg���O؈J�p�lD�7��\�?9m�0�~��?��_ro�i�d�YL��w�{p��BE���/QQ/��e��%�wT����ʏ͚/�;?5�,��s����/��_;�p�i�&���H��a��0$kl��~C�ސˡ"5"1ԙ[(�I6d���+��/B�����4_����Y���p�m��lX#7,�����*�9��s
�?h��Q�?"1��}����K}O��ĸ�Ŀ�¿�½����ü�_F�^ƐaYA�ނ�v?F�\!Q.�Id��Yeї��E>�uN�>#�Qp�(y�����U2gOY�cV������r=��p[¿+O{��<�� �¾35pTU(΁�&=��"�ZJ+sR+�PE�*;�҆���*-�r3��J*���L�t9VJ��B�D���P�\:�E%�s)L|0>h'�o;�k � d�/*��	�<K0
�#TH�/(�' |�|w����@��P4h�o x\N B�� 0A"0�(l�� �H,�#��$�@Q1X��&�8,��P"
�($%�$��ws��>WӘ��[���Z�$m�ԧ����B}���Լ��|S�5��L�Sbj��O��&�3'��'{���&����h�ljf���?RQ�[S�:͎�æf|`��`/���K�[��������ӟ�����z���_��>?7�r�@��P͉�=�����ߩ(��{?m1��D�m�����;����=f|�c��	�}�dS�Ts��=�7ӓq�`�dWj}d{��<A��dF�1�5�!��8-1N�I4���,%7��q��<?�Y�*�f���*�ŵ��\m[������Ŷ��CUa}5��*gw�����_i��mp��C@?�{�c{��֑J�P�q�T�_��󡼎fs~;�(���e��'��x�l ��v�`��1]e���M��ǋ��ƉB�D�y"b*�:��8Vv�8r�8�^K��=��v7?h�s� �X�uʬ,��/�����C�?�j�����
�Wg](M�И�FϞ��?誾S�w����[y�7�co���H����4_4j.�TWM�+ՊTp�G��1�x�e.}�C_�P�V�l�e:�2ɏ�E\���x�� �D(�FD��s���xIʸ �_R�/>�U�"�-K�煤�\�	&���$�`@�i`S���4g��'��e�<�~�FY���)<�0&x ؇�R��������w��P��^j�O�1Ɣ�!9����-!vyj	�H�M
B��P�&6i]���hYg��=R�.h�58�uv&lj��5[��P+,�
��N�p��y+�D�����(%�*Ņ��5�YG&�\:~�����׆���^��~������kK{Ϟ�Z<�wa�oyi�ʕ+���/��?���_m�tc���v��;]׮T�9�sl�|�\��B��B�����'�.�+��
(��V��J��ɔ�Ùs������>1[|�in�uz2���g���FFS��`T ��@��ѻP��� ���� �0t5��'2Md��´�V�J��H4'�a���$��L�3��Q�L��FI�R�-Q8W�seN����<8$�*S��
��R4E�g��,0�	�,�P!xZ��#�c>H�� �v?�s�);v�v����]l���"}S��+�zwn 0��<�����k8�.R�5��*���/��rv�X[�p�؆�VEL��Y�87^�8�8�_�ל��6��:��1u�P�xO���ʙ޲�������wZ(ǭ�X�6q�Y��Df����pnv8� z�`s^�i�&�&s���ʚƴ�j�x5M[�
��g��fk `˚��M��cj`� ��6��)E��~J��|������o������~���'n25`7�
�C���{tC�P`�O�P���D"���'p[}:����`SC�v;CӓSbb㢢�T(!���������$>�v�z
�����z�j�޹��'�lV�����%jIZ�bjҍ��(�p7�5ߙ�(�	n���H ��[���t��(���MTT�)��K��HH**�����o ��\%�w��bKB�+��(��Z]LDdei�`���������x��<����_�pa~~>//�`0�}U��F���OF�Q�V����&88�l@�eM�k����m۵��۟���̓bj�WE���x--��+k���KU� �^*����eU��"EU�(/N��$*J��uY�����UI��ɀ����<wi�� J�&��J�`�`m�����=1��a{�����cS��1��ݚ��lj�Y��-���|�#k��ƫf��U3[�F�lI�j�;Le��3Em�|���ފMY�=7ޕ�������u�xC�bE�r��j��+-S7�g^蘿���+���tN�l?|���zþź�3u�'k��j�Jj�*�U����8��2����y<'�=&����	�e8��vsrTdfRb~RB^LDZtXr�)�,7���(�%�dH�hSm��,��O����y15�z^/��O0�c��H�@������?���������'`��`��C#��$<�e�0\Z�CI�(!��QS�W�D!�C�	�YT���/�|����٦�=�YIR��$�lǅ��� 
:��	�c��� ��vV�6�ϿI�5���Cd���*J��-$<�5RB���#���	鼐2%�X�.��J���>e8fV.h�t��]������Wp7+{-)�]��bj|�7^�����w{��dd��/���̗i��8�+���7\���gĆ;���/N矜�?�:k1�U���ݗnW�U2�,>h�7��y��HA�#�RB^�0^W�҈>4+?0�>�h>��p�~�2��e��� ɚP�/��_9�����m�c��wN�שׁ?[u��7l��aà�Ш!5���7��rC��I�&�E$�1��	��9��k���*�W
�Wb�W"կ��_��?'q~A�����)������9��)�k��(b��cI�bIoc�0�ױ��X��8�W��{8�=,��2��2�xK��#��'����	��牄+.� ���E
���N�^`�/pYD�5	oM!XV
U(�F#8���
£pޓU0l��[�<o�Sg� ����67S��P�x�,e�+15ް��P(��kj`M�B���
�CS��@��W1
��L5N�aB���3��V9Ǫ��	���w�w��w }��x�ہ܍@{�#`����� ��� � �p�_P�o ��X��x2�H���82��P�b&KĠ�45��P	㬊�PEa��6��R�h*�7�(rd-��4(�	2��Ҏ,�u�'_&��H�h�X��w��񘚔�n��ٟ˚��Es����ǆ; �Y37���(�i�nj�GM�>�Լy��w޸��/>��/����W�x���ks��ͣ����{�k�����z�t�5�P����c�Y�gM����x ��ֱ�( <~����xS3V1� �xM�Ds�ᦨ�}�G�gi��.�U%H��+Tt-��ȶ3s��](7?��� 䅑KcX5�YS�И)o�U��i�����r��1X�j���H<�3�1T1�9�9��y��4Pc�� ��̀�`t������q4����7ۙ���xe��	i�'���4�����O�8 �{�S{�ӵ��'`��>Yn�(���&
-G���#���l�L��xY����UY�w7�p��g3C?�~���LbĈ^>eՍ����k������������ow�y���rY����傸+5�w�
_l.�Z�~�8�rn���ث�1�R��&�_�q݈r^u��ڍ7��NӊFzZ�<#d.K��bΊ��*d�
�+|�*�
Xf��
��(�l
$kX��Y�@���#��I=���]�/}[$����Y�\P�`V�4X�,��g���l�1:b���lj��@'�aB%�kj�|��<Ǣ������Sx�&�Pӏ:���t��;����.rP/�/ Q0�T�A�CS�)%6��-R|��ؠ"6�)�vN_��H��?Uw Y��舖���N��4��B��Ѫ�jP�*�12��d�)�d���_�|�ʭ�����gϝ�Y:�sq�km�}uiߥ�����������9�z����KW���ӿ|�������WoT�>�6>�8v���ٌS��N�/��[�K8s,c�l�ڹ���9�I����=w4��l��x��`�p_�`_�`_��!1Qbs���Ma�\��'�ۿnىB�D�����B�ۑ��2P�Dd9��P �� ��8�O�����D�P�an�T��T'�t6����%����<���p���TOhH\5��"��x@���0t�	 s��)� ,5K	���1di'��#��ݗ�Ӈ�s�����U�D)V����<jj O25`�V�,�ӝ��aS��Җ��*6�V�U�u�9aSS�$o�6����/]�i�pt��cǆ�5��W�4�F�M��_2Җ3�]<��h��p�+��4<-��D[E�N"T�L�1�d�;�#�C�e���,����)Sݘ��:�>ssX����15ހ����h��7[ӑ��������e�Z��yhj������4CS�%�.vky:����{���fǶ�~~P��_ ��WcMؠo���M�Je�X`�P(T*�Bl����D 0X 	�'�	|6'<ԕ���pZm�����@���k�f׿?�����������V13Rō�p�t�4=�I15���w�7�[L���r4�� ,z�7��-.��ԃqK��M]��*^�e�hXAD��1(|pH�n�]����"L��?�fRiB.O&k�*�I����,)(�x�����۷o���[����o���k�]�xq~~����h4�D� lj��^�&80�a���;�۶���ʚm?xRL���������Mթ���6z��D��"IR�5�I��6U�hJ����)K��e:�
#{*{��Ԥ �����IƢun��� w;KcG�s�e������T��A�5p�lj�r���ͦ��b�����f;���<���l���Q�g+�fI�3%PLM*�9UИ*)�V%�+Sl	�Y1���m����='[{껏����9[�>U�w�q�њ������θ�*�6S͍��\���ײq*^) i�T����d,���`�E��$�	b1Ud�m*�Mi��S��Qey�/<߽�{NO+�rwwwM*��B\�+q#!!
�8����-4д���==�3=�֮ՙ@��������z~�z�^�S��T�_�"�p�������(�<N#M�K�L�3/���41R��115��5S���(-ՙ�$R��8�ǙD֍��A@��>d��w:���2�X+"�dd��FV���!�RX"K��B:�����XzF���|��ݷ߾���&3-^���1�X���#�Ho6���g }��@)�W�����v{$�#����O�"�8�ͦ&S��cޅrB� Q�C�*���R��t�v֨�SJ�(d笐�y-'�zz�J|\����ލ�/n�ug�٧?���Z����,sy稔�D�m�3��G�}��a���)�G[���ߙL�?Z�?��_����H�׹��t�Y*�!`�>����w�迈�+ψ�5��t�w�ڻջV��v�Gv��A���Ī�Ģ�Ү�Ҫ�ʢ�Ƣ�Φ��,�� �\��Z-�A#�Q���Q��rC"q֩�ojĲ�|�/�;��W.�w���7��"цB�!Un��c��'п�Ӿ�Q��3�!2��3>B��C>�R �⠾�o!pw��7}_Eb_Aao�����@c`e�/�E?�Լ�y!�M�S�`��u2T�f�J^�S�X�5>k]�[WVU���I���VpD�_����Y?f��{�n���찱���!���M�9��:�F�1�_�ҽ9��*��
�)��Ԕ��NS�� �Z4�! S�)�c�̈́�fg��k��b���4sP2J����rH:U˧Hx6Ο���yoGz>��Q����x"�c;��#���	����2.��t4 ��~;���{�n��y���;��|�~(O�W ���C��$��"��D C���T$��A*���(3B_�l)O1T�iv�+��$U���4Nu*�!*'ܒ&iJ�I��?7\�Pڳe-'����Wbj&��O�%���L����g�L͡����"5���j94�>���WL͔�-�fS����@�_��[���Λ��w���y���_�r��ᆱ��ɾ�ъ�����93��3ÙP@T�Ɖ�N��ޤ��Ĺ���	3��}Q��=a���Й���� ��;`�3���f�=�8�p��z����<���<�q��25����d=8�4Qw�E�X��Y3Vm��_4Z:�y�=n�=q�)���֜�{�,;���RM�� ri��*I�;Q
mf�u��Buw���̰��:�~�+~C�H�c��V`�|_m��n����0�����e��"u_�f�L7T��W�.��+��j���p �`/� [N��2R��_���4ζܣ������N�� ��qg���.��<�H�vb�y8C=���1�f�S�3E!��}�<����g�G���a���#��U_���s��)��DH�+Ņ�������ͪ���T�7��Jkٙܘ�a�+3���]+L8�u"-�x��dB��Z|�����1���ˑ֧#m�BM���U�tE'Z�O˹�e�3�i1㴈zR@>�#�3	'٤�\�
��*����
�Y�SV����3`��#�	��b*`MJ;+g�U0��Y+*ֺ���`���+2�)���rJL^`"Y�# L�聇Ⱦ���T�<w}�}�<=G@!C	PKx�"��E-�1ǜ}��Y2�0s���|�^=�n(�.�O�j�t?�iH@r�[>uqP�'��������j��@틖���nH=Q�<[5�en�����>Pp��-�I�J��U�(��9X�fHe�GIv%h'�j���f�'���vN�۷<7p�X��b��%����5��կ�l^;]���=���ĉ�_����'���y�o�[}�d��X��X����������c�IG�����'_L=��rZIqFܤ�M������n��j���1������V�@��h�X�$�<�D_����I?�^�a�p,�f 2���ĀjPx+�L�Gp*F`�1��$�!Z�t�%�)�y��q��%��R]C��Il����! L$x� M�!I\��g����	$�C0g�b�^�W ��s�z��w�v�wx��A|�I��G�h�%QC����P��%¥f `uX)F�O��6jv5'������g�ld\�i ��8��S�(ܚ�mɃ�^%q�aS��PW���=ϟ|�D?��XMombCQXu^PM~𞊘���m����y#�Y{�Rs#�j���k`����lgGY�PC��`�奞��0��̰����Ҋ��P�Ƀ쎇Z8�JոL<o�P��R�ekZ3U`�>Y��̆ 4�ޫ_�O�M_"���W����-���$Mi�<%X��r���Ď'���'�p��	ݼ=ݡ����^^h_o����� �����>65l��V����S�Tp/�ǣ1�@�\��l�������
���R���'���Kn���w�twsF�@������~/�d�����?vF��6�}'�'g��OpLM�#E��P�d����'jI�ZB�����65p��Zt�^�20p��?��T/�O5��$pXǇ�$u)��dpeU����4me�2���S5,���$#��Ob�N��Pn��U{`SC#��l���׫5qQѹ�Y��`���v���3g�{�;w���{���۷O�>=;;����T*q8py�d2\>����a;o�"
�B�L�T(`N#�����r��]8gL�����'~�?ݞz���"��p#VG�Sb��x%�~Jr֦I� \j&U���4=:ÈͶ�mD�b�<�Z����7��Y���	΁Emi�8�_� �JU��rU*�X�ݝ�+J��+�c��vfQ��*��\�U���.c_cvoUJkQtI�!3T�$ �;D��m�飭y�F����OwfTEu�� Z�I��T9ܥ����-*-ܵK+��B}o�����_bl�0�m��Q�R�`��:5��.4�
�y�Ilg@�*�W'�HPDk���{VLLJx\�%�a�2��t1fu�A��:�� ���D���|�7������^<�N�I2�	k;��Az��^D�7I�KQ�Q�$�	���T~d�^�d���ߟ"m��m��x�r�ۼH�=)�=��� _;������Fn�������蛠��15VJ�����&Y����p#O�ES�;����H�{R�x�*����	�#b�,A@�Hhd!	�EҐ�.�ͣ�Yd
�@�)T<
���I4��ݻ�}��w_�]SQ���H@�#}�ܶ�/�Fxz�=�eh�@���׬�Sd�G9^�J�Qx��P�S��L."��5�&S�����"�.1�\N��J�'1�W�>dV.�
�q���Ȩ�rw�����.!�ޙٸ���{on�z�OO_�=6֩T����q�f�/���s�T����nG����#�;��+����[��;���6�]������q�I<����q��<��0�}�H�=IC]�S������o���ޱi�6��6+�3+?�*?��>6�>6J?5J>7J��H�2I>�?Qq��J��C�5?���F�ڐ�6�(����`� Y����B�"�OB��y��3hdҝ凅<�G���=��=��-��-������G�G��k�>PPd�[(�(��X�kX�,�6wi�H�ˁ�K����g���\��?��w���F�E��V X��JĮP���Y�2��UgE�9%�3��g���1���Yr�,�7���)�`���=���Fz���b�7��A�z��4��[B9Ma�Z��t'��ԇ�]��%hjԚ`J��R� ԄӫB��΢°���h�P�`rq0�$�XD,�W��mET��Tfg��:j��&D���2����'���hH%#g�$44�����Q�D��Pp���OH��/���7w �#��Q�>�!X�E���	g�t�ݾ�c'����� d$��E�t,�x.��#�H8/w��Q*V�]P�n��65���9��LaU�*�]�e?59�
�ɐ�g):sT]��=�'_۝������-���Pzv)azT}�j ld��Cq�X��+7W�F*�`���S� �!�-!c͎Ѧ`�搱���=�p�8��5�S]9{����h��4�,*<��p`br�01�d���V)3��w3�������x�������7>z���S�4������W�8^:3��K�fv0���f�7�ejf���=Ss��:��P�ؙ��+��t���ϛ��3j�!0V���>�
��:��9Cƞ�@�������z�L�o� &��:0��"��2\e�4�@�TY�+���
�@���L�W��/��)OV��R��2-�P�j�D��jj��t[�XӀ	Y�sXM�i�*R���LZG�u#ن�|�D�e�a�$���[��_����ɍK'������W{�_i�;�5i���s�处W
>���rO��u�w;��h|������y1��K���Ԑ��x۱8��D�Zr��İ�ab�.�د�]���uhW��3FɪQrZ#�Ps�(9�e�SR�i	픘zR@=%��3V��5 &+&Xy�c]L_R�� �@x�	�&���ܯAk��f�(gtX� 6k��"���B-0������Cd��,P~�5�NYs��["aaSs�^�c�����9�3E@�cG�~{�p�SG�;��	�؃��tw��:i���^	0 &��z�F���vK��jB��5���/�<ݔv쾩鈑��*MX��9P[(7�aSS��&/ZR�j�۽�<������:�7��\�/>�X��Pxt���Rى����kΜ,=��;9�~f��g_��i�ݿm��׍���q��o�_�]>��22�<>�5;�����0�zd!qi.aq���iˋ�V���/�%.����������/q�7��S����O��<�^�����#��	�x�6v'��O�b�r,KHV�(jE�"�q*�&�C�8��L3�Yf���Kթ�����Β������ڊԼH�Uϖ)����T4��!(�B�'Ƴ�X&���H�a�)>8�7�胄F/�	ɚ��m�m;I۞��xL��Q��1:B-G���I��`S�e��3r�i�"5����o�ʃ���&Wߜk�IS���,q,]Y�zae��O�[�_�^]�aʋW*2�=UqM�����������(Y����l7r}H�9?�{��������ϟ�?ٚ
6u`{	�x�	G�<H �gS�ոLaS ����iR�0�ͦ ���$Us��>IS%Ku�B5\%|0�gjv<�������������^��������B��B��ij�R�`�N$�T����15`�O��p,	�'8#k�(��l&stxDLDddh�/��n;]����4 �>��v(��ejv<��@�t���N�ljb��X�CLM����yx��!̱P��W�{?m�S�aj�K�l�U���\��T]e�2�ƏTҵl���"#��]��@?�g�m;�����0�F��%z�&*,<'#� 7���d�����ѳk�/���o�������7o�<u����lvv6lj�\A:�.�q�5�Y,��d��`\P�L�,|M�x<����Cej��\����l{����퓏��}��w6125jV����IP�\�]�v4iz��ԀI��i�e[y��b/X��/���4�/x~)���ǉ��E%��r�O�5d��Lu���i:��=3�����i����}}nhGY�޺�ᦜ���=�1eɦ�q���h�d�˚"�:���kOM֝��]�[8ڔ�W�U�g��6]U���OW�]�aMӞ��=�Yp)�8��L�3�&��45��.d ���I��8cf�&ѢM����f�Xc�,��!�PDr<W�f
4�?E�Gy�nx�A�A1yPM;��mX��䅱��H���P5
ˌ#r�p���2{ �h�F[<�w�?Z���D�h�7���q�e�y�wzp�w��x7M��0�L�T�_25�S�S��d#5H��E��J.��u#c�����'}������ţH"O����8*���MF#���C��d*�@�,�H���l�f5�x��+�^�z���~do�V!uX�����N$������Gݟ������t�'��O�����w��x�W�;����b2x��ԸLM���R9�T�-�!�D�%cB'������*�eG��멩���������O,n|��Ƈ������xy��j�K;!�^�1�w�O��U�����Q���}d��"�����?�-?��|i6��Uܑ	����Ȩ%��"��(y��\�"�20�9�b�5��E�F����A��m�����;��VŇV�G�G&��&��fٗVٗ�gFѧZ��7Z����Uӫ~�(���mH%���6D��rC���%�M��3��G&�G}���
7�����D�$��d�wd����4��4Χ8*,k�4(��yG��'��'����� n�𷐸�����끨g�W�/aP��ub�X�"V��Uz��?M'������b�9��R���hD+z�	�hI˟����ߓ�;�e�7s���NM�j�6��j��VD�����k���z5������ԇC��:�����n�� �VBIP��T�]��X����f������h�QR���a�XO!�KB�S�J&F�@��(�����!�H�n�8��� wb�������F{{���V��~��C��%���
��`�X,��F��O$��T��`�`DdX��cܷ		!*Vb�0+RV�����5��Z�5M9��LQm:�.�[�e?5��[ӥm�r8�;O�W��ݥ�MX�M�+*I� .Mpi lm�����h�/k��a�-Q��OpL�x[�Dԥ65��5.S������Wo�x���w_����ߺ{���3������w�O��/�ݟ�+�fv(in/,k�f�cg��3����P����"h\@�NNS �{���2�l��h`�ؙ����0�h�l0&��c5F'�}�l&j����j�p��^LM�x]�dC�\G���h0l����*p�e��:�`���-�����4C���j�p�L+t` &C�Ɓ
}o���\�W��-U��{����"�@�j�T���P����M��̦�l9���������g�����Uj�*1N:�	��F����y��b�h�q4�<Yd�e۟k�.=ٔ��@��+�ϟ��3+�t��G�Z<����[{�%ƌ�56뙰�s��2r�ok�pO��e�v�|�����K�)����bR�B�u!ֲk=��XO	?�q>%�Bb𕤐+I����#�!� �j�r�"Y�H�L�5�`U�YѲ�hX+*�9{E�YUr�T�u5 &��� +2�y%난y^�X�ѡR�pZ��5k]�>�� ִ�5�
�5��r�I)億|\L:&"��z���e"�`fi�n��_��,k��O��9B��j\��&a'��l� ҧ�Ջ��Ayu��:�^��5M*R�A�e���1�i�D�.1�M�kb༧�t�U�!�������"�k�⦋��eۣ%uA��fj�� ��Ra&�8UA�
;dj�'�4�[���[�ۊF'�{ƻ�����h�9P2��xq&i��#sG�O)=��;w(gz�um�����O�ol ^�q���7[Ϝ�u`&ed<��t��b����������Ź����������Ņ�������������Q3#����Fb��K�lo�$+���v;W�������q�$�'�!���h��cYz��H��B3Uh�L$���3�8r,�̓:��@"��E%w�׏���<:��6��C%��A�`G-���D�(�B.^����X�P2֓�����8�N��(L�Ő|0/�����a�i�6����X�H99NM	���dH���s�\�&I�{���4M~(�>	65 xW�lt� ./��jg���0���%Wh�R�N��w�(�����]?�������z//w(�α��	�ʹX+#3J�\֐4ؐn��ט�!�P��G�t��;}������׎�~u��٩cå�历hk�����[؝+y(U	P��a����T\����i�T�LMC*Ľ(g�ljj�p�ڪXi]��9MW��.�����Z����a��O�=��O>����y����ps�vw���@z{"|���???�ԠP(��0������j��O�Hΰ0
�<��7�s�@���섚t�p�8�����1����l�~;�Q>R�ȧ:$�h3FA����$��+
�j	�\���.a�g��T��n	��X~u<����ue�2'X�f�x!EF��L�D ;��FOt ���q�,���X3Sӊ�w����hk?v�صk��z����7n�<yrff&##C�P�p84F�.�pp@�vt:�`����:�%&���K���vP��(�wx�ع�ɧ���#O=����'`Sc���-5V��SaT�d�gG��Gä0`���J���~Q�	�e ��>�_/�q��AY,8�T$J��U���sS���8��8�2U����HQZR���d���h��C�����6�tV���G&���P%R�ȏ��T�/�o:7�sv�����ka�7o_]\wYh{!T����MMG��3�;�-._p-���48��Դ�����P��n]2��ij�o��q��4SM�5'X��fWK�*�j_��%�
{��|�;�ۼT��{�nG�y'"�r�E���}1��ظ  AH�Rs(��0��NB�"�����^�T\ &2k��x�G5b�Z^��������'W�����D;M��0�������JLM���f��Y��Q�Cn��XћL�Ƣ=�������C��Ih�F�`4*�D��"��}vx�m�ض����D��� a1T�B� ܼ�G&��|������������{��zmx��l�G{�YD�R�����q
��1����|��������o�G��n1d�,:��� p�"5�41:]�ɒb2E�<1�P�-c
��r1�QFR󧵲%�rY�X���F_O�?�=j�2wl|�������/��;Y���N�ٷ�;T��Ɵ�֍�ܿ�F�-1�OI	�K��11�/?ڂ���Ȱ/�w�;
�3|�*s��_�Q�D����5	뢜��V��Ysۦ{+��v��-��U��U���=����C��#��3����+��s��S��#�S������:��*ُr�ߤ�Ģ��Dr��V��Ӂ	X�I,����#���'.kC ��a�D��He�@g|O�Kg~À��@�O�G�GyKzC|MxCx�Hy�Hy�H~�Hz�@|�@��ǿ�ý��ncp/c�ϣ��Ш�1ȫ�%�<�F@���+�*�FǮ0	�\ƚ�}Vʿ�_�J/��M��f�q�pI˟�pj�u�)gL�ܧ�Y�FF���GOiԑ����L��Ӫ� : �5p9��j62`󇚚j�&���Ը�j�t�-���A)qPJ��`RE0aw��QlD�ZI��-�L�L��#':�Xr����!&x+i�j&�db�T�����98_6և���\2��G2�(*&���'!� `BAа�^:��`a�|"NL%�T)�&B2�G�����,��g��R�E*��hr��������`�ǩ���)��ES��%Oٜ+k��3�ͩ�4�Mӓ��bjచ���3�٬i6������S3h�M$k��	P�{?=4�f���`,k`Ssph�_55�C=�����ej>{���_8����h�x_�p{�XO��Hᯘ����١��AH���A8M�l_�Lo��3�f���5[��Ѹ4�P�m��^5��bg6�ij��Pc�6��/�L�M7�δF鎟o�>��̑J�p�~�8���|�\Fx�We3�i\���{�!G�t4=E��"Eo���P��X��D3\z��i��2�Eи�la6���aF�!�P��x�25S���b`�*'\���&����Ʊ]���*
��Nx�`���_�?�ѩC�_<���ſ]=���C��>SY|"1�xx�1{�	�����wK˾�x��⵺���j?n{����٧s����.'I�M:���ɚ����W�¯f�]Nq\����2��iφjφ���s�Y���Mt�*\��M�3Κ�X�
\���
�����/�yT��J��*���{]�9��¬h٧��S*�I9u��Y���qK<�k�C40�0��y�?��fS�L�d�$k �"z���������ލ����t�|:q>m8�V�gֳ����@�sqBb���'"v�]b��I�mc���*)�L������Ru�y���X�m(��'o
���UZ��&`|(�fRm0����+����D�v��[�w�uv��4���3{�u~n����ř�����@Αټ�����/��̘��[95���~��w76.�U�������'��&2��9��|$ma>cy)��B�� }q!sq!cn.yv&fn.rv6bf&�����ɰ���#ñ�C�M���DiB"/(����U:��DѾ���{h:���x<KE�(�"9A ��e8�Ñ YCI�ź �9DT��p�+��>�~����οt�ꝕ���$�,X�7q�
A��I�X1 �00"J@�gc�hHw2ʃ���P��'���E|1x4������Fps'��z<)���J��*R��@�(P�*d�{��I��`�"5VJv=���e�
c���M�[{�ͦ�3p(�fSӜ�n���gj�ąт�,�tg�ե�W�];5p�H��L�`SZv�ء�Ye�9+R�R
lH�I�ߒ=Ҝ�*����CJ�N���c���NN|������~rte�z�)���޾˴;Q��������>5��a�"5��sp/D�%|���K�>hj�R����S�iyr&����z�c�c;�z�}����'��i'T�{�������,M��pL�!�H�ux���.S��`�L$Q���0
�<����vXF�P�~�`���n`��������������������B?�������uj�^b
V�%�i����`~)�&Y��.ݻ��.
�j`Y�SS�IT'(��T����K�T�+�B$�Z��G��dD@��{�4.<w���\_<#��7).>:<�n��t��N�K��[��~��w�y��_<~����trr�\.�\A4M���U78��N�S�7���+x<����x@OO/���O���O<��)l�ljB��h�=S��F�h����I7``�|KXM��9����5����)�����DUI��Ɋ�I��,cGqhgI�HCr���Du��,CI�aJB������	k+K�������t�Fk��`91���Nu����|t����gO�=��yj|�䞴ފ��b;�)KӘ�n�TBE��Up�n�K�f��o��S?�SӒ.�eM]2�6�_����XIK��)ñˡ��-t��S�#e�=T�=5;�5�:O�w��i�CY}�V/��#0��J��&yⒽ�)~�d?L�*����L���h�T�n����NG�"������X�x�`E�X�7R�ӗ���O�{L�����㤬D5;��O5��t����JLM���j��Y٩A��ȡ�x86��r�������O@�YT���	2	I!����gֈ��è5�5R�ͨ�3%Dc#�E"�&�N^�x��˓���έ�������D�$�`hX2�$R�vB���\�FD�=�;%�x������r[�/�����x@��dJ�bT�	�1�P�*����^{� ?fѝ4�WMګa�R�礞ߕQ�%՘�_����o�|��7n|���V�1�#N�	������/���6�S���)#��)�$�~����?[�������Ã�6}hӽf�?��=-�>�\ъ/����u��BpQ-���_3(_־�yӦ~êz�"�e��5K߳H�7K?4K>�ʿR|��e�{
��J��j�7��Ԓ?�$���,������g!C!�P)~�K�*�]!�I&��T��X�w�`C,�	�a5¿2�?��b���d}�d~�d|�b|ŤA�}Ad���c��=��y�@y�@~�@~� �����{��������n`�/��q�gp�+�E"�<s��=���e��r����u!�J|Y-��U��YuѢ:gQ�Z�zᜎw@͚T3'4,(�F���{t�=�UGn�k��j=a��>dV٨0�fm�� �C:�2���S����f����	Rj'�S��P��� ��!��	�vJ���c���I	
r�o硤871�]��P�}�t���hX*V�@�X���Wq�jU�"IxU��<"�K@��� 8�@0�P�^!Nog��ZJ���9�&�PDƀu	�d�u|�Q�6�9`�d�@�فx����=���(AY/�HפK��9N����!T�+C֖)o�Rl�4��t���"k�Ĩ_��٢i�eh ���%��M�@k�=Y��>M�:S�:~)��`_���X�@����cL�wn���M0��O������kK#���O��r�zrg�~%�in(en_�� ,k�g��b �}�y���k	�v6ۙ��IO�5���{Ń����l��25���/��M�f��:Qc���N����]l+5��*��n��Jݾ2�`�r��W.�WY0R�5�s��R8mo�j�D�� zJ�i��B9PS�(�.��C�N��V\l1�[�|����{=�� ;X����M���E H��35'�������c��]֡<��.�haȥ����~q�����{ne��6^�����>88rwo��eE���)�rIc��lL�u�u5|���AG�'�Mߎu���p�*�|A�Zn����i�+��kik�a�I��a�2îfE\���l_�7�������Fk�E��E(΅�χH�������+zފNpF���)5�AN�٫*�.=sZN;%���Qִ�UgM�]5pW���Z�I5ㄊ~LB�E�%n��]�a`�8��#`��F0�ga��P�n��qe?A�OΘ��,aQ��1�G����^�����;;������v���W+Ϋ����B
~�4�"|��G�o����F�F�/�cvk����hIw��+�%�!�k	�6S�Xkg68856�C�2���edj���<��6-?J��mn����;0�4����T��6(�i�`y&�0 ����㳻N��\Ȝ�L=�����������������?�x>cb"al,nl4aj2ca.�ؑ��GҖ2N.�_J=2�vd>sy1��b��|��l��B��|��L�������!��ֆ:Nb�4)��a���6�H@P~��'���&�f�9LWB����$�|��� XX�Z`օ�9R��֎]~���?}�wo�����r���nu�O�E�da��E��Hj2^A��)% L�h	+áĨ > ��FJ@�=Q(� �
��g ������A�r��l�RB��"CG�1�ʟMG�@%��L�o�J��sx�� [LM����0u�2��4f)��U��LUE��8VԔk���[���^Y�:7�vt���(4BG��}L�� I�R�Y9ܜ�S7�'wKv��g"؁���z����'�/-t��g��u���jI�
�+[��ΐ
�������N��i����q��5X�MԜ�Žj�R@M��6QVg?�%�K�d��W�B�0^h��^;�p��������q�zB�gj|�|}���p�M�D�y�ϗJ�b�X$�{~*�J!��d
�A�
�<�V��M�L$��Ȩ�@h����-�N�Ϛ��/�? �������65P�ģ^O>N�� �tR��%gD�I�̯�����??��6Y�25�(C-QQ+����8��!�(H��K��;T���٥�q�	��=���n۶#�X4�D ?j�i7���888x�ʕW_}��7޸~�������dtt4�Xx<\A
E���C����h���D0¾L\���_o�O���K �x�G�?��Χp���  �(�p�86I��gL|W��9� ^�����Y�~�o�5e� qE<��**���)�=A�5��Sf�����aJ�U`��*�1FfF��<#��4��6��>��"�:7,7V�"	�����{
V��.y���s��������f�gzr�wGv��U���蚳�-Y��O٪�<mw������h�}��4�Ch[�-k��� M���~]��&IX�(���dX[3B
�5Q���ף��@��������o�A�C��0!K
C����~�HoT�'*���M���Sp�>�XD�G`�:E�!0+��B� MK ���<��m>�'ܭ^V?�= eĚ�1:o�l��h�7�;g�520�ˈ3��?Y���Lͯ��@�Fr���`fG86%M#ċ8w��v�m��� 8���4i�+/<8��-���\�%K�'F���K�b�J�:�G����Z\=�z�ev�l�����K��G���[91w�B��HQ{S�ʂ������Ĭ԰������T��+ �$X=9�F����@j�+$ ���,�S��)Ag���bd�U$���%��N9��Yv2ԴlX3k.�X^N�{�,����n�<��9�Q�����}��W_���K/���)C$�sJ�-��� ���t���R6��Z��mf������#�
w|j�&��MT��7�ڗ��,�g͊�F�9�xU!8#�ȅ�r���Eu�,բ �f��a��i��i�c�k`b��P~��2H�U��������Z�Z��Z�;���r�e������7\�w�wbX�I��ңԊ�bC!��D��P�_�w w����;�6�+6�+&�+
�2�K�s�S�#��=<�.x��{q���wj<�e�%�y<��{���B�_f/q����%9뒒}Q�{��>�p-��l���Msޢ\1�N%�FѬ�7�a���Z�~=kD��1:�X��h�U:|�_n$������J|�����N���j�2�\�3��bj`Gk�J��k�PL*���P�B��iĪ`buD��XL+��2��D6Z�q�f����g���:f���2q1FZ�Byx�f����|�A@��yK�� �k�T��Aυ���PR&���d��f�2�R8���j�D%'�adT4*&,���"�(��d5� ��d$��1��S1�����H~A4{���M#��Vo�Rud��r�����&M����|�A��AM��D��e���L�q�=S���4�{�3�bj�U��o8��	b��ɿfj��^{p��;pE��~�ε���}��F{JF:�&�w�Le����ߗ:�/���)i~0ano���XH��G`S�j��Ϙ��n��,�_�?�Ԙ'k���Ӎ���։��n�X�a�Z7Z�ݿ[3R��P�+W�)F*� X���1EJ T�c�oj�b_���T}O�l�) _�V��D7Rf+3����F��å���E��o���0����_`�������@�枬)4F��wGwY #�}��9��l�PQ���C�}�7��������7/o�|�w+K�.N��\?d���*�l������OZ�7���H�G]u�48�t��셚��*���\�K��w>+�\Z�zJ�����Ya�s".e��KZK�����gc�NY�<�8.[��9�g�%�F��A˚��i��fA�*s#g�ʡt'���I9dj�hX:6ഖuB�8���S�D�e�;�y.z���e#�q��8���9&z�����s4p��9
�@�"h��N��4b0��߇����t#=;�;ݻ��]�.�Oֻ�_@;ѷ�������WH��;��6n��"#4*�*b���[�߭'�Xh���P.��΄"e��i*��*�.����"h`�l�j#��&P�M���> �h����HUc]��������{k'�ڎ�=w���|�9���MM��y0O��_�n�����kc/]o=}"y�?~t$z|4zj<~�`��\�񥴓G�O,��ZN=���<�zd>}y!��B��l��L��b��|�ġ��	��Q��������j���$'�R��,�������~�8��i�>b ��OE����4�G�p9���p�J��ȧj%,'6(���s�w�W�/͞�կ��������׾}���㱉����:�J3Q�&<N�F)X����x�9�HQHX��<V�C�(.���`|Ph/������$�zP�v���v)�2t���r��W,k`SH1�̤L5'����a��	���&.����D(j����<�lj Y��i��U���e-����9��[�,w��4�n>�_X�����Ul�ke��)�Cz�b�S��"aSob8�\�o�������9+{n�[\9�wr���p�ds�PUx�cO��1��(�j�$�`K���5�P8� �]���N�������%���B5�r��pC��4Z��	��d(�	����I��O���	�~r�	u��q������i�Q�op��L�:{<�L�|>�Π�),�zl���;�F�\,aRiX$*��������z��i��u�Q$�B���;;UC�k�"5�}����<��6EZ6�.�D���rү����O�%15��ҪQyxd!�@�	��hi~�4Vˆ��Hh*
��:p�x�{�yy�� �+gR]ݗ�?�$XA"h$2��֨ԍ�����/���[��^����866�p8�e"��
��h��E7�Ԁ���7�@"�p8�'�7p�����=�05�bj�/	��rZ����9[�c)�	�40��"59Vb���Dv���X>��(���65�𾩁My���	�
�lO�v�EL�e���ݷ��04B����|?���K�n~��&/�cwJ_}VgUjCa4XɊR���S,Ǧ�^�8���/�?���6|ce��R��`�PmlO���2��[rt���,(��3_�Sh�/���Npޓ˳�������������9���@}�*c%���T�.�<�O���X��7 $ ���9�����{�!��� |�7&��N�Ƨ��2Ќt=%���K���'R3q�|���&�$���8j�%ʛ�m~����o����"�~h�/����x �������2��2c�D?I�S��#$HIFz����Y�`gHU+�� �Ԫ��l�B刨(,��~�ء[/����g[֎՝��?9�tf�u������o>7y�:S��O�|n��+�k��^^���~z�g������v���|������������cû���rKJ������:y�^�$�&�hY2Z���'"��`t�(�ej���l	*K�ȗ��d�"	����*�L�ŧ#�"��tW�[i1oW�z�0m.%<�P�������o|�������ā�t�~>eM���	E}�~�'�19u��b����ʂ��r7�27��7��~b��a�:��m�㫸���-��o�Y4W��s:�RtR�;!柔V%��Z�Z�M���Q��	�u����M��A��Q��U�E���W��/�����t�ϵ��Ԣ�բ�Ʌ?Ȅ_p�IP	3ȟ����_��Pz�V�w�vC���J��T�W��|�_����D?	�?
��s��2��о`S�`R��1��0���5��`7q8��y���M$�$_&n	/�	ϓ	�Q	W�g�ԧ�����g���t�kF�sfɳf��p�Ka��,φ/�5�&�I���N�h�q�T�%m���O� ��mZr����25B��Ti!W�bj�#�:=�Fr1A�_15!��i\��fjyPB�T;H��` �*�ZL+�P���x	:J��,L�0	�!�Zy3e�b�<���1�QfBH��(	�&c)� ��i�2"�N@��I 0�)`F��f���ռP�0�(�4I�uB��A�'i8x��GsX���,����B
�KIGKH<���1!~;�u�l�e�Њc�5i��LIK�3�&Sٞ����v��;s����M�/��_��qi����̓�15��{��ɚ���ֈ�=1S	�M�Cbj�VM����f�V3����05�{�6��x�ݷ^�y����}�;/�;3?49P���x��`z�xv���ތ_15��P�n���gj Y�45p������]���lj�[���q�>��s������u�M�~�^7^����l�55��Z�:��z+�@�i��0Q���5�3N�&k��U���J��n�X�q�q�� ���+�i�B�e���w�C��_��M4:+��+�
U��Ś�p2x4�x�y��:Vf-5oq+.��Ƹ�"h\l�rce[�G��n�~���F�-c�v��b�p�u �Б�+	�.uU|pe�oo_������k�?��ޭ����t��G���:옕����E�bF.z>#�ۮ�������飮������{���f}��s�-�x�(��䫹	�����C�e�^�	��z6պ�hZ�7��Wc4�њ�(���Z�t-T�"^��$kV�
x�6
O 09c�r䔆}RN=������4P��uJŀ���N�L�q5���� #-H�+��v����9CAϐ A3C@㑳x(vf�,�P X�������@�i��i�p>mh��p'ѯ��A�R�8ؽ|�+��4"\��*'6�Hps�=��Yn��F�fևp �b�AՂ���Ukg���8�:��Hj��뭴j�*�Q }:�LMZ���:gp��{bo�`O��`���S'+�犎.82��`ޑ����y��?\pr6}f4wq���R��قC�#���ӣ�3�1�b����$��O<��tz���f��/J^:��p(i�`���H��OZG-{������mS���������E�0�f�R�%z`�8�/@z�v �T� ЇF�I�,��k�-"�]��s�2�b
3ҪJ��j�:;��]z�֗�~�����������7���{�t�HLb�=�Hg�Q�3d��&U�K�(��a��,~8H���X� �͵	xJ>�� 3Ih���	Dy��=���^d?Oj����k��8���o65�� 8*�Hp��� h��`��f��`�[�"���6���A4.M�dMs��.C]��j�e�jK?3Y�v���xՙ�Ʃ��]�
��W��H5.�L��2����V�6���O1z����A<Bt��P<�G���vh�����:=V=Ւ�W�Q`[;�O�����v�]����Mm��B­���5��x^u�5�-dj�)ʺDem��)U�'�ؘ�+�U�DiC�<	A�xa�v�zl������<==��>��*
�y#�aAnp���S(���Ű�7�D"�l6�B�0�\&�"_�RY�!���`��dVJel:���"��!����l9u?��Y���0XT@`������fS�����}罓O@jX����_��������CY�uj��p�dw<x�QwU��8R�"�Ѱ�:5TT ����@��Q�Ph ��{��8�A��5��w<��G�`N%��B�J�jjj:{����?��������͍���L&p�H$�yc2�B���b��|�9M��b�`�;�i�+������܀Ҳ6e?݋����((J"ljRt�_�(�����&?��+�����?�J��=;�ZX˂{w'JaYS+.��֦��V�-��?>R]��WQw�h;�|?#�/H�����Fnf��$�^��R��P[���L��=~����ן=q����Ks/����2�©�g�;��/iH�)s�U�����Z�� ����J�p�`�Q�_�/��� `SӖ#ߓ)j��f������am��&QV��lJ3�%�r��2)��5��z�� B�?��G���|p��c�F��1Vo��gwG�w Cv�c�II�$$3��J@�R�������g�S���@f�7�C�"��16O����������S��)w��v��w�p��+���-Rʊ�	u�����6W���J�MIs�A6�� 	͎���zi��j����c�3�S���׎w\�0�ʵ�ן~�}�>;����;��_�T}�d��R��@����/�^]�}�J��S���'��=�xba���ë'&�/<qt~����|��p�ށ���̔�萂H[�U���g+X�2z���/&�I�bb����I��%�,9.[��MM��X,E�1�D�=�d��b��B��r���Ԉ�+so����es��,�Bs�Ow_���7>�x��o���.ѩϒ�/bh/�ho�E�����h��icO�Fc�Fy�Fj�FL�_"C�1d�<��I���P�kíP�5���Eu^/;����K�	���������Nt�(�c����5�-�m��}�� ��!�/����"��$�� �J'�Z#�V%�N!��\������	��������������\�B�'���Z��4�e�%��.��]"��D���w<���l��ҷt��4�wT�Wd�dH�|B�~D���'�C �M�x�H|�����r�Fy�F�M��̤�Ħ>ϡ>ǣ^3����5�̒�/��^
U��y)��b���P�3�E�f�,?�-�p@�>9e���/'()�jj��Ҧ�4�ɍ:R��Xe��*-d(^;L��~�VSL���c�Ps?�ASS��*h [Bl6SB)�����C�����!�"��O�����'�q�
B��& j@���F�ɡb|m�!�<�l���, Z�$��bSm�]zߪ(�9�,�%d�IJs�cS2��,��>c���F�C�r(�Ar�MJ�J(1�X	V0��v�$$�Y(9-@H�b>��ls(�9���Pfv(�6KV�!n̖�5m�ʶLUg��'���.gn8p62�M��h�j��R=��f����L4�L��35{�'ۢ�:�v%�RLlj`Y35����)k�ߙ�w�z�����w��ڼ~��ί�M���*��-�.��_4՗63����M��>H��&@8M��@Կaj;	�@�fϯu��%����Muj��Θ�����Z�d�i���4����C���M60�7M�/ܭ�W�5etC�P��h�i�� �Ԍ�`���B��0���5%��bexNCyO�J#��
� ��/7���/[��-��Ŗ/w�O�Xӌ��G��M��L��b�D�}�"��e��%��y��4u���W}n���g�m|���G77޿���������/�39~�j���2������cj�՘���*?���@�g�-��y�}���җ�v=�;煊��e���=]���r.+�|v蹬��T�J�y%�5g��+���H�j��L�t%Dr�!>$9�8��e��h�$^7K�Z�'5[j ����2ƪ�yV�9�����Zފ�{R�<��8�bU���9	iNH���|�,{��>�Bf Ӵ�Ct(�f��̳0��,5C��h �p�al��u�px�7�?��7���ݍ��A�vc���>p!�f���w;ſ���b ;Y�.�W���ĸ!f��"B�H��J|��P!�Ra�͔Z+��J�m��8��:��ά��*M���	P[Jc"6��mT�8�vF���c�FȲ��u�{[��u��u�w�M�W�ϔ/*^�.X8��0��8�X>�{tz׉��ى]G��\�c�:������!��4�pd6pt.��|��ĕe0�^����������N��������
?<|�20n�1��4m횆FsC� -S��-��c�L��M��C#�q(?AC!h�n�G�@�𤢉J�1-(�,)�#��/��7�b��}�{�l��Ku=Ke�S�}�㳗N]x��k߼���'�l��Ο_~�W^�bt�����-��G���o�˩;�[?&ٵ��G�3{�S��m��QY���=�A�����r}�TiesU$���b��_���ߋ�.!��$8�G
��ct��IT���X��K��`��4�n�g��96J~0=/����6�I{��Ty}��R[�LT'
k�D`S�*mH�5e( `Ҙ.��W �YJ(�%[W��mɷ�6%.=5^�4\v�@�DGvA��"�7
�,�@�P�l��h/��ΰ�4e�oʉ�R5/����n���� 1�����c��C͗�l�nM�)��diӕ{rtm�z(v|/eS��fSӖ�q�W@M}��*�˚-��!Eޘ��OV�%ɛ�5mن�TmE�"?J�����������dC]���	�K��/��i��&`����Ԁ�?��aRi\&���Q��k�*�����!`����:	�G9�O^^��P)�@� �Ec�X�G"\�f�c?�����_h�<<B����0m���w���=S�u����~������Dqm�\��xYa�0�!���u\�����q~h�RG�(�#�8���������m;��������ǟرm;��ѩ4�����u�ҥ�ׯ?��ӫ��������:�\2�B0���e�� E��]��5���i�� g�'7�k8lj ;���䣏m{�1�O�ް�	�Q#�$��qv�F8}2YsOиHu�d��yvra�8��D.
g�Fqʢ��q���K�A?4(1P^8�k,B��S�����Yy��$VT-�I��K<2�{�P��HMN������Ox:��E��'�YQ��DcY��"3�(ٜ��6��ut�?)Xttrϝ���x���3/��]?�����W�;��W�_�厞2G[�	
��մf�����.}o�yo�����^ָL� �M�rO�К!nN6���:ⵉ�:���*F��f�3	vƀB�����X�'��M �}�F�! B�-w�*�q��x��Νd�g�a��@v��@�C��0�4��N�2�A���D�)-��0�^t0|Yz���v��H��
��<��{қ���)O�;ž~f)�M3��$7E�L���CuBd�~1�&���2���Ԙ��$@���fe&Y9��MM�h١6Yx�eWSEQ_[��ުɑ�ɑ���=�Wn\k�v��ًUWV�/�*9�����'�/�ڵ~����K'��+8��K/�(9{�������+g��^k�v���\��3�'���,w�N홞h�k���[X�omkٕ����cפkYJn����H�9�{�&M��Tdjr�\&K��%Ŕ�H�2t6ë����p�����Xυ��;�/%��-��f��zu~�����mS�uri���o|��Ʒo��cs����������dw����7:6z[6�[6��������%�~f�Т{ת}צ{˦-��j����9���^����N��'�9M¸ �?��<��d��4Kn[�w��[z�+:��z��f�'A�/C�_84_ؕ_�U_[��X_�_k�_�E�(��*�?h�`|��|$b�ϧ}(`~!�'��Y��Q���R�g��
����咿����q��3>�P?e�?c��c0~Ge~Ge|M�I�}J�|B"L&@"���ޡ�ަAܥ��b�_gS�ph�pi���[|�!����~]����hް+n�jnG�oE�oF�1^1=b��П��W,��&ɢQxP�U���n1�[����v%��@m6P��P-�Z#��L�v֦����CQag]a��Ԁ̫�P��?oj`M����=S��8ev�NM����ŧ��")UGIP�#$�P!.����6.2���X�h� o�"�ML�K�AR�]�`��t��
cs�+��W6c���"x�` 
<��O�s�F~|0�C%-PJ�aw���wd�3-Eт�HVW��)CԴg)�d(�3T�Y���fS�5�4β50�S���75��{��ɚ(�i�J}:ؙ�K15S�S}5�45�:5{!M���Լw������G���˷�^9wd���ɞ��^���[/��{���!�`�7L�\��u�ӝ��4[]	P�jL�d�e��
&p-p8^k�ve3��D� ���/+�^�h�n�vd��u�`���iSЃ����
��PFv6�RW���3�Wǫ���v�Jt�J4��p�0R��_����:�d���0 �!� ���1�?Jg�a�D�u��6^j�_d����h��2�:���svj��g7>���7_�x���;77�����#�PU��O 8�1�S��(U笖wJ
�>6����w�j>���NOëm7
�We=S��tIʕ���y�r#�e���9��XO��%Y�-��Ƶ��1��h�Z�n5\{6L}!D}��8o���J�Z��,�	��Yr�"{�"�j�\��/�y������+Z�EL�5Jϫ�����:������R��J�"�,7��A�FB9$$��C|�a�0�0�&�2�ya�I8�$.��T�,	5�GLx�;������Y"p���!a�n�8�(��=�����֏��EA������h�v�O+ƻ��L�n�����]|t��J!:$�v1�M�i�bZ��IG���jt�*#��L�����������f�րwDg�)��p�]]���0fK��rV��W��w�ȳ�D��!�U��u�C]��
��k���N͌�:<�{x��X��x��T��@��tޑ��K���gOO���'�����$��%-�'--�?��r*��Z��s�G��,D/����&��&���O���	�w��wJ�;���u�:t{���mam]�jyr� 4R`b�4
70�H�p��p;<Ph����Y=\ر�Ӿ\9v�|����g�ǟ���^{���C/5̽�p�����gs{���'V^�p�÷��ۇ�m��ŏ���v奏�W_):��<��:��Tt�ZT�jĞ3�'q���V3��g��{6yϩ��c�������v�92�u�le��@rP	M� P,D �##�9��d�)G&�0�D5�k�4(?B����&�PE��e�e��9v n�������	��u�/��I�pf@��.E�:lH�5g*����j��t��ʺ4EC�f�.����ɶ���]��J�jZ*i+u�E�߆���f� �HY��,Z[��I��W$V���e����a�?B��A2¡��ϯ^��?2Rwjd�dCB_qpG��!Uؓmh���&��?�KU��8��L]2��r�kJ�4gH[2e��<5�zc���[��/�f*�9�cy�񐩩��3�J��O�5�ȝ�FQ��I����|%�@�d��q��d�SOz�{x�{y��ݸ������7�����e$��u(��%�H4g� �3�I	8�|.���pL���S���1��٭F�N��
E�.*�D�`q(4�Ǣ1h$
�B�u���Q�@w���?���S۟xr�c���x
�����1z.�."F�1JB��@�*1�86N��S����?���7���(�)�[�)��T�k6+p�j��1a_S���?/���'y�$YMxN���OV�G�v����09�(��Y(	A@B��с~<�A�s�d.�¢�HX���������\37({ܼ��q8�˷�lUUUgϞ}�W�~��K�.��������j�XL �u�R�,g[n>�����l6Xwa�Ui�L����<���U<h� �(O=��۶'����/61P��;�(5��-GEK�T�{u��Pu�T���5izd��e��
B�E���(�^�*�f�c8����u}�6��%씭��eI��,Q\�$/�Wg��d��j�vj��h���d#�P1�بm>6HN���ܴqz�$#L�.K	ƚX����O��o�*��l����/-���\X�t��2T�j��H�PC|[�}O��1Wۜ�k�����u{J�o�`EоJ�`9Y��p�-2<�r���| �;�v��j���P5�T	ܞ��B�쭢9�P.OѰ¹=�B������$h�)
O"��8����/	�J�9V�"i���f���`��5|���qPZh�[�L�I�䪴�LGV�8DG3��ZN����8�~ [�j�
-E)C�h����Ǎ�c����_�Gs(QRf�������)ff�	�H3Q�P2��l+5�N/I@�zy�X��;���6F��ge;t��$
Q�d�4����i+�?T~p�b�����X9���r�ɥ�SG�V�g���Y;	 ������N]>Ur�L�Օ��gʯ�.�x��±���痫/��|��҉�sG+W�NͶ�^l\:T=3U}h�q�`�􁆱���������]Y�ѩ��L�6ߡ)v�K�d�jf���%#gH��\��)�����"d��%F�Jѻ��B9�H�-��E�1m��|*.�zv�Z��Ŵ��v}�R�yo��¤\�w<��RO��gom|��Ɵ����,��iUs~�7ز�ɼW��L�k&��
6F:7z�7��7Z�ؕ������2��ԫ�0��hw��7,�7�ͯXu��ʋ*Ѻ�wF�=�୪���"�V��sj���]váz�,y�$�c��iV�k�|h�|f�}��bj���l��ߙd�$�jE?�$ߪ_J�_HX�����>��6��.���������������������Z�T��e��$��􏹔OYԯ��o���i����/(�Ϩ�O�ď�������ؔwY����7�7��9ě|�"�	�zSŸ�e��qn����7�կGhn:d7Bdw����oE���	5^֝��N�eG�y=F˝p�=�Ɉ\��&ŵ){4$�Ѵ�Dl��[m�� Z���`����0�A@]0��A��+ׄ�k#��H&�>��Ái�f�C |Wm�6�� ��J�*�XF�	8,w�"��t@u8DU�;�ZB)����]VB���k��j��jz�k�z�)�66"��2��B�x�k@�6f�*@�qA2�EL4K�&1�V9HIs��ZX�-RX��) ���!�I)61	 &��"$yX&v	9T��Q�_���#��W�*��Չ��XeU��)]ז�k�RC�i�Nd��� ��9*�΀	<wٙ�B�@���:!W�[��٥��W��L�O.�������N�5�H�y�n�3���4��v�]�E�^pt�}M��A3���!x��1�6�'j�-v�-~�=~b qbO2�i�3��3':�';s�;�*TL�UN�VO����zh�sf����N�� �=G�5pn�l�fA��� ~�~���� o���˗O�]>4P;�Y4�U0ѝ{x wq>A�I�d.f/f.�������Դ�Z����PS�E�����bp����WT��%��/e~px���:�A�<�\�fo������	�KF����)'��-jf�٦�5�
x��<�h`���w�/5�á|�@��=E�/,�=}��+����퍷om|xw��76n������]�;�w�t����i��X��ѯL���_-��dO�����|���^�nw�+-�ϕ��ϋ=�y>'65�A��V�Z�u=�k>m�G�#�"�C5C���첋v�e��i��Y��A��Qr�,ު|ɦ�aWߴkn�nش�h%��:���Vt� ]W����i{YB[�fyqVD=  ����|�4�t�K:�!α�s���H',�K�<=�C�`��#�sX4lj1����$�	=�Gc������=���}�>D@2�Љ��@�A��ӄ�l"����٨�K��:�a:��6	�U�l������I��7�k��3��F�o�*xϫa�8�껤���<T�4��ÙMQ��Hh���Ψ	�UG�ʢ5�!-��Ս%�C����G�g&�fƊgF��ڟsx,{v<{�@��������=��r�f2��ML&����M�[�Z>�w�L��j��Z��j��J��<���С��C�Ӈc��81z�68i�0���i;�����͝��V{}���B��*vDJ����bIx:�)$��T�JnK�-���^�\�8�5�\���i��O}!k���ɗ��(<|;v�s�S/��;��4M�9��k�i�7^��W����+�����]��9�u*n�z��@���#�bF�%�=�6�Rt�Ÿ�˱��#�VB�O���
i<ꨙ����,���K���̀Ǌ�h:G�pR"JKGڅ�9>Z���6I���"���TOԈ�4a��-ǆ˵���-�N,��S�<���AYS�po��-�����r�`�'�ek�s�{rtMY��,][���"t�9q�'wi�h�w�鉚���]�b��7H��Z�Y6aE��%3��8qoEZsND��L��v����v�o��d��j/߿����XÉ}S	{KCz
l-ڦ45SUp��L��^��x	��;�8m55�Y��E�&�i�xNI�$�Q�,�bW�@�zaY��-�>�ơH�TMN�8��S�OE�O��H�m;{�s�v�M����������P}���O`�s6~���`�/t�~�9opL���p�\&�Mgl15A+�h�*�PN��)dg?oX�0X"�4�B �9�D�@�j�=ܷ���ԶO>��'�ܶc|�8	���lBB���o65�j���j�uS�+c?����5��:���d��X�i`S�CT�$�lj��"F\�[�H�,�)9.IB�b�qHͦ����E���4"�@�y���x{y�7www///�bs-KMM͹s�n߾�25pL�@��!�H
��b����pL�F�M��B���q��l{�	�mO�y�$ ���@->s�uj��!G:_�PQ矫=hj,�{�&�Z����"Y�)���,l�������Ai���iy��:]Y������U��������ѣ��6)��xRB��w�Xh���[٩!��01 -Tõd=�O���7%�ā�[�f�/�_::p�h������=�5����_����Zdm��Z������"cW����6X4Xn(5��XX� ��C�]̃����>��M{��%Cݜ�q:>Ic2Ԥ�١V	�����T#l~8d5� @
�q|/�؇*`H)�/Ê$����P�R�E�QKb��d�.�d�2��T�8�&�lM�ܕ�V��8:>~��������]mqQEKz�)�fH�ʣd� �/��%���dc�o:�)n�?i�/�7@��q)�2F����e���If��H5S�.NPi�_05f�K�d[�VF���ĉ���F���7�e�`U|vl�@{^w����驢��兲��
WN�9�q�h�����SYgOg�;�Z_���O�]8^p��l.�,�p������GJ�A���±�K��.�>��{u���L������e3Se�&+M�>8^�������6�xWZZ\jtPV��0�T��S�hY�jz���!#eH�l)dj��h@����P�)����>�����0]L�>f|)#�ʼ�k
����d�&�#yw��]���ݍ?���᝟^8��|U(�ɕ~�W\���AY.�$3������������?֔�TV�����B�ޱ��4j_Q�o�d��T��u��/��O�EU�s*�Y��NxRF?!����xBA[Ѳ/�W�����kF�K&���-��=��c��� �6��vŷA��U�ە�Y����$��D_��_8�W��b��<ڇlһ��,�G\ڧ��"�b��T)>��!��������-����%��9ʇ��A��I|�I��C��K~�K��!��ƿ�%�&$ݔ_Ro��7���z�-#����&x%X�F���h�+a�[���c��ǙnG�i/�5�V���^����h8�P!�a�ON��aMӮ&A�OFr���b�����aY�d�4؝S4@S�ƨ����F�!��%SSI���>HM8�6�&�Q40���א��!G�2�SB.u�J��Ev|��oF�P9F\����eE������nc��
�!|T��A|d��`Ce�0%�.%�$+8_���`��u�㐒�E� �6>��E�F��A��P)��$y1����ᛮgU�i뒌ձ��uS��9EՑ���TwBIO
��dI�3%`���}S��l�&}��O�pB_���@��Ԁ�ͩO�GL�����Ԍ�æ&bjO�T[<dj�`M3њ:ޖ�45YNS�7ޙw��d��l���@��@������:��9��0���15w_���Լp�����t�hG�XG�dO�����܇�0�RLljZQ�?5�N}r�]
f�j�lj��7�K��[�u̯ ��lj����p=��Ț�vf�ep2���j��+�\̃�g����&�� x�_�5p��qg3o0)����*rT��̊P�hyċ=߽xf��6>zm�77>zk��W7n��q�������ܨ��Q*�d��rA�XԨN�nd����������C�~���t��#{��|�!-=�Y�&�\��L��T��t�i��Y�2�ur>�p)L{)Tu%�0͵H�QƗ��/��n��o�_����x7!���7�mo�:^r����Y����K:�e���}L�XQ����<<���pXH��&yD����pI��?O�/��P�'"z�8��F�M#��vv�  ����;�.�G7»�׍��rҁ�mC����4�|�	��d�=�6�S���dx@��.E��lj���F=��Dl���$��p�o"�g�t1�0 ^ܲ��n�d5E��#�P���Q̪	�UEH�R��)�����ʜ�����u�����-:�������C�PX��T���������C��3Y3���MM��������
W�w���^YI>~<�ȑ��iǁ�������щ����QKߘ�w�4���~ݞnm�mu���Z�S �M�:"���"��,�)������¦]{��O��;�:x>a�R����+1{�&=�2�\�����G��M�����y.��@�����;o�~��6.���ŷ�]y���/�9~��u:t�r�г���s>���9|�嘡��k���:׃[N5i:�p,�f.�~1�|Қգ�����9�:KK%�Et��NS1�F!DB�RSbt�x-޹s��y;gh�l����e�f[�i��`b��T��MPS}�T�%k\���������7x���f��d�luG��-�ؚ�ߓg�.��9ؑ�0Ppd������c�%	
��GNy�&�/�Qĩ)�vQI��4V���70�\3?����Q���z˞Ynm�ʙ�Ӈ�*�jH,�-�Î�)M����I����k�u�"X�4����%���{R¦ �M�W�0CI`sv��LxOEm8��-�>lj�Ի"��F���G�{���o�c;{��m'���>�  S���	@�!P@gnx<�����|�X�0�P���B�Fg�.SԘtz�B)�.��A���&�F�рxb�(8
��c�3�c���N���/��4,���c"����S��15�j�`����g���l^wQ� p>]�p�%1¢a����X�xã Hh_,��	��75"6�Ǥ2)"�E�Aa5^P�www0"Q�i4���.\�p�֭g�}�ʕ++++f����c�X
7Y�ઁ��J$���*�@����+
��W����n۞ ��9$������p9��HPa�LMM��1W_��i�7�̽������gN�?u�=9H��n�݅�f!�R|���`��-�h#X�7���d��;��߄�H�cMϝ_��zb������S�F�':3��"�� YS`l�ehݥ�車M�ePXM_)����L��ml^�8{�9�}��=Gߚ�iJS��6ljZ2mٚ�(�1^˴�H>K�`qQ�A�ө9z9K#g�d\�B`�����[P�=lWHtYDrmLVkb^wJQj�ވ������]{RK�s�z�<7t���ܕ��������w��n,=����7?�-=�.>�4<(ۢ�Q��\��艥z���H	$��(YI:v���bf�ۦ&{����0"-� �b���M�U3оk_��خ����&s��:��w�h�#i'���ZN[9��~"c�$ }�8�X=����}�X޹��g���[]�;�P��\vv��ܱ��V�[�\_*?3_v�p�ə򥩢�c�F��F�G���:[s몲�������Crc�E1֒(CY�&O���2sT�,%SF dKq���bse�<�K
Q CJ�E|l)[H��*N��7����NE֛�����\v� �M�N@m�o���߼����6n?��z�Ք�#�m��*�,�|�N�iT|���Sc���΍�ލ�ƍ��)��")��H�]�������u�:ŋ:�5��i���^rA/��战!%�SO���-�����Nx�(}լ�kռo�l�~jW|$�*X��C�m�
�5�[���R��J��Zʁd���)������������	 ��,�{l"�}	����C��K��C��C|Ʀ|aG�������vWD�%��)����_�3^1q�Z���_��"��y;N7��j���k��[7�Wғ:�1�`QŝQ�(�J����OCPR���N�SM��Q;��V3��Ji�4M��h���i!��PFc(�)�	�j��*h�b�035��(�Ci�a4�2a���ER�#Ȼ#��M�f*�iaP[��}��oa�9IJR�GO�n�y�
QR���eay[��v��M �
�-� /��C蹁 01�V1�R�E�� ��.�9$� ��1���E��^z�����bu�#'TF4нC��T�8LZ����6�����k��t�{���p�lj ���N�S��]a5����8Si�ͻix+��05��j�H�u����:5�cj"~���L�&�ԧ��f�#w�#w��h����@��������=��B515CS���YS�Λ�>��]��;7�?w�����`�Xg�x箃�sC�F��՘�_����S������M���`��:����9�M�˪l���"k��%*8
~��O>���?
�5�f��+�*h\�L L��\}TO�jw(�!N:^wy����7>c��[���x��	u󙟮�~u������[��1�hN�:f5]���S������#sS3���j�������֒��g�\�
;�|:�t"Rw*ڰoY�5�F�"���p�Z�~=�p>�p9\w5B�l��Z��8˭������G|��Qv�'�q_�%}�+�뼤OӢ�K� =�����h;MsV'<���1�HhB�,� i.n��?�'Mq	0��C"�i�٤n���%c��4��i��A��T��ab����P3M@CIO�6` �����鷳�߭�у��F�v#�;��~mH�6�oη�෇��JhcB5,�i���M�H��bj�Ŕ:�5!Ժ(pfK4,e��ù��NS�eB�&�U©	��W'JL�+*szF{�N�7O�k�+?8\|p�`j8wj_��p����Cc�3釧�fd�Lg��8t(��������ɤɃɇ�2�����<v"i�H��L���!SSA�����A��C�GC��;��������ۇ�m���^}k���M]Ӡ����i2��1�rG���֙�2�P Ó�"�%<�0��'��`V�bbױ���=��z/��]��}���#�%�=���{=��X����SgG�_���7���7޿��_.}��t�f��]�7�{�t�+��um�Y]Ǻ�uE�r��z��v��r��~ƶ紥����阵�f�V1m�R&��C�%�<�&I(v�j)["gs��YH�Ӣ4�hl�S��T-ឣ���N+�iv9H`�VBu�Ԕ�	*���4a6�����4Mc�l�`A�t9MT4W�Qd���jK��jn�����kʷ�D
L|O9��d++AOO��ҭ�D�$H��cM,�CFs���uu����ݸ4s����\���>��8�3�ܐ�W��45��}Tz���(=;W&p4�.YP��S������oU�i��(e��g�8/����G����ΝP�o���z�x�Aš�p����˗��<�;�25R�L��'X�0�4��(�2�No7[��WkT2�T(�<�	���7;0�aY�C�1$��
���A���v�@x��<�� 1�f�M\��!����<��� �����`k� D(���Y�<HM��2VR-�M�Y�S��lb ���!��8���P�|�ˠ0)�G#���~>����������.�B�h4����.]�y��k׮^����255�p8�%���DWN^��d`�b����ۯ��Z8�o�I8�65j6�*"����
��K7�_55�K>�; )�տdjj�����\}9x��k�{�.�<}|��3���6F�����e�lR����#�t@���j�������'~k��l{����L��cC��NjX.;Н;��^�h-�v��ۊ�P������9cj�KL��e ����=�]
f��y��< kt�y��l(
��hL�
��Yʶ\�@etK^X�C�94�¨iUb3�*�0�\��hOKʭ�hm:�1v�i�d������փ�f��X��y�Ů嗆V_<}c����'^�^zv�ԍ��W�Oޘ\�ӿ�\��z���������=^ٵ�7y�c�����E���iMa�<�,L@�p��%#Sul�C�r���T37��EL�i2l���6R#�L��,b�E�Q5�V8�7or,gj,mr$mz"k�p��Ŵ�P帣s	�O-%�<H<���I_Y��kV��WsN/䜚+XY*^=R��\�v�|e���\�ə�c�ʗύ�:8�7>�� g�'��5��!�vwfq^jZ\j\Hf�5/�P�ZŹNS��a�h�
R���%���x@�(�a��U �	q,tɧO/���пZ�����W
���\ˏ�,�hZx:zg:�{�����<���;?\Zٸ��=]mnnG���$�D�:y�A~͠�29v��l�{����檿U}�+����w#�_�_5k7u���ʗ��ͪkf��F�%���VxJ�8)�uʚ%	$k�e�c2ʪ�yVź��'�l��ꌬyǦy�$~�,����*D�m��0�Cu_%����h�ߩ�ߩ�+��y�ȸP��}>��\��.�C�����vO� ��y�O��Oxԏ�ԏxp�{<�{"��RƇJ��*��J���w�*|3H�V��-��0�[ʻ���Q�S��'��&�_�3݉�ߊҾ�x:Hv\�YVr�Y�~PJ�P��(���WS{Ք.�[O�61���v�-�k��&��IK"�	hg��-QЇO���v�9���l�5�ā}MS,�ed6��4ǁ S�9��HzM��Tń��f�4����u�0'ܳ6��k���edĈQ�������
i;Mw+����p��,w5m������MIީ����^@�� D��V~�M���`%D����z���$FHqabL�&�<D�2�<�܀(9!��)�RU'�+��d�L�������8�Ѳ�tco�}���K�_@7�������w�;��NgS��-�mY��2���̌bY�����2��i�f��$;�N��Nw�7�f���ڝ�I����9�Z�m�%i�O��� uW��ր��&��eP@��d@;c�5�t4PӘw0r�X�M�Y��?S�S�g�f�>p�!p�јyYL͈2\�)ӡ�1�կ�����+&��'�[&�c]ʑ�_S��oAS��矘M��b�\o�xT_4�]��_�П�]cj���S&M3���fJ ��S��	�bV-�M��ټ�1��2�>�M��l�ǁ��d�e�	Ashj����*����t.�����N���/�2k��"~o�;�ݙÜ�	(��gr[�-�����G]G���7��5_<9�������_�ݵ���O9Թ��> b�SB��yQ�;������溣�����U�}T[�yk�vB�^r�Aj�n�l#J��݈�mG	7���0�F{-����ao�qwøW"��#����I��󃂤��RS���ʼ�.�Cmѿ���"�7�?�K�aV���Y��yV�1m��B�Y��.�<�H�3��u�bfp��!LbPS~��	w�I7�	W�q��������G�)'�I�)WGDӸ؏8�:��;Yw�[�Ϩ-�PX���>��;�d����Y(m/(l�+�ε9]P�,��,^VJ_%�^M4i����f8��Nmt�V�C��4,��K� Y\/B�I��R4̙_�V�^�Mz��y�Ѵȱ�f9�)�A��4�ajC�+E���nSiRS}^��nbeZ9ԩ���-�.����4�u&w'��$O$��L�&��%��&�$��������F��G����$}=�C��^IO���+��;��;�`����ת�5�y�J^c+��4��"^N.'%��d
�,6�F��g7/[���P����lk�U����/�_����w݈�>�Pf��i^����2����[�o���/����w�����j�ފ��O��m]���y�+�U�ᐫ�㪶��m�f�մ�k]㷬r�9���%a�"�jZR>��0"��$�^:�G��Q�b�?���g�{	�4�P�G�-��J�S��o4�Tu�9C��H�h��w0m+�,GJtCS���$Q�R�0�0蘕��� �h�[�8ng�TҖ�n��"�L�z*�[�۳��n���k�5k#uu�b��?����0�3�.��z��c�>r���`Cv��{�6?tkN����/�۽�7�<�ܿ���U�_��4�2�ڙ�4�)�ј�d��Id����?	L��5�i`�h \��ͤ��S��	��?$��P���y���٦�#�l ŝ�u�u��|��|�ξ�����Ν9� 15��,l�쐚�P�@S���	#2�_�}�i?/o<ƟF"�Xl��e�X4:�$��`����� ����x�� ���YY[���S��gN�\8�js��Ś�n��qa����ԘW?�5�i�Ŧl>OUbͦ<�~*�TCKy� �@~�3�|�����鼣�i[���6\�-ݝl�Q�nN�n.����vNv�v��V�8�@��@Y�ء��4����ڵk>�{��7677��ǣ���X��)Ӑ������4t:�D"a0777p45����njΙR��?!Uޡ��C�0}�D��38�H�n��jj
C<����MY��tva4�,�:�ɺ�f|�;����Ý�ٞ�8����?��~��vVLr�����(��&��M;����������s9�d��&u����;ԫ#U���=-	����BIK�PU,Q�TEBE_��S�u%�JYoMPg���\�]!K��E���� �F��jN�5$#V�1�Ҝ�j�h�c�
b2���<(<2<%.�0-��J;Q��Uh'ʺj�6���ʇ�
�7r�7��.��m��m��n%����޿�7�]0��?�]9{�q�^�����Ռ����������՘����������Ԋ��Ҿ��Τ�6yTi�,�I�qH\.�*"B��(>!^�Mc��-��G��i̦&Y�.px�~B1�'%3%��Ty��%��=c�'e�;��#n�;iz(iq"��D��D�������������/#$m\L~&k2.-el.d��g��d�����������L�/M�/����M�d�����]�T�2Y٘�\�Q_�Z��!���K��,>�����a{CS��pˠ�2)�d�\�+ ��M�	����8�lKۧWDXe�_��qUֽ��G���R�w
����cQ����B������~wu���;��4k$��y���|w�ܯ�Q7Ѯ��|>c3~TYz�g<�6����P������"?��ޒp����7E�7%���=�:�r�E�eb�ؾ,�U��2�c��@E.R�VL5Fw>���79��<�c�m�!��M��;�b����r~-�6B�31�WbƯE�����~�E�g>���/8�?gc~���	��k���i^�Q=H�0�������+�/�K��gDo�'D��I^��1���_�_�����/$��?e~��L��4��i��h�g1�OcE?J�41��X�;Ѣ�r�@����#yN�'z��܇��}d�n�[ӳ�����h�x�y^�B��W/�S"q4P�(�}�!��0?�����kv4���H@K�S#cv4�qx ���Y�4F�B#�B�kH}�W]�o]4�>ƿ!��4���	ЂMpSm�_u��k�>����A؂ �4���h)�|U��������� P�u�&�b@8/ŝx�.����a�-#���C6��
!Y����T�H�C,x�磓��׵���&p�k?��[�ɐ�G�R��`U^PS�(���p��8$�\����Y�lIgQ�&���dk3�&� }&U�E�dѵ�Ӏ�75fM���HsX͉�������15ݕB����uO�o��Q&�(������L�򯍩���'����?|�փ;�//.��J�ڋ��+���^fj^S3�LkC�i��lj�Syj��DP��BZN����W-��w9Ήݞ�s����y�y�'Hg)�<��t�q���g'e)�@1��65����e�`��wC�k��B^O>�;�ݕ�1�1zs�å��EA�T�.K�i���`�wo����[H�/}�����G�\��;�?ZbT�e/�D��]D�a"~] ��>��:�����n������܏k
��d�q���V�`3�w)���f5����fm�q���kQ�[����OR�>Ή�ai�/�sS_����?4��T�V5U������| �(/�'�i����4;vOH�ţ��P���f�i<j���)1�?z���s�u��q��r��t�@�CM3�`5fo9jg1fk:SN�Έ��pu��f�Ѻ�����in��)��*��&Ss^�`���DLPs^�b�t�Ry�(}mT�v*����h�a��X
�sө�vnẴ�Q�"�&�[�ĭ^��i��!�j��y>�渣i��"�-&Y#�4������P��`l�Է(���HQ5�f��CF��`�T��`�Xo�0"k�:��	C]I�}I�I#CI##��#���	#�������2vI�F��C�iuu��ze=ݠ;:�@�A������EP�"�mTU�99ټ�Tn|+,�)3x�A#�x�����c����U���!�r1�};�p�qMf�.mG�`��Ю��=�����h�"j]�L�6M��<���w������>:���Q��q�
�uS>�����ƫ<��f���f*�8�K��N�*�y�Q;O����/����S�����AJl���ċ��C�ƒC�$	C!�aio.�KF�ay�r���(��m65P�75H@��l�rdQO�ܷ0ܯ$
[K�J ךj?5��Ҙ����$�qMs�S�Ci��4�l��i �5�<!Y�'�K��"��w��o��-io�w�}et}��$�D��a/нNQ�P=�lB�h9�#��^_(��?���������W&wW;O��E��Tf}"�*� &�mE&�4�0��5d0���x@�"��l��`��Av~N��y�y�ǛR����8>6��D��w��x��}�{�^����p������g-l�[9Z�~����(�0��12~�<58?�@dRi\&�t2��'@Mn��e��'������:nj,ϝ����g���15b�s�%���{�Ԙ3
W?��:��c"�8W?A}���Re�I�$RL�@���V�3S�>r���'zX�۟�����7�,Ϲ�^@; �5^���.h'D��[[�X[BS��F*�����Ry�ƍܻw�֭[���8������Mp�T*8jfS�����L���=���)���;u��W^=�ګg^w�Ŋ�� %���h������|Px�g�.@�BS����ui��Xby<u�%�Ϊ��k�]�|r0~{��6'��q�������Ѽ�	�Tt0�CFA�>�φ�>�k�=�W�������m̏>\�}�p���ȕ���9�b�*��6JUؚ/j��
Ś��P���4E����������Ёڐ����J$g��Ԙ�	���/�4�T5L�jM�uHm��fm�,E��&	
���J�m(���X(�]��_��_��,�+�8(�8��\�p7�v�̍�kq�W�/GF�����=�q��	��9�7�V�ݩ��n���ԁ�����Fj�N��~����f<�j,�j<�~*�a"�j0%_�Z+�$�!B6_¤s��B�� ��15/35Qb�`����%a��4^3<U^��K5({�=��n]TG�x_��H��p��T��L��B��b��Ť���U�����Յ���H"��B��\��t��t��ɬE����1����ɞ����Ꮄ>]�Q��kKV6���e�W&fE&�����'��0��4�W&��4L�l�{&�EER����<�3��q,���<�)��~6��6�ۨ��nm�U�7�C�.JzR��8�vqꀘ�a�j���K�������7ݻvtc羲f.T��;���s�����]w��0���J�?2��z�GC���t�Ea�	�o��hO��#뮀~�C����ӑ��[\�&�w�����Hw��f��n�5�,�u�6���Fs�Aw���|��}O��DF�a0�g!����_�X������[�w"濊��&e�������/y�_p�?��C~������c���h^?�z~E������X���_�p_0�����1�?a���|��A;�e !���P��"y_Fr?��}��"F�E��8����d�%�-zƹƾ���V����i�F�����Pݻ���v����x�ž�R�.�_�8����F)Ǩ��[�|ͦ�4&Ss\�@S5@�@�����(�M�=�qSWB�͖X��bK"�5�ԖLV�RUi4�r!:���!#kL�Ʒ<̯4S"�/�M�;���H}^	�{-�t.�f�uH������B��!�Hu|�K"�	���<S(s']�����@�� _��+������"����$U�P��m��nM,�4�^��L�$�k�ԧT�oL��2��L�LM&]s,�0�1����BLO��hS��"���}��@A�725�9���B�])2�M3�r\��e15���Qeڰ*��E��"�O����O��6��lj~���_}��O�߸4w�ؿ��:�-�BS��O�}YL͔>l�P3�	��fR%��cj���CR�r ��\Sl�7�帩9.Y �V��'8���}�rS8~���T�@Mc>���`����C��o05�è9��Kbj�JE�j��h��Zg6�+O��h3�)��pm�W�����kG��=���ї�>����o����/M�?�y��r91r�������aD�OKJ�P�����K?)-����f��0!`;J؏��Jw"��,d�Sw3��n������(��hɭ���I��f�|Q���ڂ߷T�QY����G��#Mӑ�����~_Y�ﵥG��?)N�</�㬘��5&f���4�D7�4�m��LP�)���m�>叞�u�v��tswwss�q�q���@4��儣5���n��0�L���[mϷۜ�۞�؞Q�PٟU;�S9��:[�-�����ϵ9�S�,T^Vj_[DӘ�=ii�:����f��8�j.J�qmc��r\̚I�fZ���$f��!M�/�2p��y�-h���D�±�a~���mQ�f]�,د0 SISG�jӇ�Z���F���]��څ�֙���ޒc���Ț�ឤ��ġ���AS4�`|?��	tb��#�{B:;e��� �� H��"c��]'�i�:]�V'U�%mJ~]#��AXS/���VW��J�y���VL$+<� f��,6�I#��X*�%��<	G��Y&��E��E�W�;���Ҏ�"�5a;�ʌ�:�uߖu�x�� ��j@ۊ�~�d���G������'�x��[����h5���%L�Y�C���u�t�Y�EjY#5����iM+��Uf�
�n�Z3}�l�S<���!%(|��X)h�ܓ ��8���S1�\�������yGr=�����f���ljr�!�Ea��>���0��lj�Ĭ!�ٔ���港y&k^�i `jM�4�\�6O�-��rԅm12�j�� T�CU��T����[k������{�.��;
�s��q�� �Xp�Cm*j�_kxpy���ӏn~�d�͛S��]��ݿ�1V����c�H�Ud���j"�Mӟ���ܐ��o:P��b@�<�lj�8�L�Z�E�ia�񇂏;`�"d�4Ny<7����3���Ν�_���+�;�ԅs�ϟ�p���SScJR�hmb�����������H$��4�a��	�M��������8*�ĠPi$2\�n��������@� �������# �����ZZ75g��Z|cj8~N2"*�����{�Ԙ#k��me4�h����X?Om"����I@J}!q:q��Dv��/����9�<�<��[�as���qs��p��t�ss�wu�q������h���O�PgϞ
����4ͭ[��߿����;w�lllLMM�����x
Zwww�)�8p����#������@M~@�lj.�9{���"���bᯜ~��g^w�:��l��C<H8�B�8}�>�;�sҥ�����>xC�M�����+}e��;�����~���89'�[{Y�w��Y��.��� ��\����������gsa�Ҡ����[W�nM\]�ٙn��.�k��W�)Kaz��c�J4E"U_[ h/�T�4GL)b'�bƚ#���z���b}!�h^�����yG5��ނwD�6�R�)UI��DNN4?9R,�Mʫ˩��m�,4�J��u�������������ԉkiӷ��"�{ve];B�%~�&ϸ	������K�y�vp��-e�f��a�ȕ��ˀ��+����0ݪ�e!�i!�zZV:"+���e��qռ�<aP�@��lz �,b��x)6^��15���<]�$�N
���x��|��$�)
�gD�)��T�et�ZnT���G��'��=sÑ�#ы��Y���8�8�,�Z���8�4��l��t��T��x��D��D�,��.05Ȝ����m�jO��$u(��)�����������и�� ^���#��14�*:��N��e2<���Y�l�k�%��ȥ9�ѝA�p-f��P�l�<:��PNu.����z�Y��VY򽜨���o%�]��fy����>)��|���F^�ov�������o����=u��^�q������#�O�}?�����:*�9�QMvMv#����7%Y_%G}*y$`>�3�f��˦�b�����l�6�︩����Qы47�_�yl�<���{t�������}��v��~�����y���PH�RB�Z��e �d�_���1�Y��} ��!��Q@����K1�+	�.�~&�����	��5��k)��R��t x�/���%��Ĕ�D�Od�/��_���e��Q���xɗ��/�>�� $|��IRГ��PD�"�\����~���wáFp��PC��y��={Y^�4����x��^:��^���¨B|�>m��4-��m���p�2\|"��I���,zB�z��1�U�L$�֦-�L|1�qsp�+��d�:��N�j2�L�.�՞�1�r;�x�|>��t�2�ږL��1_����+7�+� o�1�q,K��f */̳(گ,W�DT%"�k�	��2D����� @�\������(<��
:�v����Œ�Ga,	PG#%!~�Q� L��37Ч8["���"6'ѵY\m�S&�vS�=���hj�EB�B}c����?�20��P�35�9���B�mZe65#M!�͡'�[bj���c��a�ӌ������޶��d��bj>z�mhj <�u}zo�w���_U0�ɟ�+�8P2ݕ�]cj&u�fS�i�3������7�V����*c�ʚ��[L��ohj���<5"�����[0�sp8��lL�Y֘�j�ʑl�/�lj�
y�Lw�P�K�6G`����&�?P���}o�S�|����/��ӛG_��ۧ���ɭ_?������ګ5�k�Qs"�4��D�]br.��7����Ǽ���qq����+q��p�n��j|���@��`F�@g+�{)���{�\��\��#��8E�~N�We��j,�7u푾�O�����#��HY��������$�_kK~V��~Z��ў�2O��%�-P<��(hj����i��<�s�1�q��EMz9#�m?��3khj��&�l&]�Ɯ�F���\�]��lz,�����`
a�"h��(��\��ΦzO���\�+�,U>6{%��P㌬{b�j8(�hT<���j㺶�\[��!�W�5�S��k�#��@s�@IPF�hR��� ��
h�0��P$�FMh����1A>�rBY�%'��$n��aketr�cr�lu�ouҰ0����.1���:�;S��z����!I�����������ttwʺ�"�^����*�Z%Q�%J��U!jj�Ԋ�j$UU�������BIV�8%���El��f�Y4,��� c	2�çE�R���x�~En�
�ؗ�ۯ�ۯ	�W���v����t�D�+�]������Ʃ�æ�w���M�.nY��-�j�I�L�!��*�x��u��y���B���U;��e�ٺ�lY#�͓�gi�s��J�O���l����I��Pw��/��L�ߏG��1}C��B�(�w<�5����Og�H:᧦Y�d25�r��$����D
��5����9.k���S�)HI��M�YU��3�YuO�'���Ś|�I�-7��3��m¾��Ձ�'��_}��������Y|y蓇��ܞypy�������{C�ݝ�򝍟v���Ϟ�~����K�W֍��
}]L[�0�,�жe���p��L8���J�)�	Sgh�'l`���L���#��5�O��U'�cy�r�����z�W���q���Y�E&��!5 �N����L�5fS��0"�i��I6e�=�5X_?�I��D�@$���&�g���*'SF�3qutr����hj��_x�iN��p1΁d�H�G����S����h�YӘm�
hjL�3�S���sP+��nj��q��$NV 6��)$8��l��,�N�Y�q�E�>��S�r�u�������8��Y��?�	O����V��}���{�>|M���tII	�Htpp@�������QMj`{�Ԁ[��A$��煦��i�-μno���Y~��TpDb٨X��"�0L'�R���'�!�^���<�P �E�UK=%�7:�g�ޙ;�W��"2t��$d[���.o��_������v�8��?m��N���=��X@Ssm�kg�y�3��)��2T]"m����u%]��{he�ڐ���Yu&qJ;�~�� @��W��hL�5fM� M���4�Y��'S*hEq�����ؐ�PyX|fF�>�m<�a"�~2�y.X�ݳ�w޳b�l�
��	�=�ݗv�������������M�n]�>P�[1�7�g%M�M�;x=��Jd�Ad�ܰ�^�.ɚ��3�!v^� �[�k�f�ɒj���lq�#�2ib)DD����+S�(�d1�\FΑF	�3"��*"[�õ-EX�15ÝQc=�Ѯ��������~��`��H��p�� jf"zv2fn*n~:n~*~v2~f,~j4ev,ezIH�LH����6d�3�t齚䎶dmK��)SٔZW��"� �F@	��9��$�d�K�Aw7�@&�1�ℤ6��b&���Z�q�g���Yd�b�C&�5%��^y�Ò��*Ү']O
~�8���ү�����t�>y���.���j�>|��?���/��WR#z]/���ء޵C������=O�_�i�Fۏf��F�GmGm5(��ez��!���� :H�C�ǣ��1�,�K,�5��PsT�,�@w�Hw��54���6�k�����e�w�=��u��v������������u �2�OE��鿒�~��}8�wr�oBi�
"�2��_S�)�
Z���>����q,��P�|��A��P��a�����h���>�|��2Z�����A_ A42�g	2��	�$)�䐛�.f��#$�I+L�)�먿Ra�&�jh�0�p?�GGq�2���F���~�@]V�Q��,��A^�!>�ԘS7�#�+Z"0͑��y>C45��:�8�lTI ��(�m��e"N�BlϠvd1Yl���,t
{�ŀ�	h��D`���֣5�\�)�����e.�A��XlU�:_��P��+��V�����)��$JK" :`S�JoK��~s�>W������x�{4���H�?�6��ᾠ�Ol���� h�#1%�^��7[��U��0��bK
M����M��Hh65P�@S��T��(�75й��L�w���,tU ���6Լ�� ^S3�NS�����f�X:�Q6b(�W�������|l�����>���/@�ɻ��oή����Wi�':J��K�z
�zs�{��{3�3 �]�s�i��о,�f�#�\�{N�V���7����X��?S3�L֘j �e�q�[��P�����0��Ƽ���γ�_��T6����y��`7�o�]�}��Ԁ�/���+佐�t�!�ўJצ04�tU2]��hKb\�*�;����؏�,������я���G?y��/�����?ښy��]u��E�`�L�ds/�e�b�6��'ߏ��0?�n��vB�X�a�h?\ 8��DK��N(w;���0ޞ�9Bt%R|3&�Ab�;���%}U���g��<�w�ſ�,�ya���&F}��e~���2�ڙ9��<a��i��L�Y�z���H�\c���|�0n�>��>�i/�1W�A���Ո�ը�S����5N6(�W{J�is�`}F�(,_WX��fs�����������|��Y$�����J�e����b�x-��Ms�0]�lg5�E�sUPm|� ���$�*��2Y���҇�M���| ��O�hN`65�im$�%	�1�4E����Q��r~(1'�R� ��f�Ltܺ�r���쥙�����)��h�dw鈡�1ܕ>Б�ۑ�cL�KJL�H��O����������	��uw��@�!��+��]��̭���7H�e�����BY^�(=���1���Jg�do*ѓE��Ӽ�L,����^PXI[z�\�n)�k7��ZH�Y�i�M����`�5���������L��Z��-��^��n^ض!3\�u��ߤ�/U{$�E{H�P�{�6M��To����j�2�i�ٸD��Ö�����%k�bZ�"��Bʼ�hR(�_���&��T<�M�
h�R�o0�G.��z&���P�4 L�3D�L1:K���,��C�BOBJ U����AyR��,ZX�		�1}�nZ���&婡8����-�u<�F[,��ՅM�PS"R[�yM9��TZOC��D���w���}u���Ǘ�^���ss���A��w�>{��w� ?�d�˷W޻3����uc�y@�����NoN��R������1�� ��̚愩��70؜FiH&�cjN �M����mk:���|�"�ݐ�,��&��a,_������7������2�?geq��悵��N�xF��L�L&���p8��`0(
�`q8?ƴ 
��������v�psquutB;����`d����.�Nv�P��YY�XX~����y���l-�:[��r�${:���g�-yj�Y�H�!I���}p�e���l�cC�B�KñE�>�!ސ�0��p��)�����k�+�xļ�3�T�2:C+�Q6'��ŕDa�"�%��HpD�TDK"�Y��(��@��u�t�=gsᔵ��������������ꂍ�9K���ϝ����ٳ�ϟ�wp���G@�R=~����o���{�fgg���322��5�'\�F��ɦ���`�auqq�������
kpġ�����������AyV���ӯ}��k�h{�5��{%g��ሠ�ERlL��Y�@*����*ǔD�X��S�R����@<����W4�5MitdP�!�ٖ�W����\��D��Uݭ5��e݃����=��5F���=�~��u���o���o�s������:~���j{m�Ό��;+�߼x�������[#���G�/�䏩�;k�R��H�"t%b�-���b(��U��D̫��[���fM�+%h�  ��IDAT����H`V3'0���K�����r_��� �3�M��4|c�)�R�ʨJd�q3c$q�!��1Y�1%�Ȋ���aY��n��8/l�(U�ʴ�� �@Ҿ+j��鶹z^Ǯ��@�u`< �J�[R�����������÷cz���]���yY���Rl�6@����a��3
���Fa~�4GÊ*!��	�`*K �!�BF��*�G��c�>qB���(p��<�Ğb�L�G��#[�#C,�i��SS5M��;!�7=�*�%�qD'A-$10*'&�6?��:��6D�al�h�1ʇ:��u�.��S)4� b�V���k��
���������č�͎�Lf΍.ϔ�͗,��L�$c�T�������]��!�K��m�T6�5dV��f&$FIYA|j��� $'��SȈ�I��2��l�{�Eu����15����y�l&����`�T�m�(3��'U�o�']K�=̍��:����O��>�.>���zb����;��緷�~����m}p��پI���+�V�_�SX8<���!����w�G�mG+�G�3Gc�G�5(��}v�R�{|�&��x�I}�M�G�����}6��k�5���{��1Cv�̑]�I��$�	�L�n2=��U��:�i��Cv�Bs���Av��|"��(���@��2�W"��䟇0~F��� ���PH�Q ��Lȯ"X��d�)��(�Ob�_E�����4���i8�(�'��"�O�B2�|�(�*9��Ā��$��ߏ�<aߐQ��(��&���5MrC�5b�#x�5D@�$7���HE���:J�t��<u&M������
���5�	�1}��0-tj��o��*�q�X�2� ��hlC�_]�ωhS��5��H BS�L}d���hhj@�,k��>�b�ftp����A�l�*0T ��bq_�t�< �V�>Q�Q����q��ho@M<�!ߒN�K��&ak����+1	~��q��$�����@�c�+�^��n�6��pAh-�Du:]�FS�P�&���5YQ��'o�Oq�_Y�&����Y].O�c"��e���!S^�vӺ���)�v����#HpM��EO�50� ���0�����Ԉ��e�8è��Qo5�h���}�l��Ԙ�jB��["�Z�M����5)�cj`��!Mt��b��r��n��i��m�[5ޥyYL���gR��7P���\ۘYӏ꫆u%�Ʋ����f��5O�j��ƴ����mLM��z�90��I��C�h�rB����-f��2��@Ss\����jď��05�SsB�<C0X(������,]2UOn�!4F�{��V���������?t��Ǐ�~���go�䭣<�ãßo��lf��v����9w��^b27y�Y�����A�A��@�~g/������a�k�ҫQ��pវ�ƃ������	�GI$����inҗ�ig����YF����oE�ޓ��
n��9�I�˔���5�9<z��H�\����}W)�+d/ЮS1k$�E?�O�Y/�i�1g�!{���5`��Ɲl���.v��Bi��ꭟ�VZ���������3
g�ԀN��ydѓ����F�g��٫	j�����Fr�p��<�U%@�
�mB7��]!�0ke�oK�7�D�y�`�6SL�5ภ9Nk�$k�����oC�&�T*'�
�Ya�-�s}ʝK+���[������^��hɈ1w�#�G��cH��J��I��M��N�HJN���&��;��3�h�0�ww���%-���ƀƆ���BiA�$;U�/���8�<��b�X4?ŋEv�R܅4!×E'�B<��ϗ�T�t-$�_�1\���s=��V`�$��㪴�������������\f�f��]
T�s�gy���5�f_�qK�uW�q���I�\&�)�C��dj��4�.C�Cn\�4���)������lɘ� &I�݂��`�J}�i��0O���"�t"�K���@6��)\�+�J���ݾ�4B�L1�#s+��1�+t���&ޔ�#�XK��k?���qSӜɁ�fr��y!�S�5���d�M��@�/h��L�ԫT�))
͹��nW]�BO��l��U�Ko��{s����GW�߼>�����}��E���ߺ6�`����pI�9�4�Udh�k-�4g��2���q_cV3'8�i���ߥ�Їs9�Bw縝9N[��`BM�g�?ޘ�)��%��r���������W�ϼq�ԩnj�,l-Sc�S~�����M�'>35�e��3hgG(k<�n(��+
������	Sc���<w���9��g�,O{:Z754��Լ��������A~p	}a0��<oj*����@`dM�)��	SC?^fj�be���H�1SC���r���\O>΁�n��p����g;+7Gk���4��y8}����ϝ=}�ԩӧ�V����&�
�������������t2�laa"�&�H� ��������
��Q�vt^hj��>��g���3��v����[���x��m'!����,�n�715�)-xV��н�����dZS)ߖ/R�	[s�=uQ�F����zr���~�マ+K���Rmu|nKJq��"���)�޶�����9�����,=�2}w{�����F��`�|gΈ2��FW<!e��� }��]��T8P0R2�>P�]!��� �EC�м���ј5�qG9nj����,RC�>ߔNjΠBSS�GLM�<*>5:�*�TV�P9*�������-+R�z�z+@�#�!����{b��P�'��:%�W�.�CA�=@�� ��Jlύ���q]��ע􇡊���uY㪴iY�Xg��0�����N~�Q��fD�D	xv�)��!+P@"$�h�w05�2/��y��	�Ʉ\�'O��E�d1bq�T�XU �+l������F:��;�}@خ�T���Έ�����ȱ����ę���Ѥ�ᴩ�����¥��ͥ����ݵ�͋K�%sC��9���EN�*�[��k�P5e)�J4�E�5�UřY)A�P>=ZĈ����T
��/35�y\t6�%��\�r.�[����1\��J���F<̍~��8'��ʼ/�J���9���;cgq�^�޿�'��>{�ϻK�U���}��-g�|�o�����i��=��W�9G#�G�Gs�G��?�g�*.��?
���{�L���żM�|(��f.3��)��$�5��2����5�*z�b�	e�5K$�E��<�~o���]�٭����C��U��m��#.�>�=>�}>�C!�c1�!��Bi?�3~΄�0�I$��Q�Ϣ����� ?�~��,F�i� ��ŉ�Gr!D!��?K�|��ej���!%|'}/V�(�{ED���Yg��2}�^SD�ː�S��Ӏ��� �O@�P�$t�Mq뤹�np�V��j0� �2�O�����BS�� Mᯈ�)cMc65��t4�5ͱ�N�8Y�N�(	'j��8���t�z�����R�Hu�D}8`�N�	����*���d=��B�2�ҒLh������'�7�Z3(�)@C*�>_���N�j���-/�9ο) }EA�LlKă�*�Є��� �l&�A��dД��dbK"<rc�"S�_���' �3e0�9��|��Fo���Lt4�,& �<M[��~:���ojj�=�����SS-魖���`ɧ�:�!�[�
ԛMM�`K�3S�0�MWg�cj�T�#��am޸�t�X>f�7֎u6�[�=O�	;s����\]�^՝05�}��9}Y��@Y�Й�_0�~4��@�u�\�<�m�_�٪� �:��'xnu�R��4��e�,��{z�3�t�>���+���e15�E�2\&,���ن4�&���ł���pLoq�%c��y���?y�����<���~���g����/����?\Y���܏�nfoF�g8�9cG&��#]�S��%&v�G�Qwd̽@����܌	�#�%�!:� 0�fSƂlp��WBE7#dw#o�����;l�&�c���M~��5�2�g��@t_��7�~�Kt�w�& v���(��d���nH5n4R�i��r���%��9Θ#�n���M�q4��4V���֧T�g�g���:#����|�Y��a����`���QCvRS���%�I�uT�g���x�J=�d�� /U��*�W��>��B%� ���Q���Լ��F��Ah��C�b���!�\M*%�C��񢆬�ɾ��	������������H��P��X�X{�!�_�է��5d�3z:S���iCC���i#�I#CqC��=�ppQ���i�r�.��U���T/�++��M��cC�r� ���4?6՛G��<DT71�]LG��"^(`(d"G�P�X�1��>��_M�>���s]�u#�x5�p9@w ���5"����!���W�Qڭ ���mU���a�w�z�K{�����ר���L�>45t�6�i�\�L�Y�W�+g	e��E�ؼAl�]�Z���#H�z�8�Far($!����D���^���G��j�L�;�E���,
��303e�%#a5��
�3YSO2��F�(�i��-�P�
����^�ם05���T�-�iK���\�+�J��ܖ<��L��9�Lo�\.���~�j�흎��O��}s�`���އ�=�6t7�4W۶&j��{��TŲ�L�"�*
�z% �00p慜�4fS:`��r�}��i�oJ�縩Q������Tvi,;AL�{��]���;�C�^_8s�e15vH@�������𽼼��L���e��ߘ�S���Ԡ���� 0%��� ���1�{k���Vcq��չS��<.�<졩 �@o��3��,�w25P�c��y��[�k���z��鸬yfp� MMճP�,<Oe,�4w��T�j?�FQrC1</>��>�j�����mλ�Ѧhhjm,���8{������ӯ���k���ӧO����ËL&������'O��������fRR���閖�(
J,��9�Vpp]]]�~�����̹�Ϝ}�ԙ��@4���?����/'�������mJJ����#�e��8��~����y���Y^pxbCY�MC
�9�������y��8lg���hōU�u��K��.�|pk�����K�kg�����g��v>�3��ŏ�.�yy��fϝ��G#w��//j��u�C�1��`m�*]�Ԕۋ��>�O	/�;�x}�A=�FS�'hj`�����8���f�s|�?359�,BC�1�ܒIkHcV'����Y���yTRjtnuT�>��OZ=*���/�W��k2�f�j�ږ)������� ���D �\�81^�w��!Q�����+�]W���#�����m��M���+A�+m+��IF�0����c��Y*FT)V�e�|�+�eJ��)!F}���I���I��4I��b��L�!c$AdY��eʹ��PQQ��2?��:�C�6ҙ9ݟ13�:�?ޛ0ї29�6=�1=�5=�35�ԙ����幂�Œ���������噂���ƭe������%����B��X�b��`��p��`�hw�p�bl��CW�Q4+[*+��"�#E�!+�KJaz�Q���)�s���
�Kɦ��L��9-��v��������1�����f�������KJ{hԨ׾_�&_6������G��zty����q��y�{��;��v����D��"�+�������ʣ���FG�62�##&��@�.�����m�}�w��H��Dr_��.\�(n+�%� &^����D���4�v��f��j��j��zk�Bp�$���<i�W��W��(���x��E�w����?�}��2���H6������ ?��' �$^���GQ�bD�I>I�}��YR ��p.��޻�����ĉ?N�}��n��q����{7�{UB]g�Γ�3�8�e��e�ױ�˾��������؇w�Żv\�I�.2���v<����������!�|��i��"5�x �/���M1��h�h^>�T��5P�*@�
��qM���p�!�֝��+���IF�C&"f���MQ Йm�-�	(�.r��l�*��H!5�c��0��DlkI���$C��I��4b}:�!�Д�ߚ����c|�b}A_�F2dӍ�L�!�i�g9]�<Hgl��1��]]�EUgR��$E�j$Qz*�)�֜A�_M�����s9��45��L�׼��(3�mi��T�"���f
��A���qMc65E��^�y�bS�cj�jS3Ԙy��1�h
lj�n�V�&��㚴�iP�Mͨ�x��l��|��f��8��2ک5���15�W'WF����}�Tg�lo�|o���\��F�|{���UL�X��2� �k��e�1������sܶ�5��y��y!p���@T࿈���O�sB�<C8P,�/���{s��Y��t�1�bH�6�}����C���'���zk�����g��zr����>{���{����/W6�ic�7'?Ҷ�&,J�KB��P���,3i�$�Q�H�]����	["�~ �0�w;&�F��z��J��r��0\M�n+��.a,(9�Eq=4���䷀�Y�z-�|���=��G��S֙������_b��S| ׅ�+<�.醐vOʾ+a]a�ɘK�E/ԤR�i��z��b��¨�Մ�-��>�i��r�ޢ��|��9�iԖo(�ހ���N��r'��V���F�e�i�X{=�IGv�P]�4'�I�rTp�|'�i\bWe��2�[�F4�*�O��OD�����Mᄋ1sӜ$�����A��-1Ė��ʚ�8J]�<_(�Hp����`eM�Ho��J��������J�\g�dG�xG�H{�!��=��=�א�ӑ�ߟ18�5<�12�2:�04����7�����!�h�k�!m�������ڲ�����8Q\�P.�D��O���8�����dz1��.*J��r�T"�Dg�&eg�wd�&2:�R�����t_��n�ھ�ݑ����C��T�[w Ӏ��@�%pS���ԩ'Y��9������끰�!��S��=�����}�r��إ�lS6I5���yl�4�x
_2�-'�����Z��"?i6�����a�b
�Ǧ�t���ac��>�"�X�W��\�g=�:��\� �c0+�20%Cj��L��UǓ*�s�n0?��Ƭi�yBU�H[ �s������uC�HW�G4M���BД��ł�lVS�>�h.��z
vf.�(ol�����t�\�^[Q]_V�Z����n-�v�j���am9��t�:��t��L� ��慜�4�8���8��&$Z���S$��w �eж��Kb8�\͓����d�lq���Y��H���ԘM�ۃi<45`b��4����l���x�'�"�0I0�C��̲�~B99Cڗa65���/�����Ͽ�fw��n'ģC�^�L�(��w����i��8R��� :%r�2S"aHy$e��oL�Y� ��yBe�$
�Ԑ�b��1�� ����a�f�dv����v�t��x8ۢ��P��.�v��O�:��o��ܹs�@�{x��P__�޽��z�������ͨ�(hj,,,��������G��d����xooo85��L8
N�5¹So\8����YogK����Bu�b8�s\�y0}�w35e~���-x2͚Fa*�Nihj�!�֜�h�b+s��<�\��;kB�sfj�-���P=�3�s�;�ߟ���<�ye��n�ݝ��μ}}��v��U��K�`�ʊnm�zB�>Җ���Q�/�@Mc(A�:L�D������e ��D%"��A�)K�f�r����{�;�45y��bC�)�Қ���M�%rce�q�)����庠�ni���aVҸ$kZh�R\
Vn�� ��]@�	$�ư�qb8���E��Dv�:�b:��{1�{��ݴ��Ԯ����h�V�b#�m#Ju)��"�f�Y:�(�bd�Ey���D	8v��g�8B.KƧ	i�����D��|�|o��_(g�������������xmk�PW��X��L��B��|奥�����Z��Z��r�����������Œ������͋U+Vg�/NU^��[�Ul]��.o�״�K�K�Ms��s�ͳ���Ѯ�>C�@�zl��ۨ�4tt��Iq	2Q���������in�45Y�:
I*�SS�F�2����:�s٦o�$X�&�>k�~�$a'�w39佂�O�s�j����aIA�'���Y�&��������~y�������̈́�.;�q{�+�>�c����Oc#�ʊ������������裸ģ������ O|���&��E����<W�.��VH�u��*�k����DBl���y���a
g;������fc��o�Nv�$� �H{T��l�[�-��]�����»A�B��?��~͇|#�2V�A����1��%'�>M|��Q��8�pΛr6�q�̣0�5	�@@��v�M6f��1�C
<�y�u{�uy�=�: ���N���Kޥ��b$�vR�]t�N�����!�m���eH�'M0Vb"��ca(�.��Ȣ�h���:���7��9&hh�4:@��ЦR��$M
p\ٴ��=�\�঎,zO>g�X4\8Z:�	5�@S�c�a��=�,���d��BQ��d�hN�+���Lj�I�4�� P�4d ��$l[�h��4��BS�M'w�z�����۟�@GlB�&�5O}M&Y��R�s�U��{#x'�0�>nj �,�}��iK���������U&�� �b��[G�ทy����|瘚�Z450���	Gcf�!h�)x�)tȴ�	��e�.cB�9��4��Qmވ.�DF�C�m�C����9X_�@S3�]9�WM�"�?�b�7�f�+����5��2��!S�`��	N3'��x�<�@��xRa�|9����y^S�2��`������O�3X&*=ω�o(K����V�7�0&�t����hYĶ����ޟ�Y��;W�>�w�უO��[�~xy�����]Y�������پ�E��fa�J�t�I��RW��U:~��@�'z]����	���`ލH�5W#�P���5��0�V oM�\�R.2��4��@�_$�/������ˢ���ڡ����o��{�>���&;�8XpOʾ'b>�q�	=	���w���y7�	G�q+���Q;�	͔�=`��v��j��B�-��Fo}Fc�h���J�7�֧��5���T�JD��n���!�;豎�'=�EOs�1\4L'�I�qT�"g��E)qU�Ъo�ҡ�� �rV=4}}��K�Z��(�"�h�PZcI��D�WHljKAOQ�њ�(���
�H����GQksdFE��X���axA�Sj��)Cø�r��d@Wԧ+�m��3f�te�gf���'���D�u&��NdOG�A�U�(Z��u�򒠢�hAL +�˔�8���3|�N|����ey�9!lt �IJu
�{ұ\�?�D�CBRJ�k�r�i�Iƽ�N�+И���n�z+P���G�k4{ՖDu)�}?��V����j~Zw��E[?���(����끸瑨�>��Ms��:�+��}z�.�i�R�A�^�b
'�&��� b�0!E�^�-���a��8��H�2<!�)a���89�7F�'�L�z�H�3Ğ�"ϧ�\�K��|20%�^8+�15�I��DbeJMMU�&		�o0��dq[�y�\�2O�.�lN�N���������#��dj���BC��-��J�M9�,fU:�,�\�Bi��w�GkR�F�7'�.MV��U,.�V�M�n�V�V�W,u��E���m0�4}a�R�2��2�iC/��4���i3%~!��H"��8�-�_ˎ�h�|�������Y�s�O��cjN�0�3|6��b�̦�@ ��?��w��@����'����T��8��6 [3`��@�?}ɧ��+�g_E۞%��
p�P�W�=��t��_kj�}�y�� M83Ͳ愲1����eT���i\M(�� ��T���(��T�O$�]Lr������\��#U�\<Q>hG_7'���������c|<�юv.\8�<h---���=i4ZEEŭ[��y�hj���677CCC�X,�B9w��������B�����d___pp����M?���1�6-}2�Ը؞�v�d�؋��at��k"�*p3��G���	�2SS"G��gRG �	�OchjL)�a�sDPf2�lU.WU��FʔIFձ��y#�[�%�3�[S5��WVU��57/�t�{k������@�ww������.���3��cz»�C��R��Dl(!z���/D.�]%��b����o/�5�P,4��;�$�u�q�{����W�qSӖ�ḩ��Ss�M9ԖFK�.�[�(̏��'D$�g%�E�kC*:e5��ƙ���ֵ �F��R�v��
R_
�n�C�;���`�vH�$���ܰޱa܉6�Fu�Dv�ڷ� ���X�v�z#B�����
S,��y�ܢNn�N���Vr�J��"7��1Y<!�#�1��	廚D�H}Se�h��@� ߄pBh ����Jq�)���	�)iű��Iꦼ�����������妽����ʵ����ˍ�+�+K�K����.�T�ϗ.O�.MU�N׮�խ�ԯ�hV�׻�\�~��ڥ��5��as�}m�}u�}eL�<��j��N����*��Z����Ӡl��J�I�
Y\l&�#��N��2h�o75�2�{!˥�f_�tl`��0��(�J��\(��wʓ�$�?ʎ{���Uc��-�?�P�e��]ȴ9?*{Ү:�u�����~�.�|�Dic3��s���rE_���������md�QV�Qa�QV�Qr�Qh�QX�QD�Qt�QT��¾fr����gS��R��7�~[8�*�e���D#��q��\��ɮs�i��$�v��f�a�Dr]��o0<����dzm��6ɨm*j��~��sS��@zB{3��N$��(.�h�����bD�ǋ�K��� x7^�V��Q�Q�Ap/�q[F�)&]���6���B�Y��,�<�1.����N��6F;O{D�`\����[e65F*�������a:����.�_k25�P�:�
ǁQ��QF�T�xd�S^O<�2	D��Y]�:m*�i�`�g��K#��5�<5�c65�%��2�Pe�hM�Xm v&����@y@o���@ОÁ�F�Jզ��)T��5' -�$EU�AoN&`}��T��4rS*�%�2��������t�>��Q�6r��tM>CWȂh��<�*�fF�C=N{	���1#t�X�645f:�M��D��P��ZRȭ���h�Y u6�yM�Ï{������;���!�r|�j6i�`$��E>�
+�GU	���	m��&�5H@M�����>�filiH=��m/��﯀��b�b�R�7�f�+k�+��S3����S3X+~���}�qS�C���1/��M�q�r�3h�zSc��t��*�Y͜�D��3��ա����eҡB^.�7�ғJ�I&��t�8�ۑ�M�:�����o���}��э?>��O�>�_�pw�ח|}���V���ƿ�,���p;/kI,��PH�M&e����3��\$z�1q�ꁔu�=��	.˅�#DOMM�x_.��w�;��� �A��r�h_�=s��C���w���g�6��m&~���r�g�؄+\�m	�0�;�ⷂO��	��)b_�`7��ݜ'�lFl/��[�;X� F`L͔�=ha�^�3]��ڭ��NCS��>��9��?�Tzr:�t���A[�<�՞6j/[����؁s2��;H�W��D�Y(�vQ�\�W��tS��C}��9�i���7�Ț�*���(��2��Ko���ő��H�OS\c�5��#k�i�x�&����5������ ��@��(bMqh�>�g��0ܨS��5�c��!Mi������=��3��?gd8r<wz"cr4e|(q�?it a�/��3�]+W+CZ[��4VB(3B@�1�\<��G�z3Hn,�눬#��#8�\9�t�9�P܂)�2*�C!Q�\nP|dnkz�x��b�~#�}'�po؏��D�6C�끚� �.��	����)\�������z�w��~[t�g���=��<��>�<�wޡk���>Ky�l٥7l�k׈K����)|�$�i�y��d�X��8ݛ���Œ9a���JX� 9�����H���T)�t!����H��97�3/�F.T�r��<50��&�\O��t�p�LLM\���j�Ep.�2T���F���L��x�245�
���VӚ�k���d2�2��\Ei��F���Uk*�%Re�XS,5TwW�;ʃ{�����]Ł�lA[
�5�����@Y��a�5/:���ӎ�����djN
)30��i��t��-.��'�!4O�C٢���_8{����Ø(k̫�0�޳X,��	��H~fj��'" #�F����\\m�l-�l,,������ ̲����(��<��?Z�����i���d{İ��5��x/X��)ǖ����Ք�j?AYSi�l��0k��p4� ��S�b��L�&�^�L��E�݅'�����e��l����m25~��X/�M�c"�F�����]�C�5��;8����tzaa�k��}�]�Wx������x�믿�����������������E�
x�G{��A�����S��8�ګg_����ogK������r�㠑��B�T��Ӓ[|g/650I|����1U�nN��s����@�M0��ښ�l�b�r���\�����Κ@C���>eLkO���],Z)ݘ����vg���^ǵu��]��+=���*���Չa�� Ce��<��L��+�J�}!�pG�����nw)�v#!6P����������c̀� �o�7�;|�35��FC�!�ҜKk��/�)�[�$(��f%Fddf��Ŕ���;je�Ӂ��@�f�f+L�nؗw��; �q;�s'�{�g �މ�zJT�nt�^\�~|�Ab�a\�^l�n�a;B��\�+V"�뱺��bp����W\b�iC��C�T��2vp:CEcIYl��˓p�<z��-��MLMT�_H��D��L�f�*K�[�sU�⾎����������չ��������������eťu��V��N��n�����%��M���pM{yCu���vﭝ�[;����o� Fnn]]�;X��[��2��8�=?��г:۵8ٷ8;��Ң׵�5:}{kK]^^iB|a�<[����Y���Y �SS#�.纕1��i�5t�z�m�B��}�^��qqܣ���91w�"�Ǽ]��aSᣪ��%�|z�Ź��^UP�_������^��㵝Oz�G��vg�O�O�}g�[h�wq�_�GQqG�)G��G��G�IG���.
��8�(8�(4�_��?狾�s>2��R�ר�{$�m
R�i��B�@��P�.�Ss��
X��/��.RP�D�Y��S_������'�,3=ֹ>k����}��~＂wY#�.Q=v�>W��b�-)����l��0�c9�f8�I���(�Q�~�N0�f ���� ��* ׽~;t�M��*���  L�'�]{�m:\-:�V0���io�q�����C��&����#�Ew��x����e�� �1�ª��U���P�2���Ux���@M��!�b�	$U��4&G�J��S�'�1khj��g��i�d2i�T}���hj`&�����
�����@y ��Lf�"�Y 0��۟9UM�JhRi��#[�H��T�2�֘H �'��P֤�Z����A�.��[�q��Τ�r�H�LC_�n/�J���-`j��l
 ڙ���dj��R���7 E�.���Ɛ�t��"V�9LR�H�����2�
j�m���������;��@Gs<�f�T�鸠9�Pc�`s�iLK�F�q���QUҔ>sR�5��2��1]����%��M�7���]�8��W�ʡ�Y�+����@�R�SY�ؓy�;��f�	�����' ��\�4X+>.k��ϻxڝp4f^Ssܶ�ڿ���������A(WV��S��gfS3����4�1�����i]ҩ�����_lN��_l������}qu��+���^�����~|��Õ�,O|�W���:��H��/`��BŬ1q�l�&��-��Ș�A��P�a8"k@{!��m��;A���e��FD���໑���nI��n�DWE�=6������2���u��r�K�#fBM�N »�'b�m:q��m��v��z����չq;�)G�I$�fҔ�Ƽ j��z��|��)ùWScsFms����������B鈤V�,��Vj/[�����wB>�F�k'�Iw�`�lt;�M�G�h����un�@wm��&�K-7�f;����]�E�:
���C�1$u�/DCUŲ �8�"��D� _q�m1�m1H�*x@},�=�����0�#�U���`�d�[�[�'knIm�*�j[Z�z��:������.mv_w��P��D��l���s��Y��#��ؾ��vm�J���,,��E��"R / �*ݗA�b������Lq�3�Q�h�{�U�v�;�S\C�n!t��Ec3yIxPR��@��2������H�m'�㵗bT���5�b=@��E=�����,Z��n�'�{_W�|]��ô�O"F�
�{��8x�I��;�L�z�Cq�R\f��R�6�U+Ĳ���YB��x�T4M(�$�PR��BOA�/������ؼ 1O$c3�9D9����%���R�T�k��3[�m�4`���e65pbV�@@4M�&�P����@S����O�ј�yj �\�:�@Gc�4�M1W]�-bj�� ]�X]*PE��|nC.�.�S��m))J�U���dRYP�H�H$�#5��I��dj�4&�Z����Զ$�"��������FiZ*e�4��Ƥi�r*$V�y��9.kQ�#��D	1��%ģ�h;��y�s��x��/��yYFa???��4���thj�D"�@�I�O�O6�����uwEASc}�z���̑5`��x��+�`���\�N��6*�����}ט0�v��i��)S~r�Y� �%�TO�Nu,Ѭf`p��NP��py,�4��SSO�N`凑�+��oG��%�8a�\|ܝ=ݜ=\��x�`}<HX_	Ϡ	x����٧��ڂg��֞F������=��������zll,�L�b�������?`3  @*��x<����quu5��#�050O͹S�O�����
Μ7^�8(����-Y~�At�h�g�=Y��
f���Ԝ�\��M$7�
۷=��i@ې@/:8ޚ�h�dBSS�Jl��nK�&�P�Ij+di*����δ�������#�k�eK�ES=���5�KW�Z��Ǌu	퍡�� R�I�+#��T�Q&K�`�v�;
Y��Bvg�o������#�c65fG_�/15��"z}�1�
�/e.���$aQ�,79*;;;��6�\R�X��<�^�n��oGt�F��G�D�F���c���_��7z%v�r��a��a��^��. vh?i�r���̩��cW�F�$�Gwn��V�4K��m_M�-�7��������%��YB�H�Õ�1��\�H��	9L)�!��V�&D����fgE�h��:���5��m����fyN�:׺<Ӳ2Ӳ��viI�������n�w�:vw�����{�\n���qk���a�݃�k��{KڝE�΂zcZ�9�~iƸ5׽=߽=۵5ӽ5���ki��U���j:UU����I��mk���kkhP��5�f�V&������7\ �Nu�b��2��bj*x�U|��k۹���@��Þ��xEM��_���6�q~����Q�r��U$�f��_�%.���*y�T�k���7�{~qu��{�rc���JP���۬�㶕�uk��(���̓�I�'Q�q�GAQG���[���#i�d���~-�.�|(`�ã>��n���T�M��
	�LFCG0�~�Tp���':��f	N3D�	��4�y��v��9���e�����BA��=�9���=��H��n��C���d�+�e1�������l�]���c��Z��.S=�nS8�$5����fmDYݬ;�mM����~.]��.�G�����Cr�&��ҧn�G�o0�0B�
�w!�F�Qa�!��0�24�� ��qH(��Ҷ9�F	6M,'�h�;���1�ёE���Y�N&@qc�6���fwǘ�5W���+����Z��hr4�
45�d�2��H��%<��ݚLmﮉ$@S�1�Ҕ��.@rǤQ���ߎ)n��nJ��e���b���Zm!G��R�19t�2��`DS�hY ]1K_�A�M1���c!5�r̚�;]yBc��e���f)3�P�hM��59��5�q#�2�bS�cj�15 hj^V�j�g�&|DM͘:qJ�>���f"�	�Ɂ��%��󘚇�M�\o��@�qS�܏�Vs�;�bw��;�f�%�;����׊�U|���&h_�H����;�M�|1C5b�`�h�J��`��~_������)C"h�z��"�f����t�=�܁B�`{��5^Ȟ,`e���iݩt}�5���g�֦<Q}�6����O��~yk���>����͕O�.��5���ɯק~�4����i�?JI��x��<.R|ט�6a��_a`�>�i��`��Y#�7�2���%��ʐ������Jo��ץ��R�m	���}�K�.�ݖ0��JX78�[<�c�M	牔��������ø�Ǭ�:M�\��0`y0�`5�,[����f��v����NV}��^מ�~��Y���	��Y��y���e��ޓ�����ۮ�ϱ��وw6�Mc��t<�4������tbw��M's���B<�a^�0o��W)G�Ҙ5��1�mAK��H M,YKy����!k�j@<]OU�S�	$�2����#	�J{]Ko�����[S�E�� ��hRI���<R�^��Y��Y[e�.�T�*
����ւ���ѡ������ڵ����%+�EK��C=�#}�}�h�*R��P������BXL�!ıy>�W���2<��`�����DŲ�b���K$�1��EC��]��(!3P��IC�"�$������-�)ʋ)��d�v�v+Fy)\�غ�SR_
Po��F�dϽ���a����SoE?�{�{?t�|�-��;��{,�!�u�����!U.K�I%3��Z�4�h��?F�飦�bC<x�~�(2?�����<N�$g�Gq��x�Z�$B�HP�b���+�`( ?�;?��,��V��Ț�xSr�DRM�:ik)��Ks:K��3Ӗ�}���9t4hjY���])�P!���D�Ak�%�ݘì�d�e���-yܶ��D�,��s<M�P��W0�OmK�����U��Q�1L��u��Y4hm���|@���9���������L\��wפRd�0����&�٢m�ۜ=����w����g-�<���������ΎN(WOw_o?_2��b0�t�F�(HL噩�K�H8< ��q O���y��Nv��Ԙcg̚���`65�&�iq�ܙ��8��+o|�.����q($�&15�q��151L��@^fj^\�[�/����� ���Źu	�w25��hH
�H���&�RϨM`�ǲbx^l_k��%�˙���Fc���]<�M��|�Q��_K�c�<�]���A��<IV.X�h���̃����y�у���޻��������
�������~ 8XR�T$��l"�������
��^bj�!�:��膦����������/{�7��,�'pDb�>I�d�{
j����1�����x�8�A :	Ėj[&�B�i��kDW�7�K����2A[CQ�j�i��M9Ծ��eh���F�q�Cy�&K�F���b�B_�\OƘ>�j��/p$�x��DM�)FF�]&�,�K��<�.����A߈D��h�C����^慦Llڊ�M�Ԗ<*������NC�2EX�(�M�����(��/o���ª���0�B�n5�c=�{+�o7i`?ip�2��6|�9v%{⚉��c�3G��2F�҆v Y�{�WJgnV.ܭ�x�z�n���ܡ�Ԯ�D�r�a%͸����o���,�(�%����aI�����h>O&�$l��M���r�'�I@8njЈ����8O�)I�l����@��@Ll$-!I�]S�(��U�u6�'�#{���C��;+������B��r�ކq{�}����j~F5;��ʹ�Oh6:���>Ms�E=�lmc����SQޣ��4�[Ǎ���l�n�W5f��n-UՖ��*T�e�ue�����uuuUe��ʊʶ�����ԔryP�����K�y��S�MC�1 �l�S���|�K!U�FLM1ù��n�x6K�ZĞ-|Tݶ
{���\����$�g����&>̊��{�"	�/}�'�ɋ,�
_Pmk'����b���!��n�����ћ��ybtM0�Zspڳ��b�����3�h\D���@�1EG��#aБ �O<�8���#�D��������P@�K�N����7���8�%GT6�X���,�q��@rY �.PQ�	��4�y������h��i&z���"�.R=��^�l�->nGHؗ�R
�PF�@36I{b��������{B���p�����a�v��[4���
�}
�<��8��8��2��<�����0����d�1z:"15~�n�.�G'��"LAwPP����+����Ԯ`BGN�
�(�1m!�maXhj����4�8"���$"�Ƽ�	�2�4]:ㅚF�F7o�W?�dbj��9aj�4��#�v��eu�q:�E��B�1� ��	�r��,�:��H�@Y�D��iM!Z�I ��JiK�"�ya��ԌEE�E���{ xo�(B��S���1����i͠�+"8W�"�3%\M>C[���қ���Z�[���aAM��_y|d%W���s9�,�*���d�r؆|�	�X7a,�tq�T���w75ՒASM��ZY_��?45MOM͈i��3S�<ݞ5���f�M͸�`���%U�����*������� _��ӟ}��W���:ѽЯ7Ԍ�K':Jg{�.�\,X�_̅�f�T�i�#}֘����I](`Z����M͉͉V�SZd-�0X�l�� �ơ�8>� ��f�$h`���gV'�qhd���� ����������w���/���p�"J��j�H fSo5{��:=e��RNW	�����1e��yes�j�+9���Ϩ����Rދ���rQܡb��"��\Fw�=��MB4�6�b�dtf��~�5�������&:>ߝ�ŭ����:�����^��ŉt~�Q|�j���u7T�&���|'�^�t�%6n��?K���x��|A�O�$�mK�b:�,(�A��0ᖌ	69���N
�VL�[�O�%�B�w%�;b�>����f(��0�-!���@�~ f=�	9����D�%��Ź�S���z�>c���`1�h	t���ڎ�9 �������Ͻ�;����5��
[��)���)Z��:�E��M��C��� ��CDM;�I�p�3��9��Q��੓�i�u!^�0]��V�	�Q�{��}Z�~���9s0\>�qH� } :`S�b`�s��(�c���� ��� �n�t�.����2��)��fq3?�[�ZS�ܬ(�ה���6�(���kK���Ӄ�'k/NԮ�6n]��X(��߾�1hL��f��"�$9�����D�xp8(��#@�*��<�,t8�9��Kw��;�1��l3���v�c�$���X��,�h.>JH�
G���I���Yu=�k���ƃh�N�j/J9D�%W����m�R�fD�դ�Y��̾5z/���p(m�h��u;��._w�޺`��Q���uԺM^��n�^>G+���2���Y]�T>�V�����tA�@ �3�<|�3��J`�$q]S��iBt��-M�N9gIP�γ)1�I����40=�K ���R�fm�`�f"_#+�9�}E&�2@r������o��D�<�92G*�ky Mf��3�x 0a�M��<��Υ-�
�Q`��4$BX�A��wJ�L��Z]C�C��"��UY�./ �c�i�<�Φ�/}� �T���B�4�	A\l5��2x+�)A�0�����x�;Y�n�ƫV�h�g�-��X^��>����,����`g����v��������c)$2���9�:��LI��a�&�@7�����
����dg�`c��h�;� ���il-����:�ځ?�������+��μ��h;K:�#����d{�s�b�.���t�g9$���%��H�=M���sM� �
�`6���)��.}�'ha���c�j�H0�l�@!�T̲�� �� ��*�g�bHȣE⪣�1��8j]<�PNNc�(���ۑ��z�|=P�N�. 7g��zz�pX&��O(�����8���p8�SӶ/mݹu����~���f���/.���1�Wg+K_op�����,�N�hj�����
�XX�ca}�3g�-�z�ԫ�x���ٞ���,��FJv�d��s���8i|7 x�)�U����|���i�yA��`�b�WY����OWA�x 4?W�!͔� �d�'���1�൩ʥ����&���_���2U9i�SFM�c&5�M�`��U#����b.���e/L$:J�傮
aw������ �����(��e| ��|��v��8�	��#�^�Tu>�-ג�k˦�d�jҘ����8NVjpnnb~iaveUJe]|Usr�>U9�:��SO&�g�;/���n�m5�]o���<s�q�J��~��Vi�zQ�J��b�j
Pѹ\۷� �@����r�R�n.G1��<���,3,Vu��6쩜�k�kɪ�M/�'�ĥW�$DD$����A|n ��$D�I��� Z����z&�|Re�iR���A��#dB`�y�wV�_��'Y��$�L����qiQ��4IAAD~Ilq}z�����������������Pfh.R�f7��V��C�Ӣ�D�$f��t�,�r����Ť�E��O�3��?��a������N�4/�������������K�%��4&�æ��L�D��]�X��\��R�P(��s��t�t�{6�-��*���S��΀B�S�1��T�v)���|tU%DW��*D�r�k9Ϲ��XA�/�[�����ە�Te��w/9�J|��̈+�~�\�YE�^xP��W����S��������{Gׯ]9���{R(�Y��z�{�n�������1�I�x�?Q8G\)bj�#*���;����`�������;!�<�X����w�',�:�*�g��I�ջ)�y��	���0OA�Q��4���"��"��"�k��5���1��>�|�5~SJZ^iMD\S6$�M)mKB�$�n�|�&���Ư3�+T�e��"�c��m��H�����rts�s��q��C���9�y:�x9�x�����0��� Σ�覧�(��*��Q�9J����ˉ�~����>�Ǫ#��nmAKT����X�&�&��$�!���"4�\3�T�.�Л����M�cȤud�fGә�����p]�,��/�6�	�۞E3�_�!�ٞ���еYTM&E�NR�)��D|k�-� ��T�*�B����t"@�ARf��\��>�w*�~eN��w� }�y���|Ĝx ���|Vg!����,�u�qL��i�b���ͦ��=�<e~|Ё�愣1�Y��,e?����(fKX�82t1�נ ��y��;�"��y��g ��bj����1u�:uD�>�������]�XG�hG٘��~3���OC�a�zР����N�p7�_S�ɇ�|��_|��������?x�:ѽ8�<nj���穁�f�3sޘcj����1��-M�I���f�^2� ��#�"�P�`��Z�y� ���K p���������w���/���=��Z��*�H�ơ��ٳ ���cr1[�S-'x��"�f�JtBИy��<e���Bz
�]ytCY�Aԥ@�Y̑��MUٵ��m��_mO�do�ӥ��\Y����/V'�����K����cM˗ڦ�(٥Pβ�zQ@\�8�)���}��5A��<�o�G�P6��.a�K\��%�uu7�u3B�(>�I\�{���6Z�N���0���ܷ�8O�O�9�"����7�Ļ�-.�.�y�JX�@�Y��y����sv6c���(��ݨ�=`����h1�l5�b��p�h}Z�5�����Y��S4��̴�-֝�v��~�� �u��!�v0�u-�A�v�r��BT������y�C��r_}��.�O�
G��@G5.�_\@S5�hj�/7^ĉݾuɐ�5��;�E�<�&Kؚ&lL֧K����9��ʤ������ּ
MiUg]���y~H�1��Y4\�층�8X�X��Y�*��+����n���	��|"Ϗ�A���2*T�!��G�\��N��ApL`:%�8N���G
�+��\��Jr7Q����U�,V�wld�w�Ի᪽��(�~��0Z�ޑ(�D�� �N���؉{�#wB���:�&Sl�ډ���
G��V�U���j�%j��q�^�D-������IMѐ�����$�$c��b+�K��x�0P�/Of9�r�I��鷦�R��{� Ln����9D�$������g��_�*��W�'d����v��vLa�L�4W'��lO Э�=��`�/e��|p�1�����,U�s� F�M`�AhM��f0*�i���l���B��q���������?35�,��_p�`�`�4k������������!bq4��d	8\�ͦ3�T�B}��!�	`l>oj̚温�� :`���3o���3S�}��5�)c`C٘���zAL �^/NP����&e������g�L�i �QfSC����ų�BI�B� 
���D�v�{�`ܜ�\�Ў�.�����Ͽ��;x���R��xr���@p���"#%uok�ޭ��>y�wޝ���\]+/.�9�������������������䇾����}��ΌF�99�s��#H�9GQY��3�E��r�qr��9�����ؾ����W�E�`@R+�g}����W]]��B�����Z����B��~�x�mP�����پk���۞��A�	�ӣlbR����#�j	�j���Y�5�X 45�v"45Չ�Ԁ���M�W�
a�v�#�>5h��:
�Ф5�sk�@�,� ����J	�]T�@�N�/���� `z=Okjz*]e��2Qg��H��ŭ�vj���96wINUcU݁}�����m��3��2~�y�\���f/-�3{Fδ�i<�:xjO��=�'�:����>4U}p��m��u����v�h��ɺc ���1�|t�f�������X��@R^�=�^d*��\������=����������݅�9�驅����:ߦ.I�ٕ�fq����gBSSd���B�?SS�*�2]Fj���q�Bg��$��&�+˓K+S3
��,�6E.M�2�MƵJy ���0�,���SpE*>�C�"�ǒ�0��Xj��ǳ�$®����<&8240, 
I��8"��$�&�	�QĔ�	�<'ˌ��E��1�p6�����F�""X���qV�#�It�e�3
�"�%e�Ji�2
4552\�
_���(c�1���Փu�&=��Dl2�-�z+��L�3�k4�-j�a%~�ȺQ`������ⷋ��(Jyݝ�A�����ж�j�i����;���}�C*�_����ߟ=�����C�-�IL�lL�5:��������*)�4�Gj�#���H�H�x��<���/��hT��U��F�7J��
�Wj��Z�Gz��j�=��朘xZB<-#��?NI�g��
�9%���vN�\Q1O���*؞�q��-��6	�n�Yr�,9g�^�� �,��f��4�ϫ��T��
�9���yZH_�SOri'��%u�F�"b�	1cĘ	2f�����'�	q�E�`�&9�).�#$uK�=j ��qp��cI��T�'M4�.L������lФ��4��lH_����W�@S~�삭�R3Z���@hjPY��tx�p�z�j����2945]ŒN��^$t�D���YN��W�@�R��ZTY����՝H���kFV�^�Uk�k� ��+�_��*
�� ��#�:p:H��� 
�� �ů�4���Ԭ�S�?G��YL�|W�|�{�����kf az�a�kf�{��5��3����|��G�����|���~��_���_Z=;չ0�w��~a�����w�nd"a�����=P�䡦fy0�aL�ܚ���$��|��S�j�zղ�YPY��ox�Ohj���_�<]Lͦ�f�F�T)G*C岁RI	��G3}�����Ǫ_������on-����o/�����~e�./�ә��N��w����»y���m�3�דu�m�eoVF��d�i>q����N*�終�j޲�5'��3���3:��x�k�q��%���yQ��)����a�,��E���t�W�/3ퟦ[�Ȳ�b|Y/���<P
�H9we�t�tX@���y��#���E�,bF��<�A�1�����8&0�k82`$*lAz l�P�����!b���$�>2�0#z���b��q!qBD[��0���i�=L�۫���Iv�`<}0�џ��Oedp�3z29]��D���"��>��?_M"k�6�Ϲ��{<���^���L7Pi����[�ʬ]q�U��E����������ƃ�MǪ��k��컼4����7�Ϳ���{/�|s���S3���<5Uڳ�T�"O��T�`�،�x%�B�4S���l1[M�S��p|��7��zb��^bb�X8n��퐻��E)qi�ngyk�ޡ�������ײ;o�����7p?g�~z��+�K�������Ỗ����;���ց���_r��y���������]�C��;�We�H[�K[��yʹ�rT����5�S*�q"S�L����:y����������qYhn+��AA�frU<�&����@@o��j�+��T<^�t�i֏z��yJS�42@+JhL`{ů����&������������+745 �{�5 ��y����[�rW";EG�H����	
^S�*Mp1�$t�A?�Mg���D�WkL:�A��*Uj�B%�ofj@&�i�"�*_M坤 ��;�2�����hjQ�2�*g%�XijZ����&W�kj FL���zz���c7�5���UY�cjVcj��N;AF�q�2�G�ҰQ��L2�+$ |F� �	4�N��O�?�����8
�X�PT�_p���7_}�w����Μ\�}���=���bP�������[S*QSC$745QQ�E �f#S�S���`Dۥ�-5OO�ד�x��� k��t�����NU45����W�ʚ�/^S�����O
�0��ohm>�9,�*�uI�o����h&���A�x�����5;��f��?𔦦���S.꫖wU)����T�Nmy�)/��.J���lܻ�a������{�F������5u���,?��jM�oJ�m`I��x��N�Z�l3�a$�$��+�#151DI$N��`�3�"Y�>�$2�����3f�<^�I�&��J��B�%Go�����֞�HJ��e���l�S�E�kQ��B�"�,�7�L�B+����"�75�`(���,2�
͌b;���/��[˒J�\�G�Tcd�L��+��:6Sͦ+�%��dq,���R
�H��H�,�A��� ��C��c�l:]���IX
�Ʀ�ix&���m�S�J���t��Ǖ��lL$688l{p�ְ��Ỷ�o{&b�sQ�=��/��K�3��nc�
�:(�4&�@H-��*��*�FA�S��UXhj� j\�_�'���\��h$4�IMVr��\o'�[I5Z�3e���
�h�Vd~�������2^tƿ�L����������U_N�Ul���_�D����܅ou�}33��p�g�'ؔ�]["B�యә_�e߱��(T��P���m����[���
�#����V��Q��;���*�oT��t�oL�/m����ռ���w��tNN�3�ldj�+*�I5"kV4,hj.��-"�ݐs&�y��E�`��3��z��g)봄yJD_�Sãg�i�i
n��'�N�1��L�H�l/��<Χ F��N	v�L�N��~;s$�?���d��2D���t��<�٢�\!t4P�@G�����hհ |� M@�5450��S��P�48� �5�jH�r%����T�Kw���XAe�z: �ߥ��m���X��kC`u���
��� ���i�7BSA���T�f3M��bj|�~��O�@&��'���t����Όt�zzfG���z�4���?���_���/��w�����>|�E_S3�_�4R�2Z�2V��AF���s���FKWF
�=P��-e��Z���L����?d�?`E]H���45~�U$~@��v}/�{"�(��ؓ/�����15uZ L�V��+��%����:rt=�����]կ�����?�r���_��b��7KC���v���=��n��͏��m���;e�,h9s
Ƭ�>�`�Ì�Q6fAB;��P �f�3.$���t����������I��$뛢��
���M�:��}v�o�~���MV�')������Uw��k�u���B�.�"��w{Bv��LE�LF�E���������0����'t;<2��=��Q|�%j�	�DP#�)��p7�Ǐ��cR�2�eXN���x �4�6�`<}(�9��J�e����C9��l~o�'����р�CL��J��e(k�
d��\P�����t�K��I��nuw�����]j�ttפt�g�Ko��hl�i�[�x���HI١Ҏ����_���q�����|�w��K'�NL>;�2ӟ���&i%�<N&�ЭF���b�gXYZ�	�9:_Crj�^@��Xh@9M�"#��L/73�,�r;�4N\��v'[
R�2ss��U��zJ�Ow](輜y�RAߝ��{�C�2�&t_�t^6u]6v_3�\7��6ܵ=��hx������E��˺�����ޗ��/H���$�{Q�rV޼�l<���R�K;����5�SnM�j���U�k��jF�����9՘BM�K���"3��Jw[��I��jU<�8-��l�4�+��A�^�5�נ� ��f�75���� @�v�`{ vAv��aI����.p
�F�LؾYz5�
CЛ�����ǘ��
mO��#e*t�NEi
/CO1�1r(6tGخ�aA���}{lt>M��3�4�@����Yo0ju:�Z-W 635B�Z�`�Mg��p)\L,�24����jb�s0X ,Mͮm۷oy~�s�l&a��R�C�HQR�5ԟ6�Ұ6�0�1���(hP֙�Mcj��I�S�\���gb�!QA����;w�?��ག�'D,�W��!���0Q���9��Լ��;����S�ܹ{x��NϢ���x��8&�2�T*
��*��R_��55p��cj�4Lbj$�--�@-0��z�����ԬJ�rM��v�7
��P!�`g|q�yVM|j����? �G�� ST��닯��F�7��u��4Ȅ��2��35���Դ���U��:Uw��p��խ�w��L%ٶ���⊊�BwyFNIB�˞TH��HT� ��憄�v�o�l��GP�v�C�!a;H��A�	�A�H� f3�"�I.����`+�hdYl;$���sf떘m���ڎ	�G��)8��3\"�G ��d�f��M<z�����d�f��$,���l�";��BuZH��[(nbjJ�X.���,��;�v~e�I'�l�������-?��Fص;f[ f��蝻"�D���c�b1�C��r�R/�h��%zwTH@Lxr(|&K���E|���q�4�$�s���z�V���	Z�����q�� <&��'FBw�BHA���ݻi�� ^p� $H�ӄ	Ng��Rj��V�$�*I�Jb��P��֪�a5*\��P���� �A�A�j̤;��Ak��5�Q�ĽJ�S�8ȋ\L��X��vm�[U�/:�o��^)L�nͿ��C_��[�ٴ62����
�ש�T�ܯ)�zoò�ݹk�Xh�ɨ�k��t��d�WD��ŧ=�����?M���3��V��:�?j�T������W}k�~nVhV�� yAŽ)�_�P.�(�T�O�<&�fE�:�e��s�x�M�f!�n�Q��x5H�7���gռ�JDӜ��OK�+"�2���%-�Ǚ�2f����f�J3�"Mq�3<�4�:�G�Pǅ�	mDB��PF�Y���p���NL�)G�$CY�LQO2[bo���;�'O��h�ŀA�tC\�a�jf�A㇟���r�����偲jXf�	-Yjg��A��8�nPe�1%��R���- ַ����
 VkOȠw�jU��㶆�A4�:=4,�ρ�d���O��s��-�����I~��8O��p/��gn�wn٢^f=?25_~�!jj����w^�穙�o�������X��H���irOf!��W��?���`@�O���P���25�)T��=�<�w� ��Bo�X��A_ؓ��� ���F`�N�R�!�X��ߩ�q�J,�5	K�r��|s���R����Ŋ����+UWJS/�/�.e��%����9gF�Z�sN�sj渄��cG�YuQ�:�b�ȩ���5�Mr)Ay#E�J���/+r�����$�;W�S~[��g����ѕ�i��]��M��%-�
�p�{��_���§1�����i|�6t(bwg���Q� ѻ�1���@@oĎ��퀾ȝ`w:I���E�ӣ�hQz�-r�1@磊w��<b�GFUP�ԴQ-0���(CFʀ��`!ةC	��d�p*Ǔ��d�=��p�p WЗ����vf��4�F���P��;�қ/��b(~� =�#y�6��å�*�t��{ʬ��	��)���]{�6f�k��w��z���Pq�>W����KW�|�֥�_�|�Z��S�/.�?;�zr�ui��� K7�My�L'��	vV���n�g��Vz����pt$D��@?�۷1�]&B�� �efJ��Zaa�[9�v~�CZ��K0�&eg��j]G���V�;O;��u�^+쿝?p;{�NZ����붞�ޛ��ۦ����l�Wl�׬C���_2����yA�y_��@�����>�N�9A�9�3��m�q}ݴ��O�w���,�/SZӴ�V�5jqjQ����ȱJ�S��p�����n;�&���&��Kf��,���E�@M�iPG�C�PMgހr-�4�~Ssֱ�iжl� `G���!�£�$�ybS��S(	N��C�A ^y����@S!�*��EʊQ��f��I!��];���7���5��D�L<����4��bRi��3�k#� �^$��#�A%������Vhjp�"�(��e�$9)SE�icj|��MMk6�����5�Lͪ��15�15�	�B3'IA5��R:������s[H�n�Wo��3۞��; ����Xp�x���1����}���7^y�������Ο>���c�����Mg�������j�DM�L��n������Ԭ��`#��P#�S����75��w��̈w��|U��xJu"�&�ڐ�l�Dj`���P֠U���߀�� `�>z (k���5
T* 4u(��xZ� _Sς��g����z���� }�a>������ܜ�j�@���Jy�L}�T���Wf�r�*�RKr��R3��	j��G��	1M!�ȅ$)/bc��.3�͈d��b!N$ƊD�8V(�� b����r�|>E$�I$L���R�4 �ܪ����.�� ��$11��&E�	��˝�-௶�ճ�]��;p۷�v����q�&&)K+�1
�"�M�sm�B��J�0���Bq٩�	��x6��pۙ�AI��i�g��rFxl�ϣB���#�B���@�"�"��%���29D���ј`,!��&pD4
G�5%[Ɠ�*��.bah8�J�4(�"�Oc�F���,��֕��0��H,��X8*9�B�`�b�4�I�	&���ء��� f�.��팭-y�A���K�j5�FE�S��HXM�
S�ࡩi0R���F��Hl�RZ�=	��D/��#�E�ۧ��F��GN;D/Te���|�"�~��z����[�����_�{~�v`N-k�
;D%5�b�vnm��.�f���Y��<����ȉ��;.F����GyC������G�ŏ\������Դ�������F�ߨ��ɥ_��_�e_��hd� s *_ԋ器���+
�S�d��Sj�i���sV�=��7�7㜑�"�dY�t� :��VrV��r�)kED?��,�	��45f�=A�'!�Qb&��ia�K�Pf��)uRL���&et���>��M��Ǔ���ҩ�X�h$U8�.˒z���ْ�,q_��r�τ�b?G����e�t#z���@�~�$���uI`�������U��T�@�� @� i��ڠfǗ�R���`e �
�� �Z{r��c�eh�ь��I���ZhX@&�`P���~<������:��@��L��OSe���y�/>�໯?��w���_��Go�r�����X�lo�Tw�|�	O�������~:3R|r8���i��Y��)M����,��S�@ӨO���05~� h^`�cX"�Q��e=����'����ӍXf�F=\!��S��T� ]�J�x����������~�E�9�'�Y�CVΐ���,?��XxSz`��]��N:��F=�a��E= ��J��Z��v��N��uw�gu��m)��2����ߔe��4���t��mQ��D��&��:�]9�s�s��[�G/2bg�����aL� &p 6�;jWgĎ������m�Έ�]�; C��~L`o�n����'�13,�,7��L�1��Qf�0#j��È�fF��H%ţ�{�Q3�cA�2��;�G��Ɠ�� <�BO�h$O4�/����{�~Pe450ї'(�:��(Tl�_��_1?G�)�v):ݪ�R����_n�MlLh��j�lk�>��y�hٱ����-mS�o������\ﾰp�����OM:9�4ѝX��1����.3��lq��xnF++��cc�YVMM����зAM��L,7�*��J���,�rJ@{�&ʳ)
�m���E����������j��*�N��]u�,쿕�+s�vJ������>dēu�%�畸�7�7�ï��_�����zA�� ">r��r��|V�rV�zZ�g��<��Q�K3�EI5�8��h3�T�$N�OVs2��,%1[S��)�Dic��A�>ٙ���%3���A�w�v�PSe��5�^M�:ʐER֏~�k���)M���
A�) �W&�LД����9�}2�vCЖH�b�ݳڂ�i�G�Ex�<5=��)�Q$]e8������,hj��������DE��=�@�I 8|�F?	�<��0�hX�2X�<,`�nnn����;wnݶ}�s۟ǆ��x��j�Pe�%駊��K��{�i�z<���L֬35���ԧH�6~������T5&,*pG��-�۷é��oy>p�.�eB�����.�5`~L���̺~��k/�����|��G�O���NOG'���Q2�@�`�g>)�T&}O�X(��l
���㡩���/�&�;��cbj��(����"��Ƞ�]��7�D����J�:�Z�H�M���V��<�ԴK�����hC��pM�@���Cc ~5h��f�9x������Z�[�h�rM[���i(KV��݉�\�9I>f���gF�(�F0�D���!d~EJ�� ��<����c�`PD3Y!!���
u,�M���':�܉��*�����xb<[N�#/#p$8���ǐy�xNx,;,����Rvl'o�Fھ���yNh��$efh8F�jj���"e����Z��,K�Ǳ�휲x���U�!!��b�h�.$�	�cB�!Dl�Ťa�l"�Cd�	\��#QX8�@�9"Zf~���@���gl�po[J~:C̖�d�O��IX1KoP��&�d�;L:�R��l�F���d|!:�����Ȋf�1�wSwo�n�B��W�ݿ�E�LaD���j�NC�U5�5�N�Ԩ�:b���`�4i	-z�^eo}_so�5�Ւ�ڗʩ3�[���������{*��fC�M�o�g^O�_�S=̉�����G[�[��;Y)=򞘈lT6�s��?aTW�fy�q"�{�ζ���Ȗ������W(����/��HJ{�.}TY�����N������h���Z��T��X�B��V��J�I�i����V�C��sM�zژ��J�)5�4��\4J.���MsR�>!�/��'D�%!u�K�g�g�IJ�1b�>F�%#�f���b⡦�ѦŴi)}JΘR0���igZǝ0r�SA3�*OOd�&r�cY��L�'W6�#ȑ�g��r���u-�&h������?A�#����F�@F*� ���40��@;@w!`���U b=������9��=e���iQ`k3 ��փ��� �Lt(���9 ����?=��S��_:�f�`���9��*�fv�{��OOS��'���'������7_~���o���?1rx��i��f��ny������+î��K�P��,d"���W��,q�75������v����k���NB�, ��n�^��	��z�^��t15(uڱ�h��x��S��T�KU�.i2����)�� �#���ɝvj��tD�_:���Cz��H��s�E�D�8�R��T�l%Iz"^�d��.'��g2��rMWrL��-���|\��UC�U��Vf��*�o�r�X��7%i(J��3�Lӛq�����*�9�4sVDX�Ĝ����9n�=H	�%��{I!]�]��]=�ݽ� @!�O�`�x���!J(8e������?-�M�1~� /���ÏR��!#�3�pw�p"���� �4c�±\1�4�ybO���^oLMG&��g
a4� �>AS�ʚ�"������W����:e�.yW���D���t����ƾ
�@MRwubw]jWKv���������C�5�����v|������Ǉ�OMt��:�8�8t�Q�"���v��*4�yi)��xn���mgd[�yj�iui[зt��%\�քu�q�f�VZI�Vr��Vc�W��6n��ﴊ]Iƒ��
�����qoGK���k��o�a�J�����k���9�73�o%��q�ݳ��3�`~�6���e���+��WT}/˻_�u�(m(<t��|��|V����eYײ`��З�(r���*Dq.�-�b��k��jv������j(����BuT�&ڥ�u�n3�m����8&45p�軂^���ߴ����.%jjЀ��
�����
�f3��	��L�_�ηi�l� ��"l��CH�M��?���'�> ��@�vk���8���=H z�5�U�����|e��kc��rtPl(��|L>���� ]���QX��A; � ��0X�e@@���] 
�F"�6:55�P�����-�d���t񧊩�Kf��Mx����{���5OSӒ�*u�RTt+$G��B"�����7he�έ������  H�w�D�G@��県�+.������r�����ox��,V�@H'Sp1����X(���B!�áR�x<j��]
�����SCÄH�f!6EI�ђ��$ߘ�����f"�#?!C���5I��dZc:�%k�N�C����P�G�4�<8h�</�Ԡ�1/T��j�(h h�ǰ���Q9��h1��Z�^!>R,�(�v�����V��$�R�|��c�H?����BI�0�,���"�c�Z]�c�,E$IM5�Xq$��, [+�v58���Q`)J����u�jSy|���&��q%f G�1D��pn@?(B%���� �QҨAX(78��ܽ��c;+`�("��#%��yz���q�ɛ���I�DfY�8�U�.K�ċ
�=BH�G��G�~>0pKTL ��%ņRb��(.���OaqI4��E�p�F,[L�k�|���޿v����œ�#��tW!�$l9W�k�jG�=#;)''%-�n5��r�\��i,:������F�F��F��Q���@ZT ="���������ή�K���
D�*�NG�Rb��zbjj Z45�&j����L9`��gHb�K崦r�� �F;��J>�<h�6)c��c;���9�ת��i,��t\t(�%^q��]V�R~�'���{"k����GD疿n�`F��Q�ut����>���s��#c_�>6Y?4�?���6;��������M��{k��5�Ϥ����O��O��OM�/�-_%�}�d}Ӭx���Spn�8�E��e���3*�9炎wQ���Z.������H�w�Ӳ�q\H���XX�$3��L�bƩ�c��Qr�*Ԩqz�83��OISb�2)��+h�*���5m��X��6�C4�&���2�P����+��ɇ�d���~��P�8��ޱN��A��p�|=C�?8 *h�d�3Ѡ���G�� -��E�P�8�� -F�Z�d����f=}��P��W}s@���[`�Xݭ�
���j��#|���A���́
���L�@L��A�����	�$��D153�(<��}�/?25�}��W���ן��7_}�Ň�z���d������Ɖ������c�����n�J��`��P�_��<}L����C�9�5��M�o؝�j����������9�`^�����icj�T5��X�&���{�3�ơr�`�b�N?V��u���=���LvW
�+��OJ�{Y�VZ��ҫ'[�3)��t�l�h�ƙK�d���.��W������S���*�R�b9Eq9G��8ፊ��J�>����:�7u�������ߗ���(���ׅ��i_qH�8����^\b��J�#o���S҇�����W!,�K&�����Gy��̈!V�3#%��)�2��;)!��qCb��#��W�u�}��N�%�RC�<d>��`*�p:w4K0�+/���G�D��������^Y�T��/dů�����:em�B�1$!=�+9�'o/�v��{����RZs�����w�9Vv���c��k���x��ɮ�屡�s�������iei�$u\��`�t̼4UV<''�	j
LȐбq�H.��)�c��q,����Sj��z����s����2�e�&j����K�-uu{[�?�}��shp�����kUC������e�^O���m�m�~`��<��u�����W�ïk_S����yY��@x�&�在����yuӂ�a�T=�+<(O����%�L�ّ����i�Jr�
N�C(T�(#\��"M���q �Ԡ��@w_.��"]?S�55�C��+���*�~�*�'65ߘߖ
���( 4G��� �Mp�0�e�X $�5A[\d�� � x/������)��| (�Se8Rfh.�:x	V@��c�C@���15��'hj� ���b�V�2h�z�F-W(�J7�4�l�.�� �"��D,���. �N'S�.jj����hjxd��G6�H������bj���jlaX͟45P�@Sxژ��9��I������hRdpd���������;$h�nA�Vޙ�� hjb#��ۛ��y�칗����}��g�N��q����db�|@p���'� �5��!�����o ��cj���J���K��5�<ѩ���?25�M2��kj��O~�F�=���x: �IA�ԧ@������x��O�zG�c���yZS�V"訔-r	:+t�����B#'K�J���x�,#��EADq0QATE��QxmQ�!�#�j��t�$3��@�q$<�&1�F�$���Dd��yEZKkF~[aY����Y�T��N�IL�e�s�1},ހ! t18eD�,4R���޽���2v�d���X�	%W�-��AF���6���zY�$�AM��B	�������c�##��w��D��`#d,�Mf�4���ah�T!U��L2��'3H���~��oo�|w��ʭW��{����C�8� �X�,� 1/��PK[Oہ����˒�R	_�U(�b�I��bq�|��`b0���
�^Ol�\�VR�vZ�vn�V���v���=G���ӽ�_�%���VC�ӓ�Fu��~�J;�`LdL�H�BYӚ��4�)��^;�X"w��T���R�X�j*x�2�V��f��~��Av�[���6��W庑7ׇ̧���ǧVnm#�tb��>��3$�s׮��;��l{������eZ����O�ӿ���,>�������{��Z�Gr�2Ňͧ&�7���R�IO�8���^~_ι'c�U���\P1�(�g���Z.jj�i80g#��l�I󄄾  O�q��%r��"Fɑc��qj4�l�1��(-z�;��!�z5̈́�:&���h�ZƸ�=i�O;D�	��d�p� ���F�;e��y�q�j�@1�/�������@��O���J~�4 �ьVi}e*e�2Q|��]PYƻ��dx�e �em��b	:�	�hd���d%lo�VS�v����v���v�����c�Z�
�i�M fB�mȄ��� �u���<����5�f��s�U�G���/?25�~��w_Mͷ_}��+w������nB�9�:9$�uT���\T����]A@z�����C������%�C:�;T�S�����{Μ3s�����;�>c�k߹q鿿\���]&3蠤���)KT���R%�9�lgH�8V|W�`,mo�x�C���K�d�K�����
��̈́�q9.���Dth%�F��A�s��n�`٬��ʺ|�扣F�=#i�j�(���W,f�Y�SJ��Y��DN�eYg ����}���#��l�o��lON�_�fį][�*8!��c�iM��^H��K��dt��Ie��Ұ=��Ϋ�xn)�/��A�Yo?��l���i,����)������_Bryr`YSe�Tp�����}H����
�.���>�g��aܖ;oj�E������.��/N��f�R/|���Z��L�6nv��RK�R��I��E�,���8��6�v"#�jˢ�U�F"��L"�̉�i����/�r���y�>!!�O��9�%G�Z�]K���������3G�fsӌ��Ε;m�Q�9cC�v���+����xQ���=�H�+���iy��>a��Y)��ȅ�RY��*i�ctD��z�I��`���yS[�ǰ�5_v���w0��3>�˿���&���;>Ǔ�-�#�I�C�6!��iG!�!]�
f�8!��+�_�������
yHfX"9U)/QZ�1[o�Q�M;$+6�����S�if#O7�Uʷ�_���W4��9@8&V�>F��gv���mB���L��J$����'�����qX��>�iH�WPM�k��v��6�� ��>���-��&v�.W�ً�Oxv'�1Eb>2����鴸��W�"�c�|����V�����=fr�稒���b��EGE<�C�5.�F^3��,�!|�׎��9Ș��ڪ�����^v�&`<���4v0 	Mw���KS.����1N;f��L�
�~+j�����BHV.b�%��gEf��v�67�,>��
&��%+y�\���찺Z}�-b5�g�%b�'%&�<"" ���H��)����͹pY�5�x|R;��>��L7�AE�t�q�(��2=�N3(���fP�D%I+#�)?3�r���^��2<nr��M��hu��媮��JN�s2 �Ƈ7�h���^��$����d/:m+�!���e(aފ�����#��y���T����]�$�~\���2�����w�̄����Ģop��)��\.�M	7�d�����J�]c �����g�ˈ^�d�U�S�2β<����C�λ�V�X�yG��f���D��k�R��T)�MQX���U�,.\���#o����kw��N�����󎌜����֖��,b�`3���UfԎ�V,R:���
�J�D�Es
�UlDэ��p8p�pJ�&�����6�<�Z0�

ͺ��g��¬��pjGD��&1�=�X������·a�O������ttd���ǹO�P�;����-\4fq�%g�fx�w&�YN��~�SN	�Y䞶�\8��<e���4�"=}cr�9KUI�A98R���-IO��ͭA�����]q)*���5����1�fO��Q����P~�=^�j������*N�N�7�n��X�w�Q�^�3a5Z��˗���EV��rn�(AHzW���0���Gdvښ�ϭ�1�M.�����
�7�����^j�'�������o�q+y#��;�ŷ+t��k�*��L�U4f.�
�������2%���z?�"��A���O���J�8���zn��J�9}����X���_�����ݴ�����8aj"��?Z#�`+ޔs������g������s�LAQ^?v�z��+�NV9hݥ�HW���Q�yr�Q!y��A�;c-^�ezڲfq�w�%���6���X���W�/�H�YDq��U&͑	*Xq
�����ĨzقؤЕ���¡�*�?�lY�n�ݹ6)���^�I�t�z��y:(��'a���Kf�a�;(c��X7�����K��*x�E�@��̟�>���IJ�L� �#"��͇k"��(ّ��fvWbǩ�"�������	=�^�oz��]�:k��l!!�L�I/�N�"�.(�D��3^���K�?�O%�*/����(w
��֚"}_�w!Ȱ���2��wXSD~b-�Ԯ�*��(�t�i�_��R�S�<��L|;��If��~K&��>�r@^YD#��fHã����F�i��h�W��&㗙a�	O���B��0�8δnkH�=��T<#|V~���$���I
$��{��.�JHg�c���I3b07�`�����CUN�����X�� 
�C��y�D%�Xt����I�:ba+�f�;�D|?+��}��@x�V(�h���Hg�w]5e�`q� ��})��:}戽J���0ju�'�(B�V� �ff��˝��.h� +r�	�b����o��&G��7y#L��,%p�n@��ñ�:w��ɯə�ȩ�[>nX>�s�s���s�}�118�Bnc��)�n�`v����Q�=����ȡ;*�}1����:�â��?��w�ߛ�r��LzĘ��Tp\�{XeF_#�_aB��c���[���r~69Z��_��	�S�3u��qIx����pW�>K��K�~Qcrn�QA����ّ��̓��5l�5'uv�P!0�
��	g"�;�|�=�@Mcz�a�.QV-�R_P��|M4�&	"�1�m�}�u���y�M嵰�ӆ�G6a;��ފ�˩����I><���������h���̀�Rl����P!w���i��E�y4ɭ|�?�꧵5��%��[����0ԩ��o=?N�;�{d���9�ݽrb2��[�t._�۾��ZÞ|��S��=����{��`	��d��c����TE���ͳ�[��|�bR�%��TEN8�Z��qec�X�޾W���Y]��%!����ME���#��x4��@������ܧ��U�P��rrK.e�Sǡ��3�e��O�����;�g��C��#1�)�_������c�O�=f>`Yx�v����r���\�#�����OK�GD�j��ԯ���_���C��,�[��:zc�K����Ĳ?�z~��뤙W�3�������^�2��@�GpA?�x�=��Up$�$��hX�4t�@���C;xf�r��Ɣ���Ǐ�ue�kE-�8��o3�A�n`I����k]����Ѯkr|M�@�Э��
?�Y���/���-��4��6�P��d�yd���x�D�A�d�7�6kУ+3�͞�k�|�_��6Bяt�8-<�^a�B����q�^
W	GO��F�UD���� �G*�ԍ���S���W}����t�ֆ�N2U/|6 p4G����*.n��uQpḿ��!_gЁ��2��������X�(آ��$���`F�g5�q�9Ȩ)�/���i�(�����cp��Š���S�N��b�F��̭i@�� �\j�pܑ�Dď@$糐�����7�D��Q��2�Ci��(�e�����y1/�RZ�Y�J�j&Y-7��%��х��lPZJ�@��AJy�6QĈ�'�%����KS�~2��s��w�v�k�pa � 8y�A�f��o���?SA�]!w�skIA�vvQ���[x�+�b��B�5^:�o+L��7�a�Xq�y��y��dfV��"ߋA)=),���S�Phw;Uɬ��C;o�@����c�b�}x�,ҍB؋����a0��`F��ʆ�TP~V�F��xb�c��K)�r��h�5�+�.�,%�Ne���
��~�d.ͬA9��c�q�P´����:�l8M�dK����V���z��ci�cd��i��7�l���V�u��)戺fJ
?�(��d㻉w�|K�β��;vp����;=V"�ā%B dTS�H6�p���:|g[ݩc޲��#|�#,l����5y'����l��-OB`��hD1���X�#�����ND~a��;2*�g(B\07�hۦ��k��r�B�Bm(�0۞�0&�� !=n�lj̭����竉óBɻӡ��a7���~���;;�	�9�*�h�k;�Xx��|e���6c����p���r�����?��+	}��h	t5��o*TvR'/Gi3�0_��NEk1f+(H����|9e1#�Z'_�1x�Q��ՅF�h97���2��Zo���9�qzJ��C�by�e{�n�C�>���.1�F�$�.)�~`!11"�8i�QoC��ČW���"�Ӎuжd�����i?j��>zZ�f蔕���ث߫��)R��y���+GG��f�<@��q�SS������}���WX��}�闓F�5Ͱi���E�T�"�4~���o���Z�=_M=�|iJr)��`�U܆B[hMWQ����{/3zPπ��B�ض�@0�=���.B{@����oXF-��E�7�bM��ڑ>��!�	T��{�b_�n�窤Zh0ˉ	�.� 7zo�٨�̖�{;?P }��\.���^V+%`��?	���J����40=�B]`�ֱ_����Wh�t?�~K�$9���?Nah����)/_�:���8(�Et��FQr���H ���>Қ{���M��G��%m���w��uG��ǵ�X�/P�;����!�,�m�T���0���Uq�~	3q�0A
�#i��7BV��?����;��E�>�z�2!���X!N�������
���|>�M��T"�L���h�:��\�ć��!� �@5Z�B� �j$�i�5�4����:�E�����,f���ٱ�������H` ����Cp���5�:��1�;(����lh��H(����vU�Hu�C.&��d~/��Ρ���hߩ
���!G�F9��F��doD�F�^	mhRW��\��2��鈴j�:��o��o>����5���/M��o��'�u��|+�5"�2ѥ�
�8t�B���2ѿ���a��f�Nx�i����L)��W�ۥ������.����������-.B������Sv*�Ǳ|��17��,0 a�Z������Y�Oks����\;d�DH�$
ٗTc�йB
$R��m�2o��6�o|�����̆ �	r����yn��r9�l���]" 3�"�"��Q	>e�0-�D�>�B������dE����Xr���i�B*df�Xs����c�Ե��q���E|��<gL�} о�L+����WsZ�h�3A<ED�@�~ɨZڭ��\M'zb�F
Y�2��7�0B@
(����)N��~�Q���b���<P�E�/E�3��)H�ۄ��z1�Y��(��js��{��h��;( T�}�c�1����d޾_#zu"ྯ 7t�.�������B�Q��Aw�T������ګܪ-�L+�P�l_�T��R���=^����D�Jq����PCJ|�eB�p#h�ϡ��z<#��,�Q�7B�<�J�N��MҐ����@rT(B�FB�D��u$���w)��(���L&�����=u8�7�?"7�B��Ñ�uC���2�V.\��7�Dҟ��Y�ٚ�U!��	�Q�e��;	��Dtl��0aOSǕg�j]������(�F�:9z�ƾY��>�VTq<=���Xc�J��}m�
pD��击���):"�ޡG�bAoM\
�fXf!�XP
���0�)B�����Jj�V��ޒ��8�7�1�K�,ܨ�Q����D����UM��ތw�9��?�[�8����n*17�u8�-@�"A�-B��ep5 Q�[aķs�������d�l8̖�I�3G��I�f���C1G��!�.�Ȃ�2�w�����;��EXP�� 8���l�j�D� n����.Ƿy��`F� ���.=��Q�X�ԡZD�c�����rI�a/ΚE�Q�!��A45�K|���c.g%0ɡ��D�T��|�(���0��ll�����<��i
��T|��|��"#WAM�8���Qd��br9�L_�9��ߊoqd�b?��-�[�\R����QZ�#"��pF��-'�e�H�Z�)�m�IG�[�sa�^�+>)�I}f�3���6� 3%:��ء�b�1�6>S0-���g��R~ڭ��1����ie���e��Msk��A߹4�+駚��i9>�䱹@R�oi���Kk��$̇R��>
l�;T���u^������Ѷ?�" �"�邶zu��)Ӯ�������wav-��;�g���|�������G=�EG�}wbJ�d~�-���6
<�<=�2\����]s�����D=�ŝ��/T�Q��q>�c͸+����G���R�Sz��<M5�,2�f))Vx�k;�n~�i'�`s��zߔ������/�C�Z3���U7�4�4w�6��l�4,�l�V&��]�S�Y�X�B�����!d�)�*���o�b��Q^�j�K�=f�|%���=�5�D�<���-��C��d��s����+$֏EL�6�_��ѧ1>Ow����m��*����7�
�f�O�U�$�xYh��#��H��8���3���P�v�]���w.��;�Gۑq!JJ��Eؚq#����t"���٠�����<uK�Rɓ0q0�B>����;2=��Ո۰���i�S-$�AC`��seW	�O��&�Pe��Y�c�@������Ǐ��b�XD��4��^��EI�V��{�r�^%��,��@a�ߟE�>8��J���_�2�ڪ7+����/v+"�������2L���hL�"��x����}�c��.��l@J?Z�;�;�} ���z��]z�H�	~�#(h��J#�>�� a&A���$>�������L=�q�H����-���� ��vү0��h���/__�j��i[�I��~˫1ǫ�ر�����s�I�H��kK�Ӗ�����z�4@#V΅�c�2����#_��8V���>�#�QD�W�׭�H8���W^�X�%��G��h b���V�И���Ƅ���WjJ��s�k���W����i���Vap�� b����߃�o�Ɏ�ա��Z�����9��.5����i�����2�N�h��C�|��/�i?����B�m���:V�&�[���y��j(x4)+��3�/���t#�/n�6�z廃�kI��� #><Yf`�
�������
�c֯i#�l�2�y)�c����(e{�U		����*&?5E�������d�'�>���@A�+�Ȼ�;�.�ś�_��S�y6g?��5�ƭp�=~m�v"
�۱�����������ɂ���T�ZA��k����"]�"�9I�럏^g@�+F�pE85�������Tx�n)U;�pݢ��I�(�F�@�L	{c�?1�l�[KwI��'�:��C9���%��/��2Ê�<T���C���ƈMxԝ���-�`)ẙ�ݯA��븠5������t�П���������$�3N)C����$�c���%��a������y��oمT���9�VNΩ떦KC%�e�8\�.��pE��W.��R\�Ъvt��|��>�ЍJ�˝�d��)ڄ���/F������D]�"��D�c!��J�*i��.LN����g�(Wp�p2��[Q�h!�#<�;�vߚ����?H��a0A$�\.J�%��?���#����"�Lj�`�[��7��7,H�IL����
�OT���g�R��9-�����p�6��y��#�9�ۛF�;e����C�u!�������fV�<qZfןE�(G�=���''�p�W�j�<OY�yr� P���c,s�����.{I8�_�XqF.FĆ��ʤA�����q�?r��:�Ds�g�O��j�����p�<�\�̛�>��}���I哮��L�;�N�I�s����8���r�X?KDm���Qຈ�*ߒ��L`��k~�A2H�>ﹸu`�j��/b	��'��/)�R�a�tl3�`��UN��0lD� 
-��X�N�S8"I�zt�8"����fU�ɞ?ݻ�x��\6����>��^�O[*
�%�� �3"���X^1-�/:���W�����j�����|��G�+,�B�~�]�c	髯L6z	1�a�|��!�N.וV}7xa]����v������zܰ�+���ǡ5�?aW�c�5�R%Lypt�-�@�J8�t���B4��YWI���u=L�`* L�à�93�f6�"�' ������ڂ�O��ܡ[��P��>h�Uߠe��XK[0e�J������Π��}&ncJ<� 1�Ί�����Y�ħ�͋'3�^ݒ2���6=
w��S.v��$�|,�o".Ƈ��~�mu���v��^��.x�SO7}���9ug��}�����ߥӿ����3uK�����5�����\��I���Y�C�λw���	���
�[�=���#��9�ϣ�U񮓭��4r�ݷ�@�ΒS�}�w"j� �ڒhg'+Rs4I��g�Q�R/��I�H���ˊ΢"���!���N��i��|��!X(��0��/�/U�|ؼ�V*�a%�R6�����ϳ*$
��)v�R�=��
��3��5���D���������Ȉ�i<�������r���
�4���:��u�[��:١����VM�ӌ�L?��m�/˷֦>�ϲ\d�#/ɦԽ��� b�6WR�%
d5M\�.z���^E:Y lϜ>Q/������hJo�c�?#|6���w(EM�Xi[�^qn�10 M�VL��Z^��r2�0K�դNE&I��i���+�G�Xm&yJv���9��C����#)� uw���`�r���<��h{ב�خD�lYn^��Ʋ^�	!�c�QK���+ɝ���ɰ�Q�x��]�~% ����~u�� 0�/��1�G��qȑ����]l�N�̱�z�H��焠�3�Mb�;BH�y��XD�y2�`�}�o��xXye]��-"��%��	��������ɏ��[����|�i&~�R&ʔ��|[T=�\(�Y:ki#��Y��z��Y�C���>�����G�C���n��&��Bc��th������h~1Xe ��������>�-ܕ �
�+k����h{9���֩J�BB� :u��?���ФT爳#�>�U�lPӯȭ��֧/(�Zg���Zu������BS�]u�C_�g�'k��{���/ӯ�J:s�K�:L�%9x�m̻-�y]-�ٮ��Vn[�����2����ۊ��Ś�>p��t�[�Yp	O�z}^����an)�2,�UNi�b�_��XW���D�f������Op3x�Ŝ��2��;.��v��P�/��;��e9 k�{`��̽xV�ݧ���g[��� �ϵ�k:>�J�>�c+fd�<�z�c��!xq���
:�_3�=�}F*yg?�����R1�/�h
D4�"Z�]~/}ӵx�l椪��d[�o>#{	�Nm��y݀��y�3P�࠿�A�mdŪ��mo��g���G�FJԨ=����ͿL��GS0�$(o�C-jv��C���_��l���`�UE5�?�Z�:v�:+���|��
�V�n�ehUN�����TY|1�;�t-��N��Vܯ^Z�Eg��ܾto���oۜ9K����9�(.��)Ô|�$O��DMS�<�#��V�o���sQq����]��_�8���[��+G��^ꁱ��Q��X�3���f�z�h�&o�����������e�D�u�xxD+m�̡�ևg�;�+3�}G3t}AE]�Bg���,�R�̠$�E���0Ϸc�W�c�7�p�DP��,��)�7�vB>��s��Sy��O=��gf{égF��M9�9Ȋ��@i&����5jI���M
������*w(*~� �Yʁ�/��
�nw|�q]K��G6x���뿄>��H�>8%�kJ�nѝ>�z��o��o�*Έ�+�v��1�{�fT`�K�����`~��}dq��m��DU��{a
���E�
���ȉ��YxU|���r�����7����	l&�}l�u��2#�-Ǒ��FV�=��EK�n4��`�b1�n�>��*��m�q))?)�u1�����׹nO�ȅppmE��L2�<W�V]	�������lTbc�P�/r�!�~�gI�0?���Q�B��l��x ��Y5^g8�u����3��+����1��� u���w!5)�yH�j��B��� ɗ͝�j����5b����%3|}��'ℬ������^ԩ�6j7a$+N`�eO�d�[`�I�~�/̚H���h�#asd��#z�(z5��0��Z�� B��Im��{2v0�؎��]u9��'���~C	]��>�d\��:-�4�|�S�:�pz���6�4�̬��K0�Pb����wkl�"���Y/T�����T1[��;����)�=j�D���qǕQIҴ *S�j��I��^�zq��JPs0;��ʸ��u�|VCod.�벾*K���=̿�h�y���BG�I��ݢ:���rо���a�S�?��aw{�����O�}Z�;1Xj�����_�'���_�w���=�~D���
�ח���Ԭ'��ב͵�_�G�n3u������;WS)��o�õ���N�m�ʪ�?��{���ȼ�ɖg��U޴=�'D�W
�n��0���ft�c���xa̭��{�5��5g�B"o@9⤾�[J���[�P�i�`�U�k�<ی��H��sCFֹ��EB�Hl�EV�{��ۀ߆���,X8�hz��3t�a8�b�F=35��h�8�=w��=�g��;�GY����.����D\�'}��=zߗD��Ya��|�ӯȊ��!j�n�b�TBc��e+�&�����4O)C�e<|���r�t��?���l��&|m�b���kT/���K��@!��|M^�ӌN06= 6����N����:u��K�	�P�1�̗�4q���!�ټ��ֽ)���j�h�f�n��PO�,��\:8@u��R��+<�8h�G�fɘQ[�L�6b�X՞=|�濟�����=�Fi�u��#ƈMq����_3T�c�	�Л�C {�k��3-��N��F#/�����[�Z��n�,3ھz���1�f~0'8`/�fy�.�_7멇�)B&"��~�DN�\Je .������{/��c���ε�M<��2y&J����Z��f/��(8����o��_Ķ:_���Yw0�� -����V�u_�^4�Fu�R�#�N���ٷ,7����VGl1� v_À>`G��yupf���a�A��O>_FR���"!]-���c�X��v_UV�L�;��-��l��o����������ټ�J,�2��XI��8����K.J�n�����3���5z��|�^�e���|>hK03�g%P�po�_�Ųޖ�&��vғ�T,�dk���U�<��4�F8�K7� ���I���~W�]���	|���P�>�:��6�����~�V�x�˽���� Kh0��4}�������g�#~K楊f���O�zg�k〲p�ۆ��ފw�o&%Rˊ���t,e����²_�B�]|�;j[�&�Uꉅ�T��}�*O���ބ#ٞ�	�VUcx�+�4��y&o���'���7�7	�q�=�+�s��L�C�ǐ�%�#��As�A����]�^)���]>ݦ};�Mj@��3ȄB!��~�W�em��f�mq�U�]���U�C'G�N��z�ůx3eUw֞���;u��=��J*騥�{��d�C*V����H*I>2[�����MR��O����Q3�ܐ4�]�t�Aڐ˥�g�����Z�?F��@��K�87�*ܢ�vh�F
	��H�p�V�Ӟ,�����eB���?#����D���@#���E�g �:b����C_�.�2��
m�@�,5`:�?��Tiu0K���r3פ��d�x)��T�Tlɴ����**~�j��|n^ZT���P�
�d�bT>֫��K���P��て�pd0'�7�;��}o9j�z;q1}O�#4��b����1M���!j�S͏b�J�����Nq0[@�S0"Y��,���KS(f$
�k�k,�kܾ�қ�U�=���U�q�r�v����`�1�M
���i����F�{ןee���g�2�7kS�[��Hf������F�q��� !߸�壊W+%�xH��q� ��ǽz>��Uh���l}����q�	o��y���U�4Ą�s�SI��� U�:"�WS�E��]PN�htɭN��k��������5�'��xS	7M��☺��&!�O�� � �b{��JZ���������J_��+��C���ԩ-��s���C�e�ȳ�
B÷/yX��f�TR�SY�?�W���K ����v��_��v��m>�f��y>+$�U"+�M`#����d3e�kN�Հ{}zmPR��Vm7�V��%h��í"-���a7�DO��	P`�I���ϵ�+5�K�}��Hd�st��G'f��4�ˢ���Q��[����f��ˏ��
L(�'Zt�|��SЯ�+�-�S6���@����@�yg���6u;�7)�����q�_�π�_E������Ħ�B��6?��X��s�x}0����|��'�r�����Qϟ����o��K2�:�y6��J�����Z�o��������o��,��S���X��E�iȦ��ߥo�[�7��7����G�lܜ�Q��x8�9����Z����v;�+x���9:��`�ԍO��@����V���!�ZU�Ze�Z�#�K6��W��e���ʌt����7��������,�_���2�����m��E'PBՋ�쵘:q�Y�5���>����J<���/2��*On��Y����xn�K]�B�_�͂�H�(1��ڌభ���*��y�g/(�)A��dq
{����H��px �&>�?�֊;++h$��n�ؙC= �;�1!��Q/ �|����>H�!�Y��Q+��^.![\&�8� �8$��ך��M�VV�}�y�~B��N�`v̀��vüF5i�A���������}�c[Vwa�xJ��D�����g�e툦�<�!�E�GmS� äG,p�{6)�`q����k1T*� ����z����9a �f��R��=NL�4K�v�'��N��;�,�$�w��p��֪� u�3����H�%��a��!f��:�w�b!�C��"A�ON���#LI����(O�����(�[([�@<�stm|�$��^O���Yx)��DU� g܈@ rs��t�^ؽ,:3>�fV����G���6{f������rb�X	$#�ߝe��؉H��/������Hdj0���d
?`�!����Ck�*;���*F����f��C��y<������Њ��!D���(������M�$�7���S�< ��zR#ū]�4�spaצ{k���n��
<_N{�W>#��Tژ=��`b�r�.����:�#�n�m�D��e�J�٠c�u��~��W�zl�VY8�[����A�X�v�<M|�-�Q�f���}�h��wpiS.Fջo85���}��}���OȬ��:���r��e<�ͿS�1�����l���巧L��#�z����Ce^���R,���~� 	�����5H�T�s�"�G�U�Y�Ӷ��8e^�	?��z&)i�y�灨~�B7r�W�J�����<N*�2��h~`�T�9����K���|�+O;���(mz-.́2�m��J���W�	#`O��O�
��nYC9��ȾG��z\�g�ۻJ"����8gg$��WS�$ħ�f��h.���&:n_��z��8�� ��(�	�>�g����SG�7?�r�-{Qr��tH��޻Vd�GD����ܸހ.h�FDb�a[��kY$�QO�֏^�����s�s���z�e�H��ܨ��),�#d�E�3C^�D|�z-j!u��J�V��9�2N��"NmxCf����pa�ÉGF�oث�>[3R��VwC_�nG<��,���7��/ƤYt���lV�HV%8��ۈl_�pE#KG[GE.Qzr����r�8�i�
�h>V��n4�mM�@���^�F�%�V�)����2_�"g�Bԓp�N��==�哜θ�-8���2T��a�0���������@��@��X�'�C��tS�(�����i*������i��ͅs�|i�\�!m�~�H?�����L��;Ȓz+
���Jcrt���G���{Y��ld�m��Y�"�s<`4�s�S!�A��k&��uq�����#�@A-y�4|1}�t>����ߌ �'�}��d{�&��	�	u�������؄6��FJ�kL��KD̷�"��kY|�Ն���f8��WDL�jãZbt�Y�#�>�WKf������''�Y�_'��C�*�K�#b}�1;K��YQ#��\nڑeaa���G�1��o�\����O��5AhxIα����;���C� 
,1
CK��� ��� ?��ӾÞ���Au�g���<O�/��EI㞶sq�h�)=x̪��Х�?���­�\tZj��f -�M�U]�Z�P�I3gjt���
A��l���{��Ol�����M*�gR�#S8\��j��m:�(\��C��>7#M��.���Qd�uC��+nC����AHZ['��|	<���<X9?��5��}����s|����d���ѽ�߅��G5������i����w������-��{3-zב�#��~��L�g��~�����{ַ��5��(��kF�o!Fw��2�������~'�?:M�.�n������Y�;��B]���M1�^]2�0Иd_��<�~F[א�"��g8��| Jx/y��n��UI��j�m�"/ei��ɘ@M��uS��Z�J��ysƢ%2G�46��вg����Tڷ�mGˑ5$��d�9jY����d��Ԧj)�����O�d�q��*:�aD��%���?(�j�N�J�{��C'�b�/gӻ؞�
���DJ�����ꇀ�N�n���c�5���I���������G'*�%) �Yw%t��Ҭ�i%n#�����5S/�(q��^Y<x�tי`�&��K3�+���L`�A���E�]�q�7�0���B6e��~/���-3�"S� =�8kWu_���iK��}n�k����m\�؄���'&U��.����<�/㬲��TV-���H����"��ѡ�>�n�&=1���+r�&%�*A�1�PiP0�I���H��d�*lb���6p����}���AY��{���#����r0�E�7k��kW��9���,��֮B` VG�����?[NBEh�c��2��0T���a 3�"]�1�Y����ݷ�X���mN��~��v;���ǹ���?��r*k<6���_'� }��D`&</�؀��$�����Z�d��?WZD��Q>���#ܮ���A-��[�*HN�À�h z֌���2mT1����A����T�5��i����9����܊YMCgt%fS�*	� 7�����E1̟��f�L�!��H�q�{4�d�y��c�fL�'�w)��6����L,p���-��HN�F��v�D,��XW�����`�����:��ұ3a�N@�����V��fs}�BKI�\Cj�^'�U�U0
ޡ�^ G��!v�q`�Mr�*�ȿ\E�g*��u/��8��="�s~��������(^iXZ��l��r�
ܑ����n��i�?|��;>��E�5Jn��V.ҙ��f�Ut�����1��,����Q�=�����a����Y뷽;�e�g��Ov����w����qנ�|�:g���(N�l����.؅�[;IW�E��UhPb�՞��>����������&��0��0q7��J$Qp�d�5��3T��OV��f�C�+A�s�گ]�>�������<� vϘ�I��7�.y.̅|Ƅ��������3�(D���\Dˌ���/�ʹ��ӝ<_V�̀�����Պ��,٩��I������ڂ�Q"����XP������Vr B&���/��	�h�~=�Q�Zd�b�Bx�aG�̞/M��"\�ZXB�#�����3���'j��Z��^�i&��Դi���Tt�4J.*.�{A�G$�0�x���:G�K�#�
%�ЮkY"���!�
bM]�@�}��o6�Δ��v����>2�j���aXbL�$մ��G�C,6Gw��4�龧��d�=,�e�WXM��&d��0��71��@O��ņcB�w�|��O�-�������m�=ne��＋�����ܻu���|4
|�`+��R�B&�ɐ�8 
���4�f��-��������g��`���m�15:|�W��v*�4U��$f]2�>�٘�n�������N'�z[ HCM��r�,�n6O|^��_�L*<�j_8) hC��!~��O���f�Y𨯩�����@Y�,|������Q�Wɻ����l�67e�:R�����i��° ah�4"V+
��8�����V,ek,}^ΐ��Z�TAⷺ�.Ϟ~��߾��;�_�ҝ7�~b�\C��7 %�����UQS����`nZ�A� �B�JlUKlZ��ǐ!Ф .Uħ
�d�����
����CC���G>�W�-?�EZ��$#��s�D�8���v��n�2vj��Rb%�}���1���.;�G+I`��hI:b���� -,I�=Pqx����ؑs�/.5]X�<�Xu�\���ϗ\�Xz�jɃ�%o?�^���ne�Z��{�`鸣�w���?|���}��?������r:�x���ݚ��J��(�y-��U��;���n�u޸�~�����kW�o\-�}������W]7�]^�\��r����{�O��:����\��޲�*ӕ�η�,�2���l�0M�f��L�oc�c��J�J��MZ[�)� ��=�י��J�w'!�$�}bj�S�ґ��c��V_"k8�=ϙM�.���eHϤ�N:��V֩8������IxQ�:)%��#z�9�Ew���q�m��6L�1lX;>��B� ��v�Ŝ���a*�+&�=|woL�9f����D��G��`�i᳌���B�Y���qMϹa�]7pApUǾ�e]�0�!�E�qJDY��v�O�g�N�Ç1�1��w�-�5����b���L��xR@9%���1O)XM�f���Mz�.;�p�!Y�q���d�J��d�b9K��%�ɒNdK�r�cN��K9�V�.9h����ʴ0�0R��T�*���!�4ce��r�x��OР�9�f�f�Z��?��� �k�2��V����*52�p���T 	�2��]��ԃ^�3T�E�K��	�/�Fwaa$�G�@Sc[@*Y P� `�'�4��f���i��� �h�_��x��W��;��=���635�������o�ܳ8rh�U��H��������������}�������}��o���O?x����Ǧ��;jfz떆�F��G�O���+95�>�q�-<�q��.D�cE��O�:�<y+#��F����Eo�z��Y8j�;l������C_�'yژ԰��kg|�+�P�G�f�<k=p*pYp�G����������w\��� �N���'��]��|x�ͮ_����k5M�xz\���:� e��c���lDd�ډS�Z$��F3U���ROm�d�
0U���L�)&J�ɒ��:H�N�b�R9[��9^�_�6 ��s���
�L9�3]����b�A�*Qϖ�|�n&KT�Jȸ[�!�\p�\�v�\ 	������<5~�y���AAGE�������>��.8�6�>�F)]���c�Yq=�Ų̀�?�.IO��](�.�tI:�$�.$���:W��\��"u��/Oџ�,ЂmG��`��)^ܐ�h+L<�Vwy��YO���ᓞ�Ɏ=�E�Y&a��]`�T�(����iR�ElL�6$q�X���UYc�U��V�҆,g�J���֧�3%�9򽹊�,ٞL)��͖#��f�[���st�������ʔ���ꬶ��C�y-�κ������C��{竎���_��Y<|�r�W����Z�$��J��K�S3�&YHh��԰�q,��fҧX���+A첳�,dd2#�i��D�	�Li% ?��I�	��dfc�7��o���(*.� :E`$���Gݲ�b��EG���\�pz`TĬgĻ<�� @�ƚ��;x(�� �C�(�Y��[�~g�/�Z�c譒��(@1������ ���G.��b|�9�@��k��Uz�9G���;K�02��Ho���Q��S�,M��ZN=: :`G��H< $dw0 ��yjp1Ѡ�O!�D����~�D��+4
%@%�#�J�\��E|�  "�l9,.��a�Yt*�D ccqQ�a�a!��+�{g��m;�<��/����>�cklh&�F��$9)[C��S�x������fkb]&�ˈLq 	d12��J�g�; �U��\l�mH�4�q}e�:A���<�\ 
t����S� vSj�J����[2Ue��L=�"&�Qؐ]�;�l~��m�U��"�	�	
�3��������@|:=�a;sr���o����_���k����k�B�a�)B.K"��e�H$��
�,�B��D8U�k��������B����O�0�f�s�����/)*�($���0��i���F)����䆳ӫ�p.a$�fm8���������T�6h/U`m� ?`�y�sR��O|j�1�Pm�}���֙6���-o��7ly`C|=����M7V&��^@u�W-Ճ*E�Q.�P-�4���t+� e�h$I,NCD��q��8F UC����*�C�K0 �j�E��R��5%�g������W~���ܾ�ܵ��3�Ǧ]�m���愒����-��zh�q�HNA+_����	$5�m�sLu�\��Ч+�ic���m0�k5�t����Rbq,�I	�I	�ʉة���%���'s[.3��L/�3�i���*H(��Ѱ�l@U�*IP��/�cZ�yVVn?+IV䎯?XZ�Q����X��`�������KgJ.�w_>�r���׵�E�/ J�\];[z� ke����+���w���.��og>�������s��W두��%��߾�u�}���u��k ��+e�/W\���7.�o�R|�R��s�W��t������-C=����44�ʊ�Jr����8q����o�p������6�^;u_<uo2u:�@�p�H*��4α4.�3��KW��ݎ,^G6�3�ӝ������s��8é���`L&rf�y)��$�|"�D�r���Er�,:��,ɨ3B�;��O�	S�7ʎ�E�C�1��bvv�C�ɑ#��8-��
��|��0B��УF���	F�8=r��!OR����y���u���s4�ԌJ�99嬌|FJZ��,	0'��	aY�[�FO3��)A�1r�() v'i!S����|�i	���qQǹl�_2.Z��q��q�3q����8�D�`)]��!���f�g����9�\�h���Gڙ޸o������&ly�5>�M�IY�' �
hU��*�ѱj��ePS.ڱ�:pl�Q�R5:_+�ǆ� � -��o4� ���*�����D�Y,�P��6=���� ��WǠFu:  ��CQ�!��V�����*�p��S��ׂ�H-�s�ݧ)�	c:�j��f}���l�8���S�0�A�\�#�p�8\e�����C���$Ø����َ\/��Tj]ڷ0t���ᅑ���<�#�#=#}s�/#C`�kg�@���O>�ͷ_AY�����=p����پ����������US3Rp�+kά��S��Ԭg�٦f����������g�����A�~�P��bPL@�T������������¾�+�6�H��M�[@z�	��T�l(����0*g�V�Ț*�L�x�"k&�P���z�Ё����U�\�NKg&^�У>��x#S�������sAypMxYx���A-��˸7 ����������F�D�x����=
Ռ�v�I@eM�K�+k��4���s+]��Sݗ���U�穇�t����A���.i�SͶO4�Ow�8�~e����`oSiM���&-�IJ�eu���\}}�55��lhj��j�J� �H�!Agoo�t_��#M��l%`_��@��p����U�Ț�����e��%�M�M�U{���>\�6Q׻R5p�|�n��{.����o\��g�<����w>i����:�)R�@�.��ȴH�v�+�_d�XH�|�	�4Db\�X�	SlƖZ��u U�dFS:vSag��"?��QS��"�Ӛ�И�7�?GC��i4>�����C��^EM��p���^�\�-������s8����5�Ȅ���y��i0u�j������:��ˊ�	��Y�' �����FG0XM��MR����Kb���汙 H@�.�΢Q���DG�<��ٽ3`׎ݨ����Ą�b����� ��舩��TX�� �tk0�LM��Tj%V:�P����hLCfFe���AyJSv% hj�<5r�rT��d��EH����
��\ж�w=�<4�� w�B�j��Ǡ�|@L*%�a;u��û��x�ů>�$�_�p�����*1�C�Ųhd�	�
�X$�D"��45$	�z2S�m��[�?�����﫦F��5���A����vbE��A�jj��MM��Q��6 UZtUhPS��`-�D��}�����������y��AY�������M���Z�U�o/�U(��k���&�Y@�J8r*������D�.-��'h��e�(������*��ss�r���܎��k�^��{��G����{^{������V*�̖쟨n�9q�����_h�z��ly�x^ewnEWfɱ��=<]�Ԗ�Nt�Sˬ�Վ�Z[F�1�@��Iub�L	j	������d�mװpqRz�Q\d����b���*��*,�J��+�c!+!�s�I��$qu����-23
��'3^�������j�;��x�S�0�pe��̂��Y��� ��x�P~�Z����g�W�]?�rr6��ҁw_������?�|�����>�7�_|����[7�n�(���57��o]sݼ�y�u�J��+Uאm���� �}�Jɥ�U��5^8���b��X�PWM���C��u��|KQ��$]]bUY��va��{��;hCL;8��rk
yo�@�H*�h
�-�8��mO�=��, �i =>��?�1��M�L��f�si4�d�x��8�E����{\A��'X���q^��5H����03䀒�" $@�QN�7f�����`w�=M�X��^P�n�����m�����c_�0/���ThjN����8)%.�p��9n�</lg9Q3�H����E!vu9���q���h�^����x���g �S	����D��ɂ�,	�dj�d*Y%Ϋ8Z A�Rt"C&h��`)��^f=8�r5)S�C��/����$�j���,����@�h��*|�`vᥞP����������zV��.W z��=�2Hw��0l�|o
�o
o�������55P���?Y�W!�6�@5�~#<����4��6���8��$�f�� �f����ト�Y<���@L�Ȑ�a����?�`j����_����-hd 15#G���&:kg��Ox 5'=+ce��]s��Y�E��3L �P��8U����M @1(MP!��2ŏ�550��s�+���W��C�2��+���:p��Y�5k�0~�J�e��� M*k6:�k-�P�,#5_e ���3���25`d�|߰Xf�%ߐq����2��AF]��Lt1�.-�����?nl�i ��@M���Y�4�>�55H@M��?O���d(���l�=go��� �S��p��L��3�G�z�)L)IԹ��4Mm��1Gߒ�oȐ!c.�LM]�_@Nm< ��L�"]>����U{� ��i8Zdjw��K⏸��$,I�[��\V�P]�ش�~W}�Du�bE߅��{�O�}��_�����������1e����EjϐjLZ�*� �0����8v��V`%�[�fl�)�O����է0a7:���E������3��(k��Ԍ4�6�:cа@�a�3�@���A �� �]�4���Z  �\�W8�-����~��g���=9Z��t=�15���gm��MbjL�e?�ÉƆ�E�j�($�151���"e�Df��\&��XM�"Ci$R�D
:���`@�f��.�ΠQ�$���n?2CmH��ؽs׮;۷n{�g��?�?ߵ�������%�( ����&���k?��Oyz\�6�m��M8(k��،/�}M�3�Ԁ�U6�a5��ې��������l1 �ZY��9C�jj�bjB�?�{ۖm�=�s���w@S�hdMxpH�w���k�w�'��Mr�N,̾�����{o�p���k�/�Y��*rYDl�J�HX��/���<��dR�T�����՘�����@����c���fF��VdD�d���j��D45M�H�|�Zs�h= +��
�`445h��[�jc�'}F�S���fؤ�1h�_���
ߐ����.�w�r��DHLM���@�k��dt�Jd��R�Aj�J�zy��\���TT1���FK�&ʚǋ�:3K���G��^~�����W����Ͽ����'��u��������<�'�t�}e��{�h[��w�աs����Գ������嶩��W ��ϵ��?6]�ؑ�n��:��T�֤V��B�C����F>9^��6K���b��m�Z�vV����c"�s*�剼�^]��>YT�(@bǰ<#=��L��LFNEKQC_k�lo͂�ti������K�
._p^�(�z���e��+���ȗ;W
���o_ξ���<��r������w��k}�E@��;��o�߹����7J��(�}���5���U�ͫ�nTܸ^v�Z��k�W�n\+�~�u�rɥ��֟;�|r�yf�n�������5�eiy���e1�&����D{���思�/��/��7��7��?�q8��jhj:2� ��O:�3k5�����!�Ɠ�K�N��fӅY��l��lŹd��D�����\Ø��&%�	1l��D�;#'@��Qf\��Y ���)�����D�Sr�53�a���t݋��{	�6�U{����c��0Ϊhg��SJ�I�Ɯ��V�T�XV���㬞	� �ϙ��-�s6�Y;ﴝw*����-'�G�":�&^I��Ȑϓ���gf�Ȃ���k_���a�k�fU ų6|iCPA�oEV��@�
ġx#kF�4��2Yg��5��4*k� w���>n&]Ȱ�4A��Bs�L� �(kz�䨬�.��p"�45 ��;����Ԡ���3�ldj��Uঈ��UC�h��A5 ��c���@�l~�<�rGA5�*�����M�^���U���Z��#;�ƟS�cj �vT֬������O?��O����?�滯>���������4Ot���7���/��>�� ����4����*�$M�F��sw�ݙ��B�{�MUAQTPT����Sx[x���#����ȶ�NO���������~��������;{߬B�,PK�=;���g�DFFD&�2#��͈�Ѥ��č����SCW3tȄ5K�Ij�v[O���4��15����J!�R�g��55�"^3�m��)�B&�V!���vH�_;��ĺ��L���jMİ0�K��2/bjf�(�rڲ�M��5͢�H��e�F��HSC|�/ ù��0������u�Z�v�-)C�� D�@ϊ]����(F �5YC4M_�O�` K8���%��S�)~�@�oW�wS�{��-�g[-)H���Yl,Yh),ϮL�T+�3Å���%	�%J�2�oU��҇Zn&ڃ�TQ�#�4�� �8��4��kM��洀�4IK��)=�13�1;�>/�� �\�_RZYP�T�4ZоX4p�b���_��ߛ��X�����;	�;����m�i�\��7@*����<���]�d��2�T��Jf�!�M�f5q���M^��_Yx�������M�o*�f���2I�nF�,LG�LU�&���|̓Z�A�۝V�佋t� ����9�ޚԂ|<��h /�
Q�`B[֜Sӕ+�I񁷠x�c��������E��:hj�u��P�
������[���B��v��N.�l7wx����
y>�>���/��7ϓ�qwusqrvuv��������#c#C��!�fj^���?��+���]��R_?)|R]R�S��S|-���V��7ϒX�����,��ɓ����9���-�3SC�j�v�����4���x�	��O5q�8��t��q�QX±e��]9�̫��|��o���TX15(n�ԐIj�\�d�o`mnaef"������>��}������X-��f�:Y�9�Y�;;�ݜ�lۃ������mkk�65G15�_�;[��l�h?��@x�Δ9eI�ȷN��P�T팦~E����Xs:�PC��I��z&�h&�&�'�MNc���qHM�/�8��Q���q��� ��C���V�mj(�j�Nu`MF@F4?*�+D�WDFe����K��C�3�ku����4οӶ�~����+o��ݭ���j�h_۟y����Ͽ���y��?��৓��o�y�x�^��v���^8�^{�t�^���@�Ǖ���W�]�i�����ݖ��������������Ճ�%��Eq�y�2H"	}��]-l����<�%�hjrd�y2�|�KQt|GSG��ExD�
#Y%ќ�(Nq;?�-]���%q����UdT5U�̍d/�T�d��Lٹ��{+io;y�v��;i��T,��^�έ�{�Y��f��>: Rvo*6W�o������-y���{:��}p���ajT��r��ߣ�m����Tw����;y{w
��,��^��T�0Q2ܝ�Q�W[��
QF�ý2"����B�*ԫV�j
a5�]����hj��J�V����H��Vw�{o<E_����}0�}(�}L����PxLŲf�8�	�k)���~�J���N��F��� ��9_`Vh�y?�E�3 ���C��]̄���4��4TĺB�5?��A��a^�b}�N?�A�~4Gξ̺-�%q��r]��� l���Ď���U��z��f�˖��.q�4�7�=n�Y��Go��o�=�BX�CYa�k��+�ע�k1�k��%o#�g-���&XTQ,�SP�rdP1�Ԩ5K0��Q0yGꄲ's��L�p��u�T�	�g�����4�2�̔�e�=���+��Ŧ&��?:�!#��LӁL(Pe���d�ga��5hj�96[���-�.�2x.�ag�S3TM	��|AC��8 5�.kp���}-S���g7�����m�;^��d������g?��?��/���?��?�ѓ{w����z+��K��Ɓ���ɼ�bj��)^|�'��!<�34 �JLi���Q�AϢ�˚<zX�!�M.��8�MA&�V!��/kjp�+�g��w�T���)�d�68�0@&���<�����|�hQ-"15t��A��+S���h��s!0��=�O35�Z��S*^��k��Q@�7
m�ڠ��M�	��X� YP̗���T�p�h(տ?^��Y/s�t��Z�ǈǊ���r���G*��Ң�d>�I��H��(AQ�_A�wQ4�"�_�CMb��E��F8��;�9�C @ �ʣ\�c���Ƴ:����7��M�"b�1EԐМ!o�
m̉��O�-RU��%Y������i��V�һ]�����ʍ��&ދ��N���;�X���{ǈ�rY�_���d��<T2�4�m��J%�̔[f�(GCBiȟ͋#������ 5�p51��4�˚�S�����[Y �س0���Y��x��N4����N߲�{qm�#'�4$�l	������B�5�i15�ui��(vb���m�a�k�w�T�ZzM�!������USjRaH��I�1�g�{xs<�\o�7������,W7(���Bqut ���6��3
So�'��YyZ���˚I�Ͽy��W_{����_<gmx�m�/���ڧ��:PK��Qk?Q	Z�X&�L�dVY*��O�4��آ�)�qCY�r�;����~�hH��%���=�cYU
���yV+}*b��!\��mch�s�ʙW/����|M#h�Wd�Y���up�KSð`�P_�w�}��'��������������9�.���Pa5l7���p�l6.�d���W������ۙ�YV���	N�R�l�K�ܱ������:�����QXy���dj\���� :����A��������Lu��=�ceU�x�����25�����`o�T�[&k�.J��(�Q�i�9%5�U���˕}׫��O�O�K��1����U��n�ƻ��D�L-�i�y�����?������~�����w"7����O���|���{��������@5��2q'cj/g�0{� cl;�o#�3�o#�g-�oM=�Q4p-�s�r`���_UP�HH	�H�H�B�I�R�&[�#g��]B\ա�x�pg���(��(45�Tߥ�wϔ9%ڣ����䖧׌��/�-L��O�n�^_O�sS�w;~�N�ݝ�������{wU��w�3��(�ѡ��^�[��≮��pc3��V��n�������LY��f?8��(M�z@i�C8t�}�0��A��{��ô�������w����t�  ��IDATڨ�X�Z�,�)�˫�ON�ą�C8��9Gª���huo
u�u������S��)���b]��K���y�{O�З@џ�1�1����H�L(ٓ���8�l��b���T��4��$��I�ۉ~[q��H����lg��s2��`W 3��@�	��B��?`?.�E� ��A�s��!ԇH�a��H�~��a��~�߃��ថ	���ۆ�e-�i%���y9�q)�aQl[�ݐ�_e����\W�. $`Z�
c6�X��+��H�r��R$k9���u-����_O��|���.e���;�u���t��d����/�ЛL��{"M3����I4���2f�$D�S��(Ǯ��]����ж uBz�ڠ:�(�<^��բ-k �ļ�#�ɹ�<^\$�2ڜdj�Y2��SE��gP/C�Y�Jj�n���ȸ�15���^���'����?~������ŏpxgke�s��j��dq�|m�l}��9��b,mm5M2����8�eM��' 5�b3��Ӌ�W��!'%�`�}гh󲦆�3 U�:��.z�)�}��8��:$�a5�15�rY����5�P����!�X)� ��|q1��]�$�2I�s!P���Ohj��� b0�-�b��$��X���`��<��<��A��yA0�!k(_�q4T@M6�F�D@_2H�7�8���[��uR��@�<?�:E�P~�Te�TU�@IzcF�:NV��)��΋��	��`X��U�q�m�2ƽ"ڭ<ʕ�����Hbj(�s��iH�M�i�����3e�!u��ي��������|UnI^uGN�ha�j��������}�;�^B�݄��������W���|Y�,8D ���qRe���.��v��6�!69a69rjV�<�5��_��������ђ.���o�5$���K���W5&�FQ�@�9m&��Si�k����F�P��?��;�s��f칡.��F���W��A���tYsZLM��1ï(�3��ނ25��5�?�^�J�����o��g���KS3� 
gvsr<\\==X<O//.l�l�����l,,��̡
�آ�q�w �����9�F�ʑйp�x�ܙ�^�[�~���:�ƫ��Y�_�����G�R](S#������j�n�E��&[z$k`�5�!v�-
����AY�A4$��i�F��:/ij���>p��ı�Ư���*�k�
��㵟X�F�:�t�|����y啳����44����\��@��&�����f�nH����q�4����;�>��矾��$�,�e��;;���pqd�:yz�s=�p�WWW;;;+����<5���45�x1ejrC�
�(����('��l0�P�����c�	�4�G�%|b4>
�K���ܪ���F���!�$��6/�i����UsǊ�#�|��Je��ʼ�����겚�����➅�ލ���ԣ��w3�}7��w�>��[1�0|dWڳ.nY�YM_8(��ޣ�����������־�������~�̞l`S>�>���� �և�?J[y���H��(}�q�ң��{q�;��-�������������������k�m�%��mé%5�	)Ұ��PiD�4&T���$�W�͖{懰B�
��j��0���p�dM$�0ʽ8
�M�����\9�U]��E!c�	�թU������ɂ[�����܈�ێۿ��t��r��4�����xx���'ُ�߾�vp�~��·��{x/�p?��]H ����(S����4��R��)�;�
�9��:<$�n��=���z�V��Z��|��D�Xw^{UnUVR�8!�#Y�ʉ�.唆rj#��CY�aM��a���N���
�F�Ss������FO"[�� ����x���=����{�'r�yג|6�|o$���U��r�p�J��B8k1�@b.�}F�:)ur ��a�?�2%s�F�`Š0���nDr�ib�X���yK�ۉ�'�oEy�8���,sY�:/��;�ɜf���]q]s��Z
u`wA�B2W#�1^�ўkQH_�b�Ds��x�(<��gQ鵘轒�_M����f�-g�-��}4'#5�����;�/�"`R�1/�]�`PS$�-f:�D�`2��04�s�)�650�%	v���*�4P�{��� �Ao2U!������X�!kHC&C��fj r.,�3�(�ej�qHPa5$�f���+�����i�{��������S�Y%�ſ~��OS������ſ��?����\_^o�﫚�)],_� J6'
�O�S�6�h4M��p��P��15��v��7ejZ��Ubj�x^�) F�/��ߔ�A�
�R�M�rl`䐺l�8��x�*�k ���/S3��?��b&p}(`�@���uj�p�HLɚ��%u�\,Y)���|�OӚ�'@v!�40���XfJ�Y��2��Ԅ�@v!���4SC�h
i�2X�!h �5O�x�[:��<
M��ȚcM��f(Ǐ���t��l�XF`��%�U+q*p*�z6�I&J�7��7z�&j�;����SB�C��2��PVN�[Q�Rɭ��^تb�*�����.��%����`�|8��)�����^�%_#�O*�}4�Ư9Mܔ*jH��K�kL�ԦU�J����2㊳S�2ӓӳ��2��3'r���w2��$��fM�K�Y2���5�H��CBBB�A��RNz�G��9Cn�b�n�i�r��j�S9��Uƹ�E6�p��T��t�����a_��`B�@�/�|s#/oD�0@�B�!�0��PF�t$�ac��._��׆t�؅CW��>v��
��T���15hj�e�i15Ce�lqI�w��Mʱr7�jv弑Υ+�/^�H} �15FzW�t/���<5t킓
�����xz�`����bggoiicffkn	2g[[++8jillnhhx��i�_��{�"p��gϞ{�7�E��t��딩1��fq���4��&Y�
rT�P5"��@� ��@�d�Yv�5��� MM���LME�쒏���h��45�c������"�McjXu���$�r�O����sd[��L.��y��o�J���ƛȅ3g�^�ljh�-쬬�^&�������qp������w����?x�������훫K�hj�������#�͙�v��D����Ҙ�C�G�{��g�eg�#��+E�R��pu$��-�q���"kHl����5�>��~:Q���������A�A�тs�M��$lq�x�js��!nm�Ҧf\�=V�*���V����Ա���֞����ł��̑��3�3g�K�y/j������L�:�V��Ð������������Gk������<�?������w?���8�M1p3h�V��n��ه�󏓗�NY~'a�q��A��^����~.�q>�y>�u1�g5cx+{d+�oYYۗTӥ(������~A2QH�0>�7I�쭒{f�p��Xan�GOԤl��`���.�QTd�:��I
�G�养@��a�9�fǖ�W�ݸ�z�z��d��Fƍ���[��ʽ�	w�LM���@�;o��<~����)���V|�i�ǟ�~�I�{O��<<�}t�h`��G}�DM��$��n�ݻ���0�޽�{�s��+8<(��Q��,^_*]���.j�j)�,MU%��C<T���(�pNy8�.�[�n�hw�4M�CC�C�©)޹%ޥ=�?kbh��D�H��'��X��%�25	��O`Zɡ�c/*���Wy�]��&��F��@��lk*�m2��Pvg�=���1q�; ��w���Q�Q�@V�9�
��8�	���Hl�r!�W"YK�����!.��t"=�X�R4�����������Y�a����YH���{�'r瓼�S}U��t�r֑�Y�>��i�Al�Q��T�h��(��`�1']�P�G˭�5�) 1)� ��@s"����)�fH�i����84 �"P0A
$�:�,������H�.d�(!剩AkC�����A&�Ŋ9^��2P���" -P�f��[45epv��y>Xe�Ա����>u'Oo2N�S��(GC��A��F���45?�����ƻ����٘,}��!��ajVc_���W�&��+h��VL��t������g��/jj���A��(�@��쒟�`y<�i�P4ǋscaH�TP��D�R�D�̗�`���*����Ed�4hj�K����!��Z�uq1�x���� ����H�B4,ڠs��B45 &f��_����!0��j���S3�-�O�d��rdY��ߖ0VM�#ej�ܖ����w�G/�.����%֦G��R���@�,95Qb��/l�VKq��AY�D֜fjp5(���7��T�����DiqjD�J������SZ�V֒Rџ\?�и߼��q+ch�d���F��7y��<}�B�Ae7Y�ʐ��X93�!+�67Ү0�1/�M��!*��/��iJ㵤�;r|�SC��f0Pt��J"8P�|)(n �4��`��<�I�R�����%c]5v���� �K�+?�0L盚Ѳ���ж��R%��S�s�.蜻p�����CݫF�:�W/�X��Z�[ 6���6��&��b��4����渺�988�ں�ٹ��C�Sckn�|Sct�����ޥK��ŋ:�Ν'my���7.��Ի�f���b��N�w�L��6�ߊ��� �4�e�̖�H������ (h��9v�\ ��6/Sw}e�2�C�j�<�p�����u
dY{X������ޠj���ӹbij�g{��YY�s�wd����,PT\���ۏ������G��skkui>7S���hef��`�ru�,��!���x<OOOT3DּxL���oۛ^yX��8(E�2x�G���7mJ�|����Dk&er���{o�M���K��Mbjr?���`o[�^��0���X_�`p��+�z�y�}ݞ/j)
�/UV�e�4���Ne��&�̽=�į��t�}��;�cO�c�%�oɧ��L=�| ޏ��1���ѿV�����g��+'�W?��o����M܋�z1q?r�^��A��A����g;��fh�n��ø��������������������������FYR?8�W*�����'����y��^hj
BYEa�T(M�=���;kd�[A�KQ$���_ܪE.١.���P���%)5L�P<��ֿs+wj�xu�p�VҭM�΍��[���S4!03<P��~��N���|���ض���m_��㋟V|�}�[�{�ُ�Y���Z R�ށ֐��;��{i{��w���߻�>�_zxP|��zc�xi�tv�r����!�� �@��(Ju��(��.��TDr�c�"X�nS������Ԭtn�wk�;�4hjH�L_�D��������j�8SI^���J���}8�uB��C�h��T,����]H�^L���Z/)�!XrR�1㎌F��D8#��(3����t_�f-�z��{�'�$�eP[]�Fq���w)� ŋ'��kq�S����ZܽP��]?���ɿ�d&�>{]���>p`4!YZ�o��g� 0��o�=˒�����8D�I��3�U�tj\�3����/�$��4I���#���d���ҍ�B����:�.�΁�In`��؏��&
�=�>`)Q�A��6��1��SD�� ⦶l���nU;ے$f���x@ 6�oɜ��As�	;�3o�wph�h����!�
X����%8��)2}�1��vH���)^V�`]. @�|�hf@�8��γ�k��H�hf~�,{F�\}���{����:5� ��:��g��f��$̆� �_l�d�ҠZ`�R#��qB�~�������������!6�f�V��՞3$DA�R�c��k@-ѻI����.,��@��D��2;���E��Ta�@�Ou�U�����:?�V\{KV�qn=�:}>�4����DԈ�IL �I�<�37��F�:�����cĦ�r.�ԏ�V��Q�C�:�,�B#�L+��;ϲI�Д���:�o��N��ʳS���#�%F/���D�xZ�* �$��~g��g��̓$�2Qzf���ؼҧ�0y���\8�0��1��|��]
|�^�`�jk��}�V>��==��Hg��'9�灡0��e�8\�knР~��Х�:Ao9]w.��ن�m���7�d���)��'A״Oj���zO�VL���0�z���]M�T%�	(8��SATh�O�S�%��r/����^�z�jIRc����Q��F��b@��j��j,����5^�z�Pw���t��)�!3V���Z������i�?���8�����k��*�)���*� ���.��{�O7�G��H��D8�����3�
���eE�d9��\E4�`�3�b~N�'�{�wg���8�������B���]�ii�f��PU���K��C�DQ�1qC�21��n�h�Gu~�ٶ����uwr�����Q/����)����Z
X.����ʼ���CF"��R�������w�7��U��eRv����<��ttLXת�*acZjJ���WS�;��XUT�����䛬��.��3t�D�=��ͻ���V�oX�Ƴ�\n�Y�V9۾��nDtd� ��2�).@Q-�,司��R��g�%�(*'��n�̬�(�_?����#U�T��*#EG񞍿H�O��!����Zq�]�h<�E��#U��̡����{=�]f�<33P�O,���7O�26ݜC_i�!��xs�5��B���)F�Ӯw�E%M-����T@�v���`��ݓ����h��g���N�JJJ���)))�s��/V%���^��j�v����B�G���_�X���6��4�LI�2h\��̑S%kg>(�5�}և#�BG�,B�5K�P]��6�=�k)�F�k=$I��h��5di%:�h	Zj�cpG��ƈ K�&�L���I�*��	�C��~��������%�M,�y��	�E6ܴ]��|�4�
���
|�j�k���gյf�pf�4�50�8�ޟ�����N��з�M�'�{��}T7)3�����O�SF@t�����&¿i�O�ep�BO������Ģ�bywFݻ�~ҏ�Ց2l�_�Iެm��2g�����=m�R��4м<:b�\^X��
�M��Z�Y����Ik���a��a��U�=5v����g�$g�:���o���4�S�r��Y#n��\oo��X�d`����_%�Ƕ�eo����d'0����up�h�fo{@��|�O�lNPʱ��w7���{����鈨����W������b���3��r��&�+�����[�jZ��h�_�.Ǝg�Kږ���ʲ�������=Y#����yz�<A��Xr�6����վ����Vz��'3/d�4�Z�k�!���W���q7q�Hw��@<n�<XbP����y������	m��ְjLz�(zO��p�t��x��I~H�6^l� ������CV�?����lQ ����'���ɊMr��20����b���y."�%�)�$�@��m��g�d��t�`�x��ퟆ!4�w9Y���zרE�3�π�./B,u�.L�Ko��")L��rt�4�Z6��,�^ ���>z�C:����W�x�f$S����I�+[6����{��a�]�9��EUȟr�`��ƁiD�x��'��c��_��E@'�I8D���c��d�<p(7�~2.Ë���_����:��X��t{eȡl��� �$3x�����^�'��_��_�	^����(<_�=���o�__X�Vq�A�o��Y�>슾�=��4e�p;z�9v�lDV�Ϋ{�B�K�t��|�+(��L{#�st��0�hK�M��Q���&)��C�x7����UGqT�� ?(ǜ:yzq�p$\,���:��j�[$��{i_l�RZ�:{1{0Q�1;�|a J拙6�`
\toP�;X��8M� ���3ҨjP�߃$�0I�l���j�mC�ېƩ���=�PU:/���Y�E���L�}�eD?O���F.��
���Tİ��W�|>5���R�C&�xi���Y횾�i^���sV��½���5P!o<˴\jj�j�9��Q���+�Qdϱ�B'�u������4H��; �:8��]�!L.f_��YG=�T��&(��,��v��|S�Ttw��Է|��p��~f���n,�ngҿ@?�N�I��C�$�$`��-;�-�i�R*6pkTth���/��$�{5�F�~���� ����TU'�� ?)�љ8�5��O�:�I��NiVXð����S���7�u�f���s�T "��:��l,nr4���)����6���C�h����J/�/��]H���;��:f8#�w����U�o�ẗ�胁r����~bFbmK-ƿ�幩��k�n�)��>kw��m����\r:��=;-Θ��U�_Ͽ�����m�S[𱵍�����?&$vB?F߆�{ő������꿄��>\�E4��gxU�g�sU~[/�[5ܞ�&Ў'������}�KJ��� {��7�V�P D7��bv�0�%�ޖ������j�3Z-L���-��\�g�u��0�.���7G�����QG���i��k
a�A�E���;�~w�#QQ��U��oXn.��M��:����f���n�r���z�����`����B�tϬQg*����s�~EFFF[[[rrr:C؎��mL�yhK��G�:��V�A��=�j6  �U$|�a6�[���g:?�܊ ��A��=AnU�����pR:�Ӏ�z񍏦���2H����+��Bs0�S��7��G�!ʪ{<�[<��dl9�۟/�2.�5��,T뛫
�-`!�;�ך��D[gn�zGW�:c¤���)R���G�'�9g��W_�Sq�ǆ�mK�~7�[%�q�?>�d�������h��(̥������iZN>,�|˿�`���;��:��e׏�v�cG*���S|��4ԃ@��J$=����E��Et�C��J|�pk�Z\���qMr��*��g@~�Z�����������+�m�Gj���E�ߞ�{KW���;4�����J���kPm�X��D��̓*JV���d8{��u�� ;��=��ҟv�ݭ�5)Sl		I
J �/�ȗw�u$6��+�:&:΀�SsT-v�+t4�5�5���d�g����+��F������f��-��X�W�X�Y�|�hP��D��I7�Z�2-u,K�������N��(�m�!P�py��<������2�Z�f&H��>ʯe8}✇%<������;�#n͹�i1�0|6��>�Q{�d����MCk�Gw7f�C$�5Sd�5}g��7��@n�C�a|}W��s����֖$�	�i�!��{��ǐ�;��6�;f�E����y�������AQ<^��I��^P�E�v�&�T���4}H�i�a��bI]���,� ���7� ����c,bu3�m���?N��Q'����	�LI�q��@y���PEĚ�K�>!ɿ}K�"[�+ߘR������=_9�<��
���;3��K�bg���
�م���H�r��t�Aw�E_�O���_��ڔwQv�Pm	QK5�m��O�J�u�6�P�|�.Z��u��V��h��3ú��'q�4��*�l x���4���2�q�$Q
Av�����`.�LN���!��n�\$�$��Ӽ,������l^�۬N�K1(M0*E�f-$��]�@�Y�	2�c���Mb��uԋ9]��lPx��4"��ZcW~��`�g¹U�qla��� �T �	��㕕��9j�8+�����2>I޺����1��R~]Hm��	�z੃��׏��M����3�2����{����r�ϰ��j�`=�ӹ�K>��<a���M}%���I��x7��
�kY暤�ua.%�xK��B	:���X0���"���$;�{����g�d}I�����v<7�'�䔤t�4�D�r��h�$ {��Ֆ\�&�o<EV���B�{d�QQ���Jޟ.�sPM���$#^ o�(�P`�[�#�HU~^��
��t����Bb��<�s�q.�Y��ֱ��뾩��2��8��';e�L�xٮ�hOe+�)�l�4���t�WL�^2/�Z���?���(w>A�%�bi�RdR����?��QDl��σ�7�k�,���rn����u1����w�,��`��en���҃Ǐ�w�-�U���x�jf��'Zl�4��o�Z���^�5�c�MId�ۭs��+�'ew󒻤R�ᆹ#�N��{VYc��0�H�y��t��(��V����%ߨJ��?�%v`&�H��&<5'���S���x�=R�D��^Oۿ��9ӳ��B��|��{O(�g����聝1�NG��[\�����|��c�t��.*���S?]��;92��$�llyw�0QQ�1�{yy}����HK#&%Ͷ������0�����V���	�F�7UT��4v�h�D��!!i�b"%F��w����p�ЀG�6�I@���������ǭ� �#%�s(-�J������0��/��fS�2Y�NiYO5�q��F83�NT,8 �	�ywVå�6�8z<pa;~n?�U2��m!���pq�v��w���� ���-z~�s��ș�j2�����HM��E&�'�0:�7ө@�������G��(�h�����e�������Y��m��ˡ�Y��ݙ?�'ц¦c�,)�O�oV��W��b�(�+�U濂j������1��S�H����Ak��VK��~���~�WĉꚶÁI3Տ$p��V��;��{�c���(�_΋е l��?%�禱f���U�f�=�ض�㟄��1��Ή��S�O��M�ף�K��_ei����������r���	X�|'kKPp(C/��c����R>`�+��Tiq����� K�ہ�ޞ����ڜVbe9{��h�����ҎrT�f2����ۼ:`g��Y���H��M��^������[W�l�z��?����:�hGc��Z�-�$�A�� ��� ��5��/j3�qN�P%S�.D%s�1knTb�k�>5!j�t'�!̾�����&l�eY������d^v��/�b�<��}��������ܳdi_��G�J<�HD�|�U�[ug��<���n�%�R8H�:��p��}�{��g��A)
7��'���2�;p)Rf|�h��l���s;��d�1��w����of��gF�{� 9��8����Ok����o�X�k�����|��Vul�����AY`=qp����v�sԲ]0#����D]f=�t�ow��Ǯ�^�/T�EҲ�\;�_��/|���UR���ؤ��f0�J�xK화6�.0�ũ�ߗ�c�l}�`>{P�D��X�z���K�����@c��M���pQDd�a�@��s�Ä��	o|0[K��n���k#�|���s�Ƥ��k�N�.�7e&D�n�ɐ�B��8"��IW"^ƚ����d@�eQ�%�*��q�J�/정��{w�0��׋�I	�k�7�<R9��t��`�XL�I���ֈu^�i�,E��^ĕ�h��Q�\�c�`��C�'�*��GG@��>w�3L���+�@@
���Ff� �j�T�tՄY�(R��3A*iz��Z�)��фen�����m���;�����Cu?��������y���F~��h$5��<#ť���6��=�̭�����&�,�.�o?��s�xr�iM�UI 
"��5^eB��1&�F~W��K[8�G�����o���� 4�E<��o���U9�+􃃌vS�j����°����h��uBB��N��F�OWw�Hٿ4���Q�,{��_����|�d���������O�~+��?>Q��O{��F����7��8^��4:9��D��
�fE��i1-s�=;��dM-�rўC�q�tr,�P��(�p�����VLe�׏���,Nt�t��s�ӛ6`��6�wy�������גb#+�� � �l�0T�`�S?�ׄRS&������Ş=)p��˷*�F��{I.�B�~RP�V�t�v�8$�&<�+��ݛ�S]I�}Za\}��9m}�2��Y�����z�ȃ�4}F�\�W���5��������fff>>ϻi�Q�&���|>#��k�gr�(�廀įcc	-�k:�.x�� 8!&�ͥu�ذ_=���EK��U-xMN��MWk��i|c40���Č	Yֵ&��;��C꜎7�Ch%x�ã�#�´7��}�	��{`�j��Q��+���-z�:Sz���t�{vD���ZN��$���{Ť�o��pzE�ݖ,tm����}���i"y[Qwmu��V�<�~/pFUv�Y�����i��ǣ��?
�G%��O��w������u=��XKzl��{�x��1S	��a$=��;�s"-R����;7$>�@�zn�������3S�[���ZcR�g�@�y�]�RjR�R�c�j�֟F|�fB�j��#����~E.w�_{N����^��$Ѻ�^�w�jS�f�rc{z+W��ůsףK��t��'T:2���ɪ3�{R�5S7+*����j����\g�3`|j�|��x��q�
����L�s^��������p��Ɇ4D�4�^�l嵆=a��PO�Un!`}U.�t���W����M:5'�$
�&��
�~���Sp攊�7���
�����9+�:�D�[��
>FM���t~"AZ+��&L$1S��4g�ۙ����B�.{����nɲ��6��I�5!�R�9��!�Αc�C�8��)iׄk�Fc�M����o�՜,��M��,0Ǌ:�\����g�x
�9D�k�&�y3<�N󏁐�(���>�}]W�b&!Hb�8>	�K��޳�,	|�Yr����ަ�V֐'	�t(�C-+h	va�cs֐�����74�S"�[{�`��)�y����k�tbK]a�}5�����S|�S��e`˯\���ň ��|,���Y��d�FL��ƛ�BP��-$�����p��]8��`ZH<�K�����\9���;��Α{[�*Z)B�E�Z�]��f�,�d1"n���:�4?t�JQ�H�-X��t��}�ڇ}�4�W.-(���bK�����ԎB˫�@�2)&A�z$%��Ĉ�"�P]�c�> �/��(�<M��B�����i��Y+ů���.V��Ǳ�~K���.Q��=����W�ahP�� �_�+}b>)�����XJ���'�V�Xƪ��r��*�	 ���L*��L�M��-(Zq�����dY[?4d�7f�D�@ⵐ;�ݞ�Y���
N��@"��칝\o���-�T�x��}�]3Y�:v���5Q�i�&d��V@߱��6�^�/P�E�;�N��Y�ɟus�����ć�� �P� ��� �8�ԃ��ڀ�*79l��@�S�wnk�:��,��-�_�3��L�$3,�u�`.]�2A�ŋ��3ҁ����a�+����F���mE��*����>Z�������+��5��b6���(�Ų��2����I4��Z��Y�M�v�-��r{���79m��5�9>����q87�m�2���?s
���o�w�=�&I޵�t�������7������<�ea6�R�^G]W�����rϵ�~���_��a5՚~�|i�14VƍP\Ejj[��&�,:��)	���^L�}�� �F�[�CNK��m�t�꧊�*9�E:��l�+HD���Ȉ�T���a���������K���G\-��W�3�1m��^�N�7�m���S���t���W4X���kW(�)�+����}ɝX^&W��rn��n�ð��q~�[�֫|�Y̓����p��cb�h5l�/0JηY[�3Σ�+��s�/D�Ƚ^��<�g0W�Fj��Ok��#hMu4��.����I�t�����H 8G���{���2���$'{�����3IǩD���&eel�e���2K�կ�mD<w�s>ʋ�T��I8K$�����D�	���I e��U�O~��/��C�}7�>ٜ:�.�u���>�'���-բ�t9lq�&��G.��&?������k)�i*{��=+롣�a"a�U���H����Υ���2"�Π�N���E���׊��t�����)�K�+s�3k�;��q*��!��� ��ì�	�\Y�dl3��5�mn��V�@��9�e�V-��V	��X�|����h����?�G&TMTԧyI.�9�����F����`���<�T����9\�y�JG:�U��vX����3���m����'ӧ%�8N�TN�~.|ѩ_�s�����,�L/�ϫi$�&i'&��=$3��f$��2�	@<x�:m䅦 m��9�z�&1�p��C�t��;6������I7��kC�������
jd����w�T�.#+�ę} ��Yх���h�DH�4H����eu���o��q~����_tOG�шjy�49��S��$�WUϵ�$x�i8��>�Ź�ӷ$9/���3��ӧ;#gBTȘ$ ��P<�Ѵ��2��='ԃ͛����\1?�N!0��~�0ꚙȷ���]4���$I ��¿�b�x���)[(F#��Zܬs�s?��q����vZx����lS0R"	Q������h��(ֲ>1�nB��A��b�Ǭ��G��`f���ީ���a���D��^h<C�PbU~�-�5�.]k	�T�]>d�W�ֵS�vD�8��+�_/�㺵&��Ox~n�6yEcx{_�V�l�9'���ɿ=Ŀ��&��A�z{qe|�wp�'@	���j(m�Z1�.�:K5[�K.|��X�F�����9�ɫNk6Z'~��}4����S��U=⧧�
����7��������7�V��������	`ɂ$�	C�t��)�����g�i��f@�R!��t|��u ����̌���y�şms�]�M�d�KJf���?��)C(Z�m΃��Ὦ_<���p�Q<[z#ҿW��(}�o�[l�_,�_�+wb��7{����JB��gf����ʇ���(� (CLlU��2�Zk�X����O#�����g�'],.��Zƀ-Fʁi�߱���ɋ�o9�<8���Y�ɗD�?�;`֤´ D�QSeK��͝�9^%�$-���/���_?�L#!�]^��?���E=N�
�O��������iة��F,P=��i�߰�le���AhUߥ1Խ���g� E�8V�����ϦH>E�xOJ�(�'�#!��\� ��3��[���?��� g���X�����/�����i� ���|�7�tѹLV�zEc�?}��@��!�+�2K�h�~��-�B��r�w��í!�c���o��b�{@��H�4{�u]4 9]��͙��Ⱄ����b�Q��h3V������hK�M��g�:|���]:}��p���qr�Rg!@vpp���d�$g+� PB���׎����;���78~��7�bv�ip��E�G8+3Up @H�H���OH���O�f�����-!�ς���l>T�
��ͤ&��ä�q6|��JzmK�E�g��g��_Vc�l������d���X��4B��thO%����!�ษcc��F��EW`��\������>�:z��FD�r����uz�.s�Zl��{Լ��B���~�XR���{8E�:��r2���-���k�$:X��(��,3�5�a5�~5X!]g/Y_
`C%J��P{"�I,��j��4xR�ϸ=��/���OGL�JIZ�t/�I�-=�Q�V9Bs�4c��+�,�{:�)_!淋��.I��v�~{�k�9���t�Yr����7���6H#l������5�����N���(����H7_"�hQZV8$#�P?��@��=��������R՞�Z�����		b�u� ژ0�8P�xa�ff+�˒���*�8(���v�#�b֊R�J����r6vE-F�$��d�s�~���)��s�s�b�࿊_	�g��<s��aa�1�L�8Ƥ���z�"�x�1�V}��;�[|�;͟�(�P��G�M]����}u}�jN'�?4��"�n�ڣ��\�{��
��`�w�����*!֐�n8��k���b�0��� ?~o4��B8���a�.��-�o�Z���у���Bf�S��!��#?@����G5Q�gT�Ĥd�\���Ϳ�Jp�^��3"l�}��B�W��Q/"���s�Ty0'f&�a����7\ܾ�CCTӼ.����%�c�,9PF<P�P�!)���[��f�±v�y�I��:��+�.z/z,��'D�/�E3[���6Hf���`#�}��Br�������7��E�(��3��@���j��5�W%��֒Q�-��������k�0Q��[3G#d�W�CɁQ���|9�Q�^aK���@�O#��"(b�!!/�1���Qbm%�$H�M��~b���,�;����3�� eF2�٭��b����=�q:�彻�4�k�+�����&�A�,X�mv�ۣ�T�����pv1P��D����:ӑ�t��UƽSK��]�x9~l�:!�K��X.� /00��Ĺ�mdf-���"�M!�H+��a.)���/9"e>�0�@XNt�ȵ�O~i��I�V?�S�W�uj�Gbk7�R�b�E�̨�+(~+�+����z�����<�/�Ê�Z#�U�=��[7�!ͳ�6�=��=�Ri�˭�@Μ*�As�.v����E�]hQ E��7&�ƣ�0ì��@e��9�ף����!��O�W]��J����I0T{��S=�V���{<���pO���A7�����G>�}:*/?*��d�ɳDG:���8���[9��2��y�����j����E]���dĹ��
���ͽI�+���{:�vv$6�@{���;B\�D��Ȭ�٩�3`N��GO��+7� ���7_5�`�������o��<Rf���y�v���3�Ps�`��D}�Pjh���O���l�[HLJ��gte�D��;�Y�齵���P�ձ�B�a��ε�#��������P���Xpds�k�5�&&��5�]%T's8�x�m˓�h��H��t0�Ԧݷ��:�r�QP�Q`!������W#�Ù}�X��;$vv���(jYT�,9�oe�Ad1Z�l5�zc *z��hDг.��EI)`ILw^�S��_��雫 �-#���,q�����sU[œ���XVdI+$8�T����c<OO�[�I�5�C���UsM������s�D�l������.�p#����U-6/�'=n�҄`�s_�웾��1�h���S��L{�ߕ��lr��
;'Qk�8���P���^WK�GY�I�/��z�^g�uz��l�����u�K� Y���Gq��6w:a��fG� �Y���3*��%V����r��s���lU����"�u)H?~����Vƺ��8V{��B�"��U	1���L4ʜ�2�5Z��2�-��ܳ�_�u��`
f�E�t�3 �zyz�S��� �Z̆�0�ݟM}zR:���I[�s��Z�In�%-�0P�.eB�BQ�7iK�����Қ���#��a|qW|�#|ed|�����x�45A;��V;xE;�V��E	2 A��?�EH�aI�PD"z�t�Z�������䁶�F^o8��{b�r�V]��"����nqi3,���v���,J������Jh?!�A��,�~� �"i�ɒ8Ҥe��sH�$pW+\	V	�we�\e
=�ٰ,���sĄx�J����^�-���Ǌ����L�m��'h��j���a.�^�XL��|�RB�����ߚ�$�T��a������j�6�Jl���Ў��������s�#L'�%��dI��m�b>p��2���� �=��6]�T���9ɧ��A. ���*�-쏇�~��	hE�
�R2�(d��Կ�bB��˽Δ$p�ў�	���=�
�.�]Y�m��N��(��ﮡ�	�r���"���FK�q�����Y-�ٌ�G��G��٢tS�ό���b4C��h�T���`:ǅ
�%}3e��enC@�c̬J��/
��А$�oU)����Cx�|�9���Y9"0}��	o ?����|@p	�������g�Ѣ��G==iFڐ�^�w4e'@�����5F���وE�-U�gQ}(<�S<�F����jF�zK���P�G�f���vJ�Y�G*�F+3�u$�n����p�`m[3�o�FmGĝg�ü�� '&�*��
Q��0f������H,���l(�/�ƗR�ێW�Z:q�xҸ��z��h��ۓJ��7��;H�}t�!����u�]��,�|<�>�� &Ik��רd�1�4���(*��>���G���A�	���	�eq#*�^�^��T��5e����V�Vu%��pI�;�̓����K��>��Ekw"�d&���8�7�->W|z� z��ea ��?��s��
����o�5���Y������:��ߗ�P���!��d��A���'c���|�-e�;Q�>x´����z�<?ȜQ�0P�l��Y���<β���?��7QPT��W�s�ma�w���R,=Os�>�*w������=<t�+���ڶ*`]������h)pdq5�1�a��Y��(&bX������'�qι&��A.3�}�3����ȧD��$�g��B�K��K�B�s;'����������,�l,��(��6�@����$vѶ����#��ȉ���f�����d��&�f�Ն��+\�ݲ���-�"�3
�³g��V�����Y>��Ύ���G$Y����ob�,�/⧤�[�5�ڜ����E��7<~�;4������rz�H��߰<���/Q��tS�̀���}æE��ł��2D �[��X��KO.N����u��E����q��) ������Rpme�C����,_Ǳ�/�߂���(����xrO�"p�RK�c1���u%?R��:P�,�8��k�.��_N�e�����d�Ȋ��Q��S�R��/�-4�7n���q����>�3�/>���%��AC$�ҏ�Ԉ{!F��D��5@~ʦ��0�<	�b��$��@��E>=���l�[i�z��0Ym�I��ǽ�dMtܯŸ3�������ܺ�l�5��Z�������yu9"�9�%�("�����y�5��B"T���G(�������;XJ |B�Pƈ|��m,�6�
�emR��G��`Gbb$3��.���h�ĩL=}>��#��v�~��u���F�
�%?�`>K��$T:�Z2��2ͯ�DI�7[��X�q�ү���0.qd�g3q��W����]�W]UI|�D��0����j�����糰���$��aw���d75�e�Aw���&#������q��h��d��h{ie��>��)��=��5��*��'�@�H�o��R��D��l�m�3�\��5]G�U��H�� k������;@�3�T�nt������VO��VV{4�&'ae�"	_}mm� (�3b����8z�+�'&̝��Xpoz%��?�p
c[q��ī����L[��t���o��
"�q�a�-�;�g^�\��x;�U;M?̲��+���A�@�nڎo+[�m���Z�V�����ܛW@�5�z�r�`�QU(_� �7�z鴦�P�(QHAU��jU�� <�I!�*1�+CA������H�ld�|�"$��D�@%��Y_Gݛ��	E5���D��`�q!�
r74&�5�8uHĐ��U�ũ{z��qW'�:�����WO+bM�~�*,֙�Ô�L�6�%l)V���; i��P�< �'h��-Cji���~*�ʢ }�,�x�V~�W�xp�{�i���N�ޏI�?(̍ �m�8�p�i��"Va���3?ؙ�̙�ՙ��Ӈ�Ƈ�ć�ׇ����͌ʲ�϶�ѻMл6մM�J jYh�[N��60il�aѳNak�U��1�tؾK�Y�-4d�
c�����mFsV��"��tOqO�a�Ј`yY��L35�������ȼɰA�5�����}�[���q.�;�Q�,�&�fm�l��cZ(p���БWɷ��ݦ�CWH}PL�S"�@��7L�N���,ȥ�E����\�����+L�gΟ�!slD�
�ؚHb��aU�<�tH3NN����ݦ�ƛ�ֿjtj��Q�Ǘ�0v��qt�}�~�P9*�>.�n�"�%��(���/�� #�ĉ�x��\��H��F�=	�H���~h��\L��V��=?��,�v�\u����.g7�a�+49k]�hn�@��H�Hq�����o��c�EC�2	pT�-*p@а�"s掺r�(����s�[���g�邋Je�b9���w�Q0v�ru����۫+@��\�K�M���olE�My��`??Qʦ�Ҹ� ���Bߌ�ƪ��}� VIPd�f�+Kf�Z�YV馾�j�|0%�d>ux�<��ߒ�������zN4A��9�8H�ɘ$t�D<�d��=����P	��(k�� ���ǿ�d��6��JH�__�Q�'���$�p6��ERa	���#+���d_���=��%w��L���DX�� 9�ai��tN:ݙ�a�#�#$�"$D��i�mH!|�%
�e�W�OI�p,��jL��������p�z�n��u��{�WQV�:��N悖�G���Wv��f��D�'�q6�}_�ؼ����>�Z�C�ƨ�;Ȭ�m�3�N����ʉs�)���J�TWi�^f��R{�\�ߤ�5�D�(�.M�6-�x��n�#"qG�z�T>T�-Q(�TT�O_����6����M���;Y��`  �AHi�T��f�~�"�!��3��r����a#8�[�]o�@�"����=d�������!F���I����F�x��fH��>���¼��+C=�La��^���v�β��5���|���5��	��&T:�!*݌���e�*�O��Xh,���L,��?m#C݁�1|g��G�l#�ll��B�_V��u�p�nv�����iDqrF�g]U�Y�����s����E!
����4�Vd���Gצ�x���Q����m�"�aBqꈃ��ùB����00r!Yjasd�,�8ڽ�
���<N���T�1����u���/\?�*u$1��u&�Χ�+(ܙ���Y������i�]�����*�2aǤ���?�@���5X�ٽW���ȗ �&�&z�\.�
�y
u��,
���݉���_�{�������Py�����[�T&E|���(̘Q�ô֕�s��k��(�j2'����Q�~^م�PH��P�l<5���/c������e�հ�51��/��/L��gW˝���q;��/�9'䪏��汥n��n�;�>�>B�#/[�mb����Ww�:�K�
�"q#���}k�s�&�Tt��Y���I63�Ag̪N߃ݥ2�-ʴ��|c��b�9�����ȉ�k+L�('����"\Y#]rON��\�R�4���	��h��C�Q#i�uSs�s%M���`��y>�s{���š��t�G��6T�[ʝe၅�-�;�ff��׺K.{*jFV;b2]b�o~f�zR_�,%M��j�đ0F��̼��?����N��/<\�ޛ��3	�������T�eP\]��'��<H`pKp����	���w�����y�s�ԩZ5U�o�U����]��V-�|,�L�����3���y���('����W���5ɲ�Bީɛ��Y���n�9��Z�������q�p�ӆ/r~��O�Ln�3����;�J7�3h���d�"��G�	��-�C����^1佽����8��Cţ
{]�I7��{�Ԩ\���ug���n��Ӵ�Q���������h�b ����8U�ɹ��jB8�����"`�̎�:"�N;��!�)!�x3J��i���¥|$8���M�nBty�~�����n�F�*r&O�?C���A'<�+�}g�������1��m8��OV���=�j�ޭ�H��Am�цN�ͷ�s�S��!?n�F��~�L��ɏh��l�XR�g���,Lzs2�ޖ.�.�@��}hF"~j�S������P��ɼ��e������m����54z�fg���3a'��uD]cD���J�%��*#:�b|���ܔ�� �)���Ջ�U28V�`,C�N1��`ӃC{" ���3���0�����8��n4�~5Px����y��#�1�?D��z�H�͜�D����$}{�o8��':Rm ���})9S���(�mTbʢ���������yЁu������X�X�NJj(�B�̭�U�^Q��<������J�f��fa��aNR�Ƌ/[���E��Js�J�/-��E���	X�]N5/�]�C�>{~�7��>/w[^,�+��V����'1]*A����~H��Cй�ݕ���:>O4��Km�Pl��C}��J^��*ơ�@V�1����
͡`΍��m���Y&KW���^��층���Xe��VX^X__��gPdg_a�Ω�����Rg�>&L*��cD��W*����:�A�؍�6@�����;�����w��-=���Uq�$���e&���+x�vPE�5�_x�3  L�f�I�c�e��ҿ��-)�X�X��?�۷�,����l�m�-!vF�#��	�-���L�F2$�(\��,�DrN���l��1��S#b�7�PF��Ɨ����׋z��i�痶�ǉ�صE�_��GKے�
FEiG{��N�n�0'�_�n��7�D���B��7���y�QH��z��U{��v���\K���ڰ�-���nW�rmh*aoɰտ9��\�)8��^��K�s{��:廡4$t�&
�_謀Bole6��D��2��o;E����XU��)��x�w�w��ٚ-������y��c�7��h�PO �X����^�~Å��)����	�A�񛵦��fǪ����y�ב�(�e���a="i/+2s/�Nſl)� ��_!Ř���bhzǠ�w����� ����������ן�4_9O���x>��ԟ��k�ҿ$
�|ϋW��+U��ܠ�A^l�1��x�H���ҙRsw��|��ķ*C����{�;����}7]q}���!��f���)�R��������e��H0]t�tq�퀎9]�b���T�D��J� �s�.Na���oiQ���;n�2�����9��w<:�P���y�y�9���E/��c5��>fϋ0f��/k��}uя�o����Y|e��p���۟vS��|��~�\';y�;�1/��e!�� �6t
� ���سUګjpR\j����z�N��k�;_��:��*mC���Rۃ���:�� !80�4�{#<nc�T黷���O���j=0"4�^�d����¢C-l�{�#M�C?���zmd�\L�K6�3NF�H9���'�ͣ�!d����:��eg�C����+2z�,F:��$�%�9N��ƃ9�����f��2�5�Vew���ߑ�{�[�[lt�SS;����x~0�K)�S�]iy^]W%M=��0�'=Rʝj�[D��g��to����9���ޤu��W��V���Cu��/�3snWt�D��*��V�(Ł 1�#�*��s�I���P���%J<����d@�׭LC��P����A���V�C��؏��gGt�ǰ���,$p@(\HE����u�����oo�=K���vo�W�2�LGG%�>�J�� 5�ppj&�p@A Á=��N�)�,�nJ�PB:P(x�+��� ���l�"���V1����z �J
��1�sj9۔�	)!�vJ�27��	�]�@�8���CB(���[P>��^�<?����L����e�Ϡ��{���葋��ڬd��%F�q���8�Vz#�^?��v��k���ܦ4�8�s�3�����G��9M%��N�:8�K�qZ�/�5D�F���$�zJϘ}�����U�UDc�@pL�|�H��l�j� �ܹ�����0��h��2�xT�w�.�!(Q*| �I�-���$�C�c
ϒKϙ�3h/��_���йE@�t	}�|<�VNP�2��������l��[����)o�����R�2��ai jl����x������2�ם�Im����$Z��!��=�72���2{�6O)�]�ɿ>��p��H!T��2���h�c:7c_�baa�ƀ0c0&L�|h�(d�)��B�̓�v�=��g92�H��i3x���x �F��Zh��(���>5vMl�C+�!=M��*ś�Sj�ܩ�>ǵ�[5�mIȧ͋�Ϲ j�u4����e�� ���Z唥��0�g�a�|��%�f��@ Ǡp�X�i�(�۷0941<02�1�:1�2�����Z�Z���l��?����đ�j��P�⽚�e��V�Ұ�^׆����~v�닢�۹z���������o���x�����SG%�n ܗ��ӎ���e&����;���F��}��q���W'�|��/AP�bβ!��A)h�dt?�����0�pM��(�1c$PJ���&2�&v��g�r/%���E9�1� @̑`N�R8�����i��p�ಿ�f�=�iQ�Bv���Nt�/�\��
M�wf���y �緓P���E����_�A ����{V�|n;������?��<�#S~�����!�DGxFx�y��}�ׯ*I��H�h��������'e���[@��jFM���HW5_�_��˕����q�КU�����ߢ�,�?L¦�L)U�r�ƭ���k="�&�E�[���\�w�K؎����C ��T�����T@e\���r��r�z��ɸ�M�3UȐ����8̂�^�P5HkmW:F�zf��j��	e��R�I?�M,Wģ��H���ۭ,P�uL����m�^��(�n��>Gl.�l��t�h�2�K���/<�8��w���r��g����G0w�ƧH���K��AS���l��Un�q�I��R#ފ���m���J��<�u�U%�n���r�&<�K��w�GNe��$���I�2j���Ō�Lcт�@RP�҈-�͛|[�����yx�F�Ď���7���݈GtC��dl��hs�T4s��dc���7�����S)/���ƽ���	�ɳA�A͚��ke]��]:|��\��3C����~bc��� ܞ�������j+P�ɜXMR�P�+UV7e�E�E��TP��ӐoǛ`���`v�}�*Σ˙?i��5#���Ԝ��ۢ�r���������(/�A�!_���-�K��#@8(��J�r�Y g�Xwơ�2]e3�J���!�IH�#O�X-mD�OɅvn/m�ZH�`mq�ީZ�1Jd�t3�o|�G�"�ms����a�`���!�M��Rr��o��H;ȝ�%ƱB�j�F*�F���E:�0��6�����	� πP�6�q���g!��ϼ������#Z��z'C������:��tRNC̓�q6ߛ���]�׫!6�S�����ʐ���������qh�W��1�ODK62��52�J�QOsT �����
���Q���SwG�G:,�z���Q~��܄Cr����=�~��u��E�z���B�3�	���ׄ�s���su���1��T�V�=�Qk��0�oa���`Q�i����us����\]h��T�����+���X/!��Q��y&�5!�I��#�ۂ~�X>��b�#.ܨ���+�´�eV��R���<�z���	?�(
���k����uz�ma�4���1�!o��}K�*��z,N¸�T��J��� �8�)Jߤ���N�Z�'L6��*���Lb������
�L�̜�ᑝ����v�C��T�]��1�I��ߌ�¡L%/ie��[��>���A���>��?cF��a���b>d�y,���[\��SbV����6���2d ��I�I1UP��n�;��c�`"�ͯC�D٘׺ ����c�!E���-(��a���aH_���A�h뒔���?}P��j���=C+N�)("�������$�y������e��n���e:,�r��oy�i7�F��2?��o}pd�ci���5�����G�ǟ��dĕ�ׇV���Q�8s�,?�	7�����-Jy.Jz|�����t	̵����/��Gp���O �$0��3L��T4��Ҿ_8�W�Zo�
O�7eW�Z�ŵj���w��{�] �S<T�/����'L��.�ͱb'�?�0V�� ��b���h;X���P�A)��x6E�����ښש��ՙ���5�Qr1�QE씟A�m��[��F.�w��;���,�L���_�bN"2�z����%o˦�G=S-!R{�~��^s�#�+C�Lݟ��Ao�����&���x�ǂ�ע���O(	3^_�-��^-ń;���Z�R�e��Y�*W"�>�孔Lc�^ �)"rϖi�j�r}����@��c������Isi}�g#�P��N��_������%n�h$T���`)'?;�B��7J���W�����پ?�m��͉ ;��&��S$���S�&�`,�wd��'�"���̧/4��%P�S��5�laT�.��D,�ᇛi��@�i6o1��X�|?��z���00Ro���z���^��6z-u򊱸��}���4�x��ڄO�y�?�����)���o@�1	� n(-��91��f�@�x�i����>��{n`�=��D�������i���@;���^�H2��$)4<�DR�g�+�`s���~u[��å��ueo%�u���j��� ��WqJ��mٍ�O�j� ���v����-9.<G#�-�"�Iv~^:�$����{����A�țyf��O韭�r�JN����Ĵin��R�R����_5q�j�����@���ߡ=Ο_%����A\��c���_6E��<������8G�Ϭ�����D"�X!1�P�{�S�:F�r\ؙ�8��d:�X�����;��v~��g��69+�D���H��Gy��f��m`�E����JP�ǃ�"ĩ�P���S�L�FP���FaSs�	7�l �9�!p\���;[�2�s�vr��;ۻ⠆g�]���g˹/T~7C"OW��9�u�1Y� �o�p��j՗i f/7�
�_�|e�1�V�V7]g4�]�n��z$;#��p]B}XS��x�הX�%U�֞�>c����1���C���0��.�gV�[Ti��<�6/�W!v�����X�!�P�~D�Q�(\E�+��ȷ�K�7R�d�kj�զ����P�����D���Ћ����E08>ǟ��-�7�sv�3(T�q^u�ً�Xs����~���]O����/�����[oX�YZ_�ǽAe�X_$^�4d�}���?i�y� 73TΐJ���!~W�r��N܇q9�r�q�#��l��i�Y��$TT�Y9*�E^߅b����K?��0�-IW�1k������6eA.�/< ��C?��߃1M�kh�ߘ�R� �b��ߤ�����LB�F�zYg�+�.?n�^%Fv|��9��ԕ��	<�\ΠS�U�QW/���g所¢o�%�R���*3�pW_D���F�}�pO'5����I?���nq��JG�vS6_�An�CP��#�2[0s�u"����eH��
��i[���[��n���T/�����gqF'�����azO0�A �����]���kE�䣇�}��}��}���Ͽ>�M�#F�#���e�!1��c�\�����h��߹�FG!w��oGmd+��� �a���eOUv�,�:�-�w�K	��V �0���~�`��P�c�6���f��z�e�@��2�b�g�rx }������,K�s���.pj�	��kn`'<�jThk�]�8zY�=��83���{,o�lh��s���ޭ�͠�nE��З�5�Nl���m������r@�˕�x���1:< ��0ت�9�����^�����>�v6�9�|$!���FmcJ{!���4�Bx�1 1"6�;����]��~�Ll&1�에A�<�ev[ߎ�3�	#/�s����w�,�錫_��\��}c��W������F�:N�&�*a�&���8h'ϩ1P�X�4��^����BA��q8��c�ʡnN��������ԓ�Pc������M���e�/n�nAKn�muka��n*�","w��%K���l|�Z*�Z�EL�_x^y{�J�1^�Z0e����%��9�U�����SZ��_���X��]*����I��,NB��e4<q{e�!��	m��q��� G�^I�[�V0�07����)G�l.����s�7����\D���L[�}W�3�i�j��+��Z=�y�~�!�k R'sJj>���W���Õ�ƃ�g��f��9Ͳ��r^��<?�V;;t��6���=wD>gg�.'k[.���$A.�i��U����!g�2�2�"��I�ob�B]t�9ǫ)���,��,�I�(ޜ����#��)���\W�;ɝ��Z�;v��u��m��_�%�t���)�(���̻Z̄�ɞ<� wDwԛv
�#��B��'�i� �*7���t'���/�0��6gQ1�f����`�HhVr�w&�I�|�gj%���h.{'�d\�������I" by�4�<c����% c0�w'kpgOu.�Ӹ��}��E���Y��ùv3�/�.�B �x�:���@�sá��D�V���AySb%��*�\!�8F�?�ľHg�&�aqV�,�\	�G8�/�n�||��_h>��N�(���:Av��I��$��7>W���YMs��\X]S�}d��N�o̐7]1 ��x�'}�
qf/�EpG�Q�NQ�uOq��Z4+V%�k���m�/Q�hHJ23��{�p���j�ׅ���x��ݧ���N����������X���D�N����l^ �eG���	`����J$�+A�;��^Iz�g1�H���B$5F멾���,9��2�y/s~���U��f������]������엕�����������ٙ���<��zDH��r���>[����;4ڮ�>o�A؟-~H(�ۥ7���Ah�� �/S��&	���y���wV�,�e$/P(S���ݹ��Qɋ�z�8���AM����c�MK�m#\�mIT!��,��0��o�{4�n��!��;G�,9�D�y(��9�����p7pg읗�u��-����v�+�q5����������������u���t�-�ڏ��!��^��q��=i���n�?�ɣt�$����d���R~����`pԼ��`z"O6J���5���4��3�`�]5�p���Ld(�Lc�cZ'�q�[oZ6���o���6bA1�4���a1�Ա��pmZ	9��W?�d�I��Q��f`�-n�k��@];��k��O�Ѥ��_�����tKp ]��On��].�6=U>zQu>�%J�)R�����y��������l�% ల@i��M��.�mr(v���ލ��vj���qvCdlabf`QV�e^����ZW�l
��*�����@��An��v���� ��}c�w��S6�lB� ��Gic��dn� #�ј��.�����$A�J�YtI���*Z�M�b�y�%�^�Fg�w'�Q'�Z�-�*��B�e|d^��7������/o76I�Z6V�8�Ơ�#�0��uL����#�~4�=�՘}Ѣ�լ&Ѽ�x*ys<�v�&=>��.�=A�	�"��~Y>࿝�&DqX� 7�.���$.�s�%�ܼ&����f�=��ԔV�W�1}�f,���N#7��P*n������/�Qw����4Oj�n�}��=��EF��a�t��%1H�2�{��=��,�yO��C����u�S�O{��Z3p��.���T�N]Vx��mS�\6]t�v�ǓiKC`h�Ys�ٮf]�T�ϲ�S�ҩ\��f�hv�O���|{�fg7g�[�����8�d�2j��������%��s���L�a�ч�/����&I_i�j����A�VCQ]��V��>?���ed�5��t�d|7��^4Ђt!D��ȩ_2�	�Ex�b��Kxߨ!]�1W��N��5C�.�OD.�'Vӧ&��3	�U�Y j�{��FH��fݥ
���������:�εz
���H
���W�i��XE�br���~�lB��n��L�FVu���(%Ĥ�.��zV��X��nNaN��D)D2_��Y����]�{�ȏ�XP��].�?�Ǿ�*�����i07���uyn�2ߑ�1X�Uj��Ğ1bє�'1��?�[j��׹)�9~��|�/�^q��&������.A�,��2���D�%|U[��.P �t	#�8[�e0C��1U��\�������li�\H( �P�&2�Ja�Fj|��ɼ������}�=������zu�����޿�w���4��;8g�"��c��ǥ8W=)FLú�md\E.`!�X��{<M������L�Y��6J�u�|I���R�i�y��l�ʷ�|���5;�v.�&���t��(�~�c��w�O���^�P�&��ť@4�'�� �n�x4��JO����}�8�<����iY`��7t��3ow�<A:��I̍�!�˄m�t��ob��uz�t��j��*�(go�(Zd��c�`��h���f�^��!LԴ�D��tTBک�o~�m'������<L�m,^���^W@�����1�{����oA�g<��
�6��$��b�ھ��*U>���iVx���h�tB^-S�:۔���="�Jb�_��Һď	��#.�G��Y����-k���������>S���v�����޿>Q=?��z_�ݬ=􏷼�C�V�w�a��i�t�w����3��������uT��Fh��2~:.�A�{|��9�8��a��y��Ϡ�8ʍ8:�	LבĶݰ��>����J���p_�`K&%����D w|�N�0tFCmC��NV���\�H�Iw4�QfvV��T s�G�4h�o\�5(���v"��txYIGߛ,��xN���+��k�Ϋ�����/L�[��g��𱿽	;�>y���g//�V�^^,r�	[x����z:Tv��D�,W����X�k��o�����0[k#3k4b�t%bR+�i��'�߰������ٮƙ/�n�I�C�6ꆟ[�\���Ca8 cN�&F����3���H��䟱�2I(���dQ���y+x���b����忈"�6�F��J�0g�Au���u6=���U����.a�!��k}ŝA�-�%���4�Z�0C)�)�F��os�����v�sŀ$��O����GN�nv�@�6]�f]vm`;�r3�t#��j�'��R��z4��Px�������Y����p;�����V[YOW��@[Y���e��?�݇����rY�TI�L#�)�m٭FPaxT�;Y��?F�[�޿{A~'�'s��׺��[�4��e��')(qw�����N�5�e!V�ZY�׿��	��*n_m�j��փ�[_��g���#�B���
����F?-jm��sR�k�v�]�����G7���+Uk:����Z-����3�������-�N�0YE�l���%4��x!�I�]Ϳ ��j�U���N4�����y ��'2c�7j��q��p1��p���t
a�N�BL�G0(���������2О2��J���#}��� �|�&$�?�K��	F2�~>�#���P���{�����嬏��Du3Ju�6�D"y�rfI����!�	�߄G;&ȥ-�L&r�i�My����tv64i�<H�8o�σ��~��*iY1Y�ĉ]��za�C�B}�BC
�W��j���濽͗t4��n��֌�_T����xM�fҞ>�+ϙ��C`��L*ߋ�-m��#.��o��C0��r�j����������A�O���BžAv����1P9��"�_�@�j����I԰<���F||��F�0��y$���eAl;�SpqRс
HZO�@,8H� �u.yF:�Q�[*�J�8�ه��`�{p#. 'H���ÅԲ��
!�N����0�{`��\j��ΎQ�dE��/��<�11���$0�d��p@��~`P��k�w?��ʑA��Ɨ�I,��B7���gl*��{�ۮۻ���	�GMCi_w�4mݺ<�x�j�l��9|[�['y�x`M(�b�����>&*���I4������j�0���������Z~��L�*����*��l��3������G����q���i���Dio�����0��şP��3��~4o2�-�-6�<h��x����?1�&AGn������a׮<�VsC�+r��c���ONͶ�l?�e~�����D�І�?d/� �:�$��Av����=����<)7ll�������x�_�p�������]���S��
6.oE�&����E�V�k��ֵ�3HIz�.j��\8㝬��&��ώ�����o�}�j�-�Fe�.�;��w٨�K,��'�4�a�c8�����E�[�I#���
e��/"܋q��?�i�G��ѧ)���Q�A��Y�c
&*� �il�H鬪J4Y��/�Y��7*4�G�j����Z;��n��9���#��KM6]X�����E�O���}⣣t�}����A)�]zri/^����dG�>G�a��C(���>������@3~�}���f�!�v�E��[�3�_XnI��"!�ۅЧ@ ���f��􃃃R�~���j��6��E��M������9�jxm������+tl1���P����]T�q�H��r�h�,I�讽�Ǔ��<�ȢT�����f#c�k6wD�&D��W*��ӝtrq�� 1�Ŀ��] �财�S�ɀz䧑:�o=�ԙ��s+1�����>��ɤ�\:%�E�|o��~��.ЊD�릺]�d��>��Hmb1o�<�x�s���d;�E�PK����}�j�j�%��>^l>Oն��HxdT��<J��e��ze�;����Vc1$6��Ym�Q["_ %���P�*��C�~rd�u=���*#t���h�B��==_�%g��&=q��)��Ƨ�[�M<]��T��Ly?֐�'�_LF9�(�B"��.,e}^�/��+����*y�\V:���Jn{|�W�Y���6{���U��T*`��(%c��%2#�E&����m��+�[H`��YF\���ȶ�i�i� ɱ!ɂ8��6�q ?�IZ"�����M0^���*�>�P��8����*�� Ћᇹ~�&����5H���H�:��P�%�8>�u˓�����?e����OY��Go�y�.p�%�W'���F��bRbKCJ�>���U��v��R1\U�0�5�r���Ē�w�l(��1���H8V����a�Oh��L��渫ل����6���?�?�o ���������6�I���g�$V��JE������Xs��!N���1�h���O �-�'͜����we�C`g�~�d���!�lY^�wpʴ���67q�g����E�J4|�A$��^��P�8'� s��� �g�EQm���S�߻����$��P)��eSC�v#���&����|=�P>�?&'܃%��&��{bP��E�Y=��?��������1J(�á�k�k�����C�y�NQc���XF!�1m&�����3;q*&�gРĭ�çC̭A̧�ϭ�H9~K5qM�k�����*,��]�˭����|5���H���>����v5,S�dL�]�Ӫգ����#D��*��0�`����J�&њV��4覘��S�`pL	���Q�Z�ȔO7ah�]��,���9��'B3�?hӱ30�����t�m �Bǲ�������mE[ag;��=����$�E�Oݶ-��{SU���U�<#SY�����(�)�KOVU��GS�#�/Cܒ�1�#�`g�\?�C��;L)�O�W$��b<���S�e���B�"m�����l����T1�DG洧��\��
�d����X��G��R��i2چ��{�\�(�����C�_#�se�ǀL�tzǥ�Q�E��C��M��ĩZÅ�c�#�J��Ӎ�z��6�K�\�������.�u(���
[�qc^��1u��|r�a���g��َmm=+�J9���9��q3b+/מ��5�YÀ��!�Q��gN`b^����Q�!��_2>��uf5m7����_�M=��G�o��@r�#�8���gl72����E*���=ɓ>��5!��jQvss��E��@)Wc��򗏠��7��i��G���_V��^D�Y��?�;�lD��GMt�9�������gI�8<̚��V:���!X'}o6�I��?�Jy�����P:P���jz>"�>����z�m�� o��i������6�c���ż����1��{Dwv����ki�/#C����X��_K	��j$�UP�����\���`�s;?}�w���O\�H��P�"csI0�E(��P��lH����C����@����AWJ�k�z*^�t_��ۖ��}	�:W��J��Ա(Hq˟�H�v15>k�����+װ��o�h�h3�ENf����	]م�������g�r��ֱ�i�Ff��a�ny�P$�sKOr����I
�m�#���ޗ_�m���yF"��?��}�'u=&����ç�p�ť���W�3~Q،��%�������r&2�B����<��d�jh��5t>(CP�萂�d%�7��,"�y>�p���)��*�O��O��;!�`$��$pRh��m+�E�N����0��9����Si�5�D8�2l+g�XR��e#{i���r���Մ�{Za�����/� �y�0;����[[;y�2�_�gD���M����g�V��	�#��wLC���a��V���9�9���J�kڡ��xr�钬�;Țs֐�o�-��,���c@����
L�����#���v���W��W���J���Έ�L������%w�=.�&s:�oD���D{���\&�*N�o"DX�����	�9�fC�P�dK���~�S'���P\�õ����/�~�FR���n��{����(����g0O[��R�|(�4!��\Bd�?dc��x23�����ͺ�B&k�r��
���=�
��y��%��{:�g2�C��m�Qh��kg�]��d�+�����;�s���&�2���w�/�����9\���I�����'-���l �B��+��1{����a��֩��e��E�W��:�:⎜�^2�jb=�s��"�t�S&��/E���&��\�2�wJe��~dj�U>�G�o���h$����I�y3E�J�����ځ����o�$���Px\���L+�!�#`�,^n
At2���Lz��]��;��P/�\�g�}�8���.� �$��	DN��`_!1����6��:^����*�:��|�Y|�z}Ȝ�}r�}���n�\��עXȰH��9�Y�����1;ബ.����.�&��f�W� i�B���w��i�k�]C��mT<T�~�����2�����E4=5�B#�25WGWO^�Ƹ�����r5�6�����`�1�xCUхܘ�@E�F�:�)
@�����$I�c��X���QM�� �E�1d����8#63p�jД�;��5<�΃iy̹���Ù[����">?Y#Y�U%��S�2hr�k��"g�u���:w��~���e����L��11�Z�?f;f�*E�B�T�fj��������+a�d��d���_���z���������e+��u��U����$����h�o�v�V�%�XJ�O]g�d�ɨ?^��ڧ�[#�%p�~zR�g��gA�^�)᫆h�`�f�a$~�*3�s|ɤ?a�H�����Ǉgr� �Ds���$h  ��GV��&s��AiM�:�ߔc;�	��ƶCC牓C��T��/�e'!��s���=�u���Vx_�T}��k����p���4p:4��yϝ���l�k0ΛAN�[��O^��Wo�=��c�_��N��I((���"#��.�٨c����lsn4\w�� �R)��&,����P�] ���T�駨�qr�k��/[��C���n��ڐ"f�b���%,R�GJtT���%����j
�ʂ���gf���j��Z�����A�+*�|��������.U�~2��A��������B���ꃩИ'�qtT��(E��4�#Vv��c>d�sv�8N�1��s���e������_F]�v�i8�@�L+�mߏ,_�5�u�;8�ܭ�Ζ�[G�j�C����qtxmvx"���bR�E������y�Uyۿ)���v���Gw���/}�>��>.)9�d�[��N��I��ZK��@n�Yඃ촃��������xl�x{���*o�㶩��4 �v�k���V�H2��c$>��{Y���v�G���2[��R~�ؿ��.f)b���C]u��{�hh
�U���e�ʸ�$4��~�f�$f�d3��]\�l/.��s��N�v�Y
qĄ�3��u:Voٶ�hTQ�	k�F`0qC������1��������6�
�e��5��J�塈S��U@La� �x�?J��%�e�\]�h��9Z���;���:����H7�:+�2/�/�P������V��Z��>W#$ P���A
�����:V�]���F�Hr3p�BG�9��,?!��B��mVtQ fF?�2���4��q�� ������Q��h��Wtۈ���t��U_�oE���@O#���� j :- a�S����lj���bѱph�>{wݭwyk NKϧ̀��;b�t1O���ǜ��md�拂�@e)���i��s�J���")UD�R���0Ĭ��3^��m[���^��&����(d�3�z��sA�w�[�/'ŵ���J���/��8�\3)�vt����Z�������SvHh:`C{8�����Tup�2}�5����Bm�.y���ފ��}cp�����R�%�6&����6?7�M"��1;��^�G��`K4��Y9_�'uw��o�L���Z?�Am���V����|m���K�7UY����ŗ~�+��u=�Xf�|��.�[w�ٽ���q����o5�$�}�(��"qרG
�H�h�br 	�'`pc����b<�쇱i�wM��e�9_O��4�������OQ6�(���Q@��?enfEu%�*%+���{ۨ�j��􄎱��b�:ˉbKQ�VD��Zq�|�o���K��(��)ƞ��f�zrP&5j7Ƭ�x~R��<&����3T�(�$� ���P����)�3���V?����r߀��������(�fa�$��ƞ�3�M�W
YT�o��tu��:��A��I��M��ӽ��	��䰗�����۝JO��N�b@N[+�T]�׫�Tk��7��lv���7�3�����6m(dh"��e;������Et7"��Z�o�� �-f��V!�Jbt'���S��N���|*�&]�1P1�6��l�,	4I-P�=��,4�h�2U�M�	�\n����2˩����|(��45����Jh�B���� #��ơ�-���k����.���㐟����2��K��˼H��hW��6Y����g�En�8{�Ǣ��`�b�'?����f�b�ϭ���ln�G3������7�ͧ:]7�g���:�9�y�˦�<|�7���j^���@��|͒�_�{���8����h[�i��t�	�X���xpw!X��`�ݝ������{�O{?֨]5�7��^׌}���!��#6T7��7a��8Jw�l4�>]�TXn^LK�Z+�d�?1ȝ+��>R������Y�n]Dj��P�R'�Y��%�+F��x���([��1��a��a�ar��N��1���ѵ����y���TP��j���u�B޴�V$�`z��Jd��W��Q���L,h>�
���L{/1H��)Rw仿���,[:ŗ�bi�xM5�Et�U�J@����K����v-��z"P���w�����k:/��]GC_�o�v1i��}Γ��lE�
AD=�W�+dO�b��}������c0���Wn�D�v.��S��2?�������V������EA�J�%��X��;��׮�綹����P}8!�/��H����U�8A �^�Z�8-瞭a�KaNzG��*��_<�y�c�)�Ɩ���0毫',Dg�t\���k3D��Sh�w��g	�}v���C��ҚR�����hU� ,S��f��BrP�A�3T��8���j��lkC���z~9�xNiC ��L���.i$V�w5ŷ�Q����W�^ �w���:@�E�1ΰ��b$:��,V�q��+K���s�
Z}�*���n��^h_bhѶ�CqO��W/���b�S��^�q)�]�l�hu�~~�}:D����9�
 ���:�2�o���29��ɥ!���%V	<��7n��5��AUS�i)t�vMLSCF㪝{���UHfM����w��ǽ�D�5ݽ�����V�\���./���-D�)��zx?��q�Y��M�u����%�(N���[iA�7��Za����W�q'�v�̈N��X�If��%�N�67��@�uхBzɮ(<g� �6~�sh�b=�ǜ��?��E�D�rq�mC��0��79j2�:9��w���y����
z{�V�dHk"t�M���f+f����}l�8Ч�`$�4oI����:iu�N��x���v?<?��0Zk���k,p�-7���̀w���K;D(r�Jn/��������kBy_^)ԅ�*�\y��q���= Tp,����錔���~���u��>?�.���]�1��d�M����7P5�,�����c0�
�`7�|)6ZK��߀��5���uU����7H���9
�H>�f���~��.;�S�>��V�0��aŹ�8r���������vg%YӾ�Sc�yإ��'���7zMjP�����l}��T�\�0�D٘��q~��{��*z{F���o�_�T�L�}�]�$�9aUw�M�$����Օ���������|�j���ް%N��ˢ�{?7�����]㪀ʚ��5�S;�S;f�˗[Z��s����H�K�W���hթq@�A�k&Ք����|QtJ�3���$Bb��,~���: 4*��Y�C65���֔��ǎ��??Ro�N8ptϱ���q��һ��g������J������"Q�?��uϟ��oq? FR�P^�ܠ����!2�&]������/z��I�F/B*!u����z#ҡ��II4�鹯L�e#>F�o��.�Jt~e*�tj�9�S�O�#S�5�`�y��-���(�\Ӄ�d����Mg}�ri�\�|j�g�ZXCƻ4�BGv�4�J'e��i�?�֧�g��w�F�Ȁŕ9�O3v���^\���1@Ts,�ߥ|���i�,4�����od�7�)W'�-���6|�s����X��j5��D1|��'W��^h:���:I�0��=��B�,��ѕ�:���\M��LG�֞���M�&`�6���fw���T�_�U3�k���?:5���ze��$�������<�Y&wI�������⟅u2�>�]{�����w���7��}�LG������`��δ�К��e��J�l��)�}e='C	��V�d��<L�o�Q�X �o��~ң�r?^�HEnY6��������pΈ���		a�ZD�1�����o����a�c�=S����w�#��t",�B4�	=�1}����X��)�M�p��8;��=�P-<�����yy�����s���+V��1�D�:yr�e��=��7,��ş\�\?;����ꧮ�y����#�����M/���s������KR̉���2�p8��І:��V~sP��xC�����:Q����� ��R�I!�|�!��8$��ic5��㫉�]5W�C���ɻ�rOkU�鴹����bhg�kM���$Ё�ܧ��R��k=���E� B+��oC��-��v^���t ��H���NR��$��H��H���g�?��\��0r�v�x�@�Pz����֙��<E�< �(�	��2`툲����F�A�s?�j2��]�Kl��)m�>��|���^m�	V��35�g�m���<FmLT0�Ψ��YYkZ�T����l��b�1�l&�t2�&dd�����<��wF�%���Kl�}$�窍����c��<1	Qʑ�8���E �4z]��]�����³��҉2�!�4��L�1��dC���ٕ��!fa_�����S��=�́�p�/:S��7���ǜ=�P���G�rҤ׾ň$�ŧ����i���~r�0���p�mh����/'�����BV���?�4��+)�Qe�Z�FVZ��-�aHl� �9q���1����l�yf�a~ԥ���~F
��=�*�3�8�O�n�}���0�
>�\I��:��_)����H�9���F�%ۡ�������[r�M!J�=ڿi�@�d:��vƓ��x%r�c��Ф#�G� G9P'G�\xZ{��%��e�?�$1���$��QDߐ�{
���}�T�h�����&���z�����s����}�a��]$o��QT���siR�*_�n�0M.��wj��"��i$���^�C����ʚ��&i֡�xKO���(��&�aՙ5��-��C����d$BW�L�1�9$�.5b���>ߚr�� A{%A��HQ���� ����V����e]�v�}1��ƃV��Uʬ5	�_�e��x��_}�ޡ���ϊ�f0��I�.�,��n�<(��Dz[X�w���%22\�����r�V�O�GE�Z��w�ڞ��Z��O�W|�VGZ�����>
����^�`]9��|�q�&_�sU�]<P.������H]h�k:ݕc��������D~H�xH�3�H�ф�~�'��|�bOg���O�#o�"!�3�=��e�.b����uٮ	е���q��^~xҢjGe�x���l�O队=Z�Iv��cS�d����;�	�������N���w�\����~=K�O0�1�����h�0#˽+�1��塓��C8{]�loB����C>Z7s9U����������*���n|�)D�K<o�8;��'#���m��f����X�p)kƙ�y�����њ��ME=�	�Z�Z����"�x#}�	W��2O��=3E�ƌ�i]*�S�`C��Mg�/ɭ��{P�K��2���Ok(�Xz�!���&xmZ[�L���2[�3{?�zjS���otj�U�Ϋ1䗆6��/
��>�0��C������!���Љ��XF�î��4��Q_Xe���v�6���-}Q���egһG	p������v�'���&D�֐��醛8"lKo\M,3M.s/�T	��ο� �����⣮Ϙ)���rd�86����O�hU�T[}�05*c,�@��D��
a�����5�ǳ_׊�h�[4�{�=l=(6�S9����륑��CJ�B[��}�C��I׿Y�����Ddh��҄��XǸ#B�e�����p8&��:����TZ����m��ST%��A��Z�O5
 ��1n����'��KMeh<�Y��Vf�j
���۶ʅ�6���ɦ˃�CV�qw��ȵ��a������Q[��d�Ҭ=R+�����K3r��C�C�kJ�TS���5��z�yE�NA�q#J���I�5��V�7請��=z�l�b_��ʏxH���/�qM�;K�C/D������)k����N��O���\�:1��m�B�u��=˄EpS���cG:O��KF����0\�d��z6܅4X��
���:�b3��y���z�h�V^�k�V[}�rG)R��-K�_�&�s�"�$e�d�E�:xz�X��uB2���h_��-�0���:��N6�`�E�_oE��2��RLıEl�Ǚ6��=�!؈�� Κ��������uūx���h�P�����3`޿-,�U�=�B�#S����ޕI��x�'��n�Oa����� f'a|��/�A�f
s�
)e�F�[�\@A�t���S��0$Y�iӋ�*��	ۼ�><��(���=�*](���(8+Q��PM���,�P�_3Q'�����t7{�B6�TF�@��E�ul6����9����lje�����yB�A���3���LrY���ż/	�"��DC~Kuo2c�������[�z���{\c"���8CW"cW�Z�(�M�~g�>Mb�/M�?#t���p��I�9:�3۫[|,ܒ��\W�����_,;;Q9w��F�U�����i�eX��3Fy��$m7�'�L�F;�F��ٳ���* B������b�ϳ4�J�|�퍫�U������һ��Q��پ�㍣�f�џ)�yj�s��}T�mO���U�O��u��g�Y�m�ź�G�B��1�?��?�:%�}MZ�MZ�7o�8WpTM|f�o�y��Q�(�����z՜��ZJ��$>0S!��7�G�u\qJ��c��[zZ�?I��f�RAٝ��FE6X��C%����g{Sӗ�����A9�v\.�J��o�ʟ`g8�l�T�uآ~~�j?���4s���?��|��?C�ǿq��`{�꜑ ��t�J_��ƿ�_$��
$ ��M�"��MC"�nM�������f�*�\[���٪�y0�ǳ>���t˃t���⍙!λ�(�RRA�#A�U/�"O����kI�]�n�����4p�:aU(S���2��Y�4m���i.a���Tl:v�D�{�X�`!�`�Ԛ�#Qc·�o�+�$q���U;��0R*��Qa#�e뀗���P�lZ�`����a�f�P����������z��_5�΂u5jߋ���]r2l,�~��q�Vt�~������C�����vr�%�r!��W�h�tR��0����"[��<����r1��M��+{���2�]�6}N����l�Ue���\q�d> �蛊�dB)W6#���
n�iW6�kN5��z׭��F~Lو�AA�[�m%xX�L��ֵ�����}��ߣ8�����n�XQ��Xb<ic�d���*�����M��K�����x3��c��Q&�11��1ND��ye�1j-Lg�;Z��|[ba v=2q�o6Y���ë:�1�M*IM�>I�<�4ة��r
�J�ؼVai
���|���>  ��xX��Mi�A��NF�l�~2��2�
�x��j�;�LNa
��(�U"z�ۂ�8�*�  �OY5��8�I�6�_�P46��4܍tx���2��&�`� �B�݄�EK�yX��AfF+M�x;�';���oZ�Q.Ls�����VV�zyvh��h{u#>���6��a�Vo���({qs2�o�R���S- .=�ac�mZ@�y�F��y�cA����hœŉ��~^�����q^�	t�z@�ge��w��eL9��!�x�k�J=3�.Pmdff��������N�m�$�N�8�����P<,d��N]j涝CPpY=kK��[��� x��B����a�x�[��0�������T�>��b�?�͜�8�3� ��*��;�b���
�\��ؽ;!��(��Ϻ��`x����6 j粒���I$#J�d#����>J�N7̉j/ ���1s|����KNa�7��l�PK�s�i�V�A��r�Q��n,���%�������,��{Mg����e��;4�՘/���MR��X=~;
~��g�KS����6����\/���\4�	��,��#ns�<M��?���/';���$Dm�n�;7d�Ճc����c����`j���S%:�)p�YL NҀ=&��-S��W2��TN�e�DP�h<�/��]VZ	��.���ɲ���G�D`��B��{g(�|����M��&׋�#Zq�v��z�`FX0�m��U)�$�$ե͕�����$һ���(�o/h��
9v��y����g��G�����G�c^�n��I��(��##F�>�E~��LN=�G�{>��u��վ=	�:��e��5�H�Xhԩb4dR���G���՟�����C����<��	e��ר���{Rz��4��8K�Ӂ�~���5�G�G��%u�YX�������k=INn� ���7|b�k��<�]����W��e�
[��q˲{��)�@��qq�7�4��$-n�܃��`6�TI�44�/�w`�Vk�m`�m��� ?�%�<(�b�9�04�YaS=�į`��y��;��!>p�{��[�~٧=v%`�Y)5vb��NX��&��q��(��S��K��OX��%}��b#Ƕ���j�������Y��%w��e�(���N:�B Z�3�����j]=���D�		�itQQ�{�'UqwbV>�U !�r���(3�04$~��nƯPj�N���V���Kn��gЧ�^ LIW,ws5�D��x��aM}%��a���?h�D����g�;s݂��:�c�yW��k�b��2A8O�?2��}��2�b��'�r��ٟ��b���� ��D�2�@�����I�s�DT����w߁��Q�·c�����Tm��ɻv �d9r�u�y�[����Jޒc6&�fG�}����MEk_�!9�x�*�{�:�XV9�@z誦�4%�4�#n��"9�3�(�t��*�j����!5���7;<��+j�7���U8+�-���Q\
�}8F���9��f�m88%��P���Y���*������c�'c��)ñD\`��ʄ�V�����p`�|��Ǘ��)�
ON=�ekv�Y(��"��]����i��N��Z�̸[T��! c8Th�c�1��a?
|qGaxI�1�k���ۦ6y�3�k)N�z|B;�[���klbr����)7"*(�T�˩�3��~AV A���������%��y�Zd��1v�љ�d��"9%���vzfĻ�Xߒ5#Ćk�J�kU�s��N�as���u�W�B���%6t�1�&2}����#�V|�械��(�4�W4�k�l_��3�?E1�Ff%��'̡7ƀ��r[�­a�~�V) Ц��V��*Ὁ��h�Km�E>6��D�Y�,�E�Q�~�M���#�M�씤"MM��WZ���K�eW�������?�9�,.1N"�չt��@~��Ƥ�����IxI��n���Y����T� ��O4
��@*�'�ۇJ����>��������V��{�nd�:�	���*O0���έ��C-����ҕi�P,}���X�~V���C*5]�/j��Ѥ���<�P���qP��瀪s�jK�6��g��5z�F��,�<��X�
��4��F��	6�>� o���9X��cP���c0�7���l{�����[2I��ub�rj�v����a�?������.���i�OR�3V�@g����Ԡ���˙�����V���+�8��9m>�)��*~�MБ���ѣy��DTO��!��Q�k0C7㊩v��1�i�(��c��7�uỘc�gٶ��>�F8�]�~(�vA�yo��䣋�ux����,��ED��sU��u�"�a���m������Gu�1��=��	�	d^3�R�PA�_��h*��F9򆑷�Vߜy���73�<���Bd����U-I���|ד��iR�A0��_�t�J ;\~k&u����h��K������1p7�7�!?��KL8~��4�T��w9c��|���0LGc�EnS9�4[��Fq'
�M��V�����g3�k�*Ä�E��<�E��эuĥT9�,R�
?�'����n���@λ��&���;�����0E^Q�L/mN��Z
��ɵ4V��Twi^��i%:��`��t\�B����m-�J�<b���Z��Z����9mvo�ڞ��wb�'B�DvaN*Z�7�j�Y��y Z�X^$xa�xR@���;�
�ݺrY���(�vD��s[z�q=u;��9�*k�G�#o.6¯����n����[**:�Wzv��Hnf���Q�7�P�|�`��Jq��RA=s���y��l��X��ռS����o���A���adʒ�4�
�u�!��tb[�gt���j�'J����d͇����S������bv��h�L�^��h��c/�l�>@��9����
��tI����R}��%��z�:�YQ|#Q뗔y�ޫX�Z�_�����U�0k�rBW2�!�dz�KT�����`W������O��C�������|A�j6�g�e| T2l�+�((D�wطH����z�k�>���'��g��LU97���7�)���m&\�,�\�\&}+����P������#,zP���-�\�&�g��X�՜�՜7f�!�Qg�j�B@2�����Ǉ�^~�I���+�~���
��A�ߢF��ݶ���й�����E���7�����7��=Ͳ%2c�e��Gj
�N�aw����VȂ_������0��6�C���w��e)$o8n����RbV�ѕ,o"�S��p�A� }Z���1����������˴'k4�`�W��e%��\����^�R ��\���:��ҙ!����3�6K8Wtf7s�>xGln�а֞����j��#��q�t��[_ڰ���;0��9��6�����kA͜�>VOaK�ޝ����E_¨��1����.�������]��}���	4(�$�	�`:��,&X>p�(xP:>��\ۈ�0:����7�ס�g�r=��*�)+�U"��%�@I ���K�pH��fK�rG��{Bj`�i�40�U=,ڌ<�ͮ6��at�0mƆ��Tdd&-�i�S��n�#�����yL�l�/�Z�^0��Q!��H�=T��-�w��w�xx?��g4�֜��-iqV�ؠ�m�)��f Z)�W��keB���y�&)���.�l�����N��')K���2t��2�~�w���{4����=s�ι�m�O����\�5Ƹ���JL]���)g���������c>��ڧ#�i�m�n4�ťӢ�����h#�uS��h���"�LDގ���ȫ�:~���q�[(Z���������ZQk"��N��m�@V	BfQ&�<���yю��%�hx݈6\-�tM�x��}��`��c���ԨkN43��ݗ@�ӓZ/�5I�'O.'����.ã�-Y%��'+~7�I׶+<���P�LV�#d�a���7�~O�
�`h sH������J���ɲ�>~�٥���,+���1u��G_�$��G�x��E�}����L�&{����+����Ɍ!��T.$K�iX�L�y�aVРԃ16[�_$����	��R�}��ڃ������R�G�J&Ā���h�=q�D��|�v%���H;+�5����=�������y��7�kF�Ck�
+��4�]|9�/��y\n����YGC8��(`+d������S9�B2���i��	�a�T�=؞��J[�x�Ru��uz����`�Ǜ��c�y���[f.�j_�<t�-�*��)��ͣ/0�;䦁�u��ڏ�ڛY�Y΋�%5+�sն������4��0��M��\)�ǧV��Tٟր�L��h=yx�B��c�o��3]��t���eo��,1F���J��I��k��p�܅δ��*���v�(
�9�Ч��l���?�x��8�M��T����ۓ\e3*%--��!�N=�+{��Yq&�܉E�R�B����3{UOp�'B^�F�RZ4n��o�z���%)2� " �:m�c�"�������mPKv�l�Z��}=��_r�k�_Op�/zR��ăy��csp$K�hs!Ȥ��Y�/�g�n����5���R�
=��яsN�@�/��0ݘo��B�G\�r���c�*�/�,�(�Kڸ�
�%���X��c���r�c�RO�#[,��N7ctG*b���=�/.�-��U+s5�t�@��	(�&�2��'���W����(;��k��i(K��|U������}��6��S��W��jr�]�f Ҽt�����@�oi�F���O�:o�L`"7W��hl�5���V���m��)��9iG�J76�h�p-H�U�<h���8��|JC.������������D2��>������)ۢ0�75���]�?���T#��d:��-�̐~L~�Z�.M,��������6��i���c&p�!S��ooc�s %�%�?.<���PCRb����@xK\9N�L6�Ama:S�1���=YzS1 �+��r�Gp}��Y�6;=�F�-�:+�d�j���us���IY������3&�Y\b�^9}DZ���p>:"aP3V�����҂
��o,�ں2ߏ&�����@ZgG����+�P?�Y�5���>��]�#��*Ě��/3s�M�'T��k�����X��?�����Hj�)Z(�s��$�գma��h�iƷ1�t#��}\_�L
��'G̊����׃�P�{ч 4����ʸ�"�_�+�`��hJ,�����=az���d6Ȧ�޾�˾��c��Sn��I�L`��6�f��yt��׶=/�����U�Y��x_7�X�y>T��-�:oˇg�T\��<�?��RRV�+���� �}gj���kDmمq��9�Z91�ȑP�p6��n��~�d0���k܁���
 �?�C�:���bn2 ����<0��=���ɢ+	�~?s�Ax6�*��^SR%�a��Q� �!�||���+�n-�j�Ay�����4	�$�m(o�x�dYy�\��W�R�y�8Yi�}��if^�wB��>_�+�|J��~5�s����N����<���98I^B�Sp֏p���H�s�!.�ǁ����ËIB˸=�s8}�e�DZP*�;��3��5{쯟P���I{��&�?�	֫f�	�i�����@�4Vʷ���&s��3�ֹ��5>S:����Y��@l�qD�D�����Xb@:ʎ9N�#��ة��V��z	��r�@�ξ!�9��=#4�[�z~�����p� ������ɍg�Գ�����螚wJG��N�"_�ޱ��ڔ����?z�>�Ӱ�UR�erQ�h:����(�>9�em��o�n���RS(�_��� W��Z�zK��QXt	���A�'Y�{�ď���˒��2#�e�5�\䗓�b��خm��ُ�3WƝΗ.Hp��//�F(ڞ��ߡ�{�01��H��)�����lX	e��Pΐ�y�5a�Ҧ�l��z_?���ԈLM��>�NX_�7* �Ց�5r� �1�@$ p�{���y�*�@��a�#qn1v�i�IAem1n�6s.�N7��ǻ����+[=<:�2v3O1�J�:t���$c��2�09{D��lİ�E}>~IK����>0���б� �Z3!4��U�e ß̗�R���|����*{������"OEx���]������y1�Xֆ"�~ۭ<X�s�!3i��䬴�H9	�?�vl��5N��_�H����N�)Q��<5���Q�HT����\��>��G�~�CcF6�oX��3�A	Q�2�v�A�C�m=]���Ku�
Z�V��2/�Z��N����wF�ƝY�y�-��/%�%r%�[�#Y��Xv��4�*i�B��V�RiT�R��,��l�~�.��!�{���^̧ɥ�Gr���A���s��S��xa����xr T�k��/��P���Y:�'�;�vW�i-��I:S��C�����'���B���=]q�35Q<���c�k����W�a~UCMG��gß��>zY`�����(�]�F���-o�җo/3;r�-lqߩὄ��M\�-�־�hi�`�$��qP�L�K���q���P|k��Y���P.����p�SГlz�mU���i�!N�ТU���@r����Gdy�ڄ�WP�����B�P���4C�E�[�`U�ȹ*������%2������O�]�'"�O�-�T��O��Y��=����GU��|���c�WJ��v֙C��ߚ�+o�����"��^��Yn1n�dJ%�M	|���G:Νh@��1��y�h��	��)#u�r�[�o��3k�$�p��x�JX�rh�̟IY�1YA+�ߝ3���E��Qod��"?,�n�=�G��=�a"�������/��9�J��ާ7��1LN�\�MrwXiq������b����&��'�S��R�\bKv%�K�@�C��[��9�����獃�+�}�H�w������Y���i�&�:-Ć�^�GȨ!�3�8�.}5cgv!�����m��y�O�����T;��O�o뱩r����[?0��&�|�>�ԇE����<4n�1�����1α�h`ǋƻ�~ޮ8b1T��VM7���B�r����ΦvrOv��2���/��_e~��G�\�n��,�=��ՙ�)�����#�AJ�-q_rij/�l�,j��{������m���#����}� �d�)1`�󞜭�
��#1j����ߗ���Ȯ�$�2�:4��x|�y���;M��^3{��L�����s��L���Ậ��gKC���n�>:Zx�a�QC�緷�t좃B�!�?����h�tjP��k�Oe�[&)��?���.����gL3Rd���t{#x� ������<��1��Oa1�|��=��@�oC�'X�o^i;2%�Fؘ+���]jf,��BӍ�g7��$	KX32d&,�1�L�W|vS�wx�3�ׅz�No{�܁c܉�uل��ׂ뭂�?����kOS��P�C:?Aέ��|{=���UP�Oa�
qp�Ԍ���%yZj�,���悮;I&� �X�k�[�8h�6�}i&�*_��T��F�څǉe�;���z�"qD~@�I��æ	&;�����w�P}�[J��G��Z{�f���"&�r�K�P�\�P���ef�E��uIrɿ�K��Y�o�X�EA4�t�AЇ�v�\a�`���([,�$���{h��C�j�N��B0��Ͽ�)r$��b�4W�<E�]�,�x�ͫ�T�R��O&��Q�H�8��Ղ�!��N�Ms���XW1A\9~���v��\�+.J^�=��{y�3�c ���[��=�`_&=����}'2��-q��M���6-�q��,�b��!��-8jQ���~Z�Vf֚Z�N�rʎVJmuF�ޏuT��5I%u��"��ϒ���c]�U�+�"�.��s�ӂun���l��@��T��<,!*hu���N�g��v���r�Z�yzF�� �`*�r���3x�p��*4�+��a�p�'Av�ԧ�W)�|ڟ�/Mn��?Jr�{�IX,Ko�p�]��UT\n��Y��m�[ۦm�_��׌���*�.��J����L���>x�Cْ�>%``��3�!ݜI!�QDKe�����Dƒ#�O�Ne$�Rq���J8-n���Z+�ڧ8�`h�i��)X��cX��[�T������S�۹č�_�9'�Ra��bx��ci��}�
<�T�򹘾���(*�f�����T���炬�����Sh�R�\�A��B.t��{�WA}%ۣ<p���$OvI�5ll�x��������t��8���#��x�U�d?t�1��2y����Te���ؼ��4hH�M�Drk�@*j@F_nw �����B:�����S躰������1:�ri2���c(��N"̔�lU��	��z�?�JE빤�j�)O��-���e+�~����ջ����0RŁ��4��Ѝ��-
�_����0�M��%�)�Oj��_�JVU���8\f'�o�0a��f��S��BfZ��g�|�g�&P^�i}j֦vd��A�m����!�� �y�VM@�$�tq�ľ���O�'K��m����߳F8�\�^'���\jM�K�4`=G)w�K��\���Z(.�5r��6��W������i�6�T��a)�]G[�Yŉ��[_��wjI@l�����JN�{wGUa(������o���ʂ�/��df]Y�2�S *�b%�Q/���8kh�j��3F�����9 (���Z{̿cS�r��$[��s�QJ�Î/
�K��e}0�wPE%�lD��[���i���O1˦�6Y��j�V�������W��i��ֳ�;IV+��Nezd������+���O/&�^�.:������0A��f�qA� k=%gUfq�l��C���$<��/����ķ������$����{��il�|��%��f~���|��9���#0�ɒ���u������,^�C3ߴ>!�p�H�[v�dW�A)F5�@�Fmۖh��r�`��5P �3m�T�IN}����� 	癦H�	��q�%2P3��M��cj;F�(��mhws|t�Х
�R<�uԱ�y"�^�D2�����uY���L��)��ʼ*,K�
T��Y=��2n�E8J5��V)4�#�.#�#ey�R�W�W�K��Ո�����F��X>���;~r��DH ��&�1OQ��G�kta����������o^��&� �5 �C��H��%�n��ϷӽQ�}� �$��M`�S�ǳ/�@�o4����7!�t_��,$-�w��E���
�,�^���c,O|�e�V<�5��g�ٹ� ׌~���1\	��>�y��^$�n��r�\$��C�W$h�ɩݐ#E}��B��]a�tXY?�m,��Rhm�	�Ø��O��� ��mA?� �W���9�I����K����df~��o�n�	!�G�Dh��D-���|��C���ᶸ�y�!-�aB�A���~D!#oтS�����)-Ik��ށ���'>o��b�LaO���)#��v �2eĐk���C��C��R�VX��������/��8����m"5}�F�~�q���O!�-,��4Vjz�O�ر	�r�,F��	��d(�oˏĦ1ŭ����Ʌ�ߕ���Gǣ|�9�{�B3�Zn��*��7fW�y?��r��ǀ�O��d"��7I�U[2U%�*�l�2��j�t5{�ql-��2�d��vK��%��O��3r
kZ����]"_!�GF�bJ�a�V��+'�!4;$���7�M����:���q������0;��3c��i�~�cj#�2A�S�2�`7h	�`p�o�R���ϵ،��Hv��D�� ����a,�����B��Aw��K8�E;�3G�L��7�&f��R�	~� f��DV��{��軂���AχX� ��v��f6���42�JIg�w${l��4���|����As{G���&�'�g��w
P`�2�L�F>3=��ń�Rx���?2�<n.<4�j�����뤫Άp���#�s);�tO�E!�Ƨ�"M�����X���f{���ӹ=�&����a���G[�T��w Q� v�"�J�zq�B^��9�3�����#O����p��s�W񧰣1��{rJ�Ʀ�~˟�L�W��ՅD��Ά0YO�e�X�^�0T���U5�h�����o���<åTE�C��0[�[hW�T��>���Y���S�=ֳ�>����e5ʈ�m.s��#k�p�C9m6����$��4H�٤N{���}E��L��}���f�R���k?�wR۹��ؚM޳&�5M�pQ�jv��eR�\lW_��W���l~"qU��Q]��[�|wG����XJ�B{�Z�ov�&;�1+�NTXٚO���GE����;�^�*�i�Q���XցG��v�@�k�����hS�(er���b���E�/�c��-�55��v���;hD{�8���.�8��2٤p��q�V����p��^�Z���ҙG��aR����ǉ�����d`I:�m�61Z<�%�yHj6a�:T���%���T��$>�XpkHTHA[G��Rb�+_d0X�6@L`~��#���Y�~w�	X�#�^�������>�׻7onVR�.{4�ۜ�f#����i|k�H��E�I��<0"�_k&��QgUۆk����n��f�Ρ[�AD@@j���C����n��~����k֏g]�y���YV)}vG���h��	��؊�����u���h�ހp�8��P�dp�E�%)�$�Z���	K�+×?_fuͬ�� p�.$��K�|��0�kAP�/"Z����}�p��'�ӕ��3��g�bX���u��%�i2�u���.f��r��A����N&Bc�_�L��C��Iɠa6��Գ�0�gL�r:/3`�њ�H���o�"i�۽�F-��]�o�����`�~�\r&��җRP�3�Q�*L����^�b֩F�lC]��ʄ �������q�5|��c�BI�X)�cIz��]gC�V�K�g̫и8w�MZ�EV�V��� �1��F��8����xo��xwrCo�x���|:Kh� ��+�1�7�r�\����C"V+ӚI�C�N�G�8 E9=(&�Y�*Kp��� @�9�4�'K�`�菝��ʧ+!��|G�"j���������6`�L@ȶ��]ʃ�M۟��YC�^�h�����Ɣc��(�y��7��J޼Ԯj�U/�yY���6��
L
	[�^X�^�E� q/����!PQ6�w�?�=��N�~e�ҽ-��{�}$�dla4c�w�f�e\���x˲S����m�{���4������66>�hL�
m�d��2h�珑2�@�
�_���C�#�O�O`��)��%	B�_~W���� =z�Iڠ�#�xm� ^�)��B����?�r�2_��Tޗ�d�l-�U�{�*ҕ�[�jv�4�;3Q$+nۛx��k�z$��u6�kò��.ײ
׿��J}�S��/�>B��|_9	��|����js���$l֑��`̛g��!�j[������%�[�P���ժh��G=�
�%����l8<
H'�o1�A��=��y��ƃ�������ң��s�E!�@9Ap|#�k�z�ꎾcH��k�c�Ym(�$������Ν�1�Z/����}�[n{k2`6��fMK����5avҒ8�I�{�23+�J�NJ�IHe"��)_?7#�b���׿��S��8|���6�z��`���E����t����k��Г�"jX�����l���I�d��giE���w������_W5�0�զ�:W�����L@�L ђESfS��+��� ku=c�K0`Ͻ[鳚$�k�Q��^�8����p�m�
B�q${^�1�oNP�$NX�[7�i�~TIW��Y[Yt������U��v$�?}}�@p#��{}x�w�5K�m�g���m4�z�K1/x0�w��m�~�:z��v��<f�{=լ��w�>�Bm)����/�-uuG��f�^�U��Tv�s6̊6�'/�Fj�Ҏ�+X'*7��Rc&�!�����0��H���6`�"�=Ĉ�b�E4`��Kh2I�v�XS�X}x{�:fE"Y�,� <�������2"���;N��:=}��p�r���|u�T�E�wg�$=4���c��v�y`E��e��h>�e��,��E��V�_������5/g���	�����ӷ�?d ����4����bl���DqS�����P?BP�L�Q2���g� *{0�:1�['jI6=�!�Se���-��������+������>�ܘ�̿^���QC%��O�87�6�F'E���]��`��sI
�5E����ٔEP����/�����Ӹ��ErN���J,cm�yާAN����Ʈ�F���\k���5N�r	p�����zl�2:K�TAB��l!��c}�ϑ:\-�>G��~*�ޓ:�_|e;�����%�,g�wc�U��t�"�F��8��eăE�J���}-�n�����~��T�F�g�����Z���/�q�+q�H�T˯��^#���@��j��(a5��T�	¢��ڈ%����V��{u�8:ݏ����B(����ކ</<��bgu�$u��	~!]�1Lp4>�"���?�q1~f!Fy�^��pA���@�T�A���|��V8 1�Sq�2_�NC0�ы�u̷�4O�V��Ǆu"��Y��2��Y�3`��#c�iB`_�A�\���%���fQnq�c��}^n`y������V�"U��a#v����E���8�%ە-���Z�v_����'t��tH!�k+������v<2v:|��:?S8׺5��c[��+1���Kd^�����WA~yfw.���7,�����w�����<Z��X#Q�2�E��P'���&B(,p��xQ��*J�y�����}�q6Q�eY�(P��7��-2�30�}Ď�[�"�b^�u�Q��bjf�q�!�0�*m|HҺ��e?蚙�.�8��uI�rq�.0���*�s������)�HtQ�/ʹ��1���7��T~^D�ק�#?^�̀�v�%��P����pE7]�Mz��Q?�u�206�s��
1{,±�j�l�+�X/�ǾT���^7�M�kȂ~����NJ���]�~�
���L3ga��7XCa�:(�2�f]^����f�<�v ��*eZ_f���=��Z�y�&�42v���:s�m�m,�۽�m��2�ۏϮc-��D�^�T�@_�rq=|p0��?! ����庯���k7u��A�����K>��h�>ו��S�I�L]������)M!�3�
2� |��Y�����pxp �Z��Z��V؆�
{+ɰ)�%�j(�h�J,-?�Y߶}&�[�e:d�BW�N�
,�����KI�T<x��<<�zo���r�)�,֯6�>o��Ĝ@��`�r����T����ry�+��̢h.��3�;�ßu(�BD�=�<�2�v��3��-�Ys[�൅��'��(T��i�(0��%�N^�w�p]s��Y-8)�b�=�=!!�"(�I�s�����@���S�Xe�({e���:�(
��u�7z*���%��"�!����/�W��u�����$F+����/~s�BA�{qI�ե�M�!�X����èp�t?�-��3?�Z_��vn�h�o��Xjy��Ah�.�5=捤�? e��r��3wme҃�E��� ��:�-����;�*�� }�_�
x*@�2����8�Ya�|�m��ϱ2�q�"�x���?X��T(�������[o/'@�unoWVj�8�r5ɦ1ʉn5��� Pi�P��!��J�W�b�?���C  �`:)3�.gU4p�����oh�A�·�/��j~�B�1z��fm�����𳱻
I�����q���*�Uړ$3�W�ӛ(�Ե2ì�U=E��;���
}��n��H�с�o�ox�B�/GS�żc�pt������ԻUU��?��˗~�`^i��<!�]�<��>m�ځ�7����D�n���	T�-��&����R������T�2`�O&74�G�S�j���A�m�"��g�1�_��EOz��q�[���4=0�_~��x��� C@����ʟ���lGZ�0O^��+�z���ѭ��-���%�Y��!4 ��~��F�܄#� �����:`�UvS��}�-?;r�WT�1xL��6s?x	<ӡs�Rmp�oyyS���U�l@^U|y��I�'��*���}k��t��t���b�}�q|�r�7���D��)����z!�>W��:�o�/��bs	�!�����a	�m	M��Vn.,�g��M��#���d#�sjJ�{����i�N�ka.��Y Y�{�
/�z�����ͦ-q�/�(��v��4z��h���Q)�פdw�)4_�@_�^��U�\�/��ȥ���4�JPK����V��� l���=��������H�}�v�2 ��֔��	@e��Ȳ��l� �@YN_��>;5a2�6A�d�M��f"GObw	���EmM�^�� ��Q����J1[8i����h��'O&���#n���}<]��f���H�$	j�t)�<eC��sv��k ���wF�+x7��{�����r�2U���(�$��Ew����i���V]z��ݼ��'��Ȏ��ǿ�Q��1:��as�{�������&��ݨQ84V<���o��?dF'��9;�A�*��� ���V��瑦¶ xv�pF˖��v�x�%�+��:�0�i�}f=�f���&����2�]P������ ��S�BQf0CM����g�����g���ߛ���۩��jQ�]����-�/".e SP����]���=��KC�#/�%�/G �a�ۑ<h�Q�,���BZ�\^;!����;�o��#
�����**Wܦ�w6���Dօ<=��NP��Wc�7d�Ύ�Z��R��gz-�����P�M���%���*PqCW�ִ�Fq6+0�C:�W,έg��VK���Q^�6%UЩOP�I��}j��J��)�Y��r&��-v�JI6_���������S,��-s�u�t�ZTN�%�H8���J�Tj�M2�b!|г�OIM���}a��������Q(�G�$��6J^�܄��	��E%���7B�ă�*�; �^cu�*xߠG���g5�����W��	�_�e5��������}�,�@�O�86,��̎9������2���˺�^aE^�}�W���r���%�Z����,4cb���ܠ�����ixVle�_��4�N��x����n�8��G�7�A%f��o��+��9�5��2��)��(ǣ�[�y��Y���B*xI��{��i\�x2���8EБ����p����:2�v>g�g$�`�N�W�R�<�tjfs\��,%=8V�M�mv�+��kݓk,��?Wv�h~�n�B렮��I�,l�3�["vq�So[���+�� ^�d���ostOcj�*�8�A��v��ܨWV�%:�3%Tv+jյ��E�oD����7�R��K>|�i2g�B�˙��zC���O3�Y�k3��O��.1�b�͙\I&���^���I8�����0�a�7���G�Z�*)"8�����*]��-�K6�H��ґ�j���C���ge�T�<XL�<�m��ë�
�mOD]��EI4yhU.6@�5/ǛĦ"��H� �r��G��!�Y|C=�J�kI�R7/�Il��?�}!�~�Isw6`�������G������m� 8����%�)!�m?�RIkj�$!4�s�Tv'%���s+�d��V��q�� �	�|Z�uv8����Z�4O�=K�hj���w�F�`���W6�}�+��4��Doע��u���/���ػ7��<�Χ=0�xK<[�����l�(�%�c���CʎE�ꖍ��� �DDTi��G�Y�m���a�½��ߴ�8v0o�.#J�u�=�(�RD�&#��h�x����*�Rw�f�ک3H?�[᭏���[�P�9d0�m_(ʓ)�6UH�6���\��n�4#��B�H���cy�[}�g�^6V?�/.�?���������s���z[�<�9�<���P���2ѱQ�,	��@a�{���i�0��Q�r��Mf7�*Q4�9h�Ż�B�Ȉ����gUԂm�!��������@�y܎O�MZ)��ϋ5B\�7��9�?������V�%^$��u�1���x)����Y'�j��'����~ɰ
�|h��=?�(��9]�R�<]�!;ͧ�w��1���wCl-5����maUB:&e�ɶq��~�o�~T-�J��S�뾹�cʂ~Z�gt��H��ʧ$��[���Y�����9v�r��h�$#��I�#�O�։D�ʼ.a�	�w�?Z�3�K��a����j��ٗ���nҗ�hՊ�X��,rh(�ޚ���u?����(�$�?(�/K��1�*03:�����tك���d�\P�iv��a}�Wעi���k���ɫA�1>*����6�((I���^��q���ȕ�_pW�������y���N� 0���V������Up����;"ޒ��2"@+���2��B?�ӆ�8sn��0_r֐����Z��#zz�21z���כڜ MGP��D�*��b�+���w!�=��&p�L�3��q�C��3�5�^�Qyd{�[)��0�B���45��!m
�E	���@���`i�2���!dj�A��On1�ݡ��%�������gu�.9��DSz�$�q�M%K:���Y�h{�7�k�K8V5>�r(�!'_MU��԰ �6~a�!\f5��DYn.1�H�i��<8�t���+��G\��'�H�9�?`derT�R� F=���`����4gz��̞dD��x>��E�s+p��'mN�3Q$��ϓ�e"�7�ǹ����R�T�s���}��+�gJ�j��r�N�������Tv\�ژ���K�G���.�`7���ߔE����%�؄�c�� ��,��4�C	��1ƹds2Ѝ:����l&�c@ ���H<U�ݓ�_J�L~����&�{9�� /.����~r1�G]����B,�a�3���`��]��]U��T�ҕ_�2����@�;f
�^��L�q���E&�8���ue;���삝�j�S%��>����zy)m�F���X�;v�便WZli๾u�|��W����J�*=��m�$=u:Ne�ǔ�.�b�S��d��	��^��s�>J����$L���=��
vx�`��$� ��qy����oe&�:R��U��H�>e�kGܭx ���;��Λ�Y&�
��t�H�`��=ZDy�v��S���d�3�+;����㷛�7�)���3�s��|�w�__��v����6���q�Zf�C��P�3�������Л�n���ָ��<������|��Q�E�������@5�ld �&_d=7�S���:RV��s*�_A�W��Lr?�/IT��}�tY�5`��S�����êH�!��?c	Y#0�Y���͈gN|�#1�{���6aS��u�<c6��ufLo����-��>���Ge[� *�w�3}���k�Y����1���o>m�Z� �hu}~̰ӳ���dY���|g='�t&/5�5�,y�r�(Fޮ�� M i0a����Y����Hҽ7;���|w@��>�D���{�YR4D?�2��W�JcR�����л�ap��}������E}DZ$ O�=���տ�}��NYĀ*M�g蜺�	=L�3�e����}#���뉈gE���oN�/�"y���k9U��ia}������G0W((���w&�7���L/��8�t�!Ѩ|�<V�U#�K���*�:��K��_M+��_״x%X&,�~>�x���)���˘�6������)�rs>��z��=I�!�0W.��mU`�(���YF첑-Υ3�e�0����g5.6�v�����Ɨ�uN���u�;r/bڊ����z¦���2�]�u��#c/���ٺM�&M�{�UYk�#���h����A	QLy�o�
\��u�^ǧ����p)�㉹�ca)����_�H%�A�ʦz���@�WF<���t�yw:bJM�H�&of�u�*^c�fYW���Q���!�ߓ��#�%P�V�]���>���+�Bi�t.�i�v*�(���!d���{U\�v�h�˶��t#�.���-/hU�ζ�u4��Y�K�����L������;/:BW :߹*���:�K���0u��ҧl�Y�o�`^`�q ���t���B���G�M!��m,Ble�ՙQ��1&i��Ӵ
tHB7æ�9gʊd��|�/r�:c�
I���S�\�#���a��_*�;^�:��d)�p1Q�65�jd��RIX+�����(8c�Bi���"-ߜ��05	q~a&;ڷ����H����h��K�0���.�n3��d��nӐ����X��E�N��*z��H��B�������X��M~�����v�Xƒ��n��覞`S�=�K�LJG9_o�҆Z¾�C��K%�O����~�O�#�d��7��~�1�M�T�V����k4RkB*y��\ ��OF)�iJ6��Q}$�縣�TF�����.���G)�x�j'��t���C��/,�L]�d���f���'��l��'{��������l����7'B���c(H[//GIƎ�\�\o�v'�MV����Ё�K�oǥ�1�y~&j[�Պ�7F� ��+p�@T �d��4(����On�v��=J��z��uz�S�Kh�+I�& _G����u>}ґ�HF��@M7�
�����B7��eȆ�P��#)�L�z^�{��a���剄��}�0?����v��˖�}?�e�n��89.a�Ƣv�1�U}���H^�Ke�ѩ��:��X�} ����UaE��C`��zv��N�{�8\��e��}������_@�n��#\�}w�G��hl��/}�o�Mw�T���q��+�HLVc;ER�c�vI�j�]�9��xFU%��<f��l�^'w0�Wo�[�̍��<w�ʙ����̛�	�7`�����?�rN1��e{^��
���Ndch�Ɣ6(j	��r����ʨ�W �L�#����>=L��p�~��D�K�ɇ�9ә��>>)� �Ƭ"�-<g%T[�w�)<�i����rGrQ�/W��e�udG��~������8\���1��9�
�P�w9AW$N3Q	�ٕt�#�X�#t�
��.,��(f�v�!eM��	�=��A�7�	i4�aU�6�q k>���o�0	�D�����Hckv\4
�=-B������g��awǑ`����Ǹ��q���Y�+FFT��&!���̲\���Q]�,�}! G�C��6.ߞ$tq��\��Y��6N����O�yJB��>��յ=0��HF�����uP͓#;-!?�Y�Ȏ�POR!���j.�QLt1�"�&yN%,-�x�O�\f+@H�`�٪)���c��~�C�ec��8��*��E�U�{?�/1U��¬wn����U�,�B*�b��#���8T��f�sݹ�,�S"��8��F�VH�?� �3���*���4�\I���kS0D�TA��z<����L�����^���s��f/{�]��$��%�O�b*Yɓ�SM�n��es�ŨH�0�~lӧYYl��	��j�Pn���Z��S���^�L������w�7���u�C���]�H��m�ݵr�
����C�T�w����h���[��ҏZ`|�� \�é. �̬��^�K�w������:p�E�� �xb���`w�Iu'V
�M���J-W���`E�*������iy�D�O(u�ޓD+#����Ӎ��U��S����H_}���՘�����>��t!!���?�(<@��R�2 0�
�K���'��@��������P,�dA*���-gC��IhH���D�������I_���@s�_V��E�:��!�]�+��-5ei�^�|���>Ӟ)��nTd����
!Ɲ5\8��ܤU:0Z&�7{��'#|��&��Z�١��7$C��"}������(�/�pQߑ��vq_̖!�r��O ȣlKqrP8�e&e������M2��{��ᇓΟ�(L9á�����2�A�+�T�Z��k A�t�9�2Y���Zo/Z{��������Z}{:L����FX�C��K`�'r)�3˼_)�ws�VTn���X1C�4�AQԐ&m��<XK���}��cϾ�.[4�p˩�f���ʈ����c�`zbY),�|�_a��-C[b�>HH/�>��#��E�@��0k�; c�tm�~�Z�>I
@ѱ�����j��Y�E� a9�<�U���r_��%��a>c�kƖ�J��n.&�_-x��r޵r�F��l=��^WL�H��6�L�XՔ�m�(��Ӡ�c����g&:��/�Z�QcE*_	�)�c��5�K:r��s�p�C�|^XF�u�Uwy�p#Aj�\����l[]/E\�lk�1�_p���}����N&�l��(��%�|(��un$��f�����+bfM���t��ey�R���k�����P��A�'lI��(	\3�L�s�&P��"�m���>S4�>�
�#���Au:�(=qd�MQ�kb���st�Tp����������q�2�j���\]����ҟ�;�)�F.ɝ�\���)��h���Q)�-��K�Y�ޔ��I!�1k�W�B_g�����d��vMEܙ��t�n����[�Z1��+wIb�^�X��x�H{���(���;/�mM
2�Q��1���B��D=Lsߴ3���D'�cD��4��cV�BXޅs��c�ՒJ�L@B/1��&컌	�(c�!�Vv!:�����p�mڄS�+� ��e��P���E����1������lF�W�ӈ`��#J�*߳3�!�F]�����b�}��u���ڑ�ٍl
f�ZD;sjR���5v�R��5�ؘ�[f���!�"k���~ɀ�zW��Z�W��h�]h��U�L}�O��&����LۨJzL&�a?��D�u2�k��
2���)$eꮕ]�c�f�.�_����=�*m���-k�����"x��_wo[o��xF����̒��/�з����ޠj���;�B���;�
ʣ��d>ο���F0��ԝ:"w@�uL�Yv����S�UQ?����=���R��K1F�l�B��Z��VOV��q�w�5� bV<,������Bh��6%1��tgD���vu�Y��ޫmnn����u"O����>����'����K�V`�t�`����%)�|�S��q�q:����AR|��(ӻ�g��%Alס>lRE%�v�xHmBհƖ�m L7xsY�i��FW�D�Y;(���p�6��M�EGBt�e��Z����-�l�'��A�@�誁�Q��,|��uܺ��I	�>�B7�U�G��,��8��ݖ<���9�y���霙)�@�d������s;� �� ��Z�;��m-}k,m�G7~�_�˝u��E���f�n���$�+���e44�<�*���I�U-���=��R�5]o Ԍ��.�w,=S��ڷO��1}2����!�P�Q�ң��`�-n`)�?������[���7��PqD�5)6�۟���2)稺Ӭ^�w�r��w1������P�M��U;ch|�f����^��kE��c�~����2BČ�ժ
�`kV�I����$6�~�s�-��2v., V�'+�'8o�LF]��I���������P����A�c]e�?; a�]�߻e��z�k,�y;bnw�Ƒ1(���>`N��,�n�y�,Ȥd�u��O�!`��ji,w�AÞ.�ڼj�V[\�J�g��.�z<��.�&�U����Q�G�O�7��� �I#Lʪ�v�n���F�oJ��d�ud�Fs��|�ؿ���G���/�t
����+��{��h����6��vΔ��� ��+�  ;���Г_�ɀ�k��Q<m�<�J6F�^N���{�0Տ��?��1G�1��1��&k΁���Ԏa�dwq7N˃��j�;Wv�%�aLp������~��x*6{|�^Wt���M=m;��a˼�Z��{�_.mu��V��wJ7�˾��A�"+0�5��!�>�[���:z��B`" ������ةqQ�?��c��(��8�
ѰlIbv�*LE�p���I��,���$�G�4|~{
�>�\SM�(a�1xE�x➛~�A�;�2�ӫ�O1ν���aza��a��s��ˇ�.�������ڽ����z�ߤ	p��ɜ^i8Զ����Ld�t��>ș���ʉ�$M٘-���u����>R�AJ�z��l�`��ߒ<:W�^ɑ��o��)7��>��&
�Gk�XJݢO�����t����r���%'�ӆ��ܜ��&��091�[��,���+ iD0}��/�<Y݄�>�ۥ}�������������n�覤2��L��r^ï�p���F7�E+e-P����4Q���vVA'_�A����ix���|��� �
ͻ����6i�F�w�Ǳ{h�_��hy{��UapN�1 f,������$�����)�}��v�Zf%	��ͷ{�5��ίh�m��] /��"6+�}#�ĥU�����&m�bC�ǖZ<O��3��.�O�+ѱ�ׁ&
�J��U%�⟳���0GoR a|0�;�U�r����FԼ��M"���Ƀ�`�\����֗��?���<iJ�e�m��_����0ԤkD,ux�)�篇a�l��w��%l8��	\p�֌�����u��%x���'H��Uն�U�(������(�-/(�n���DO\cF�������]V��Y����	3,��q,:����=S��W��������7_x��=m�K<(�ur��p�����Fv#1�e/�-Ef
d�xVQv[X�f��Bk���*t	�НG������X�0��3rt>��O\!���-�ܒP	P&����gSc�=���g�a�U���d��䎄і�3��~���!�2')dKKd���v\�W��@�b�e�����ݹA�_�ҳ=�x�U���J�Xl����p�ъcە�2<8('�0��>�0U���W�xE��西�IX�XoYԦ�1��h�d��p�/^�J�lb9�n� �X�p��~id�o-r|y�	~2�T�/9�iG	�[�I:�NЂ��aN�@Ҡ���Q
�guʇ����:��Np���g��M?z���׵>\���(Ʋ���{;�S<���N�Zԗ���M���7I����qׄ�[��q-F-)�\��S��'!]Y��*F�=���R��'�
J����c`F}������P������o��_���8�̔-~���p�9�9�h�l��u���P�}��� �V���a���%v|�A�!%���<������ʺ�-���OWļ�j��ݦ�H�վ��j����Ĉ�����B�K��_0����N�@%߇�SX�;�-i�t?�Z�VF~�HaI6؂҃Ftڍ�&��D���]��!�E#�2/��?1�k�H�u����G�U�(g̥ר:�,nd�ae�t���S�^.�@�
�_�{�ք�~@��{�a�hO.*y�Pٷ�w:�1:2f#-�	i���%#��)�����o{�'(R3}��bV�n�ID}�
�Z��|�;���Άa�ci�N��z}u1ח3;��oh�/�E�^�9�+�)�:(�E<r�]FI�D��!��^�N.g]���@���ט2��� I�#��T�V1ۮ�7^W��)C�v�cNE�I>[��M��0��NP���;eV�y�G�����w�a���T*��L9{n�'=w���B����$���i��*��zWtn�L��A��̤����ԕ�:����iT9n͔�H���n�Z�0��+r-'[q���Ϟm��3g,�֌Jr��-/0L��;"��|������:*GX�T���,���4f�{��������_]�K1�"��n�$�(Ű�����K*��ۉ�Ī�>���Ք��IN���qH���2`�q�
K41�2�N`���Ee�,H�-���
�bS�'�0}$��������d���}M6��C��/^5��� �H�	=����Pq�?&gE�╢cB pzm�#�$�rv��GY�m뭯:�@���}�vv[0W�eyF�u�5_�!p�t���ē�������t��h*���2�_����δ�h��B�n�������K��]����#��;��S �`z$1��s�+h��J7���$C�	�F�R�xxigzA��ѳ��8�I�C��j8	E�>���8~԰ongwh�`t���7��l2V��e��b}�2|ˤ�g�b�MI�N�Y|+�^-[A�V0�c�/�B�d��j�d7��]b �[�'$�e2�\~^�^۪���m]�(�]���;�	�AYY:�
�� ���+q��y����]�����Rl���H.��Ύ4U����ie�}�x�S&F�cX��O���G�Q:c�&�z.N�f�V1u��ѹ���2Ѧ��������ReQ����/ƪ�����آ�S^m��3K��JJ�H�v�1kF��а^9ߠ���Km��.zTCf!�i��,�jؑ��(����<5���� `���U�����v�M�����m[��K^�GW�}'B�&���IՓ���G\Ydu�u!�m̦�	W���L��S��0�wQ�NPX�(7΃`	54��`��Uس��!�E�șX����.Y�0��`㕆����F���^Ǿ0\?�/���[�8�diOb�{�;��)-l��+�.�4��Ƶ׻P��+2�漳|\��c�Ҽ�}�0�WЈ�NL=��\^���-7�67��o.��<uy��>t��.?'�6]]b+��	L��6��9���<b��
Tj����m��݅�g�s��|���n�����>�3~KlK�IM5���g_�f�]A��N_�v"���k�sTə�ð\X+Y��N�Z�PK�0o%H1���#E����q�8'"��ߓ�G5����B�S�S/�p"к���#"�Ͻ��$�?H4k3=|V&�V�<��$��*}%��N[	r�ƸY���d�1"��}���ܠK�/�wܿHMx�f$g��fwhΣ0E�V��]od���H�(�^L3e����=;Q^m�ZO?,o�N�Tns|ޚ����#����TI5���lr�����|-8B�M3�"���k�-h$��[���пM��ž����kcf�����dx��嶻�B��;I.���K�<N�Ϻla�ż��0JWh>=�y3�ڢ��� �vύ�vP؀���#*�o��r���M%���7k;K_���Y��v�ZrO;�S�F��"��O~;����ɴLU���6�ˍ�C�T�n7O�l��w\j�����S��U��4\��fS)��aۑ]�y��)�Q��_>���d A��)ޥ]���y;�bh{�6��p����6ٱ�73t���֯B�^�B?u4c��2%8�~W"�4;f@^U�)FMK�����jC`�γ2�Oxq���~��ӬM��JS��-%��y��La�6�����bm$�"%
͏��_�ߖ�O�8�9���V���J�%�~L����G��G���������MR��F5���q��:O@�������O�R_Z�{0v�y}��+�Z�aɿ"1�`����N�;:t�l���V����B�Q��T�9%�zw�+���%�N��jsR>p�-�s���n�Z�:���F�Wv6����v������!	��d������l����$Yq�}UQ��#����K��5zxՠ�ee�Zl�cD��?.�]F�7 ���'˺g�d�!����(�����+�/R+�
s��v:�b�>�p7��6Ӂ��n�W����?+;��9��ީ�����l�4�H�E[</�w��|�V}�g"$��!/SG�x�=`��X8�� �=plH���,�P5�)��X�)�
(�H�¥C�D�z$�oa�`Ym�y���D���]���ΌO�⥒�>U��D��q,;�1 �=��G���]0X������W�U<�".�TI�{	��\���q/��E�j���#HA<�r�Xe!p�n�ƺ��7/7�|fi����S}�6�B5���h�-q��q�x�q;� �i#9(�@�Y�� �"8��B��  ��<�����>p:�*�ƽ��{<O�Y�ٽߞ�|�]-s}��./{+f��c
�h��3m�1�H��ܟ+Iz����(YL3T����0�K�F�~�f��#����*�Zlx\Qĝ����2~���=�A�(w�1�Q&1�k��G��-[��l��~����Dz�X�� o�Ƀ��S�g��!�:0"-V�.�n��4Jp���w/��u����u��`p���X]M��p=jy�z;�Ŗ�.�3�f���4�z��AKB�G��=oo�ɎA�'� @v�K����Hx�W��3MA�ࣄrq��6���[$� �*�"oq}'�o�vU��׻Y��t| |�ea4��U�	/I'}��޶�epSk�������۔ר���V���r�Z~�꥓A ��&4�	���8���:C���Y+�Yk^f�/8N<�S�~�2�7'!�4�Z�������:���^���)���`l��8^��D���i#�d,��~mEO� 	���y��X�����F�9tʅ����$d�&�(ҽ�� �ʼ~U5�"WOu:�~�^�Z6�݉��%���IJZ9z�c"l�N��@�'j1̚��f_�Ǽv����;� ���:ECve|.�S�U��i^�����Y�6ף�짗�v��ZF�1�>a"7ը�H;�K�[��,K�?L�e\So��AE(�(1@�Q����c�ҍHI7������Iwww������fۋ����yv�����<�1�H}c�� A���Q�E5�`�����}̶�$Uv�d�) [�%�*��9�R����R_�7,N$!�#4�w�Hn��W�o���v�F(��^^������Mf�_D��_�ӝ��$VU����w�m+������b=u��r�������D�7����nt�o��܅a��U%֐߲���p�C�T��T��6��L�;X�7���	J��Y�pѦ0��0��|��?�hdKZӅ��]D�!���-p���-&6l��6�P �������D�Hp<�ѥXBy�q ]F ��v�I�_����P�,�)o�6���q�N�6�u�������\������/w.���Ki�b���=�\;�2ꉶ�\`1�A�B��ș�0F�2�&	�!~'�h	���}ג�ѡ/�<p�ڛD���������T��V�����������j���w�UZXB,�_\����`Az�,�{���<��	BO�V�@LK&?������c�~R-<���׷ln��ė�����`IN��yJ��qI6�B/�$��s��	����c7@���{�D�i����ӏ%c,M0����ٯ�_�����~W���p�;�fg�S��6��<u�^�f���&����I��\�l����8�����3X?}N0+��}+ǒ�pn(�ߞ��@�y��}qQ�
���w�QP�;&{��u]�/Ja�Ĳ�ۉ>R�'����&T�P&����m>$���J�BL�LǑ��Q3L�в��?H��F� �m虖���d ����VN�H��T�[��vvؒRq�.Sn��"`�pf���?TQ��娧��B��$u.��}ACA��c���pmB���(�m�Ƕ�#=��0���1�=������������^�����]���<6-b��[��Ej�D8#z>����h<w�ۡ�����)�Xe���-c�pL����`�����ҋ?�2ތIƑ���L�?6;,w���Sn��rw���u��j���~�M3������S_�l(�$T�z��+;P9f#0��/@-]�~�ҵ�����T�,o�E5�\�E-6^�͕tlm5#�(\���gq�X�����|������b���w���
��'b�����a�4<aV�k*��u�x�Ur������s�f�����=X����KM�T}�����P}�U��S��93�ry�VQa04�s���}�W�d����j���9WĕZ�h'f�������s6��N�@>"�e�6'@ ��
�a`F��Z�ov��l7dB9�?yd��ԝ������a��g���y'�[27��F���J�h��a��,s���f���ek�ĭ�a�Lz?�+2�!������m��i��aIV�:4�Q�Ҳwо�����O��Q���m���׎�"'L����?so�y^�����y�����ο֧E6��?G	?�3f?�;�b�'��i�-YKa���䆞���e͑ɴ�¾ӥ��,�V.�Dg���/��Q��Z�$���.:X�U�E�u��j��Ia�XwyAqPX�����)C��`)���m����H�`!LٗL�49�ɬ��b��wӑXF��ϋ0��F�UR�A�=��7�&�Ʒ�m�E�+��Ro��(t��+r��9o1� ߪ�����V",��l�����7�y�� �(���sl�i< 1&>	z���3��]Y���r+�f^
�� ����R2p����;�%qVJ�-v�����g0Fq��h�i�L�e"��O�����������k��N�h*���D��n|vU����i� �+�2�� �����s�ڊ��1��zan])��)�C��������D��ߛ���\٪b:o���ޣ}uH�����9������%�w[�M��m��_O��8��>YGx�����{���h�R.ym�ڙ��
=�ghR����3�yX�v��]'�}\B�?h�Su������%8�58'8��aB���,z��4DgP�����a�zʧ�P��=���m��G�=K���T�1<!����N��m�A����p�30����pv�o��vwր�����%�˿�I
��Mw��gNZ�eE�DF!'���o6�	��í>�J�m[V*"^1�,O�laf��x���4E�:U�zf�X��^xF�����A��������~���K�4 ���H����n����K3)0�8=+#�$�]o�������c�$��kR̓�=�7"I�_�	l���f�9g��X�"�{�d״����U��[Q�ԓ����푵B3#�bIl=aT+h5T�!9(T��o2�:o'�Z,պ��p�{�S�&-!�/Q�t���R����܍�U�����Ħ���{�{������3u�m�:1L���{phZ��:�S��Ɵ�N��Ni 9ֈ�n[�%`��=6p���!�w��N��r��+'/��?�"j*o�Uұ�`�ZCѻP+��s� #�Y6���5�0�b�K6�ܢ����K���f������=0�su�:�e�c�K�s��66<�Z�j�B�g^=
�Y��D��u0������
\1Y!�6�Q��zY�5w=�!@w��^�MZi������#���@*��0o��x~��h����9]}�A0q�g��'����WX��F2:h�o��?����b���S* �ӺeQ�G��F'�rl���)F�ΏA�N���->��(�Y����+���R�T�ۓȭd��!/���G�ҩ9j�� ����0S�wԏx��
�T���8��A��0�W�Rx��B?�����3k���F���/5C��4+��Y[�z�1�����^i���_CJ3��9��W}#����{�C(�u��):��'U씯i��4���v��m�g�{�-(��(�۹��O�g�E��QXs����!U��2��PZ����e~NYl-"��nĮL���c����x�����6?�aZ�����/$��Q3�+�h�	�=|V>hga�5��j����5�9E���PrY��i�r�ͥ8����� s�p�+�\aR��m�(���.�u���5�U���U�]K�e,��8�Arl�4Q� I�Կ��d�p��+�l 4�v�^4�7�?��ϿXmK�.�	�ycb�أ��WS����#�����Gs�-�E��q�	������R�
co4�>��$�o���S��N��#���B�PL��6gw�Σ�o�>�c��~� ���w?1�P>]=�GwP���i�~��K/�.�A~������ͩի���+9��]
�hh��IQQ�����?�~ȗ�+�p��md��G1E���'*w*��O�F���:W�)��4�;s�3���
�3>�mtFfP�M��I��8���nv�n��[��H²D�1�sy��h�<������[���ݻwmQ�k�@0堕±���"�ު��9�T��-d��#oR���&�R}�;(}Ɲ{M{���F�(�iV�r�#�+��F������C��?�"�:o���1=`O��a�v��v����'��0�5x7�<x6�!B�>j1+�ٯ��X�6��)������ƣ���Ŋ�냉:�XCݻ������yT��	u��y�dr/�	�/�;B�Z��p��ySqu�u3����I�y���$ϕ�F���#Ģ�]��^�Q1��jh����8軩yӭF��y��FU�B��~'sL��4?Z��ʓ�W��}%kQ �svb�܋_�&A�G�uF�*�2S���t���0Ӿ���M��r�X����^o ��G�r�tsc����f0���3O�\�(�-���Xj0������~�����Ւ/�P'*��?��o�8�����5x�Le�$��n���➱�+l:�
r|u�J��:g��l'��l_sN��'
.��YՇ���Nf������<wtX(��B^wW���t��w��D�>_����(aU�E�W+���	�L)����:�B��b���_���r�O�'�~�q9�zۿ�~���_����V�.��r�{/1^���+C�3��.���kq�q�D���mF�����H"��D�dپ���r����A�z���kk��Hb����5��L�a^~����.��@�TC�i�������5���m��m����-���Fg��ly&��a(A����̓rq���UH�´ ���s�b��V�ݯ"tFSjO�9hZ<�F3��s�.n�.���y�T[�̅+��X`�It�ɬ�auљ��JU	L�]'ZA��ɔ�XT��M��[����ӳ?���ݶ�z��>sq�������*�ͨZ�������9à�l�.H+ĵ�SI��Q���vsk���Ga[,�Ku����Pۋ0td��T\���)�����B��W�X��|���lEj��Y���X�L�9��L�^�Nծ�s�F�#JR���#'�X�*X��u�rN6�Hoۼ�}E�'��Ʋ��iQ�.ے�+��jZI��DX���e��9>[���B[CA�H�L9, /M^8Sic����_��E�&� �4��$�!��޽�r�d֣�<�}J�u�Q�26A��b:���Á��*_X������S���8���Gu���&ԍ\Rb�F��$�;��^3[ #z��Җ�&���4n"R�ʉ�n'A7e6�c��
`";`�+Rw��3��\e���	@��0��>����%��W�g�{�E������S#ǹ��zrˣoko�mH����k�� +����Q��&�F�T[8�R�����x�r����{������������˄�HE��IKc�VY�cnKB���Ye��h	O�X)a�.EE<������?<m�_̿ܬbK�"�.�]�^���3�ܿ����t��Y����Z����z^�`��OM<������ֺ���認)��#���=�:����Z�����@e�"#K��#��D��JS���V	�:T��Wc\�����>.^xw$Ѵoi�,6y>�2�*,�{������4�}�]m5R��R[(����n��\߰�[[*'��W!�@2s��92Q�׏�6V@����*?!7�����ʀ������,x[W6��;���p�v��+ԛo�9}��F��|����܂h�J-J�8zh�M��l��̈��I�}���Vf��������0�Ff���ޖ��Ľ����c4�w@�R��b�X��X_|���`Y�Y@��@���i����ʅ=y����_��;)�_Ͼ0C ����Ӡ�	3��7kK���(o����fɘ�0lD�j^��W�R*}�)H<�6ӟ�4T_��g	h�	Pލ��a�LI$�YB?K��XN��y�=k�?l�f���O:q>�����$FZ3����L�C
B����Ǻ��t�T�Z�֫.k��r'�a�:�� ��z�b��VbA31M;�We�ɼ�"�1��}a�Pj�ߋ�9�;���lѳK��h�p#(����1$Y�SJ�sh"�X��e3G>@�4u:V/W	���3�R���P",��l��F,dԖ�y�ܝ���iqCv���z�X��s�*�=���.��-��f@������T'���m��pn�rw*{���I}���( 3��c!P?	��ocx �@1� �߈ԫ���\�D��Ȍuc����0F���Aj�0�1u#�:���	lr`���U�����˖�P�tL<$Ѣ]/si	I�E3�݂�hƳh�^LY�������/nM�qY|�L�)���\D��R���� 6���$�[mR8���nY��"i��,�TT2�9�ޏ�\��ݢi�>�x�Z7?�w|�bɜ���k]�Nl�Z�6�I(A#�K��Q!StXk��ā,!��U_�����U\��V����C���l)�D���g�ZJM ��]����)�T3EZѥ��8͇���~Q؎[[X:R"^�E��}ʐ�w�6�<{��<y��{�xH�	�!@�{>��u+��6����*x5����n;��33QE�M=c�a��iI��n7b��>�fxd�ū�ES]$��L{<�޹���urZB�&о��{��Dq���R�=@{X*���z@0wB����`s�7��(�Os�d��B��؇)��F�1��鏱�{ɝ�X��i��T&�i&�鿚�����6�b�mD��_X���������x�[|�뻚�x#�<z<eyly�jA<�d"�-fZ���V����>�eX2���>D�S�bV��FO�X/����u�|'�t���5P���-^#Y�&V� YT���T�;(>T�;�⥾�����>�7h�<J�Z.�|��9����׫;���`1�q��xC��@_��VE�(�.���⩪��i�V��7���9p��TX���x�����E��>Vׅ{@����}��q�ӱm���y]��Oc�ʔ�v��!E;�g{��'Z�����ŧ̉���H�^�L��Ilc���#��>|�GqG�~�7a%-�Gk�vK�'��hf�M��+A-u�J^+��>�o���j,��a��K������mCfL��Z�a�Q���}
��Q�_����|2,�2|���;��F玴&3�aus��\���.�����4�4R���v�r���|죻2L���Yd�¡�< ��F=osLp��|�x�Ҵz����W���� ���+`�s��,z�M��]��E�Zr��KG*è�+��H���Z,��dEs�i���,L��sۤ�8pԏ`�?������lg��)��b�(�ϯɑ��b6O���D��+��0"fO(V�!��|�s��Y:�XT�c�3�-�/���m�U�sJ���Fevm�\����k �r��{]-?�Ȓv�\���%܊Ғ=�u]�e#�y��3B�4��j.�Ӊ�����Ձ[���
�\�4�-�.�B��φa�p�uh�V�g�tӅq���*�P�U>|g��BW35��"#�8	�G����0^&�t��t#l>F͛�>����4�+�� ��?x^h�<a��+�%�}Q�����������0q�;O?�~�2Z6��0�Ԭ����bG��P �n�X�{ٖ]�<�	�U�p�u�[��5_��xF�EP. 8�`����y��Ͻ�8
7�~%��k}�	���,{��ˤ�Z5~��g	C��}kr����.�0�b������x�:�h�����:<c�b��ʇg�f]L�4_�w���Կ�?5c�>(0�9k���"�(����n`�4^#����bb��Jޅ�jq쮝�3N��>�)6y�Q\c ۜ�*�6]��O�V���f�����ܠ�o�A;���EP|��NQEK536��:"�a $඗r�9����}���#���h`��c���m�������Ƿ�g}�W���1-��'�Ȯo]&v�};e���y�:g��Z7%���( �ϕ��eF==����^�<^��p��h��A�		\
!/B}o�Z�ׄ�|oX�}��B��G�Ǘ�������&�M<��ϣվ��bɞ�5��M��ײ��$�z�P�_�x���e�WTn^�6Y� ^���l�?��zU��) #�PAF\�6zW��3�~ӈEˣ��VI����D����f�O�c�7ɨ�t>N�z�Fkp^n�����<�	t���a�>�yG�W��K^���om��$�[7v�[�{l���~�B8��N(ܨ9�B�h�>;/j4CN'�A�v֚�\-rNu�+j/|�Ҧo��{�Y���V�A�4"��}���$+�S���2��.<헚�n��lE��d�̱i.�+��ǘ}!0W�=��G���%���mb,녉�.�؁��0����-��euC �����&N����j-� s~���I�6hy��'-�9��O���;r��s5�cmQsD_�0`�d�ua�vep�'� 7s/��L}���<�"��^�c@�+
��^e�/|A�V�u��Jس`my�Eܿ�J;N��&t�Rc�n6��y~PzZ�]���`���n:
�����?��WJ�qSh�,Ղu���>$��La0�~c�zqu�*�yFfM�V�#\G�Ɏ	�����P`-����O����,(p �8NQ���i�4,�s\Dh����"��Ya�Y|J���
�5ε�3t6ೕԚ�z��J�a:�g���$Ǥ���%D���j)\�{&7�|t��~b%�ٜ�Xr����&�'8�4�qc���ON�}>z�R�� �*w���ʴ�S�jhKH6*��Ot�0k�Ȯa%)Z%b�����C�4�$��/�按�	���y�{5'j��m,B�߶�Rb�a`�*��dpk�<f6=�ٯ����4�4-z���ꑎ��J�~����]�� ���/���4��DS��r����f�Q=&�KV��]�*���x��Ǫ����`ߴ?���۹۬���d�w����/�e�౏m�J�"����ˣ�J?�
�R�d ��xԗf�~�N���ԯ�~Kl���Ifޗ
�����:��:���Z�2rj=��uՋ�Uơ*�}=�"+ ���v	s1��{)��4��f�7'"���@;.��!��/�f��
��H����R�;�U��͌�5`��0{�_:z�=.>'>�����G�\�����Q����}�M�w΁Ey.u�[��[�*�|8ae�d?�22�^�`��}R�rUQ+,��ؖ�<�����-|�'ӵ-�頙v|�6v��M�3,�����z��U��� ���)-��U����t=�����_*�{�>����P#���k&`2�k���g�`qB��W�^[���wa�a��Y���\����Ȑ�0�j�П!��>;�C����D���MhOh���>�F�PUs���N�@��f��]Q��sc�RB�u�6S�u������(N��C���k�߭��3��6�ל
�IڽKd4�ts_xƴD�),g����F��]��fT��Myǳ3Z��Y�"��]]�9B�o��	6���r{bQ���6?��}áF1�X�Ǚ�д�N�e���c��qO�ْ����=�~���}��{�ʼ;��x�8�x|��|<�G�zh��8��Q������Ը��HE^��^t/=n����v�Qb`�F��VH'�Z�:�զ*���ox�rϘdŔ��3ˮ�3ʅ+�e2ʑ-:� 
2N�Zխ���-�T�6(�*0o��/�^��g�`+�6#z��>���!f��Y��<����5�͍V��� b����f��l����*���aY���ֽ��R�ҧ<I��D�'D�(���K�
�DRc��F:$&���T�O�<���Tuq����Hؐc �'?�Xo�'�$�����]D�W���f�T��w��|��N�`/�R��=���A�~w�?����n������I��w��qxU�#|.�nZ����'��н<�뽎s���y��/E��Wx�����i	`8�g��rl췜;��v+�]�zw�̈�Q/6w���	�_����C��שt!����ؼ�evC�,!s�}��.�M>�@���'�����@����<d+��F��o�oq��Nt���}�r�v+���b�0^�l�N�ۑ����v�����ds��l��6q����_�9��*B)��r�@��)L�c�ы6F���"|��U4�����&J����B2���bTϚ���8�d~`��d��ޓ��T�Ѻ-�����|�I�!�����z�V8�$�ńcŊ��r�Ip+f����@��϶a���K,܄%��f�� �����2L�>)��NoL�X��]�m��p�O(���67݅F��C�'y�k��p�����4>`浢1�xx��a�r��S��va�"+2�d��`�P�y�i����/.�6�+�'��eA�+�<��l�	�����.�:{={=��=��=w:ݷP�;m%8��-:��Y4��!��j��,	6�k@IE���}�P�m9Uc�J��I��2��ng2c�6��,@�����L���l��4Jl�Z�Q�Q�5
`|%�F1��0�(��d�_�a��+���G�'�cY�ơo�P=���C 
�6d�O��g��̒�>J��i�~4@a{�&.	�'>˨Cz����?"e O���|mr�b��&>�`Y��ȤS��(b�>���e4���*�NE�1���@~S����x�$�Xԅ����b���	 V�AT�n;��V����k՟M���X`aV��$:�BZ�{3������9�G%��z,�K��gR����;�zd�"�A����o�M���Մt2��{�ε�~ؚ�"��8=K�F'X>\�;�qxݝ��?1�
U!!r˿���)<QH�qx�i�w�#�HwU(��em��˳��z�rkR�2�>�R♱Z��=b��%�X*�B�H����.�������t�i΂��f�b���9Zt>
H�_�ٔ�`�?J�02�]ɝT�����j�,0Ux�:dB��ކI_M&yl���N���G�]Q>�[H�.���V�<��]��YJ���Z�����98���;H-bP��t�$J���fH-�A�5*Xw��A��AÍ<�y��&j�{�D��B����ܒ�C���=RqD�b?�b���#�}��[��[��	������}؂��Gi3Ğ@�v��k���C���<fؼ��D�r�Iא��5�$��!U24�W'���Z!"���/�e��ia`E�f ��ջ���P+�nl�GVm�|�t�
���m%X����E�k��V��m(,i���ms#N҅z���c��l�I�A>({��w�� 7RǤ%q�ݼ�&���j�/�TuK�J�M29�?�M$`j5����N¼�ta�;g���,@di�����8�&�v�4�L*sD�֘60-�Ç������Kk!�q�>W���Y���E�g{�˱\������xC��D�j�+Mo'�y��� �Ts����Y7�7��K(��
�!�3����e���#��g�N"���_*q�?���U&�5��'>�v+����`�Y�18F��ps�5�s�����J���� i��z�����\�s8S.��^��6��gH��B�%�_�/����U;�q�R��ܙ�����m\.[��x�X���
�J >=?A[�~��RWi5Ro�v��i.֬�v��
aR�k���h���Y�BQǱM
���*�<�����&�1`z����}��>X�yt@����T����āWֆvߥ_�s� ���e���J����U��P�!�������M� ��c�q�*V����I�l��I-^�5��I�[�q�T���O����y��\�>�u���S�8�m	���P	��r{q��&��7Y���"U����<�� Yj����
�p�����D��$������7�O����P�EO/;uIZs�����Dm��سZD>����V�O~��0������S��}���C�h��֨A,]���@��N��5R�C
�:i�*s���a�W��(���Lă���w���7o�6���@���|�����U����1d��+cv��}��VY)���r�>w�ۉ���O�>��׎+I4>��q�[����{�Tk`[�t����RC���!���ȭDIm�.�@R��$����C[�G�D`'���*�>픫߅z�&2v��O4��wY 
ݧ�"���*��jI���4B	z����ro�qE�b�(�=_L`�@e���Z��������!�Ɏ���.�	-!W�¦���<F8J���W�D�>ͬ��*0dLh���2��q*�8�?�t�����Ȝ�[˽���Aq��e�o_yRO�o��͎g��������ד�HoϫgG���v���V�K}�c�cb=RFͫtU#��kG�|{�q�"���U��2�������>M��핯�.�������;f�����,/C�1X�����|���^�b�q�1?G��"��?��9T?w�xA�z#�y�4��rE|e����v��2z#@�'�C�^7���*�1��S�&G��Q��Mμ�\�o��;�;�N����zHF���ZÔ�>ﷵq��o�7/�|�R�.��!q�U7��`t]I�7�ia7�是&sǸeu��m�����F��W���f�;�g�������|T:�
�T�l�b���g�Ķ�$� ����$R��3q�G�gN�)��c�g�5���9a������9���a�|��j[���v���jtM��y��B���v�>��uX�d�}9�Q�b�M'�<5�̎Sɼ�����T�օ'�)�H9��u_p�x=.��	�8�M�l6};]���sw><�Y8�%�WI��T>yK��`}���aiD%w��h��|���R��S蛖o�ɫJ����\:2�Y��Hj����/��h��ߨE���]�Q
���'N|���DArg{A嬄�<^�a�T��~-ezrc��m0�ȉy<Z� �,�6��M��p��Õ��C����њiJrC���ރޔ���E���D�����:Bc`�I�Sc��b��M��E��Qs�w�oQ��O��R��Z�F[k��y����:�Nzbp��T�P��=!/;��C��m�����g�7��d�~Ef�{�m����׻!M��g��A�	�[y=F�� ���#nQ���/_�E��4?�0��U%Ӷ���\NM�s>���^?�!���䖊�v��V
ζ2�\��ˣ>�C��k�λ����R`�t����_֡9N��[�z��r��_���Lib���v*��p-��Nts�3�y���9rM��!�;H%3���Yr�IB>;�T���q���-�;�Zyȗ4��.̱n}�9��S��x���_�&{3}�oJ�4U��%B?.`�� p���7�Y�QՍ(5��΄-�&6vDѱ\%`�7�]��.��{hY[�(�����?�<_���|����u�~�MX����{jD>���<�n��}���o�.̋���<��i,9�$�al�;f0�%�=��	������:$����G~�8�;x��8��56��{����o���Z�6�w�Ҍ���o�GY�<��.X�	��;S��0ls�pA����o����xJ}�w�cS�q�����7�)����F�8X�� �3������UbP㾆%�S �w[(�U�,b�6���n���˂bӜ�n���N�cxէ'?E�*���jG�|1����M�P�8�ї%� CI��.!q
�q.@�ʘ]@��k�q�2�y�2.T.e�&����Z�CՁ#4��yYI�G9��M˯N(�G��D�]��p�u�����㘞I�hă3��r��i?-�h�pq#"��bZ�*QFtP���;�0[MW��0y.� 1(:�
Dw�~F��"�O�QB&�_*��m'|6[�K���4��!#(]�@��C�w�	�WMdV9��Oʨ��s����#�+V��V�"�����^ɂ��~��>�����i��簡�������S���_|��$ s�ku�<�U�� <x�#�=�C�H<T"7Q�6QfYI��3�&�4�o�)T���J^)򾭽���x�Aà��U�����t�~yY���~�,�gQ�x��)e�r�*&Q�8%�H��'h�d?��^ѝ���8�IC�s4�>�f����Y�;olO���kA���^͸T&�q�o{�U�u9���[aBA%�sm.�|:E���]h�~�&,ߏ�8��¯X;�\�1I��_lg�|�Vg��� i�GyrX���\�'?(�:�K۶v�O���5����]�,�!�;m��Ҿ��b�N��J������/-�[�AB�:xt�� 1Vho&��o| �ݿIc� �p|���iک���Ya��_w���&0��J�<�� ����1f�A¢Y5+"�jy����='�D^o<�N��2�6��1��2	=ĳ��P��2pS�u�*��I��w��-PB��;�Δ�g5A�?�y?1�keB}R�Pv��?e#Zi�2�)b(?��}9�%X�����xl�;B�.׸[�/�2����<M�:��'?Z����(%41�>�D� ��rm�ǝ�Jj�N���x��/b;"v��h~ =&!^����`���H���/�|���G���u��r9�����6����S�J%O#͉�S�Ke���߈x�9�����+n|��Ѧ5����͢�f��~M����F^�����J�����-|��noaQm<�&n�'����y�	���C,xF���-���5�|���锃��?0Om�|'���T������)R����RG����v
!_��
�˅Z��a��5Q�A����ҙ� �D��NUL��rr g���9�p����Bw�UJV�@OT,����*<2���$%��:�45Q��^
�dc/e��`CTsLn���j������{S�=���N5�ѕ�<��G��0�ћ���9��h͑��,#"�yĽS��O㕊BI�:C@+ĄbE�W�ٚo���e���D��Y���X�t����e�1�a�s�7�XZ��/���"�N�
6����f�0�	�U_��%�L��Qi�Ni�N�#�&:��c�V�6O��r�i��r�`�_gW.ܨ?�o���8��Ro��!^Og�04%d�	I�ə�5��rU&b�4���I,t)�'����G\�����7p|�PSq�sd�u���y������p��qvVBE='�ʵϮ�j,cC�j$`7�ʔ��Ups�|c�6fi�p�P�*w2{��ֿF���匡��8l�pk
��4d�񧼼���k���m�I�r���)I��9:I�p������Mŵk�O�b���F���1�Pc�K]9���|\Z	�ڌ�!�}������F�ُ�ϲ�9�6#��>��X5���(�1��C�bŀ�Q���5�u�B�PU�~���"D!��(�4�؝�3�5q���;"��R�XL+�>4e%��F��v�����=M����"��Ε���O"�#���uƻ�J�����4X���v����b�E��� �#���tkREo����xL���� ���8�y?�w�~����T�v+CY�(S(9�]����Tu���'z5 ��H�A�����OQ�Ll��^����i#�Z6�8�c���Y�?2�
�G�򹷶��q��M�j����jC�����k_���ފL�o��M|�|�p*��,�7����X��/���p�lR'���R����FU��U*[ub���w����U��X@�~�Ӟ���j���{���؄<<�V"��7$|/W���/��=��Ǒe�c���Zp}��,����|��,�׼kD{ ��k�-(�h���t6��@<�VuCv��^��{aQF�y�2��8��)hT��~��4k%����a�O�1ާ�x�\y�?6j�����υ��f����m��}�X)��oj>��E�9#4��5O�O�L86��<�.�[l9���Xn�9�in�9
<,����C���]/~I��wXB��iІWd�����?k�a>:��8]��>p5H�>���j8�����c�r��>�EB���Y{|�')Tۼu�sSS�����g�����������T�ef����<�3|�O������[WNml�>ل�3��F����$?�Dkd136�0j�)#��9f��cNW-��T�k�#أ4�0�: 1eB��4ĩ�]�D$R�GW���"�37�{RLYqW����C"iC�����!����/��&�4����@��|���/���_��;.$Y�z�-p�,ֹ#�)X2��u�p$�*�����E:-$��&g����?��|�|���0�`zH���(��M3�sz�:De�O��B���>����@ƄwH`���=
j
��m)�Ũ��)2mFw��:V[�}Jһ�)Sl`�@Egn����W�h�,�u�ȍ����զ���گ��7K�w�8Mq�u1�V�x����rWkE��)���
t��J���`U���kճ
�^�r/'����g@b�i�N>1�KEW����@����Ͼ7��I4���'�sy�Ts�n��kՑ��3�������ƹc_��+7�� (�i����8���d?qя�Q(0���wS�_L�S�@�ڲ#!j����tZ���j��z�����A>��4L0��im��h�?(bK�G]� ��IV�]]�Fn-Q�:E�>�o��t�/��-�6�ה�����C()�14�%CHK�tw7������)xx���}]{������'���j ���f�����3�hs�U�����CٯFzEPFem#.F#�E��B���G��F�YD�Ƈ�jD:��aj��@��{u��?﯈����)D�D��^��Q\���^��%
�%��+F�p��'�/A�[A������`�f�����ˠ*������?D�����w0(u�%Kɷ��1)S�MXw�u.-D#W`�g-�1��Kd8�K�=q ��|(L,�k��5fc��a\��5��� �����e��y��E�������>RD����P�0ͱ�j��[� &�����u��n�d�4@1Tc0�ȹ'Q�^�V�U ^ ��-D�?��Z���M�؊���Y��y����2����>����JG�|k;����w�]hRY�(�Ȃ��z5�Hל�e��HDz��e!��=�o���6��_����������_�b��<x9j�tJ�=�`3��A��$�dkD�h�6^�5vb�MD9�Dď�*V������Sq�X�B>g2_NU�_���>?�2Xln��{_�~Y��:�bo�z��$h0n��W�����y�y\1���6�B�B�1|S�iM/ zF��\����j�n���z�Jwϊ��g���_�@��?�L{<8z=����gFGOb��W������r������q��l10p���ȕ�8����l
��_
~'hI��!�1����5�w�qC��]�ky^��Z��T����������T�HW�������6'wMM冮�R*��ѱ�����1��g]�#9�>]gWy�H�jQ�yф�������ī���v�Ph|�kI윰��QIj�i��r�ӈ�6��gX��{�����w4MGt-,��P:���n�('�>m�����,��Cg���A��/ǆ�v	R̮���=o;#J,���m��VABz?�������\����R��t�~����������@.h_.�R5�Z��4���D��_<���6^�:[�_��+��l@]O���x���:� o�ZS��h#���ms�?�ۅ��scČA��e�ӿ���,,+/���Y�ngwZ�"n�'�J��"ӂ�lQ���k+���ߝ����p���xeV�)�⧴���	��wY

 է�a�sSp�Z���bB��2��<T�@^i��C���f��=�ewxy���4���C��+Y��ښ�����Myh5$��8�Bw��m�_aX�[L�f/��7�}�:X�RH|�Ę�:D�}�lcR�bт�!F�X�Њ%��~q+e�� ���#
� ���*�T�?��2,�ɪ_�!G��7d����J>�SßD5n�8�濗�L@7}u�	����p.1�i#����8����,�~�C��\���L6�C�	X�*�:�ڔ���^A|�����\���P��`�l�:k��}s�꾼����m���P\�N�*���Դ��_gڋq9(90V+���W_���N��k���2��������T��?���qU]��|3�W��q��%A<E3o�}qd2�mPpJP�j(��"U�����Ol�"�Q+�3F��Ni�y�@!��,��<�z����e��v�����[�@Kww	�S���Щ�Q���V����}�M�X|*��ٶ���ts�tK�LS$~N�p�t���w�Bڔe&��	l�{N�#s�Ɗ$�l�ɤf8������7SkM�c���'%�dޏk�_,蟿H/7������	��)���9,x��籺���Dj°�d39��y��I�j:���(A!~2���%�-T��7�j#�ѮS3U�Կ�a.�ҥ�Zt�u�J3���B��ŋ�Da:K�Ƚ\��D���.����=�
ڔ{_5�~XhU�"��WxZ"�20�3����<����f�j���6����X��֟n�	5(�/����OW��J'��n2�Qn��Q
<gq$t�S�~������MjP+��A\�J/nS]#＝���j@�ʐ�ۧ�������$����5�����f׃#�m����Ĺ$�� �_�MT�8��/���	m	MM!e�w�s}~֘��]"l㝪;_>/.:��� Yo���JKGF�#00��o���Z���zzF::$�P8f'�ӓ�7$�4kgA�G%h
<+6�=��=�	�Y�s����"����:���n�y�|j���G�J��)�݅΢J���!(��WLcK\�2�� �ֻߕ�Q�#T����G7fk�{?MF����~S�ׇz�ǳ5�{�o^ǳZ�I��m���B_�K7J��BT���|U�+e���3��\�|�բ����9څ�Եo|�`�!j�o�}&�����-�/ҍo���ل�*4��|j�����d\�Q��MU=�� �;ly3��DӧC�,ñ���P�HI��T�?����O��Qޏ�sAʆm�;]�mJ���W7���^!���/Pc�wފ�b��5��5�K���C1�g��UaV�6��|���D��U��3s3,}�@��5�3�C�Q\�AM@�hr۸�=l��!g����3��g�DZ^vW]��_���m�[w�UG�^�]�Q+�d����8#q̢�a��ҙ�)'��O��?D�fD�ȫ_j^d�r��%lz�T����*�V���j�g�̰S�!�B�IfG7Q�4�2��qVp���vo<h�����QNK{T�����S�\�P[� &%9Ƨuwd�[����p��?��#;��������_�i)�ۊ�(o�����<L��R,yMy��t�t.�tޕlƍb\s韗҅f�yVt9�T%���7¶
��v^�s%v�O����ҩRK?�>�H-�58Yڐf��dE���LFn)8W���_�:,7S78!^�;f�HT�X}H��ʂ�$����o�A�� g�0W��;��N��nV��1�
�2���.�ޢ�	�iUVxg�S��=VJW��n�q�����*�)�.��Af<f�L�h÷J��PiG-F����Е,nH0������/L��WR�j�#dh�~ry�Kf޹��62?l��}����0��>���d0��_&u?�|R�P�����E"������D������;hA��zc�%G{:�p!��`���� �\#��&�ǼmI�U܇X3
/��k�f����_�FbI�w��[ƅ0��,>�.>j~���@���8I2���G���*����~�"Ծ�"S_�\��s�љ{��o�'M�Ҳlki��~]�;[�enng��z�l����2���^�b�F�"���\��T�������=�,]�?��G��*ʋ��c0}�tE0S�0��U���#c-�<I ٯL���/֓�����b��4�S�]�@�?�L─�+�"d,����˄Q�v�+�W��Y���_�=���6��6,�f*0x�,���" �/��"��:�+4��c%��� ��es��o�)\���9�]�$5��z��4n�<[��_l�c��o���/�ߔ���y�f(�^}1-}���bm��P_��j.��^�6�;7͡:M,4Ƞ��6u���0�o#��'�L�%�T�G��o����*��ԧ��3����v�;hdJښ'��D^_�u�4�dI@�w&S'���GO`�x���	�1�2=?�35���Q	��_t��D��Y��w���lhh��������㙘���������҇�BYY�pS���ŹHE%��VŠϑ�!���U��紇դս�s��0p_�[6� �1�
_��,��*\6ܥ�\U�]T�^4h}����8�C�6�e%<C�K�:�*Z["&�+�.�����wz�#Vc�M���I�6�U8�H�A~�������4��cC�|���âk���Μ�y���m�c�Yڊ�r����XU���N���R��.�,��c!�&�f���Ȇ���� .6�T֘���T�dd�%��#+Z$�H4���P��1��Q��Q��R6���I���=�[�S�nyQ��?�>mN7�	Z�q���Wb?$��ty�H<�����0x��U�L�k=�$[s5zQ��X%d|7�/��O{�<8t��ڔ�86���p�]ħ����o����b% �Y�$�s��gs�M�s)oUE�Uyȶ��.h�Y>>�W<��������&���$O�^�����k���_��sĎhMY�TSK"�i�U�����ֱ�xIL���s4��W]S�i+�7ѷ��"�I㰗�?���l�^Ge���_���y[X�kgkĨ�6h��p�xa�S����>��^8�V�F���g�RV��	d����'bA�vW�/�_��k!����͒�f7.@�Y���<���� �:�
�7�bL�a#�!i�7煭1��$�t$'��:hB琺'i�:jl�k�Ȯ�t`�?�aY���~����BbV�Tn)D}?�ZBɛ�`yo����[����@D5'J�h�h�����'��s�П�ў�_'==9�Մ�,�ǫr�w��k<&�7&�¨�Ω�ͦ�ͳV\+l����Ji�O��'#E<ݗ�ݧ{v��
m�x��BvlEtf�L��i�%���{^:da��{]����:�L%�%��<!�_�ʨ��[�r@�鍟+�
�-da9fD�3#�c��ǝ�T��L�"`�{��/��/�)�C{��5�fT�Э�	���x͊LD�q�%
��wc���ESނ��7�3��0�>A���b�o��32,2E|�7/���S��
����f���/;�N��QF���S41M?PsOT[j
�M&��!։eX��}Q�E�$� ��z3�L6��-����m�WVu�k�L��\�HK:�P���� ���K3�-�������<�%�S̱RL�%w'_���[�qJ���k��}5 �_�:r�K*��*T�咬'-{W�G�p�_�_��<\,kkC)(�F;�1������)CJ��<��x1�@3O3�H=UW��J1�L+OO�`Opٌ��&9��lV�K����8��Is��Ő������*�n���;�"B��/͍�7��S������8x��uL�3m�Ŝ�M
yAx��?B�q%޷�mE)8x���7��><����q=װ.��x���S?��QH��Zs1�!����~���bpW��dQ-��:����Hv �,��iK��P�f��zb��Wy^�� �)�`��a��u~�x�`���yy��~�
M�g3����$��98ĺ�.�<�u��(��0�`5���(�gD�文6�5'���E��[����o
�h�#��h����B�)))111�9~�~�~'Q�`'gg'�ں:��
����)h�oN�,��o��Ll�K�E6��e��3����<)'���t��SX��vD�/i��_��c^C]uE�8i��B£"B���Ut�d��Fs��sɶs?��l����]�a�2�h�s�M+N&��p~]�od��O��..����5!���ERŹ����������q��^�$� ����f �������d�.���^J�S�6�NT5����雹�Kt�Mc@W�z�"�ą�����*ׅ�}T����%�@�w
�V�˹�9o�\s�\�i��q��f������e�xE��q�a���Vb�Y���B&�GYy�	a�aq���]E�L�}I,�J����u���{��**� ����+E#Q��Y��BQhs�|L�N��Nn9M�W �����0�o�ĸ��@���� ]��~��|��bo�o��q�S��T��9>w¡>*�R�,�Q�����j�/DP�d6�����c*P��M��?�D#�����09h?���rI8;�u���&栳�I4 +r��Q"
��M��r��16�u&;���(��"���ڗWFAJ1\�On�9��E�>��i���
� a�eh�F��z�~+9cTډʥb���2�aCQ0��V��k���
�j�T p��5�%Ly kz+��<�{;8SU0R��zy�cE�S��P���F���(�_`�:X���,���ym�o�����+ww�"!N��6�,�P�e�E;=�y�b����@|���Hc|(c�w#��x�[+EN�U�D>!�D����'�?�Wpv	�S��D	�0,R�
9��,6{��E�������*5��=���� %<ةЬ^Ų1���AIlRY�(�u�F���S��瑯U���C8��J&���Ă�t�p��}:\�ep^�r�����O�Q�8�$� 02�*�#���*S�8��^���ޭ��B�83��UQED`a�گ�����c"���{�)F��������PUژ���U�����U�Pd݅�-݄�D��Kuh�������}��;eeL@k���������(�-��=�C��8r3=,��>���Gc}2[�0��/YL�X�˚�{����ׁ̑��3�X�γ�=��a�
�~�&A��Φ�I!�lgW�l�iD�3Kt|2����Cݒg>(��dw���ږ�L��`�G�ĀOyBD�7^��x�X*�d��tХrIZ@	"eف��X]5���)׷98���Wxz_G`Vd>^,'���X1۱y���tݻx?=��{<W��;ؔ����i:Gy�R������Z#boL3�2Ի2���Q�������Wv\?x�;�ߟ��KK�{��7�bzzz=��ѱe��[im�e�l&���$V7���3�`J��p�3��ķ7�< `���k���(kS���GdB �pr�\�����	����9:[[[[Y��������ggW�ޡ���-ԐTԠ� iI�ͽ ��@1q���ޟ�g>���u���������y�/�������#�
���GE�g���3�	�C���0 ۑ*[����o�(R-��-9y�
�B�&�~=4�}����r̆��z՜�l/+�y�;l�j�x�n')�|q6z�E�F�{j��hH���Z�})��j«j]�&y�%�k�g�� ~Z.	Q�Їw�޸� ��8A�*��_�:1^-�gD�"}���\�Hm�#ӃU�'&��K@6��"t�c�����b��Z]7{�S�m�S�H�;>3���#��q��K:�M�^�U:�����<�v�:d�D��
,�gCG���㔏�y�8�l&�N[�8*�����Wt��SP�wo�xS�pG���/Ȫ��ݖ�����7����5���K�k�tVc����џgi��h�yd!��]&���W�Q:=�\WNQ��C������[X�ωN��Cp�<�V��L_��bi�'lh�9�'�L>+��?x���a윮����}�%�x��mr1Mݡ�8a_,.(O�)<�n�'40?/xU�w���<zI%�s,��'.p�L1�+^�W�K��m�&����D����In�Q�H�-���|�Z�b�Y� �e)�(��e3.!*�',O���ݟJHem�(�	w�c+��+�xc��X��g��t�� ��G�8q�z��{A��AS�ϱ� ��0X�q�hJ`.�Y�Pr�������{��};'�h�E'Щ.��x6%������n7����D�\%.q���2&/&F0����?Ň��r�=#:�fN����*��v�W5����v��i�Q���>�e�y������QAg�6�#�P� �jD�
�M���X��m��NݗИ�k�/�2nC.���C[��D4�͠�� ��<6ȽV��~��o��a��f��e�@���e��e)}	!O���(ыѷe����b���ͬ�i��������.�Mi�3O����sZ�#6�`�	 g�$4����A?���Z�5b�Tx�%!%�u$�� Q��� 9x0�^��ȒlC�w���^�w�9%�
�I�b\4����o�eF:�hV�0{�`Z��]�|o�o,	��-����@��ʑ����/{�� U�O�(~�����O7�{��ӗgy<�A��I�E֖���@Z�֥�%zv��ϯ(���Ok�z�`(�[�{�=5�cmKDX�UjCU�0ǚ��l������5��Gs��e�B��ڗ�c�?�����^g5i�N��e|�/O=�^�-�DD��2�`�{�C��F�.X�ʦ~b8�Sp��j����F�ɥN�O��2�#�Y+���䔖������䖖�f��$����
��_
D��+���ٻ��e������	��{L�_l���y��(=�8��~�ʠ�:�%�"B]K4�\4��5�5"U�\z��蛏i��U	Y�W�9'���H6��-�69e0�؄�}�V�-�4�^�y𝭺�^���/x�]�4�-�׳��Z�ע���ܴx���[�;�wY�oܰ�c �H���1Ő�g�����qOe�R�/
�;y�H�*k�����E���[��[��w���>a����V8Xp4�a��o�S��P��Q���L�L��9�\WR�𹭄�\�/�KI��B�t�h��Z��x�븇�	�Yy��cQ�E;��C�&��QB��i����ޯo�M��]!��Q��U�&U%IYE�*�{�&���uϿ�m����GI�=w/n�H���t�&4>�'�-Go-%oѴ�,Z$�������KG�����ى�|�9B�����%6�\����u��k�O���ɓi딚� $���!�?þ�6nu��/��S7����r@d�����'���~
<z�,a��F|H���S���|��$+q�힂�W���~�/���t�RNc$y��?����?�ɓ+�ʒ�&d�qO�s�i�. ��D�J7<o��w2�zѣA�~���ͮ� �sU��eA�S�:K!݄׈��+�^3�JA�a��Q=+����F�Z!��R���;���_H��ӥ�_.Efa�$�ĨxG`�	k�wf�Ɨ)����p	�$�&꽗��Ђ�w�!�&$1D�/����s��*F?h�b1���"����� ���+��F�3��^����Q�f��ef&g3�;�DG���;��!���\��vm�q�򘴞�H�S6�ZS���@�,�d)j\8��\w��Q���1����X�!�[Q�"�
��z�!.��=���x�T�4�JB`�Hx�A�l����d�o������R?�!�jrP��uiM�f��GKH�UQR-�7.rv����aU�.[$k|���Y���b�:Q�&'�M��1Yp+�K�>�(=�l�y%�初AaC��R,�USl��g�4�:6�E�&9q� �xu��l&[u|�E)n�)Q�=+m�s&)����d�_T�h?�<��B�GQ�P���s۫���}B�7��n���	ynP��Sw����/��-$I?���j2/#���]j]�"Y[�PZ#��d�Z!Y��bW�g�µƲ�O9$�;�xtQH����@���9o�Ż��d��������ml��r?#�ZKYـ_�n�/3��R��Y�#�����ݟ�+$��'7e��3x�NE߉p BԊ�B VR @Q�Ӏ(��1���
�á"�Ŭ����P�P��=͆J�R�����*H~Bs1��"}�����F��,��v�������Yg3w	��Kܵ����BVA_��tߊB��㎼��t����5��$��$��4�e짡��Iƕ�?b�����2֫8TM�`bc�'�qq��Us<�����s��Wq&�a���J���L��˨�!����^���|�9���Ɯ���@U5�f�T`�1�l�F|vq�퍌�I��-��5-~��0���F��n6оf�n��#\[�?K��\��Yoz�q<
���+������~��jVZ}������S��EZ���Q�_^F��E���(��&���p���w�_^Ƥ�F��� mi��uI:Ѫ�C�e_>�D=.g��[�����|.w:�1�/��<\ <���:��y9�cZ6E��e���xɔ���� r��M9��H��(�Q9P �D����[,�����}3�l�ƟLp���#�@�`�Z
�`c����o\�Y�`QWi�n��o�&�Сq�����������O��	A��������A�,A�Y����-��@5�DEػ*\�Z��Pmp�Jxd��'5�x7l(f<�C��֍���F�R�bEm1Xʁ�(�"?,֊�� �`�D��qxί�-ڱ�7q��{�W�����e�E=��jA#p�뿾���wqa�KmA2Q���*I�G(N6�{�c[����Qp�e 2n�H~�ܠV���w�=�Q�[�,�Lj���|��.$�:j$�����J
�_�ym�,r��,����1;�_��V�d����}����tFzs&�9rg�C;�Ba��5B�+1��)��q�P�[Q����v}�:���o��~V�"�c�,S���j3�ˉR�	�˹� |��"��W�-���� ^�@�u��q[��P��X�d���hir1�x���)x=UU�����}~,݆u<���j?��QONpt����r��U����v3�
���>mJ%,�f
k�&�K��j�rw���L*l&m 26�-��m��e(Aԓ�(�P	m:��>��B���s�����8����_��������o�mv<��T�Q�Oc��LsG:8s>�����$I�I{�C�$47��B�H���D����S�`���������!����8�������=������1u[	 HQQ�Nr�dȗ\sd��g�e�}�K���u30��n?���Z�L}�d?{�������o�7]X(��1}�l�Vw:�$m ��c�w|6����
ј���)W���c7���F�[�[���?{�t�a�����i�-e7c�0��U�(�0�|/.�V˃��T�X__g�y�����h���+Ŀ�UԨ~/޳����d���͸"��Do���>�A-Y<I�G!UJD���s�_{��&��z>K�D�zh&�#���H�d_�H�6ia�5:]�̷?l,��n�9�_V:Y�y7���j��N�_ݺ�돼��6��fIJ���� ��x�e�d ��d/	,;���V��+t�ǳZR"2�z�$>or���4��� ���^�S�@�<g��f�;��9A�=�/�@@�Җ(��M���Bz�.�wd��k_��t�4(!�aEq?��.���#9(x��q#��tfyr.q#��]��#�D� <�7����hP�ͨ���d�����U�ko���lQd*������&Pn��:�n��v8�Uq����=̼Lo������5�7"��9uc�PD��U0��0�-�$�tt��{����9�g=WZ���=�Hy�ݳ����wp��vLP�ޞ��
����p���N�EH���+�S5*[�������Y���~?��Wǜ2�,���+�(�үc�s��e	��-`-��2�KN�O������I����k<9� �L�I�5�C\wu�gV�+�x+�!��ޙ�Yz��Y���TL�Ф�rQHf�����K|V�S����ˍ�c�,���Iڠ���F��"��2'��?L�-]�)g�ovZ �6Y$8����`,�h��9��U�� ���g%n��
=�=ô��񃿸OVs�	�q ��T��r�hqV\jؙH���5��I�('�h�Я��� �Ǜ�B�)m֗ W1:�hf��_��7�[��j�qG2*�i%7V|@wИ=s�O��'����M�Tʰ��a{[EW���w���f�E�$Pv,�>u}8~�l+d{ut[_�����UDOR;IB'IR/ODd���ޒ`^���nT݆vR{�;�֢ϋ%c5�ؼ���ף5l�>�+M%�c�.;eז�C?���6��e3�1�aI�Y�J��o\�Bj�"�2�6a[�����P�Ce�mj�R�����,3~�?E*	<����l�D�|�X������|R��j �6Z��O�	�B�JrVנ_a�Ǳf����!InH��S'	�����6Z(���G��O�T���pH���3VI*�!����!�_!5�'S��̠���F��f��Z���_���7O=I&�^�j�0\< � �U�=��
;��ݱ��}i��:$J1|�E�~v^n��cE�]J|��eܤdv��IN��Q���c����UA�x��E���v�t���~5mi�zuyLn `��c��r?^ksʞuR���)����ϱ}JwR������[u>��zU1�������$`BEU�0�8�v)+�+�U���Oh1X.�gc:�f ��tT���6��TnN��=�&�n�_UhZ]dCFyR�&�"��/-H�B^��b��"�ҏ%��8������Ys��µ��*�m�V��ߟ���L=Xt}Z*î��{1�.=�M�����Ϡ��xj5��-������ݏ޴5Z۸9�̮�S�M?� `�J�o9����u�x�ͳN5T,�<����%�5`�Ӱ�'�f	RN`]�$����ᰓ1g�-p���A��aU�û��@�%4�]��W��}�ebl[�^䗥D8���ܔ�4���y_Z��I�N
���6E��U`f�\˚��1,��>������L���MO��YM܇�bG$Rm:��v�+��(#ɧN]5]X0��j#D�_k�4�h�Y��x����]X�A��Q��G}�u��c�T�kT�2�e���zo�Q\�.(�L�L#A�\͟�O��c�}�o��g;Fj's�t�~������#�}�I�g`��-�0�\�^Ŀ�	�;N�:�z��(ɳ��v�C��D\�'�q]��hѦ�NXRʝJH)�Ƣ�7�܂�;�)$�3��84����;b�x02�Z~�*1�t!���/L����������捵��1O�S��S/Ϟ���8�<н�NR����ۀ���A���������Ax ��F��[���qߠ>�$7j��]6ہ��)Y4E��A�)��wS���մrҿ�L@�9�=�F$�	YЈvg�mq����}����[N�X&`'ck�c����Nngm����ƢH_�L��4ҁfʊ�"��gdo�z������2��)���Y5�&������1&?�H�1O؂$|��AjG}� �X����T4"M���vJV<�O��!���i��{f�W�@/Wy��y�tK��/�_D�ݯ_J��\^M��&����{,��"���_��Q�W�x����1����f��&�$�X����5Y�����i��L�۰d*( R�>�K����M3-�@��������ۭy��@�q���f���F�yb��W�'�7*e� ���`qkc'CE�Fi��L��녵����C�S�刱p̱p�@�]R��u�u�4���Vӑ{�����C�6�M��9���X*��W�@3��\�"#O�+���n����Yo7�Hk���l�]�j��Ý�����g�U�,�LR��^������g��ֈB� 0��7y��ʫJ���h�k��5:L������?�����+	����V�$^&����21�h�.4��kL����g���!q�':�:�\*1)F�J��'i8���+�6�n"ǌ�O�HT�G��G5�f��`�N���M��n"(�V�fտ���i��H<��,��HE��YK���^O����HW8� �ֶE��sgm�B��Dz�8�[+h������qS*ry�����JZ`��ܠَ�ߤ$�Djq�OYO'��\�pũEWɥ�K�� Q�ZE�@޷�.�֯.JN�y~r�uF�z�肝��˺�[��m>{[UmA�����
�|�N������37��yj Bz9�����\����wp�Ӌ��#�8뺝"��p>�K��R�ݫ� x�7�U֕��cel���Rc��a�	��v�>1�|��q�l[�:�L9�N>�����0��`�x<tu��H���6u��D ��3	/^�q  ��o�Lj�ìל�B���{v.�}�S�܊����A�,k����|�{
��gSÅg"���E��BM�z���Z@���Am���	���?P-*�F+Y)��03ҋ�)x#I	�&z��6+1z�HH�Dq��Dn�o��W�E�����d��R�=3+-��q_慛�v�Z�*�CK�*�O�9u�V��YWyӫ�y��9�����]�{m�xU-?m�yl~Aw
�&�g�"���/�*��^��|�"'��k�_��Ƿ3�dN��78���<JGMr]6��A���*5��_�H/e���m��H$�E��p�Ӑ�F�d1Ux�+x�K].a ,�;��bgIń����'f%JT�.����9�8�'�s�1ׯ��3h����!@1|j��S4��U�}[S����]��ihco��l�
�Z������:����h������n�d1+��j��k�B�Yê$S
X�Z-.?��Q]تn��>�H����\��~�Ȃ>C'�NŌ�!{�:F�I�sZG���<�L��v�Yf���r�6��u�#n$Kxn!&T��7m�2��2���,�`������QnO.ϛjO���P�Q��I��l��VE�Ŷ��+�&R8����\�4���&�i)荟��<m��h�Qp2t�]3��Th<�E�HA�htJ���ɚ9��J)"�%P*�k{�T*5��$���s,a!Ma�f��B��6
�Hohq�<�_Bi����F/N��鯘�h'#ߩ�jep�t�*��k�l�n� _l��v?ax�?��$t�iwcSm�|UڣB0�#5+��ì��t~����WJ�&�T�b+ve8��$��#I�!���~����L�M˧���Z�IO�VH��ªFrlI�g�q�
g�jی�r����l}������A�I��(Pm��xo��B���'�ٸf*Pѷ+0"m�n���R����;��x�b������w�Q|�n�LUSS]m%X."��B�Y�b�(�������h^���.#iVp��B
��'[ǿ/�'��"�:�c���4DU���9�upQZf���X�{6:��B��5�TJn��ѧP�X��QśLO��&{�����u�"7�Ț���Τ>�p�V�'1ڶ�8)���ߦq��B�W�0�pΟ�,]$��:4ـHu���O�VI����tp���[�d�UP���{r���.�.���D��&���)�dw��1߭����g��А:Dc��~��r۵W~Y�a[N�>t<r=ٮ߳O�&=�nr�I�RM�t��[$_"�bB�yg>���/��5[D�	iXi��	E�o6�Gi��M�I�v����$�cGF�c��5��G��@�`�J��	����i�����.fM������H�.AN�)�ܯ�}(x^��u�nZN(�V��i�pz��~v�S��_�Z�A�!�'��Y���=�B�:J�-�XE���m�W���G�`rC3)cC0�N��d 4�;������="���i�<F���G��}SR�Y�t'h�=��)t,9'l��hU�k,ΫM1����i��C �=�5~n��M��k�f]�߬�GHT�b�1+�E�-�[�I���d4a2q�@C�u���瀕QF>b8?����&�6�FTD)gMt��2�r*r8�L_�X�0X��|��x0��,�S�QI�=�w7����BXǬi���L:&��;���в:���eoo�Z'��a��"��@k��ĳϋt���PsP�_g9r�����Y��E��Y��U��e޵y��u�	s"_5���y�L����_b{jdq��Y�)5��:��s�Am�r�"��*��yV�e��fA�OHec��ľ�31����;Ȕ������V�Lҷ�)�"�o;9��)1���	��,�ȝ jA��8"[4�A�d$�ƿd:���U�D��������#>�����vO}��7S�����F������J���v��P�S6��}���A(s��Q����Q���岆�%������7^����r�Š�pĵ�[���C?����?��6"	����q��_o��8�'_ovٟ"�ku��X]D���%K�f�֖�^R>�������ڱ9�+cYӴ�<���]��\K9��Jڄu���D����6� ?�Ua1�_��y�����DH��:��vmbQ�O6�c�=���7w�D�]:�=�5�ċ��?z�=̡����)��;���������8���X>��Z��	^5��$���>�v����4]�SzX[&�@�Ԓ]����ߟ	{���Z������,>~E$��r|W�HW�URW��:�m�SeR�C��3�v�r����I�Y�G�=dA3�.���1�M8	$��I�/5Pw�f���B��W�$���N��WZuK��D�Z͕yx���QL㝤M���R��V3-��sJl�*l-��&��9Tr���w͔�L�{>X�)	���5��j^� �EH���r|��C�Yp��Dk�P� ��%�w�n��Ci���KqPܭ�;�ݥ�)�G�s��~@��&�\������v`L�#�O<$�#~|\���� l�T���α��v�?�1/���M!�&gO�Ώ���J1^V%
@�Z��[vT.FLcM�h�v!̴��ӭc>�m�v����t�Ψޒ+�[\�b$�8H$|"	����I)֣��A%���z�F� ͡����Ԁ�����$+�%��Np�2WR֣���.'�m�yڀ⶗Z?gY#g���-.�	M8�I-�����N[�I�2��j!���.x3���jn�0�m{[�
��3?H
u�\����њ����C�K��,�C�͂%�
d!b�]�4F��/;ݓ���~v�M}7�t�Dg��L��i�iC���<E-��R�8��y"�l��4�m-+Eտ�n�n�o�0���A����Z���H��~�X�{�/��S��(,_\�1c��Bl�Q�-զ��`�.?q�*�C�6q(p�
h�߰���J���"���LK�"K�-) ��L g]�w�}���`����wbv|0	�4���m�A}�ե�4Y2��eC_��.B�ty�T9h��e_��DD��W X��~U���3�l�]��~�ds��p;9ϧJ�&�,2c�n�ŵ��-����g_g (��/'�J�'&N�^�sC�%��]tI>
LI����H����$��d��J�I�(ڿ6�O�����{g,�sp��g�_���0��ݏ�Q��C<G�ӆ�- p<s���[!���q[)������5�e-"�T�`j��6*J:��R���uiF�>��VЮW���e�m`��c�h`�(⅚1����5P[x�L�XMr2�������SeV�a�>���o� V��:>=�t�=�"�����لߕ��_�R<XA�k�UA�VC�kQ�q��v%�b?�5�,崵��Fb�~[3�G���h ��� H�8Z�ZS,Ed�q��j�k����-�|�� ���"�!�٘�5⃱r�\���wl�k��~hz�<����02�b�[T�(.��Jxb�:��n+Z<���^c(���u��1Ywf�ݯ���3�P���mB�A_�6 $r���w?������#=7>	��ʳl�ce�ec=�
F�7�+%H�r�!�S/|gP�
�y2�?)4��5=1݇2}�w��^�2��c�}l{���p������ɞ��{mPcm�*��-��Z+�0U���9h��'~�Q�q�G�7�8�	�V_��n~�L}/���B��`�������[���n�༠��s�i��_m�mE�����L�k�b���|%�mk�m��ݼ�>�="f�2aB��Z�Ͽ�����d��ލq��6c:d;��A�.��+&�T�q����$O?�\)G}P"D�X* �ݖ�>� O`g1u(b��m�#<p�%z`���t`h���Q&��=��	.�����	| H=&;���y��-5��Qº�6X-�)^<���&Q�X�N�9P����}�VUy	�����^��U��r���׼W�XN���J���T��1������K~�URZ�3�E-&O�O�+:)���������}�ӼC$���X-���%���>ߗ��r���/
,nv5ַ�rҲׁ�Z(���AZ0:�&E�Ư*�?4N���w��@-{�|�S�9h�Daq���������X@���^��0�I-����I����	���V{�"W�93�+�W���9���1\�����B)���3�'�����=I}7%n�t�o�j�-?��M"U#�V�"<��E��fs@?	� ����	T���>�S�^�?m�6�\��b��v�Q7��v��E�7��]�U��&�	��mG�O'��t5!�O�7�]�]-��� �6�	��))M�qMH���"{��uU�@( {:��6�Sq\uO���R���ʆ�3|�&J��gLI��}�E�]9�?2��1�Ϲ>M�g�n0SR��T��Q P�� �#���q�Ύw�0�xT�����x��ڇ����OE�t-}�%�%��U��0��Ud�4��{q�@5��	�0&��z5!p��s	g��,P�+x�F{(�{d��9?�Eo��w�������|6�c�Xɺ��_�%�X�_5�xpF�s��ڣ,W<�:]6�lY?��l>艒�,�>���j��)�C��l�n�6>�����+;@�V9�O�`�J�q��K3���56��y�A�����{D.I�7����}��xUk/9�]��Eq^�vb�<d+��B�?�o�n���#9�s�؞Z$�	���G/��\�t;����uDr�XŪp�����*Vf����>�E)m�I�ط�<!�t������˽����Ed�@h����C�O�Ş���H�{ͽgÕ��a��5�'ą�O�6B�6U!1����S�R��#͠fޙ�y5�r�������X�v�!�����d�z�u߀a��_�7S�Ï�%Q M�]���n�W,�(d�k�ؕ��,��	���=�C�)C�S+ݪx3v�@�6�.�Of(�^8($g���I��t�me��P�s�r���7�d�8>u���������������U�V���^������������7��/�
�)���Ň)j,�Z����0�D�:[��}ί��MJԫE�O�`�>\��L�=�\:�/��vP��׀6�A��[zr�𻉎��U1㨦�S2�I�,ڌr`M�9��e
�i�ֈz��4�u���M����'=u��k��G��LP�H�DEe����T���/�kxV������L-[�_�A��:��ی٢K�y�d����v�=i?Z����fm<��N���=KYYgyg-7c�X���B��L��l*݉��|N�Ԣ9y1��/2�Sy?�em&��e�kd�&<�՚��sD������|��l\4�܌=�#\��z���+�R����LA��~-QiD�,�`�3%�Xp�!j\5lkBM��0�
�e����$���B�a(^��v�:?���Α���B>���o%�3 ��ۇ�Ɵ�j^�n�q_����@���:_I�?�;�)2���jP�����X��3��� ʿ]�B"��+Z�	͍�^m�^��~�|�m�VM�vm|�Ub�a���UK��˓����?�#Њ���L8A\����Dq��G~/.Ql���\��Qn�v!�mDh};򖞆���6T�6#������2$H�����:xrأifj`Ц������� 9i�xohp,n���T��ؖWVN����=ԃ=\��\������[d�w��~��X��;� n$���v[�_�^K��3b��"�}�G����E�O])����gy�B�r��[��@�w��h�L��ٛN����cAٜ�Ȼ�݋O�o&�^r�3EVS�΍�󱠕~v0�W\��t��b���b���EqFM,5�W�F�N'T��y��J>
5H�� ���/�0�{�8fij�)F�RuL��X}��v�T�L��(.��Væ��N���#�u״t w�����$��:��?'=)c�RƼ��O����C�����b�|uכc�6�YB7��23'�3ƴ1�4�G5:��d�3�w[��V��Z��R����>�Qi`�N�`0�:��P1�80���?��dj��\boQiQP��ky�f�1��;��i�b&F�:�>�ީ����O[��p��L�� �p*�m�+���-�c�Z�`t���;�Am��K��K�%��%,ނ�rѰwʘV5u��t��������*�$�so�siDs�r�!ЃD:�)7��D
���4���'�Y��0�o���5�J���;�l�p4��l��n��ȧ���Q\5�ߋbq�a�b{���
y1��G�k��@Kf�	�N���gcn�.��+���֟������4p��8�3��xdw7��v{���B�ZY(Y���Sp��ٹ����2���N^�h����'�ܭ7")����Mɘ�"6� ��9��1R�R�qB�1���P*���",������)����Xp]��GAI�ɝ�`��q��=����+�� �i�;��_g�]c渓�Ȍ�iɬfW��#i�FiK0~-�޻�ʶ�p+/�0���{����a��'uYK��#���Km�^����Գ�9��4:j��u��O���Gȅ����΅�Q}K#GǨ�4�M�/�۟L���Wnlf!GqP������w�.X03}���]�6��Q��2GϹ��Wk�i�!�[�S�K�_�˄�,!����KZ���E��ѵX��_��}��p7t {C�-�^�P�o�Jr��ks��Mk�*J��*��{+�ml�_')5^������Z��_O[��=��s=�k.��Pl�Dh�ˤ$�(ܠL-V�3��2�[\/��,N��HV@Rp��&'�t��4"�_�F��mg�ݏ5��2�@_{�&b0>B(q�U
!8>P���_`�6��+������ɿb��oM��qyz�@�!�}EX���K�d��P�Rϕ�R�6����4-���<���.D�Z�����o�Ut�=E}�A��2F4T�7V����C��bٍ�)�s�,�k`Ԗ0m41mt��/e�|���3����8�+k,r�;"ag)/E����=6#�uJڲ"94#���<��3`Fwϭ[����7���U���Fo�^�׀+���̮��5�o�I���?,���_>�/�������=�c�C���<�a��a�JU��x�����=�����_���V�����dXlW�5 [k)#^?Z 50�A��81��F�(�|�K�۟�]5��֔Yp��B��+1eA&6�ͦ��1{�3ѱ��uSmL��[�/�ue]xv@������YšC>-�"~�q�Q�p��'��c��-��ʏ�l���T�����+K$�+Ia�n��1�"�K(�Lɨ�m�Mm�-}���Y��_=z�����?۩�����Zs3mr���3����,|�Yk	d �0ea���5+ݵ�`�#ꐯ����RL�>4��Xe�ҿ�KT��f����8�n���0K�1 �����9n��>���C�����9m~z��R!_q��RR��˥)b*����X䝜S�q�ܶ�����l��4�:}�G�'�º���@�C���W�ь�}8A�d�����b�ڭԿ����� �Jk�-�q���O'�ո��~TÅ�*@�&�Gv�*�<�c���vt�<�<����;6#�::�?�4�+K�C|��eܕ=�dt���%3����$=xJE7�y?_��! �7��f�e������p�鮉�Į�
�#���'ф YB��e��a��u����9�������b;���&��W6F���&����M���J�X\�F�ͽ@��#̀{B��Z���t������>S���6��q�j}մ2��r�/7�q:��Ϳx�&S��&�� Dok2��8:���-��qFdm�����C�1�aë�-��8s�:Dm�X���0���� �-H��\�&���M��5��p��Gq���eY@KR�b�x
�N{@�P�h�� ����a8
�'}<����ty𓽋cf�cM�W�P@H�wBB�||�9��c�쳸��(�b�&!H��o	�u�S	����X���"��ri�шߴ/���������*��{1�*g	��=q|9ѫ�M��w<��%۰�5¶Z� ���{[#�I�� �~�3�ǟDJ�W��P��~<�9��r�� eN;��o,�7��p*��C���~���,�	�ݢ
�΂]�e�َ�{�\�Qȑp��6 b����ݼu�C�S�H�Ǝ��*`b�o;����>6�iro>�"D�w!Q������;���;_^�%v��K9�#�3�Э�oN����#��˞;���ˮ�S)\�ݻ�����pI���+ə�F9=&�.�{�"��~��ŗ-eU�ɤ�Q?�tB3��D:l~K
���|�w����C#�˃A�V��o�O0�m��ֿE�q}Óx+�r�W=~PuP:X�Z��f�E*vU���]�uu�sv6�42��5���B�g��k���Q\�G�
$?a��k�ը�]i��_� �bP)�
�96��gaE�ޠ��c�f�O�������,����.�P����,�N�K�����P�;8�~j	{�~l�B1
�z��q~�DpI���!ZY���#y>y�q�r�M
��\x�v���z�D���M�l��u��n�y�A�uWp_��&>�m���ǌ6עV*����<�^9{��v�z��L-ݸ<H��Z�*U�ZbI4�c<XK��_k�=,<��6$�.n9R���3 .se�����vwMb�����>m���I���72������к�����ۚS�)9�v�p/n�;�a ���j�隉U�:� �c��+�U]�
H�S�JdX�]v���"��U Xd��;Uײ����	����ZD ��TSP>���&���}.ǕR��<cS#�c���y�e�d��%��^�|��K����ZA>(k� {>u9m�L=�H'�L+�`>���o/R�-(D�c��'^"�O�u��wㄋ�)�{�z,��U0��,pv�	6�b����)^��(b��o�;7�{ZA/�|���ꧥ��������D/�D7�6��Z#&�s��Ny���	2�&d������������U�!r"
���:P��K�Hh&����U����R�T�=�Z�J�VR�f.Af%���	j�|��e ]�V�����3٭����cViek�S��vȩ���<{�iڿ˫�u�g�/���&�����^�Y+�?�U��w�(h��b�Ht�ސ���wJ��_!�3��- e6뉠�>`NPa'u�D��	����Ğ)a���9̛����ox�U]u=m�&�Y̻Is���I>�H.s��4��5�y�Ї����GfGg���g_D�_�e���9�K�l�O�\�.�.�pR��S��y0Q | _�E�����G���|�j��\��1�w���%�0#D&UO3���3E��! {{�TV�L�rv�%q�2��)^�;7^�%D{�%��GVW�<�Sώ���&���r��SO�w^�7QT>3�3�x����8geߞM'v�=�{xZ:��b6�gnii &�na5���$Z5�|��j�̎&�P�ʍ�d��p�3��]��y%+�EU��J���c���g̑�k0�.��/����`n c����y�(V�E!�8�#�c(�)K�5g��F�x�?|�;Gi���"��<og>���R�:�1�Od.	D���p�>����}o�������e���X����? �D��~4Vd�\n���*K�עH@�R��a���,m�p����]D�K��폥�����o.ݚM�l��C���Sۂ��<�#K�d ��B	�\p�DPȁ��EBqlg~��ܶ��̐���]����9aAACÿ>�<F"�WQy��]�F�1��4����Q�9w�ͻ=�($�>5U;T�	r2J����~0%\o�~j�R=��}gX��6%����笝����������FTƜ�ꞔ����{�H`s��=� p�	��� ��$�!P�(I"9�6+O컌���k�{_��~���:~� ��u!6�O�7S�m>��(^N>O�����L�'Tƣo���'�?��q�u�� ���;�G$J	5H-���~..q;6S��jB��Mu�p�$V1�����ܔ�e\	�p��G����/�>>��%� >�!���o�z���L�"@F�M�U��������:��&�#Q�	߲p�>�O��X<ǝ/q���s�4S߭��S���9��l�R�"�,H��I���t%�o�&����T���+�P �ף:��gt���hӱ����-P��x��Q�HT��Uбr�h�%ոu\t2^t��u2���~��NauT6�j՚�pQ���fӃ%�'�y�5k�N����U��z��?M%�5�k���h�o��$�P��	����#���p��z����)�j�o�DMa��H#hp�T%�uJӻ�;4��M?���y�!���a���Z���|��B)s��J�� S��yY�mo�����9)�Ё�"��a�ݓ!�T�_5tŌ�!YJ	+r ��[e9S�nd� DC$6��$�{�r�	������P&�+:ҁ%���0/�V��]/�.W�M9��5ۗ��Q�>in��$�?p�3�Y�d2��⛲0�_��܋�"������Z~�z=L�FV]��寮H�A3�0�J�~�_��Ԁ��$px��2�p4(�=�R����f ҂̠A�o�R���.}�5�38�w�=5����ױ|u�BbD*�mJ` ��8��\|��_ �������!}�2`�6���5W�DH+M�5=��ϟ�aMg.��zP�~���@��i��H��^�9\i(ZH�J��Os�������,i!���#��"������0���F���Fhq]/Y�[gɈh:������\�0�ͯ�����y����u�y��0XV҉ŷ��S��-�t2�,�,r'���
x,��ZNIMb�mh]:O� H�Q�	�h��~2�}>����B��~���s��|��i��X��HMc	a���5'��U��\6S����WT�?���XM�jJQ+��zT�s�r�[v�2�ހ��^h�ۇ�D���<���r�:!�WߜBU�t��v�i��g;��X�w[�9yS\y��2���p\t�[h�)��X��ɳ�L,�|{A�������me�}r7�M�Ls�I��1O��=V�� F�H��W�;�F,�p�/�KgC֒�fTa���<�����YZL ]�O���yOK0�[�\��7^4��˿�Y��;�5@�V@�.j4)[1�(+� ��'8���l�*0����eJP���q���̟Is!�;�rU!�����e��P�,���_�~��!��A�LZ?:?zo=Y�%Ĩ��>�T$�Ł��Ъ��`�
�䊅Ր�_�<�ysa*�b�t���/�;��]�o(�Y���`?}�">w�����0ʲ�ړ�If��Bւ����^do��נȯ��uu��%$���,{L	ߌ�����3���YN�C�T%̒wd>��3(�CkaZ3{@��J�lV�uGw��;KN��G��� }̳��P\}�,�e6��,"ÈL%B�]aΝ$Yc�`U���.᜜.���� 7�{=������Uþ�xi��d����u/�����siVe��U�#����E8v�*�a4��okT�땮y���o�0g���1���x�b9�U�E��z�G6VF4W��V��|�WB<�-%�X#쎕����L|����(�����Vc�J�bLO�C⊋H�;&�9��$� NCBW\�@��?�1�=t>��w<��n���?�8Z��Z��.�^p_Z�2��l�t>f�ɗ���k���T̵�Y�)�8�&�g�?h������3Ey�Gz�V�8V���^�[���P�M+�U���e5�~��h�gh�
�!��$�U����n�g�蒆��N�-hƞV���-(��˳i��j�t���'�ϖS��&7�ج���z��.����>����z��������Y��G�Wa���Z]ɹ���� ��,�@����X���R��d�{���\^K)��*��r-	ˀu���nݱ g1��:1�< �z�7s��j���☆�RU\�X�����h��̣lp4[�\�u
��u�D
�]l��|RY�/�"Qa������>�<�lf�2ob}qe/&��\�/�OA�N&:����F�Px��F��D*.b<��l~���S�q���ky+�}kp|��,�%{�F����`��f�b���0{"U�'bp%g���\�G8��X=������z��dfѸ�����n��ì��L���\��J����`�[�N<⒥X����[�v����@ȫ�fDO�Js��dL�ډ�2gr������;����s��l٪�ݪM��\��nh��/lTBs�3�D;"�r��vR���ڡ�������O�h���h�]�� ��BU��KSZ�WJ�0����#bi`Id��d�3�߃��;/Z��WZq46tc��#\&q`��רD*�a���Jg���u���o�Dn��TC�yD�	_���y��z����@��oQ�B:�{s������/s{��;��73�f&���#�c�4���*�<���S�W����+�ES�:�)+=H��N�r*�c�V¥Tp廭�oI�>S���:w#�ȝeͶ�wĒ��O��4r�?�3ׄ��J8{���]0�C��̊;Zr�?���>e� d޼YU��I�����s��b#��IGS�׵Sh��;�K��h�I���ҵ�/�
4&��e{)'Ь3gCku|��ί`H�����_��19%���X�!-�S��[e��Aqo��BN]�j����l���\���ۋ�X����$�������ri��!cF,���l��R����iyXg���5�{80t<hnݯ��}6����'UI��Y(��2�3⏌�b�@�B�I����w�%3��`�mG�݇�L[�UlB����hgGkk����P�B;�2gk��ڏn{-h��E��>��8���s#�n��o�0�"�.���������:>�I�|2�G�ĕd5b��*��$Ydt,�OS���R�W�'6N�uܸ�=x7U�wo��f�^�'��@cB����-gt2���Z��T�RU�[�SU�fM����P�+)�DjD��3NéA#p�d�<
�}�`�BǡQ����91��tN�"_l�ו7����l(�>;�Pt^�������M������R�縮���b��0D��F �K�%y!���-�K�Z�W��D��k���z��fv?4��L��CqIFS�~
���{@5_[mh�~2�M9>�J�Y�k�a%-0�R����E�?�H8� 8��m�>��s����,� ����\�N�	h��f�(��W	�`�������4�N����&ՅC�v�������u���}!ҜlV�U3��'�._jS����[���t$�Y23A��i[��;˨4-��� qG��M���`�km���`?k3VK��(�-еj���?$�"�H?���%��_����7y8�P���kp_�m����^�D�H�е���WT���,-�+2L-n�I��~�&h�5m�$ �Gm�}�<z�M�:E��(\��梋("?n��P���׶�T��|D$�������<p���p*X�SXX�y�������z�8R��!��:�a:�{12DX_�>�B�}��u=l#�١�T~�Z��/,���U�b!���0M�Ę7����y�M:y��֑���e|>,:Y�ʽAp���-���PR>��8�u�AS��g6�_8�H��s�n�����~�&�n�͐���"K�'2OƲ�����6yӛ�r���!�Z��prf�cl|#+J���fBD��E�Э?=j�s������u�x��$�߂+G�D^܊�L�G$t�Z���6�'��7jز>�r=V=�A�����.��
\rM%U����S�,cț�
�n���6��LE�Q�"+��V��GL����w"�Y��&��'SO��|b�P���VƜ�'����+ݜ@�,e��'\5=�G����� z)B*2�"⤝K�Of��6M�g5�2/�ӏ��Ɲ�QO��*v���l�P&���P�Jז���r/B�L�X!cx�c��L\�m��
1xKuR*�o�?�,����8�cB�Ѫ��*FnYS|��Kd�h);����T �VP�EE��)> ���Qpw
u3�M��1�Mш-u��6Qb��w[Op�r����\�¸�Iw�q�!�HrJ�Q�R%�3Ӭ�_��X��<G�j1�b���4�u���k�����1�6�0��������l梪}0��Ϟ4Ȋ<�x�s�Φ�y�E�eb��plBy�� d*�B̾�Y޲�ܺ�x�x�i�:/�H/�"����ӌҳr�Gz���v�f�Յ��N�0�����4u���Z�X^\P^�yݺ�<��"�M�s��s��h���mQxrK<,�&zo��ek�BK>������!�{qUQI���ReyY^IQeU�k9�f���4�
�����y􏋬ك��RQ��|IU���t Ґ��ڵEY�g띉�Gf���*�@xT�h���������Wؙ�'�.u���7n>f��΄7��.�d�v�9	q+mr$i�1pvӒQ2���R���Oざ�o9R���Id3	�3�e�4����a��U^��y:�yZ}>���d|!��}n�YɗA�Z�ܔ$%iV�o��[�S��������?V�/��=��c��Kx΄��������aw^���In��R���8c/�|7��zT�2�K맧����MA�����V��gVv!o�,�T���M��ZY��'�V��}����՟�<?�'YH��7�Nh�Ȱ ���{��I�τ���2 �r� (l�L��2�6ڐ��#^?����H9:���p���/t�/�/|�&"_���K�;96W��4��FiGsTWim��!9�ϥ�|��.�	[�ң�"��[Z�64˘���JQ�uꯈW�(�H���mnG��$6Aź�9JX䔘�a�əP���Vn88��2>�w�C��܊����~��̃M�rA) 0cW3Tm��l8�:��Z�f.�Lb ���c׾��۹l+k~���eC_�P�����Z�U�}}t�����S�oT�g�'g��G�E�<�τ���U�2�#b��?D@�C��e�_GJf;_�'��^��N��ә�ܓ�ܺ�،�q�y4��t��鿶��7�/a��7	v	߉��?�g���t�J�4�j@�LEP�W���8�}��T���L5,P�
�:.z�c7F���~���A�O��I����茒�
�45$����E�k@���>�(侍+�ſK�������x^Ų XF�^o�ep����Ͳlb�V�w�U˜h1ޝ��d�0�_��.�3�2��wΰ�'l9e��g�8��S�5�)�ʶUZ[H]L�Z��%^I�Vz�aԀ0���S���њB�&�Z��]X����2��T
�o_zW1l�`	�P�?�������20s)��);����y��J��~pMp�x��d�h�%{V��P���Dp���&�A<�e�i��ֻ>�b�N�I�C��cq(\Xw�kM�������B�A��M�!�x�@���ϲ����҇Y�a��-Wsr�2���5���[h�­A]'%�p#`�8`	����V��FމB��v��BQ��
&�!�ݦ��Ǆ�Nn��b�+�퍐�KO1�}G�q����c�ܠ�E����z�a���jBpD�i�Sqȳh�Wu��]��L���k�33H�I�!�?�~�����@�m��Qڮ�߬���s�!�f����;�A��E��,�&H3=��7�Q�\��[T_�ց����h&�45ա�k-vs7$|���K�H�;��0��U�FGG/#{@���%�_S�r�
JFG9A���j�^��w�xR��*�6u�N�u�|��%ԔL�]�Z��a]���In��Uw��;�������sS��������q[d��)��n:��it6��7�Mw�]z���7��7^Z&^^�L�.�J���*ZO���1{��� ^�HSK-�K{I	�����a2���F��W�Aģ��g��P+�_�؊-��/I��\�Ad��=q�̫�[Ӡ9a�[��O[��;���)��	WP�/W��� 6��h��Bk��o������e�rmU�ZUd�=�]O�$��J1�B+M(�F�#��V�Ȧ9B���4O�Q4��k�cGH_IYI�S�<�î-����{X	x��R"ty�� C5��$�_h\�f����g�!)Ʋ_t6_�a��y��~�.�8��g,x�t�3� ͖Ezk��&���ɔ�- �1���e��Z��B���OY����&�|%��{�nR� G��|��Ba#p��C�`t|���g#_
��t�����	��^8�X�Y��T�jl���DLh o?���(:A��8Y$�� GC:���P��sο�N�a!=�
-E7c��,�|B૭��(rQ��)�`�z�H��ـ�n���4�������K�;�(+`8�8pf������]l���X@kS�h�h .����
C���O�dC'�&�'ǒ3��ERvE�&�q��5�3܂�܂�W��R2X)�
d�꿂�~���[��%�?���t��Am�!NrM9|/����8N{[,D3k�VBH�h��b�]���;��pf���+߃�6/pu �X>��p�������U���V"���l��![*Gb��e8���'t4�[�R����r��n�|�l�'0������]H�@~Nw�M�,��hF��cO����8��__!�k:�t�e����K��N�l��nҖ�;{f\{�R3�/�����I�'�����I��G;���)%o�eF+TݘTwW��H�"��65)�
�D}8�{�J\��I"K������L��c9��p\M©EC�^(]��zkw/d� X?Mڭ�I	_�,��	P���7�F�XU�Ę��\�f�Ja�.Hr,�����i5R�˥�6>4�pA����:td�=_7(tY���w�V.5F&Z����v����2��(TֱD�1�D������@o��d�i��u��;yڅ� ���0� sra%�z4�4k��b�Ox0��q#
��P�%����\Y*�b� �w,�J��,���g��F�]��8����|r���A�
�F`�x���X��L<m+��%�7���.�J��\�\�W�51@��Q{��XcQM�Va��p!)���M~���Ɛl���赖�EFF֝�JK�K�)*�(��^T���Ӫ��j��W�;�ֆw�ah�+�*#� ��d.��V��
�17`��L��ڜ����6��:3�|7������/�����;�g���ܜ2&�4�:$+���0~�`����0}������A��!=�AX�ƿV�0'�b��S�A<ګ'��\XV�~���*��Ql��$Ki��r7弰���%Ih[�o�5L����
��o��+�g�+t O�R��6㴡������[�-�-��x��P1ź��yG�K)B�D���p�bP�������OV�IQ���QY[*������f�;KO1��[��mZ�cx�
���>����-�Q�cm��ui���=���X h�l�0���@�ߌ�n��7�1wS�h���<��d�7C]��WQSF?<��d7=��P죘hʹ"^�ucb�܈�����KC�����,�C�؆`ڈ����*$a�����(��*B���U��pL0�����:6=V�%�	��`�ݠF����1��+޷�a�S�5�2���c�H*R-`X^����I�l�^�fh��K䊜n	c�W�>#���K�͡�gJf,f�Fz(U\lK���n���x� �~r�D��Б�.�Q���Hϼd�<S��+|�Y^��_6�S���G>R p͎�l�K�73߽D[>o'���e�i	��.Q�9��&g������o�e��v�Lǭ��!k�hH�9l�L+��j�}�~�!���F�~;�)�%5��_��<)���bt�����$����?e��ϋ�p�{}��A��l�5Y?�菱 B��0���#���t:೹C�pf2��ļ�T�����>p�S�p�z�=��yp�gl������ݾ\��z����1�Ue�SÁ,�bIȲ�@*e��m�!C����Sduc�k7��b��Ѵ�@��J�ME�kօR�S4	�[�)w��B��6���F�P�����Q;�ï��Q6;�ƒ�"��6_��3L�F(��*���O�[� �ڌɴ�*ۘ�n$�]m��#e��Yo�i O@�(������w�'�CME���N�}�����|`�?�QS��w�X��~%��D~ �T�UdH��.���t��㭢����J
�Ѵ��$ӛ�*7��G
�Mp�us&[_�@���<�jHz������sF@������:�:AE�ٶ��zP;��Ah���?B���[^H�$�;({\S��Q2G٢��n��Ȅ����H��y�kb�|$_1��wU�oY��O0�L�G�S� �.��I�:���mp%3��\F���^CU�s^��w���O�
�R�������ʑ�S�x
�
u?+���n�F8��l�������s*p.��**�^����Z�����A_�"7I$���鎄ϩ�$_KS��'/����-�TU#�ɝG������IQn���U��^#���w	�[²��y8<{*K3лd�"rZ�pw^�b:%<*Tw.��EW7�}[�����4<�5���Cr�_/:_���i��f���ON}{SlZ==��� ��T��c�-��h�m�7h��BN�E�w��8w�స���[��,�	� ��u��U}�{j��k�8�s��F�z#dG��.(�ľZ���}��R]#�R��d�8_x�y��]�]#蟽�2�z�[c%�5�c�+p�=��#	��+ݲlªm�ö�6�XMƉ������Y"�f3*��?���`�����4���,B�g!�ZS��_y�¯���(�`0y�o_��~o���<#!?���,��h{��=�E��x�H~�u��\�O�I�Y�6r��"�Γ&�����
��z����q�l�~{�d!�h!Pw0��M�q��V�7�M��xL�a���ֿۂ�&�2�!T�+��o�Sh�I��2��q�O`�o�ߢ���O:[����|�l����$�1S���e�v�)8i&4jލ��S�h��`n�r� ���ˠ�%�K���a���x�9����އ�K�7x�V�UV�|ƏF��(Пr��NԸ�N�fB*��b"��˜W��2K�����ŀY0�YҸ��GW��)	�i \:m���n�X���������5�C\p��7q��易�J(��� �� ��]����up��me��
�u��lx ���n���#������m��^���,�hJL\r�� ӛ�?c�&���㥙V��;��x<����Z���il4�ڧ��HaI�}�2i!�!�٦�Vv'EM�C~��n��P;����!I!I8�
s�e��o�#x�fd�Z��s=����|�O
"�銒��Iz�����i��HG��(h����?�T�KX>���)Z���bÞ�7��QE��G� 6H�D�2[g��R\�'+" F�l�6��[#���Т�޿�_J}�Ws��t(V��Gl蹫"�p�X�vŹ^ 2W����ަE~JN�̢b�y�����?&�&1�o~�ͺ�F��a�f+�/kӞ�V�]��d���>��9|��EjZ�μ��D@�#�_���L���1��c�c��㇙T��[��΅�Q��9���I��D�{9S�k�?{]T���{~s@���/a�C28U3�D7��&?��P�]I�P%4���:�}�V�\r�T����������dl��o��)P�t`ॣ1�}�.�Z<9K �����J�[��"p�:�j<ݥ����0�Ag���ĕ�y,�,ZA{�xv��vQAo�q�,o�&�j�Sۮπ�Vt҈��v�G9UfW>4�����u�0�J�;��^�kq���s��2���/�$J����z!䅱�z�'�º���fI��G6��0�>#�5�S�R��g�<�H���	�1�ۡ���T�C4�X-�w���v��,�>H�Ԧ��%���f~�=�*b2����*x���p�����z��Kf�f�����D��AU�!3l{f���q�H�a_� �;x��L,c̜~dLÒ9�0)�K�����pMxvv�[����cR���������M���P�ǿ�ۊ����7�������mng���3�|/gKT���������Ӟ�svFN�I����x��� �����y:��+�髜��7W�y
<l�8T����V���&�G#�)����4�Ճ�pQ��$�9�����������8����	�QW��̄t�B��u�p��$�;k�]�ug��4�&��E'��ZL��Ao?�n�8� �e�2��|�4��]��	2�Uw��}t�b<�S�f}�����/a�VG�S�SAgW�S1	�N�Y�����Ւ��'!ߕǢ�}p/�Y�r��HA�n�U�vE[��J:Z��T�u�����aO���9f5#�:�_����ꗛ��ٔ�����`�C>��$�"[��+�d��"$�Ҍ���9�c%qZr���v�D�˖�쬧��Rx��l]��68���^E-��uD��ZC���q���<�u��_&_n��/�r�~���~J�e{����r�_�]�'fȨ�#�F��q�9�r�1�p>Wq��D\��Β)=�"�_1f����HM�����al@�M��x�������8��:���<�j�3��M��aT�PK�� *D2� ����p, ��̅���4�` 9�t���C���i�w�] �����H������\XGQȒ�.��6R4�:���ྫiw�f?��I}����U�	˜�4���_K�_0]rV=rVW�V��Bxe�Y�IdJ�3D@k�X�v�96σpu\p���|p+���|�|PE��2����	pd��Y��Xrw��͐�L�F��޷^��˒�}�,A�C[�Z���9�(�ɠj����HM��}_��[�LdL �&]a��xyԅ��.8�����
�s �v�3{�4����}'�"�Oף2�j�H�f?�`AH���_����7f���ָ�J��i�d�5�ȬW2GB��,լk��z_���\Lm̃!���@>uy�#6�e�g<�uǨ��&f��F=ͻ���"h�VtQ/2���IW3�� Oכ�j��F���zW��;��J��Yq�h�-����TiPW.NP�.�{��3�3��9xڝ�f�<�r|� ���`��������4�G_�bϞ��W�lE�\�U^�N18S����h���56�a~c�(��0�NU��c�x�bd=���xkci�B��
�m�Z�,�4U�-K�.�G"=pِ �7�o��XqH�x���e*��4�{'�\ϓ��z�$��q&�є���U �F�k�}<�����)U�UU�T�ى��7( ���a�
a#c��
�,sU
~4����s��ޯ����'�h�L���P�g3K
��D��(3H�B�?�^HIDMLJ$n�o����jrTz`$��7��r�b�m,�-��R��l����!e�U��r����_�g��P��$����B<0!��H@EAtL-��t��3k�p��2��ZMd^\]a���`a{h��#��RP�B�#O��Qă�1���L�Y4�Ų�
�J��@��O��Y��@ٸwY����fig�G��нW�����>?w?��=m<Z���d�kW�e���ݗd1u���k��>��Z e��X;Ew�J�%)2�����u�l��	�	b�e�n	�%z�dañ4��7�����\3Cd% ����U�$ę�UM~J�P�?2p�z�ۿN3��ݲ��r�	-�A���Z����[��JuL ����H�6ZZ������3G
�7����ˬ9Ȯor_�|^�Ĕ��2���&a�8��1��i0ϭ��"晹�ܱ+�-�](Գ��-��CU�[$aδ�lC��1b�3�蜧�IKBb	�������D�o_��_R���˫�\�����NF�լ�i�a"�s�:���v�v���$'�Ri������b��~>�r
���Ȅ>q� B��3��kp�L�~���r���:�V���}K
��0(F[�e	Ҭ���*��`�����l�J��$���R���)�{��j����?B:ŵ���b�6�J[�&��Gd�?ԯǣ�̀�
��b_�d�����D�:F ���}��_k�-M�ڋpiF��#�w�ft
��@�У����F���h~�[���Y@�R�HpO)|;`w%�O'/���?7��F�%�v*�c�vO���n|)w��l�llil�_2��'4��,���}��6mN����>�^����	\�އ	�	��L`�~�W�D%n��6��DG�f��f/�]5;$�T�S ���b�1�k�����"=�2 SL;��گK�G�/�
� !�&z���î⾦��-F(m�V�xJm
�H6̌�Ho�YUQ����Y�P�����9��I���hG�j���h�~W��zխ������MgAإG"��6�zZ�Y�����o]�x��Ӟ�8;s��������ި8�$��x]},�W*:�?h��.����-���j�ꚍ(0�@i~X�Ϥ^3��x��%��o0��j�RY6ud��K�
va�'�`���X<;��
VO1�wquH�	�|JjJ�g���֬�]�V�:Ƽ����V���̏}%V�����>��Ml�2�0i�]*����)��	���B%�d-G���rzZ.��s֠�9��M����c&u�>-�A�p��u�x�5\����Rk�)��J,�iqpD������5X�}Q���)Guz�k���P���ĘC�Ա<$��2�b���8Mqt=	���Ҭ5��m�)��c�1�T�/k��:�����s�:�~0$ӡE��~�ھ�/3p�d�m����Y�����J1��"��h�5���&乬	.�8�L��C<{ҧr�§6�68Dsr���D^��:E����������/گ���q.���}�;��(�\-
�E�q5��5C����1/�1(M����$��^��_����w��O/�W���6NMJJJ@@�돊�������)���M���i�kM�1��������}?a�9_�a���[� h����.|sN�S��W��?���"�;4gN���ZGߢ�z�*es�U|O`D��5��������V��t�]��l��t#�h}M����KGM�0�����<���L�{��1�5�[���2jv�R2���w����C�D�����DQ�ǝ�vGuɪ���9d��Q�?�lt��(����{|�?��5�3��*� :.��$l>���������(�WG��$9jJ��w&Uڝ+�;�$����a!�J���Q����,K��u� ��K��UZ'(-�P�=��j��a���jӷ����O�]?�\zZETV�U,�ڀ��Y��fb��6a�{4�N�RqD�)�u�`8�ɼ��4�<�f�Q��zG| Qn7�g�#�nץ$�����o��q&���P�k!?�"U��q��j7����`Ӵj�9����*�fD�]E�z�-ȩҫ�M���������!�)c��&Y�om���z�yY��P�MY�'�!�XA�une_'�u��Ƚ%" �}��20�>�Z�j���	Dab�Ŝ�	��p��u��9%��F��SF��H���C�~D$6:	tt&���?H��ߣ�E
X3լu
�Rs�Vޭ��%����ߏ��՚��ǰ����$��C�	�'�� 	>&���	���.���K:��]<����wO��3��pu�9��f.!����O&�	%��TH/��P�S���tn]���e�C�(y �b�����W�i�ܺo��ccP�8�v@����/._vFm���[ֻ�:f�A��&�>�D��B�%�:�૗{��%���7���w]��<�g_C�.�>:�:5�=��ز��c�ɦ����<�zs!�� ����\XC��T>A�'"�^��`��l�Iy�@+��e�a`�!�S^٧~��>���H)�JCk�\�`il�;0�v*�["=@��m�TX��e5%B��W�/�1b^��	BFCMH�uPE�7��O	N�4�"��/��`dF>Q��ʅ!:�!ɷd<U@\�����t�p372�0�_ʸu=͛>Eq��,�2[��x�ȇ����C;���e�j�Qd>����|�Z��}���]��������^[����.��{��	���U��#����S�Ӏ�=�(m��s���"�!߈�y髇�p�.���ó��u`�b�۸f" /��E=[�x�տߠ�@ǉ-2.B��<h!�`���/�����	}�U����[e^�ttd͒�� N"NТ_e@��<gs��en��UQE/~����% ���<��=V�j���3���!����S��1�w4߆�q�͕�De��vUN&=Bw��<�2�v�-N����l��g�Vi���!J�'�ޒ�6�_�)Xc�25?p@�Y@���ǖjȐkģ���Zє;2x8�_W_h�S�S�,>bWb����^��${���Tsz�e
�ӧ�v��&+�7���pj&�	�b��V�Y����$�4|��s1���б6���Q�B���/�*9~�?U^�2���L
߮��%��GG�wwwy�111qqqQQX���A�A]cs*y�"���_s��$(����3�IW���P��9=���8������2`�4R o����W�:�'_?�).���1!ƺ������+`�����KH�Y���r�	��q1�C���wѐ��}^a��]F�%�{/�X)�L��B�?���N�BA�z�+�<p0 $��+�JsE�"ȩ����Pax�mr�4g ���H�+�Sp����{��\��a�]L���
q�V!�h�S����re|�>��k�~;<?�q�+�?��1���J�]��7;��Z�����F>r��kEv�$|I�<��B,�m�R��j�r{���p����e$jqh�����X#��Xm�T�}�;ꤷ此 ���Xޗ&�:sw0�
+d�Q�0;{٤9��P�˖�������Pl;����vdɸ�F*��N�PZxYfErt�W̄)P��5Pz���A�:�+�1�~�q��q:�M\n�ɢUH>(ҏa�w+XA%�����l�WF8�ID}�'y�{Z���:��odi
�i8މ�-K��e�+/Cj�a*��<��૥�P
Nz����$�C\ 7gL����ē��o?O���'�xf��޴�+�em~n>�@R��ׯW�Y*Ɩ3�*��{��ʻ��3������Ƨ����Wg/���������8�Js���k*�l~m->6�8�2��u��V��< ���L`�1��gF[^��&t�w���$�����("W�x@)F�w�����hǡ� oz(�Sy�Z�6����\�aoM@����`<�d��.����9��;����(�f��X�Uu������<��w���g����� �,��_�aZ1q��,��6SwI��h�Oto�@��T�|����iu��r�1��	�o�&M�9�����-�
��A���[a�o���Z߅�S��sֳwl]s�����u�4���$q���y�խ(.��{��.&M6a��]d�ʧ��������WI��7�껣��$�~�n&�ާ·K�u���T����\�@�:�;��oa[স��q�j��@ܑ���ިB�.1 �E���K^Pݮ�\q��g@_0Q�ր�Ӯ�9�|���,�6=�]z�L���k���Q*7(��M�g4�0���ҕ�K��yݿ����cD<���a.��E�;�� ���9z�W/7��h�%6�S����?�#=I�u��f����K�U�4l����Z���Cn�n�e$��LC����Q�	3��k̭�h�ǵ�,$�E5d'@IS�)����	��{g���'En���=����������dzFFF~~�>

��򊈈�� ���������A�D~�y|/�d*���ԝ�	%p�M���V��<�$}�Σ��~��X
ëV�l�����:u��mr�	�!6w���	����"n��ǆ�h�Au��o��0~X����4.�Nk�jecf2>sY�reJ>�T���R�s.�R�&
l��֦qB.����x��4	���_�kB	A"N�y��ysA*i܅����, ��D	�6�.yG@��PO�A� 08=�WԾj��w�i��z���Hi�ܪ����W]�u���%a^c�U���Ļ���L�`?���h�!�]r��k�Z�ĵB�a�:)��M���r�k|qj>���v�5���T�D�.�'���s��(����N����Ȉvx�y����Vf�uv���4u���%�5�������~�;����]r�7��+ ��چs�*]��C,�4nC�&�S�|��߭Q׋�}��{d~z�$�G-��$s\�a҈_�
� ��<�wcHKJ�:ö\0��zx���$&�����o�?�5�����#���uL��|�޷�M>hF֬�ײ��"L?bdɛ�f���8˴�cqQn:�T�od4�*��-6� ��L�L�ͥ6/������W���^nr�o#�׻ݼ���<��A&kiM\��_�$$G�Glup��`y���W@n��U7E~�6����ci(l�!bd�k�@6�p?��$�9�2�����ÐNh�diӷ",�[��ɱ�s/!۠i�̰m�r�l��U��&,��Chc���^��! �*�^���D]|��S�g�J�J�c'��kS	�b��V�-�V���c��~mS�+�NC�T���OG�<R�9t���^����Ca�0FVnQ�N���������s�G<��>�zC�ݾ���ۍ�r�)J ���˶:n��]�#C�y,��]�+u4ҩ>D  ����,���#�7{�/3���,�K������2��m�m��J�t]:1`�#��t����r8�`�Q�[�,6?����̈Qu��t��'�_c������'��SR��C2��Vt�ʛŁ���+*-	�-�_0�]�4􍸹Ht�`�ꂨ���
m�e42�v��p���=���*��0�R�i]��G:k�D������<]�N���Sѧ�\�J�����
@����V��\����7���� z���ӠNS�%!iI��򊖒�>`[���ւ�Ƽi���y!%�!��<$���������vFb����_�Fy6�K��D��?�%$����E@�OI�����¿w�{{{MLL�O�%$$LMMPQ�@��5��~��N���䶜��������hnaή������ֳ|?Kgr�"��A:W�g*M�h�B�~j��hEy����r>tޞu?�?iiu�8뻿|�	��nRO�Ϊ�T����V��7J���~C{��nޤ�iC����3F�&S��:ppcC1��(
��<Q�Ay0]���v������Z�n~G������r������W�V���H��cz��c.޵^��I5�F�H��)�>t��#A��vp+3��L权Dt5C_���ګ�6n|i��������h�Y�Ahy��2e��V�ٚ]��]ޞ�L�U?st�F�3k�,� �+UP�IԒ;λ�n\}U�__�XZx� �{׃CEq}��I\��K�1��l̃X�t�Փ�ش�\��P�N//}�:n'�O\ۏʅ�aϧZ
R�r���VtA����qs#��36,��~�%�S��!�}��oo"�e��?i4��� ��~g�x�[��u�Tns����
,ԹQb� ���)�~J�|}�}�sn\i_B�������c�Ig��گ<(I���	�����	VK��2��v��ni��9z�&LN�s��
�xs}��W���J�Z՚�+����:��h��7o���4־�*ߡ��ۭ��8����]��Ѐ��������?Y�����~$��)?��g糊�X �)'$�ip_� �P�||�k� ����wǮ�����/�=�7uoh�c�0��f��m�>�ODn�g���8 ,���x��%Qp�]4��@���F���u��CwX��͖�{['z�b��/&����mU;w�,s�_��=���+S�ť�R��a�(�������ʐ/�����+􃮐�w�g����V�珦ұgˮH�l��<���ׇd���|��.OZ��[��=+͇���dO�?��D(�p�@��i�w�q�]��1�K��i�k;���yՋ��n/׃h��n��+�[�C!��l=MǬ���G�ڕb�:h,4\��0r@-ϺBN��0�y�=0�������C����J�y���Թ=���%�;�+й1�X�=����'zx��X}1"��+F"�*f��
U1!�d��!���p�V�D��[���G*�>ꬂ�#���W�a)���M�� ����
�r<q����ð�
�`�8aI��]�@��"/����l#s�4��|��e�N��i8ܜ�dd���}�	lZ��Gs���w̰{�����J�WYF*<�3RH^]Q���������������rTX���M" p��H�����t�j���l��"?��WBW�;	�-��y��8�K�V��9:"'""���z��-%%%!a�w,2666..&#2#6�m0�{dB�Gj�4�t��Ye�׉I��g��O.�)��MK�(Rb��L"[�t@�gc'�.&o &���8	�=�}~j^���3j�;Z��_V��(ʯy�b�6ڐ
9�*�7��́�Ⱥka�̀���y��H�Z�dJ�:OpM�n��)�	�;��m���aǿ���\���B�3~8�	�K7X��/c�d��w�C�u���,�@J�@��J%�E
�����i��3����6��h�g
���+�yK�I���?f^���d4�*R��������VyW�����&�q��e��e��}�h��޲����mT���~ �H�Pb���!&+��y��ԉ�_�m<��^+f�t>ܻ���M�����e?��=�,I��eX�斐l���`�owN�ٻ��}�f®��G��
�ݭ쥪<��]��]*�Dw�&xa$���F4���N����D�,L,߉i����nʫ�>��!����<� ���s:�1R��뿬����?X�[.vYVr|D�J�$F~����H��Z[N񫪿�k������0�3�6�yV���cr�����ƙ3����"������Lt$���hY�	���s�<��x}�����Wdn�s�O[Jk22pXշom�n�Q�q^�mÍ�0R�,be�W�� ĉA��%��<�a���������ߣ`��\Ъ�n�<I�d�"�nRd�O����|!�,yg��#)�o	�mX.�;ԲXn��wO=���M4v��_Bl]eFP[�����������e�i��V���%=�c0'��5^��K/�<HB���i��}f���At����O��k��j���N]�i:"��)h���ȤQ8"�-I�r������&ϔ_.[7�=:=��j���2�-�˓��+����c��m*G�J��e����؆��"0�܉��Hu�ȶ�p+�=)���ll���\��'Cu�Hr��8A�g{����|�$u�]�[�o�`VPA�+�!��~���h�Ҽ�C��ׄU�ؼ{��
����J�k�zĀ��i�toK_�������P�����vca�޺~hƀk�hIS���:��[�'@��EX1q{��!��7�d|�3Z�HʣGQR���ˏ��+�M��q�F�G��b��M�����=��R_��Lm64$�����|q<:<$��|e��1<��]H_?�x�j�n���Vݨ:S��%դ���%ȑ���jӿ����>#"�t���������YZ:�W!���53�����-):LMM�.��/�L�L50��
v����?<��cy�yȟȶT�R>O�ZnzE�!���.�V@�������,�����!�j���|c��<��~Y�%��r[�j�KV���U�5@w��58�z?�M;hk��
x��^Qo��N��߇�9�h�8�I����gMӁ��R���5��ս���w��X����]X����Z�D��Ǎ�.|�Ϭ��� |�slGx���/e�Þ�c�*�o쬼��j���m�WG�����u�Qg���F#�ܒ�~%�uE�B*� �/�8��G�����ERd燊P�i� �
SI�$�M�M�r�I{�t��"	Cy�؊����Y����������O`������Y{��!C��y�$nc�3����Vo//���v��AUG*��&-%�qw-�ƷcM;_�+����F�y_#̓*��eƭw;��0������^,%�T��L��t�o�/��*�%hkXboY3)n��ެtgf2�CΫx�tC�r�*��+�mR�De�2|�1b���A���_'��C����0r'�i E�^�S[�+��!�v	t��b<3����Ul٪�8<OԱ���hv����rw��x���Xy�ng��fk��zF~�Y������j�w|��*�I��B�J	0��V�$�y~3{�J�F�S4�8�O��l2�����J��š�e��En3;��鎍��PO�=T{ҏ�p�7E�>" M�=�4���Z����:?4h3�/�w4����N9��j��Kc9_����/5�#% ��گM�vu�Nc��Ѝ��F��!��ja����P������NW�uÀ���T���*�qk(��P�1��f��M�,�j�P����a�_̌��Fp�1a�-IG���He�FG�ߕ�*}�Jd��s���:��9�ei���0�iƔ<��xlA �,��!K��U��6!��Ux{�D�����۽��q�k�"�Z�Z��o�ɻ<���a���} ��)L��M؜����=�	JE�A�X@$�s�oFhy��`(-z�] ��m�LCUI�?oÁei2�͑uZڤ�Λ����Yػ]�"/�	��f�%��E'�a��fY�z���������ޜ��;Z�u#�~��r.|������@B��
L�t�r�\R3�����֤������RGTC���,�
5L�������e�K����m����Wd����Λ8�۝/�/޽�'�ѯ�l�]�]Z��be!),�E�X$�s��uV��ďWˋ7�����������,''��lllNS��m^ݑ���*����ACC[B��,�.�}+ܟ(͕��.�2��ٕ
n���I��L軨�^q��7�V�l~	�o?.%�`��r����z�g��#>g�/�'B|l�v�Ė�+�Jw�}h���p��Qt��L�%�߻��_H����y#�p�rj�"��#��`C�;H"�����~,��]�l}Qc*iY��H�Hi�Tg��j��5�~�9��юQM"�c������&%�O�ִz�]���aBkf~,����!��_�oI"�&2��e��_5R��G��O��hc�Q*q��X���O�<z�BF��|d'kg�����W��5]�i?7��l4g����Z�O�o~,�,V�Y`�+��1\�}^j�Y&g{��	W ���;5I2���*_�\t=��+�`�I�Ӌ;�7t�8�&=u�����+s�ӻ�N�K��'�KFW�bף56~��s��)���6��ߨ�K�c.e�Â�6�s6)�;���D��+��p�霁"�����ӫ��GW�@3
� V�h���v�~o�&�+˃HRn-�ĕHB�K�iA(U�c�&Ӷ M|x�Z�����*-�v���ఘ>�"������{�����F�(]����d-Md��ף�OW��e��۵���}�~��}��M��t�<��rWD�j���ud��B�⚒������R��'7�$�-U��Q � �|/�m�"��d�q �%3���o2RҌ��jS����nJ��3�yZ��&>:]��NpC��'Nhrݾ4����&�s�G�3/�eE�L��B/-�'��qW�ݮ�gQ�����6����ѺXϧŭVζ� �����r�>�7P����`J��%�1�Sg\�(��^��VN�y�IDZ:�:�ü�f������y���Y�q�"P`�*�V�?8d��3eC����rj���nux{V��;���.h��R$a<� �-����i>�����z_�^�/z���-*zY�Ի�����u��=�ʷ|f�����\H8^�mSM���>���ͻ沠�����5J����]��Þ*�(�Kr$85(���!X��X+�#�QuJ��n�"�4G���$�"�c��5$�c�3�H[ӻ9����zFA["��1*���$Lѷ!"\B�+U�u*�}ċع��2� �Ө��=2e�k`����� TO��	Zb�8,��5�� �N6J)
�;&n�O�TTi�0���{)�!��Ͼa�U��l��=N�,e@�3���i@j�C�3k[;kk(&�u\��r�ѱ-e��E!z&���cLa�����@��m",��ȋZgLL�}k�O�b��>D갆#������)S�����D�Q��:W��U�����;?mԅs����A�x�P����
��Q�0�+Y�Fil}�ה��g�~T����ǅ[�Ź�_����6����ݿ���j�	E��;��q�[�W%(l��qC�]y�J�+e�2�
m�P���r,�?��Uv�m��z��wLP?H�I�9d%�*����GMe��׏DE�ӆ�,�5O��6w@���.�I���S��L�l���8��D�#�*%Z�����Yb^��(
�p���v{���.�*��ΘRMZ6`��?������w5�T���u�cۖ��0n-a%R�EZC���H�ꬠ�����hd�Z�zE�y��^}�qE�DU�X�M�R�Hj�II��Qe����k��c����n)�MzŇ!�v�Ĩf�.��kkS�`u���=L������FH�vjEdݒܶ�f���p�8s���a��کD��`�x^f;�r�W�y�\N/Pz�b�pC�s��u�1/�ۀ���PA�s�W�^��V?
���1�֦��r{�T�p;��\��P��wX���n��93��y� ���=���;:��N�P�:[D'��b�\������s���%h���J����jϾ@n���g3kl�͉�̍�U�
|��9R@��;"�����hΫ�<f|y�w}���s[eZ�0�oh�r��PUNv�o7]�o:[8fKs')��-�!fv���6�|:�r:��l��t�� st%}ս���
�m�����^ �?��jnD1�|L-pTG�K�����<�ԍ��â��<Y��r���@z+������He����FĻ��,�Fw��F��@/�xTR�H-��ʅ&#�rLaiQm�PJ�k!���܉�o�b�%	���nM7R�˼ݢO�3�qv;����fDD��~/�ܰu:٭�o�h��y���~�����������o�K���������KΏ���}P}�zT��WLm2����=͘ӄ�B���!����Ng�6;N&y����V�m��,��ѿSr4+���5H�����v�p?��fŏ�M�>����ؔ��ގM�����d������ST�t4��T�{e�Z�v%ɲ|�[h��ԧ�����hϚ	9?;��,�O��ۧ|L:���~�&>�9�{��'��G���`��-���x@�1����|t�*�jm��܉�^�����AZ�Fÿ���4T�_�`T$�3���p���L�{�4�,��|85�)����� !G]�����7$4M\�mw�<\��	�������,����:�d9���з��Xt4�3�ι"�2�g�yQ5�[G��aLMz~�tBC���?�F�v
�l	��0Ղ�9��sr}���������H<H�&��d�\QQQZ-gREN.�׎�����99���JFF77wgggee囈�������vWSӱ=*jj)��{quu����?~dg�G�����*($�~�O�(JaJ"`�n�B4�IK��J�L��H�HM#�H��"��'"�&%O ��$}��� ��w"�;3ݣ�р��_]�1]����*���Ǯ����4Lj���>�9;Zn.~Df��g�$�ݱ��O&fye���?-K"��i��`}ۥ������/$9��&2n���ɵ�S���3Nb��,�f*�	4���)�_��]5G�4Ɍ6�+�>`P�^.�2�g�$c��,�i�x�1����	-�o�Yy�R�
�]�l�<�/��E�:)��Z<���<��$���?4�d���]��kb�O�$�dlnHla*�5s8����p�D��c�CG���e�#���롢�����,X��N^�&�=���O����Uа�i����X�|Y���4�7�h��T^=�8j�)�UkʹݲJ�kO,#lk��W(=-͞@��h�Y`�ꐧ�<k�Hj;�rԫ�K?���4�u�-�;�R�y�w�W`M@�9��,y�`�����%�$�aTJl_3¿r��n`@�K����z�����>�)��6�l%Y��M{�z��)Z�G�m5��a9A�a�cL�3.��*i�k���5���Ы�o0o�dS�|L�9	�E4z0�3޴���hxd*��ݒ!X�Q�PC^F�cq0ts���5er���L��?�V#�qP��#�x:�,����:���0��L.v�-�N�&�S�ɨh�Rp�LY)��Q<��e$�������2`
�5X������=$DsW��"�ȹ�?���Xr���sc���]�Vfk�}.�=��Xּ{�2�g2�g��\�����$��jW�%�Fc-���O���q����~�pEֿ
ѿ��#��%j"�)&���ɱ{v���gx��yz��|�aw;��k�m��\mkʯ����I��>�Ռ��,vQ����M����Y��͛�޿��u�n�<z�%�i�F���wXo=3	s�Xe
��	�C G~�.��c�/�b��	���u�l��lZ;��'��7���r;�	��Du8���l�eP[����x[4Xq-(R(P��w(ܝ��xqP<��)�%��@p/P�<���s�3s2�=�U��-�u]��J������fA�?-���A|7�'-���V�ʘ�����	�;��xnBπ�5�e��NY��`�ۻ
nm���=�Q����f'𱢿�ݨ�N�̧���p�����w��<̱yI�vt��|��o��Z�L��"��,Pl�x�u�N&�UmTii�^V�i������]=�H��,n8��)����e-;��gmҋ|�cL�Ë�/�=�G�6W��b{�#e=�䧌�-e�@!+�ȷ ���z��C�x�?EA��U·hO�Âd��Sq��>^�=2�5ɼ���R�
ʘ�\'5��f"�����p�j����@a�J8J���|#e0@a���W���w`��\y��T��v� 0R��hGg~�	\z)��#��B�"��GH���8�ا���8x��	�#���N�Ŕ�'&훜����:������mw�
m;���w�O����A�uo�T�Zzj*�R�>�d��ޞ�:i�P�F�͌�i����S+�wڰ���;L�0&�`1�@!�lc�`D�w���b�g0���lB��x�X�9��݃9%��th]8��&�s�(�<�_<�R�l7�=y�w��E��l�~����T�(WFtZ�-�}P�Ve���V��γ6�hlW��5Ob{��u%/�)�h��u�f7r�z���L��6Z��\;Kd ����*�SƧ��Y�h�?Cw��$	��~�O��F��7�a{�Py?�	�O�qpV��hZ�Y�|{\�~!��&.�����T����~9�}��[|ы7i:~��G-"�B��Ţ
����
�-V%��mHX`�?LKb=�h��j�\�5�6�e�L��Y%���X����ʸT��l�g�w벇��a�4=���J�E���?95�#�F���~-�!*R��F�*[�e�?Z��ψ����k�Q�q� *[x:�&13���+<v��{���6��ѱ��Е>��!@��qʔbύ!���a�K�K,��H���Z0�?��Xo#���&�����f5Y0��Z�Q��X%��p��iK������4����H�_a��w�B7�$<.K��N��ia툠Lz|Gx� �3*��?�}k�eB;GR�BSP�s��Y;V�ӈf��`8�ؿ�2 ��c�����Y���NB��
e�7������}1��ъm���n�k�`�qR2�s/��ʶtb=�E,z�
�!77;�,>z�H�A�H	�P`ږ�~���TH��Jc��\׍bO�M3��%1�0���\��h�{�x�CZ�G�B��W.tP,���~^1���|�h�gD��Q�꺽����<$�bdlGh�II�v\��,*�X��䋂���q-�u�P������#����g��B��>[�m�7�֔ٔ�ξ��c���R����)�#���l�G�C6�f�k���[��zu::�V�v2VRj�Gq%ʑ:/L���>R.��W�N��M�������R��)1˜��z@�r��H���bb%AD�+�����؃�SZ��(�Y N�.�~�èA�4<Ix���g���Ğ��?1tsǆQ�C7]���&�n&�m���J
���R���S92w �*��&z�6YX��%RkiAC�C�[V�>n��*U���{���E8e��B�Esd�m����,���m�ˣy%�h�K�XRl73���W�$[��DD��ϪP>w�v�VO}�rjq�%�IN��X�564���+���*)���njjZ>��BӺ��f<����uuuO4��^��x�GAA!**��յ^�A�mڊ��}���kv����"[��X�Ӳ�����E��Y��Im﹙�s��3�=��l/�Ы^L|�49�k�=)�:��G".0�HV,(%�I-�����%�s�1Ǎ+h���YʺJ�4�~e�oW��w6
H����̬;5����aw��$�ݫ�?3���.�1�ms�ka�R��w�儰�#�/�^	���C��@���
Lҥ������WT�	�ά��J��&�q>T0�� �/��d�Ƅs^�+�T�����c}�l�t���n]��G�E�VO|����=��)��5�|��ؒ%��ϳnm�Y�0	tP5d@�t�F6��i���$?3�U����Ɋ�f�K�;� �}(L�a�X�P܅x^�;��S&���+�lS&�HE꣍B���8�=ENN.�)�3s^�($��wt7���J�1=��Ŝ�FP�Z!ش�.����f�W�8	^	j_	���S{>X�L��%,[kM[Z��k�ӭ��5ә]?:J�RRP~�ؤ�<����W���������"�؉ʝG�������#J�Z���N�w;�@�^DY���у�� �}�j³��F
�2�e_@ޫ��ߧD�@O.7{V������������OH�`鉷���;F�O0T�,°�荸�-�+�p:m_�Q��[����t44��TF���0G��{�er�Z%q��W�^��Y��,8]�k�V���<��7�Rg���r�����-4�� V�߈�q:�O���%��٦�^ݎ~C���\���E�XY�!� ��/^bY��xEvIh=�Bg[��C�o�?��p^|� ��������}�8���52[*��y}n?^��(Ԩ/�&��l�'g�<��|�sYAu����B�Q;N��֧ᎇ�j���7Uv��.7M��x�}����p�0� |�ധ�Hp���f!�O-魍�9M�BT�uM����E�(�8I*<TM�0}b~����c���V�2e?�ˋwE����ia��|ULA6T`�I�s�41�N��w��/	�nSmu^k���|Z�ܳӜg�!���q�#&�w)�%�*V`�:޿��hG(i�)�PL.�L�31�6l���_e�%6�M���P�^z���F�=f�@����C��sE� ��6O-�@a����-�sLT'���r�)���Jd��g�����&����%@���)�� �����*�)ǲ�.f���-<�Ɩ�1�C����p �20�|�RCC-x��%N8�s��_�������L���rj����������֖�s���=�  \
��GOMMMW����V�=E�blb���ݢw���+���H	ó�RV��K�SL[���������[�Ai�ф����~�����i����so	���VQ]\�:7p;�'o�B?���$KQ��n��]b�Q�J-N�Sn@r�M�^zx���\�2�&R��dq�[�k���a���ܸG��'8�e�q��JE[p���~@yUX�XN�1M�]-XHO�?��F� Ά�g(�^b���IOT٘m�V�3�>�Km◊dF$qO�5��t�%�6o,���f��W�ޟ��D\�@��~!��:x�f8#��`M`KD����ĕ�R=	� :���
�/�J������.�]>�vO� n&�a�1��K�$�/0a`Em��+�m\���o�	�v�w~���m<f��q��3o�#��ui���5e��������&8�/AS�\Vj�m��_�L��ľ�Hm_h��Ŭ�A�%d�2v>̭��xIV��s"�J���9������گ�X�S�9�]�#Ǝ[O��X�`�;^'���C\8ԲqަF�Å�<T����75>S�6���\Bɺ����M�w3VnI'����M�aǎ�:&��}E��˥��ú�����Q�mX���;�� zá��߃�fٻ_�t���KO�\�/�X���9�:��Ӹ�@�����U�o"L�/�N���3O�b�ٙ���K-͇��D���3�c���1��	�\8j�(\�Tl(\d��-7��4%vݱ�,�L�W���O6��Ƞ9�W[�KJ�c��(�Je�%h��H�I�Du�'��=�0�AXKf_�������#[P�E2-����.�I���Vi��L�qǶ7I��9�,�\s_v��v:~���d�sQ7��������nM��VL�lJɭ�K�:��C�˕å�(8�\��>�W��8���y��"	�MU��Z.%Mc���q=cW`�k��\���U�RH���Z_�&u�)V����*<ibhӘ(L�)ާ�=1�$�ǫl'���� �9����l�ӟ���������~ep/xB��.��\���f�%<��F|E�����=e4�g�B���('(�2��+�F{CF6�U:��LJ�ʘU�b-Ƀ1+���	����l{7��d�aP�����r5�����B`�Ϧ:�������Q� /VQ�$B�X�<CJ�x�؎����:k��?n�00����d�e>��
?2�|�G5V>��)		�I�}i�U�^]<&X��ħ�,%i�yA	�!!�����ʁ�*.��.4�i�$R�9���t�5F�`��ŌOT�4HJ�fQ��0��}���陈\���wr �$�3$Ճ�Mڿ�3��'�9T�0F&k}V�fo9�k`�yc[�i��j�"�*sج�Zk� ���'�X#;�q�{�h���3���A�<í���s��`�)Յ^��F�0P`�D����tA+;_����ޤ���?���0h�����q�sO�gFa�Zni�+�O�h���H�����Y�r�ï�.� g���7�ΦwRcg��\"��I�N�[�إj�;�#�)<!���Dea^Yee����eư�^����������Ӭ�iu.��͆�tG��*�V���K��d�匐ܒ{L�@��|>����Y�!�ȉ�R��Lݶ?f�؅s�ՒW;��%\�h��kѻ;�_m�n58 �X�O���t�Z�!����K�m����$�����'$�bX��Y����5^A8o�(�/�$z*�ҭd���:i�f-�E�����R@�Y�(I�Ő��o|v��<�J�4B A��oC �E[��bȘ7��:Q�p-M�{FK0i&�H���'����ک��<,=�uurK�#��rw0�`��[�ߧV� ,�����d�*���@u�3�.�`E���c_x8�a���hS�Jq���r�8��@e|B�m�1z�h_�Pv�h�؟��, �d�	���z�ۀ�*���;+��4����%� ������"���J�ِK�>�}�3���U������|�r�ߓ�(ݟƂ_U!���Xw���!vm 2i��w�zD^nO:Nv|�]K�l#�X�����}���sW9y�����̋�����[��%�j�.dku�^�G�9bl�/��p����:����t흔� �P�*���;]� `�pҨ��l�y�P�Tu�[ՋX�"���W��Y�~�K�^a��4�����������8	0�g�觝b��m'@2�7t���������?�[U��r%�����(� ��Q�6Ѵ��l���zn�R�:��?��f,Ƣ�'ҋ �]����3r�̴��� L���Iͯ�Mn���(�+U�I��e^[K&�`��.�բ?���]�xE���3�Q!�8�B�fn�ME����#M1Y�BR/��/`�'���?a���Q���B���B_`�6i���N56���R����Ѐ��<����pm�*-�cO\�H�>��i��3��bS�d�'�v���i�2@�W�:�E������@��1~���<�a�\:��!�w���S&��GG�f���~q9��0��̾����Q���J�����������^s��p�=� ��yȫ*%5��⬬��!����0w�Vi��ط{&F~Ñ�sO�=n�8'e��O�N ���1��D i|��"�i��M"�E��w�z|�Q�\^H����)��_<f��kJ��8���ӛ���q��Qox�Jw��	̻:?���*��M�^�㆛R�FjZ���m�͜.����|�8|Nf��G7}I��8�YV����*��Ec�UY��~Ƌ��a9�1L�ɨ[�<���4�߾���Z�}��tC�c�X#[jk}�C�Π����5?[�+���fQ���:�����5$�EKC
YE�:&l�s������^�I=�Z�Ĺ4|u���
��@t���[u�l3p��S����h�$)�u�h�2~�;�������M�mn)�T5��Ô$G�J.��wCГa��̢/��-^�=�}��71؀������{��h���6���d��������A�J�O���}jx�X��Ы�d}��&�2|>�i���滀i�KF/�tI=~���X����P<��z܎�i�8@�f��ݮ�4�eN�5�xŎ�r4r�5>��;	�bÊ/ȕ�u�L��[{	��=k��K�}~m��F\��п
�ɱ��1g�f`[��N�����zI�6�_ǣ���c�>Čq��1��hK-�X���&'��pdGe�e-k�qU�d�aq_��֋�3��|��Q�}��|�����M�������*���lQW��]�I��vf�ɺ��MY�?�Y��3[,�hP|�V.i��`a��O��,b�~����
��ڗ��F;�N4���b
(�n^�[&g�w[�@6���\-r�
5�JC2&~�X��t���4j_J�[����?o�sc��Sc�u�Հ�Eˋ�\�%���ʨ��-I���%��AXV��1��c�b�Y�9�ST�\ͳ����/ID��IAgz����rb �³o�R�eU�l� ]�� H��d|?I�g�����{c�_\-m�s~'��JY��<��N���7k��jo��~������
SZr����ME~��_�s��j~��٢{�G"�	��z]`�8��_:�`�y...�5����K��y�omY�3�H(R�D������ss_KH�*�~1#11�{�<�k���O���7@R�X���R�6>b!�b=�k��m��Y<::�Ŋ@W���7hr�$E���'���eь*�(�])bK�P�5��!�z��\�O�z�*�4o�e��G�)~����$�S�d&-i2:�%cg���kԷI�(�E��}��(é���������V��s��T�-�4G�=�-�߸lH�I��V��|�=CpSh$�ǁae߫'���o�3!��X0-�~.���aJTz��6���	,D�dX�2ۋ�d��z�F��n�1�x�;Y��C��U�5{X� �z�_����drnN��]n�흦�����dU��M��A�ָ將�4d�Z��;�����T��Uw<9Z�β��K�:�W�r��rTQg�@��L8j�{����Uu����=����Fŝ�������JɫK��'E�B^~\���>>�37�&n�ښ��ʁ!E�-��:&t��d!J u�
�]�%_&8}�J{���Jg���im;�n�ۭ��~��/��Z��	��iΑ'f���a=A+~�� ��բ셤A�x�ȥ{��K�7sE���a=)� >
����t�ɳ�Θ-h��BAC ]�J�y�h�]5��ٸrSD6r��p��[�頹���C3SK��x��~./�'a���}�1E�"-
���S��C��}�LY=~��'�F�)�O�#5�{s>�L�OxW4��P��P�y�+�(�^���o���D�1�:y�,����(�2���@�@P�*��v�#�,��T/�;)٭ �𻥷�=���%éq5ot,�%ӥ���+���B��m	T�ư��
��2���4YE���B��'F�w����Mhnn�#M���W�/�G��<���$�6���ީ�
��/v:���ܲ�[�����|���x��3_�)h1:ᒡn/A�y\��ð��D	^��6`Q`� ��)�Ʃ�v��M�j�ߗ9s���}��L�s�:h�1����x+��{�������<�Zѵ���u� �Ёyh1�eoG��th�mGڃ�R�OIYt�Ȉ�)z��oy��c��0��鮥�W�D�E�,{+�wl��\��|�$�~Ad�&��~�Lд�����N��)d����gd��Zʲ��$F��T+	%A~ײ5W��m���1��vR-�r�^_|���9���NU�(,���~���˩�J�2�L�����-p��=??�W^QT�����}7�ɞ�#1�2�t�[������"����sl����'�$�ɛWS�煚���Z����� {��
"0���р*�\Q?SD�2���+s��ls�րz���tP/Pk�DA�"�o _ё��!e�@��_㓠j�6�*�l��s�Z���O\9��a�D�M��?/m�3k�����,!^7ޙg�ۆe�y@���zE���e�OD8n�%�o�6�`jk(�v�r	�_���5�%Ãy�#;��xM/2@�O��X���fSOx:T�O��������z��a��̖��K����R P%AB���������Z/R�Nq<xL��P�$����k��2�q�a�S5�$��n(�軎��R �i��dvT
͛O`fEGǅ� �I�5��ɥJ�>;��e�K�"�ެ'�fl2\V5T�v�PD/^�X���'��쐌
��/���M�/�nG/`���}:)��:�Ӂ2Wf��L�1�TM��?N�~�M�3����5���B����l�[��Q5-?:X^a��UZ�4s�c<:禿!eP�I�O1ҼɷX�#�r���OJ�����5�2~G0�i�N|?��T	��0���\f^��I9���@	_��Il��wG���� �$�I~�i�9����W�*G�a�#�	�ޓ�����??D�w~>Yz�܉X{��^�d���i�D�oz}Z�A�bN*�]w��y�����5�Ny�N��N�a�o��|��(N���a�<�%��D���a	�����I7-F�_��K�ԋ��r>�~�?��q������y��j�a	�ZIR��'?���D�0T�L\��Ϻ%�/�B��>`~~�����y"��9�3�6.L�	6��K��KP5Gm^o\�V�vtC�s`�k�n���d��E-�ś��!�W�}�i"�͂�+"M:Zno(9$��~_���UM|v�Fnfn�t�������T���:u'ϙ$��-�M�z$�L�H hs1�?��3�Ql�+t���Wd�z�+�������?�g8u�?�pK������[k8���}@�g�	4"��� ��c
e���h�����X�ÃK������Q�Cd}��o�gT�n�ěZ�?�i/=`�@���7��N�i����J����5��a
�=�lT�|�?�p2# ��ί�?}���ݔ?Ias��q�w*�3�/;S�V���m�#�L]��	 x��<�f� ��y��g���]}������T$7>�a,���G��f�5�P;��5(�h��v1�5Vr�	�KO�j�J��N�1{a4����ד��]ut=��IP�KP���Qe%��@/�ChI,��et�\�B�����������5h�I���C�98�-fl��''&<3�ŢZ'�ߜl@$�yM��y�^��~�T����^�� &��o�F��h?�U2����;qV�_�
��ɧd �UB?��v���E�4��ld��;���X��[�+iƿE?��*ВG�8�̞"�&I{F�Ն#�A�y�\kL�'��^�޳�~L2�W��b"��?�G���k��:T�~���#V��L��t�+�V��~V���wv����T�*~r��15B7�s��4"~]��ES���Sw��9/;�%��ٔ0Р#��W��*���T��3:����n�|[���|����o���Q���!<�<�/����M�o�3qiשVi��\���^�E[
��f�/�G6�-�|���Ր�Ig��c�I��v�x�����cߜ�ƚ>��HS᷒;���w
�'�`-(0�P.��4L�e�&�y��5T�=L�����t5���tt�*���?
�8Ė���C���צ0i�Q�PĦ$6<�%�t˧������*f�GҚ�L�����7�E3��FS;��&>�9��u�S(^z�r��l�`���]�2�x�^'xߊ
W3l�������x͞@�=�_�Ϫ���+	�5����Q	Ͽ�vN_�HM�~3	p#a�T�z�3�8o�P�5s�4Q���o��ͤ�%�0�l��u��R)F/��<����:��޼��W���ֺy�6n��*���P������c$���}M�l�����7Cb��µ�"<����!�p�b�\f.J��JCS��'6�G�_vs�\D��r��T�$��x�4���-��V�6���6����˿vU]����uu;`9P_����Iv�f5��Sc����K���� ��m#Ğ�B�X�z޿�gF���@���t��q�����o�C,� ,�e��j�ՙY���?�oiI�n���'&��f�������L7�>"W�j6_Ժ������|H�i������� c��FWCBOgWS�0x�t�߹&����n��l	-Y��U��+Zc�֟�Nx�qKL�zI�ۯ��b4U�S�\�p/�g�H�_�*#���\Mk�����\���w�A�	�������e��#�.����2��W��t`�M����^kͯ��t0a���
l_+M>�b���d$����|�!���X�W�,��>Az�>Q-ЇڮA�m�7;��x6��W"B��
)��
�F���F�C��@#�t��3rO�.��},��B���J��b}%�-u��d��o"=�e(�*��?�Y���Ѓy�%!��l�TQ��6ja\� ��7g@�X	�凄�b��2��#q�΢��ƿ��u�t��	�Kj�#�)�Ryj��mU!�c�ԙe�Dį�XZ[�5�#{���B�a�<�:R�H�I|ɼ���_��N�*���ה3�K h�BY�V�΍I3P�ERE��ӥSЀ#��{q?��f��MQX�
~ p��~j��'���	�D8�	V�8���BcO�����@ f�'��#��*"��;�i_�G,+Hp��Rr�q_��~��b|v�1�oG���=JF���H��*���n
��o�xw��J
ϔ@K�P�=�땕����bP@���΁�qυgl̑�t`HH	N�i_##��OW�h�F�
���ʉܻ���Y�Ho�'�_����@�ӬN�:�֯�N���-m6Ɋ7��;_��Zv)�*�'b+�dHʤq�%1�Q^��
ʝ�+{z��m�s��5r���Z�T5����aX�%�+ɖ�����U��#�;A-SE�H����p�v����HU��Κ�f�i�h��y���}�R���:�?�8�������d��iL�k�����s�G��ZJ����PW�~�����q�pr�RZ�������Y�Դy&�4�+�����Y�Z�0í��k��;�,8�X٫���!�2����5�d�$�Q��J�E��(FK(����~��麖G�,QE?�0V�[ �zp�12M��j�>���̪\�^w9Թ�1
��'G��[km��͜P&rf�<n����a��\G���=�ދp�����s��7�^�<�/�b0�`��o�Μ�=�c�g�`xr�󰲞���y��p����f�h p�f��|�3zM�pf܋�d0����j⦂/���D��كy
-{�&_���!*��[���aK���	�6~q�=��m_����(��u��qsf��5x�r8NP�����g�1-MB��>���m�`>��@���}~����[ Y������oV�b;i�r�� �OlĖq�RI��Y�Ĕ��L7ѯ��Y�j��Xo�=�Yq�����O�÷y���V7f��Z����@14ip�G�d�`����4ߊ��s�)O�2x[u�&���EY�B8��˅�˟�7P��z����eϵ	���P�ǎ�c�a��z8Hy�KZ�M��j=�W	�A^�@S�B	�Al �V(|�E�[Q�H��/A��\���Q�&�4��kOd�ژ�X�{�`��TC�fޓpI�P~Ա�8Yl�7�����)����Yhknc{ѻ
���2���0�F��~d�$-E'e3���eўEVNơ~�bg|������ۑ��+�l��^��2�W�9���=�+)t�^��>�{����ЂUa����7���
\@�;C-ut[��t\10�ӸjrdD����;��Xb��&�SK��e��\ףo�F[�eDM[]�	ge�/��(��pp��`e��'W(���?����e�:tW�W�r{�3Ɍ��	ܲ����XS<)���w�L��8WaKP�'" gzi����ÎϚ�[3�1�#,��ac(N#�1K��uK4uب��5���u��9{X���N�����'�*�Z�F�r+��\g~�:��堄'�.�$]��E�U���RF��3��{�a�:Z���V��{6zZ�2H��W���d��\]�2��ʀ����'M��g�
{�� "s�!O���V:�sn���'J��*i�.O@�3 ���u�+~]�om�i�h�쇬�f�~e��>�bz��y�[-�ܲ��H��6p�#��<d���F�qS �a&�7*�f_*S�xcp���>[f�?�}��ZK�{d����w�s�&���c�7�M��-l��K���-9\s����vuhk��D�а2��Ci5��q+��Qymu��/��*u�h���dz��8.�RPd�]/|#���,�<ÅQ�,䝐w��'�74������#W3��}?,8�u�~cTq=�W.q|d���v�+���n�T@^+`�Lm@�(�y�?xڏN��剄`�X%C��`�*��.~a�.�M�Y��EI"j_a���j��j�Z���j�yO���w�.��7=ZR�C��_�o#�ur��h�Ħ5"�w��,�\�� y O*+�[��A���E���,�C�(.���߅L�[8^�d�9�ْp��+�y�+	
�|m&�E[37�WJ;
����j���i��=#����Q�t��T�Z���0*am�Z-��Gȸ�߳�nL�wR�����J~�	��������ݙ�1��0�~��F����8���ȮS�Ȍ>b�L(����s�����mW�U���Ĉ�^�Гov-��ӵ��䥛�?"8m��������y�Q��"��;��#<Jϱ4��|3~�rm�����cM�H�d�
�:�Rak��ׄB���跣�����G�}iAT�Wx��+G�?�\P�0�����|���6���L9��2\���ɻ�K֗�,�I��;S6�;�kz��(bMrTҟ�.Bj�(���%���*�e�_�8x�༼JQ������`7��~ZH�d;�)�����v� ?�vy�HDyT���eQ��=!ߘ�c�)�ok�Y+�d�Xk�n�P+�]�d�w�����RG��n~B�y|̛Y�����.�7����Z���`/��F^^��@<gR[Pm@�g��tZE��(��<M���-slL����(? �.�^���7��C�C1b�y�͛�Z������`
Ɏ]�^M�u���;j�S{�n~���B��W�o���?�j�Ӡ�O�soqGe7R�r��3S[@��iKִ�w�f��|Q��V��X? ��.��Nv�Jmi�̺�*���L���V�T�������@��Dة�����eF�3���
r��<!g"�A^Ĳrn�fs$�W�v����]�c�as�Xُ�?��9�����Ͻ�� `!�Y��Gk/r�=|�Io�X%�u*/��ۊN;ת�v�[o�GW����*Ͽ����97����4���x9t���M'�?�ŕ���� ��9�oT)L�=V�]К�2+�f��r��Hp��f-f�����4��;�E����d�L�mo��>�u$���]������@s�v�G��U��9��K\m�m"b)�p����]�S���r~��}\��S�l���\21n�ѩ�W#��O4���˅r�]���袶���$g�{_�{��ұ��c�	�|N<�{6)���R($���y����`e�3>F�^~�P���O�7��:��
`������*9� 6D=� /'��{��`o�J�zh^��|עb��PW��b׽(7�u\�-CwE�f������E���o����-9�l��f���`=��x���X��M���`�i&7�P����v����l��WPh?7p<�ǹl�6�A�\7|���,"'�z��o3$�%�4�39�����V[ �%���pj���?�Ogy�E��!�=E�sL�P�4��Dn�'[��cx�Z|f��t��w ���Y�3�r+q�1B�t/!F�)��	�	+�k������e����L�aS!�ޏ�v[h���H�7�S�� ��������̦Xh�D��@���V��VpE�iV�[���W���p������Wt��^��_������x�݅?x�_�4��~�f�Z/@�#Ͼ�z� �%=ռC�33��MO7��)dk��Y
;ٌ��+��듳[�#�}�����z�$�cr���2J>ڦY��gV�0쀄A{�ZF�"%�6pM�ꒁ�`��mb�zY���ɔ�Yd3�D�N԰ ����	A���,�	�O�Z��*��*5�Y,3ʿ������zO狞N����	���y��	���ggglll{{{�׸�hL�&x�'��fڙG�f�xP@�!�[W��R"����$���أSZ�Ft�ԍ�5��	�S�j�k>y����������؈Ft|�,���$�F�d�Z3�Q��7���3*(@9��) ;s���I>50M$z�p��6��p��E|��h�A��Qw�Ba�w�&F*�e5R��6��:C��a��|�^>�&> �ؒy��v�'}�$DT��2��, F�l���M�N�B��Zw�o��:�g5����4"�V�ﳲQ�ډ-�C[�6�z���:S���t���F�SZ|���U�a�a��=�序��v��niH��a�C�ȳ�Tq�[N�$�v���nvm�ڴ|38�$#���Cl�
-�. w{���G.w��p7�a�*�N/:ˤ���C�zW���A�I���A�κ��@9�Tz�ѱRɞS՞U���I���b
���xΪ��ˇB�oޟ�Ҧ2�������f�MЖ�R��]�}�(�����jt�wD�ŨS$��]�"�ą��<�_�~�H�B��j��x�*����i`	rb/�r�ŋt3|�mm�[!�#��=��_�1<�m�0x� �Q��罻��G�B�`��'5s���"�c�Q���Ϻ�fS¯��#p�L�l^kl�m�h����������W��]k�
n��H�L������(���M��$7��!�~����zs�� �fb�Q;W۵T�5f��aۉ��)�_�Ү�c9=�q���28�	u�*�d)��#z� �� �0��]j����[H��V�֋|+�鴊	���Ԙ��0ޣCȟ�b?G_PL���9<�6����?B!m�M�����l��K���ܠu�T*�z�=:�a����FOY+A<:����_���dg8�Sb`{Nw�	/��Y~�R�6�!.
ۯ*����I�#/ڪ�ŭ6�A�����d?��Py�{ŀ}fL���G�W	��v�T��jnr!�Jx3�K%Ef�WO�}s �EF�u4!�T@bS��9ݗK�TK��Ӷ_��T�nc��g���xI�aq�űs��@|�8%)�W`S!���0p�,���������M����c^MP���U�i�9[�Ks2mФfhK_-2��.���6�C���J�}@�$�reAu�OB
��fsR������uF���gc�� .�L]e������7_��ï��Ð���f���+���q���5Eǃ���.�a%����ׇ^�u�83�1��s�%& ###�A�\AR ���Y���s��2�c�kw���Zق቉���7��2z�OvL���C���{(�}T@���YU&�m���E�p�7@f&���cB�'-_Aq�7��'�HT�b��ou��l��v��]�g
�e�����&��Ge����Bh��M#xl�QDO�/K�i�I�.i�\g��{ݟ����|Xc#�4PXM���"���Сwu��	�T�� O��	��"WN����D(�?�JA�9�0Bh����}�<g�"��z��_�y��D���"��4�Y7<S3� �s���ϡ �=�ش��0���I^����(�F�sm[D{����-�/�,��c���韸vT��ϳ����C��(ڈ;�km���Rc�cu�N����c������~����=�m�gP�Un�;G���H2&~��E�<��u���B��r����;¹'G��X:�\��t}�Ͳ|�"�^�B�Ѡ0�S��f��f��BG��m�ۿ�w#�M�W��-]jB:>�hX­���R�h��_y�y�S��_o���ҽt.!J���% ]� ���tJ� %"))��tH�.ݹ�t,"]g�>�s�y��9�0�0;�|>��u�����}��y�U�D��ҭ���l�U�Ԯ�.�e�7���±݈�M��	�W�1��5���/�U���P�~bO`-C��B�W���x �y�����t����#h*��K�2J"�g��;�^z�U�#�����k��j6n<����pn�8u*w��}�t��_�~��|)s!�+Ǳ�IEs3���eO������6q�@��*1s/ם)����!ô�
���LEp�t��[tp���D*bT�셪Jmt�����(=�gs~����:2�L�`���3ñ�4��<���<�SXH���ǰ�vsh3��d�چG���;
�DI������?��z���( =�z^��Er�<N��_?��]�wP�]$�:%0�Z����l?�<��(b0��L,����?�}'�{�,��Mre-t��j�sxfl\����"X�ҭd�T��jm�9%s��H���	A$x��q��Ώ�gD�!U�BР��dXx�z�&�xF�Bc�H����ӧ�l�h����qg��Gw���� d����oq�^�	"�=B16�e�7��4j[,�7ɓ^Oԧf�x�$�L��y�/HQY���neç�������f�j���}�xZ�����^��戶�J3s��{5]{5�ύ�3/�l�Eu���$q�}RO�p�tb�)�\+G]F}�Vy�R��˞�n�'O�/���hSU9�Wq=��2ޔ�@ꌍ��!z0����+��{If����s?��OQ�m�y�
����4�F��C3�!����B��E��O:�?��us��t]عd'�O7�������[v�#*0�ܓk�ye�|ۺ�̃q�_��^h�9$�8|u�Ҳ(��JQ���#�y���j��Z���[gw+K��w��V��
�63$bԚ�)�4$R�x��p��◢o؁%��u���_[Q���T��x���4��t�� [\�O!�x�~чږ�<�3vr�â
��,:�G��'~�����a���u垉T�P��.ΰ��`�~)���\nؼ��t�|���N�fHf��eD�ֺո^��u��ǧ��z�4:[I��m�;��7x����\��1��X��a��������51��Rz۔8�\����1S�	��������	�z�(B���"��~�Z�~pT'����(�e���/��N�ǣ�����'%�7?-�}��_���I)L5=����@WY��x�Bl*����̾�z�Q�m�ě*�t�
�G˺v��s�~��IE0;)(�6��*_j�VU3*���%����M �b(��]���^g��_��G����'�Hk�j)Eǧ�g`��&ٙ 
3�
���mrPx2�3��8k���},{����(���'�����Vܩ4t���Ǆ�_{d7�/��4�nYrҩyx�t�����_�JP��� ��l��5r&w��~�[)�!��y��Sΰ�dܗshi^��W~���-9lP��w}q
�tċ�.>h�hw�!��ڲB�I�Q3v��.P\����"�Q�N�ư�W�1Y[b��uI�7�so�/���5ί�3R��=|9V�����5}��k�����漸�>*y�=�|j,��v�<qU��s��g�����Xk����³|�)ڢj���R�z�X���1��ވ�o�d1��c#�|K���q��P<b�� ^Ľ�jő����?��-����c�m|V>4��N*��(r�7���e�Y�=�]g�|�Iy]Bu�H�?2�^� �,�'���$�
;i2� y�� fi7 ET���X����/��B�3��U�E|���P�i�A(=������Z�C�����º@j���8�*�I�g`�R᧎=V�/�_�w<nk�+e�k*c�-F��V$ԅ���at��0�4P_t�'�+H�4Z��v�S��'AG�����
I�j���OT���)�����0xF�z�T-HQ-���M�6�.I�/mК�ڈ+��J��%1��k�"-���	{�r<-�$��?=�%9tv����򲩧'R�,GVX�PW��=I��h��+ݬ�!�U�W �{s�A��;���e�����,e�bςE���vQ��8�������c�ę�*(A����G���3�;LP����<4��)l8\4׆�a�%��5M�[eĪe�p��~��eN�>C����8�c�����)��M���:a�oY����a%J��Ē�$3"�������e�� U���큷n�­5m<��������!���n'!��?iL����c��k�.U��=]�� ���ȕ���3�k�PW����~�H��A�5��pO��.�vNҬ���ί��}b��(�������S�G��L�IJvBCi��=cZ�^���O�w���Ҳ���֕���(�"��{�^���v�y�hr�A�4�������^�&�+D<���'�5����Sm��P����i����]VL����3ҭ��[^�k�ؚ,;����Li�le"1ڵ�����r�"��T��� �<E/a�9��0�Hϟ�TS��q��a�2�<x�L�kyK]ݥ;�� �H��%���$�ʯ"������/�u �ay�Ėf}�����"�<�%���r,�	\�&2���J6"�hz8X�� C���4��҄t��\����nd�K��t��� �Mh�7(�=�D'�|���ט쇓�[�)F�o̥�uR�k�r�R-��-P�4���X��o�o���[D���6K���s�I^B��H`���`��R�1�L�:���f�<����'e}Gh�����2f�g�I���ݓђ���M�@<���jҦ�ޝ�Yނ*�yҍ���a��	Yƒ����O�7��t��Ǵ�"	�+M���LX-i!��UltS֯`���L�/q؛V��/<ȱÂ��c0	�8["#Z�r�,���4>^�.�:��!�9 v�Kl�o�B_ԙ�Ϧ[���x�T���F.���I�P	��������E{ =f�����-���p/c�~ԢO!fԈiNs<�$�*΍����7j�9���1��;�7������Py\܄�*D�����j���U�x�����՚�˓]I�-(�p���H�Ě-��mŊ��8�*!)����1y���ߗ���}Y2j�)�Y�)b�����[Z�_B�}�T��`�{}�,_��l:jr�4�\|�e�Wۉ_c�hc��0�4��_2_����O-5K߃�R)���F2��l"Ta���7W�����B"ܝ��ܧ)Bu�1���G/�9��������i��NKNNNKK��%;��&]Ǽ�;/��9���oN���4C��0~0p���4"\JA�ү[{±��D�B^�ޗ�4?N�T�u�	�E��c;��b]GA�V|��. �����k"}�vc�yn;w=쫟�����k]@�<�MC�3~��ahT����닐W�X��
�"�a.��?��E��5 �:�ܪ��=R�$�.�h:�|��_ҕ�Q��#NF!(6�2��Q6���p��ϋ9��i�8.��,�,�5�s�"���x��Bt�c��{*`�i&���0Kξo������U���2�O>?2�x�)���O�����+�0���&3g����M8���8��3�h�	
,�Z�0u�qi��k3vs�����ob���H�EE-�"R	~�m0|b��Po�<F�Im���&�w��#>M��M�.�����$���ͷ��C��\Y�F[Zl�:��/��;��@��nGd�ooIWG�Fż��:6[}�o����Ę�F��h��|v{��\�������k�����&-����y��{�p)��mo׮s�m(\i�F��G��x�.��c��FE�Yɋ�
�a��6�<z�z����s���-��c������kD�Ф�R��U��.��q�%�|B�;�R@h2vI�0����:����@GR ����
�Þ&�eV��sG�4���L]�QgA4cT��ұ~cG�NP�s�~�ְQ�Jڀ�@iߏ9���k��x�$���B���g��wau����ݑ�f��m�_��^9�~sY���qqbw#7K��H	�ٕ��&Icˉꆅ�E}�B�ີO�A.��9�?����ۥ�{�3�'�)��b$�^�w��N=7�A��Jr���Ϭ�E�Η�~�"^�aAи��5�OS���m�Խ��Q��'��at��n�ϭH�b�?6瞹E��E�F�k���V;�'�n�QK�QU����a�E�b�q�g`�"8ۿ�`<7:X�U��\,t���WG�pM.�A�v���ka�"<�<GBV����u�V] �W0d�f�f/�h"T�O������l `�� �VS��"�	�K��T�xDMdhF�*��*W�Lb�%V�'U�|��愰%G�g�8�8���L��7i�5�5M�Rs�%>������T�	/��X��1wk6�jPi{ǃ�e�ɖ��4���s��sO�p��tj�s��r�p�*u+G(�]�\����f�� R����/s>��n�|��M)��	AQq�w��m��t0�Z��LB��C>)�Cԕ��C�c�#������`'AtHA�]�3(f��ߘ~5�[���4�с�k�pi��������*wuo�$�71���A7���l֎��d�x�m�ZӁ��'��
H\^�/�P���s�7@M�W5}��'�K_��m|b��X��A>���"V���'�.G՗����z��o��[�aZ�âB1Y?����ȼ2�h���@>�x�Q�/]����"pK���:����Mà�0N̰��	�<_�"cx?X������si����Ԭ� �Y4Zە}����8���V|��8U���ai1�?���{X�~�<v��q-��MR|AK�`��?<�K�EZ`��M��˰������"�g�|IZ�@Bz�.�V!dYZ��w����ٮ��l(q���8�[.P��^�v�
=��p�o���߯��C*����dzj��#�3��E�+��M�i����s��5qT[�6�^��HJ @�F��,T�%c҉�{5+Y��;�E����DM�^U�@��7X~	Z��-J�D��ؾwA�K���8�0�(uMq(�������C1x-z�$��y%��������f*Y7���jϓ4�%������$=�������hP
�6޶S4��#ϡLzjɉ���QA���ڳ��E^-��0���o���2�y�@�N ��K$����~\.~P��n>;����i���A�ױy�c�Nq��f�f$��8�+Lat#$@M�^M��2V�a?i��9�rd,1R:���h,UQ�Qr��@5��'=���H�Q�+��.�'C}$O�F��S�j�{��Q�4$E�Јw��_UK+2����z�P�f��'!��E������ϟ?���e~�Pա���3кy��^�xO�f��d;rJ��!_�S��C�8��}$+~�l�R�%<������xw�J.�	�sJm!)�(D�iT�-��� :�>բ��|c�o�-2��c?�Y����x� �
"��,f��{�,=*@�ޥ����e��tX,�&�$q]L�e�W�tq�f�����į����3W��=�҅D��~ˤ?�o�I��Ii[ή�(X�Y����%�z�!��25,�l;�P�����$��|.;x��A�4���ե]�0�T���Tӕc�����`|������Vӧ!�C��
>.��]@ρ�|�Η��o�Mwe=Χe`Y���(^#g*AR�N�7A�F���_yڶ��׏v8,�㈍#ڔ�=����δu�y�����������N����zz�q*`�f@8�j��'�*�b��#т�v�e���kh��%ZQ!�s}�>��,Uܒ��?ɚ����yaY��?ϖe3:ت3���8�,��˱��y��)Bu�������v�����6��/����R�������AP,j(�|0�MByFz'h��`5I��mm�'��e`L^Ң���Y�b,�v�S+?	����)]�kMY^x�X/۷k+��7�S����P�:�]��	r�"�C����2O�)%�7,F�A^s$����3��N��g�?��d�Vm�z\\���YF|��Y{yY����rU}|hU�8!!��}�ӆ�?λ���E�g�m�$�q��'��R��Ri�*I+x�a�WZ��W�5/�?��q����,��v	(��9�,�@��A��2�gé��H5!���2�5�/�c��u�#�j��Nn�>�-Bʕ+�U���ԭ�����J��ʮfk�Ə��C�tϟu�~�#�:��bN"�ʠ���c 2������m�P���wZ����a&Ɏ)�J^�	�t�p�8	�͘�n��x̀�S_U��{0m����a/���/����ݚ��Z+�ej1�
�^�V(˨!4��Kx�-B��l�0vN)@�J$޾5d��@�$�������N�/�*�$B7��(W�2q�П7��N�?�C.m�>	S1�h�;��a1-��#^��߽�|��ڌ��X1 ��jj5�]h:0="�2
�~�(�"�cy{fw拈��{�A$������ce�!��6��4W���;�s�v�✞?<Ϸ�BW�~o ���/��BB���e���R&���Gb��A�3��E��* А�p�{U�+
����]���K������6 �>ma-��z���0
3f����D�2���f��u��r�p|��鞘wZ���^�v*̡�ӊ������y�>�7>~ ?��~!�mp{@p�?�m�*[�"�j���ɏ�DZ2� �|J�z˹�+�p�/��$П+�*����1�),����A��;���s"�.��D0�O�Ϝy�5�STA;�����A��wb�PC�HO���+ ��ءw�B�g&�K�#��X&^�6f������7��n��z�RX�4tF� �8~H�~G�8�`�N!U�w�b��O��@Xd�*�Sr���$�6>���������6�d�F�YO۽f��B�~8OU{$6�9k�9���T�k9���׍;�-n��vL'N-1v�rQ�K�e^�l"�|�����eeee%%%���DD���OOe���w��t�%Ok�f�f�>Vv\,�������[���zԩ-�q�3UdFp$��M�LK�HA�*X���I�]�S���=�$h��4���NX.����đ1ʻ��_����J��р����
������ħ��j��{S��E~?J��9Q�)_�������𰨑��j��E��g�e�e�8�e,�� �U1����t^��	���鶅$��_[FlVIG�Di�/�y�PP�&:Ś�]��R�j���4Z���(tH�{Z#��wR��|�=0ͷ�����W��e1�!8��aT���x���W�0�KәUv����Ƥ-ch)�G{Z�;�7��;�Z������:^��?,��:���9���Y�[֩@�ϋ��h���e�<,Z����/oo���H��Dߜh���~B0�D�j[��"��J���2k'�.K	�t�Bf$=[shb=P	:�R����]���n�������z2��A���P��ggKO��l��lN��D	�N�t$�P��AXl�DGP<C��2��W��Htײ�b��d��K+�a	%b��B&��Ε�*Y�V�Bĳ�8��8���U}���w��V�Ԇ�=�m���w����m;#]�A������H8`y=��=4�\(���m�%I�-�G��}�A�o�%����z�'Gh�<�X�{</�E5�
�b�2�v`ѐ>w2P\����٘@"Q�vO_�}q���|S\<��b����5�*�(�X>��^�����Im��u�#�ۂG7�r7�%��V�.���k;.�����o;�ɂ/ӂ/o����.�M�r��s�W{�'�ir��g��g+w��k��/r����n��ݔ����c�NQ ��Ֆ�I/d����0��Yiju��F��������SL�+V�=Q�<A�T��Tѕ�0���s��C&\H��.����B�J�Ĝ$��z��<N�~�����1T�������)�����~�Y@&��4��D���m4b��H�#~H�ͨ±�۳�.�/^P�7������ڀ<�/�4���!�oW0�_��ӿ׭A�#��zv��EkjiA	H�m6ؓ�`<|�3�q"��6�߬��5�T�v�d�.$('ҝ�	8Ǆ�3�� �D��{rS��֌ȑ?;Զ�%�^ة�����M��B4�v+ȧ��Ajn�N��x�G��	Ґo.^NB�$�NF&�(�t`�V"S8\;���
]�4�P��Z,$fΔ/V�-G��X#%փ�L�QD��53����y��5b`%���]�w�-���]�%��	���_.�|�4\+4��\���3�M1��\s*T���F?�f���\��W�g���3�5#�!�����oƆ1�cdO˜d��f�/������UM�
�qa%ALU?�-�A!�Z34�������m��*jbr�����&dt$ت��
`�[�s������C�hQF,��zoɋß�̑so$��*mL�Dc�����x��N�0�R�J4TE[׃4��!�G�-H<��h�f�u0c�}�I� *6}����7�t��z{�FrM�{�ji>�����M��vY���df��DT�p�]�tߙ�0�ˇ�E)1���u�22��ҏ�-���3�^�R<rYS���XZp��>r\xW�~j;��6��2�v:��/�s���\O���wu�ܑu��� ����^|��l�>�>G{�����1"�/�G��dO���7�O�`�{���#�[��Ì*��hԲ��]H4��U����E��y@�a�����w���??�]��������VTwlW�x2�� )M	@�i������������Z �E��~8P���̓<[g�Qt%��,����)���	fA�wR�����@,gx	�:��
5c8�S���wԧ_C75_�6��lKv�.���-ϭ�٠x��ܗc8����
����_Ɖ�1�-e���d侶M���L��BĮjE�=1�J�*�O�� �p7�?5���{�$
�AA�f��P��T063}�C��eEkw�|2(�uNJ����Vf_���U�G!����v�t������5�&����T�6�@U�|�G������YE!�7�Lk����˟��!�zU�.���9S�'+�ǇA��+���T�Lc������3�^��zC�6{�6�3&f%ͭ�陑���R|�8g�Ӷ�`[�9�a��<~�g>y>�Ǜ�q/)��ا�5�5j�yvA��Wg��0YͩqE�tCxt�fB��\�R�㭢X)�ì������i�f�{�t�Ω,Ⱥ�����UL��
B
���w�Xxn�==B������=Pp��o E�2�g�L�]@�cl�@Q�3��-���w��<��~5pyow(�ǮV��^����N�M9ɀ�����e}����6������.#�E��㦫x���R��KS?��ﺖLa�56rcB}��h��tF�[mIh\?����FW�N����LMt�E��ʕ���k]�׮]��3�b�Gr(Kܭ6RX,g�g�9��|������C^��T�w�'M+7�vA{>9����w�'�����5��>~�c�v�����;H�55Gx�d��@���5">�U���U՞?����vL�F����)g�(���N-�ggXᣬ�\���K"Sl������ᒜ�g$`EBP_fo�`�xo�_��U�ڨx*}m���l�V�]�g�H:A���Z��n7AG�d:P�XB�1NL�kӺ� ����$@]��9דּ�!bs�8�7O��rX��ZO"b�i�h*��Mg&�F�J~���݆V�2�F=�!u��Д߯ F���䏖h�?R���-�Ë՘o��h�ӳ��Y��g�[��_�?�N{��m"?c��h��˾���t��˛L��JP\�{6"h��!��B_��^i��*I�Y��]^w\l��^~tikv	|�j�d�d�#3赴T8�k���L�����)1528�0V$�u'C��#���0U�3�7v����ľ�pa����+SY�,[^Z��ZbJ�#��7:�*�p�u��o�	R!R�ҥ�P���B�b9�^8�gK>�d�^��z�'�v��'�.���4]���?�?V�ϣf�pR���||��X�2�r�9A���`�}3q��*��o>J�zz�Mj��1O\�	+$C�\3n��U�L��_���%��j�q@�u��d��1;휿Y~��l"&!m=�������X���P��VL2*X2 �0�h(�;gX��C��OSV�ػ�v8�/.��`ŏ̷�_
i*���)sŭ�7݋�e��v�ŭz��71���%�ѽ0]3��yB?�(K�La/"��7°q��G 3
W<�»���㮵G{�;� f?�ߎ����}P�)f��3��c��3H�ߊ���C�`C�����Uh����o���#��z������-��m��=�}G{ǣ���ʹo&��f[�w���-.O�nz�/']nP�v�bb"��޷�)����o
5�*�;�߽{���lii��n1=7gD.�>����s�$�k���3�	�ޣg�!�m�U[��5�?;�[N{�vΎ�V���q�6�;n���p�tZ^MkKqV�z�9�9�����B���c:�������d3��f���*�Y(qq�a�3O���],O��\K�:M�SxJ�GJ͍�iMN?j�Sė@����'�BQ)��g���_�u ڬ""x\~�^n��w"�]'Fo�ቷ%�煮t�]g�q�h�H��4�Պ��!�/6	gy���;�ӹ"��8A�7q���?��0�m�h������K����#&�q9il{ e�#Z�so�դ�`-�G|�*S���9gbp��V�"iW����>�
r�{�_��k�Ďj~5'H��h���99O��Q籛�{��+;���c��"�b|g��r[����pOXA��4�`v|鿧&��6y8�Num��j��?�׼ʉ7IpZ�E�79��^p��ց0{��p��ޝ���b)Â�rR�_X��$Z՟�}>����b�c�
��v�Ī�(jT���/6RWҍOK�l�3:�+�Q\sW�F!� �ed� �
R�⫩���ُ'�[���_������O�^����x�)�����jE�ۤ�T@��ȼ�y���L��T�z��7M;9ߓB�٧bi8��Z��"gJJ�̛s�y��YZ�Y�3��~z�9
�\��Y0��A�,�)���8�ڊ��v�~?���G�/f��}����x������M�S�c�u��{?f,����<��:�+�H����	�|K�aA3{�[�K�e�ks��X���-��V��n�F��p���������W+�hik�CL}�f;,gk�+xs����^���*�I/`0T�@��k�K�����=߼V�z%��&b~��n" 墳��ER��)�Z�4��,!�9�jl�UC&��Y��~T���3�ZZV��V�:���a��Z�.�[*��}�!���g�5]��e�ò�ߖ��:)J?o}`�ϭ��,���Z����SW�;f.p��8&��wh����.,,��ᑼ�v|L<���@>=!�xoc�b�am h���[=i�5ް�As��j�������{G�U�2OR7Q�	�eZ�,j��v���9���#���R��
�����U+;U*�U�\jj[%���zA' �goN�Ҋ#��uPY%�k�q���Jr�s���yiL"A��#�h�?$ĎvFG�U�n�(0�t���~V�NB�u���w?�BD�2J+�pE؈���g�ͱ�����C%@��k;��ū&)B~s�U�G}�� s��ae��� �3� ����#M��n�3��lIG�t`q��?-@�2��>�O���(r��E��<6;H�FZh��P������T�'B�m,���v|��s��JD�a.�� m���*H�]����zt�������`w�W�~���L�ki+*|:5|�r%cpZ�W״�E{���"� ꊱ�>�z����3��s�m3QĪ3��c��4�Ph?ˬ��b�����(�B��S0����$�H�&�wL�[�o"	���ǏF�N^=�{�&7��������7��L	�-£�X�DͺJ�a~.C�(��×�3qM"���IT��s��e�Vv=޿g&� ")L��b z�P�����F���i֋�B��z�y�o'�����Ȃ_1�yK��?U�0���N$�������@� &R.�))��bg�g�i��G����p���@���j�I�y����oG�9�w�{������23�����;�M,����
�" _ïM\�eϙޗ�hm8�;��XD�rD���s��>���{��Mk���D���<���)닌�h?l�0.@�U�q�j�bULb*�|��Zr�c*�H� 65�FP�����;�l1�R� ���i�gF��z�,�X��;�G��RHK�i�0�x��������qA�I��S�3N����~kF;!�f������i�6=�A��ӄ�c�� t?����d+B9	�n/ �$@�!�8ga�R�*��t�6އv!Ӆ��-R�S�A��\|'���63V�8C�e����h�,�V4˹�T�������4+������m�u?��1N�дG����E0&z{���ş��Հ��Iۍė+�g*���zs<����̞]d�"�+����K�Hr�P/���q}�u�*����)c�p���⿮S0mIн�m	��I�@��U+y�>����,�<�3'�	C����̼1^MЮ�f�T*�x�?M|��l2�U%-�+{l�%�Ie���5�f3�8 �zWf(9L��{���a��;$jcgY������E,�Ģ=5�,�`�C7v�R�fB�x$�����\��l�㻎'_�Y_��L��vڷb��jk�Ɲ!B2�ߔ�E�3� �I���Rp`H	G�_߱L���M��Nd.�����w�/����.�FZ��$f�rm�����/���}��O���J���pp9dt6oWi����wr�F�s�8k��a�����*L[l�}�������3�#3S=�>�� q5t�ty�.�.�5nl��k�
���RPB��oxkn���@�S��<�/�C���$��Xк&@J0�A-s#�pUG^��C�«y�V�B�"K�oJ��y��af�D��F#ўk���~��B�Z�1�t���@H�u���_4�du�S\�0t\�a|�]yL,	��Ad�%@�/�R7q*����K�8���Rߔ������Z��bI��l��#������c̙�iH��p߄�����iǿ�
��R�Cfp��k%���2�,g�t��z��;����[��=����"���᝿�^)L��/�|�����K��Ψq���C���iP�g�=�� l��*~��w�T7�!R%�ԕ	�zO�Y:^�����'�
�g�T;�`���km����{^嘺::�D��_�:�����9x���#J�*jq�9n �WҪ��l���m�V�m��Ķ��?�^>��\��@�d���Vΐ9�zwRn�X?VĬ��	=�yV�"F?̋|O197��r4��g\���n���}'|C$��쿢�ӧ����?��iN�2�m���ע� >qn��~5~�����������-�g�>���y�Dg'��{n�K#C�cb����?3�s�sD�	��Dx�c�o��x@Q��� �������gO�l�I93n���g1����S;����;�܎�C	MfL��-����х*l»�zM+dƢ�mQ��Z#V�c
^p}�ۦ�f�X��1�~�7:�z��<:A39<!jZ�^Y5ڕNhLv�kq-�7�6���7� uu�-�px�Q���:9��J����J
4
���4�~�x셺/I{�d�9�����$���凷G��q� ��J��lɡo�7Yq|�3l�P�x?h��,y�Q�M}*����XЗL�Wp*���747���M��V�GK=�R�a���G�Y#�Fz��	ˡQ��H���;�����PR-�Y�2�u��@w�8r?�0	6!��)hsy�%�`t��`	W�x�a��.����i������ٺ�a(u#���,b��N���m�K��/1"�>���0������A�+��������"����&�����|_H F�CD������t��~�8�*�SXɐ۩>�B�.=��t�R7~��5��wr	�j)�}��4�f��Ml̬2̟߀k0��
-��Vs�|	�n��mB�=�Z@_���i�M��r�}χ%>��9�Q{wr�|���|�2}T��c��f�����ԓ'Æk��}''+K:l�����̈���v�22�f�5Z�͍s+Z)
���Zr�G�h�0i�hC�+Pf�1�g�wgܲ3�zvX�'R��g� ��Z]˷��0��5ؘO�&��h2C�75G������k)�(b�T�=�P�8�lo�˖詴���e-cHbCõ��-�]�ѧ��|�n�nt����M\y������OkK�o|M�ޢ�Z���O���H���N�ެ4X�"�t©�"�hӥY�PZ�+���,�|]��}�W�L�|��?�@��c^�w���!M����J����c���ǈ�����:Z^�v�Щ𒸌�9���G�r���c�p�$�ʭHs9�}[[jڜ[O�tm#�*Y	�y���)��Q���=N��eK���Xy\�A�b�V�ܣCwJ���Bg����AwL�p��j�H��x�6�#��&��i�ի{��x��������l��Հ��o�& 5��ddUf�s�V������ȭ������&�|�?U${���V^k^Es�]fLW���C�U1�����-�S81{�@�/�;}W/cV3�#�g�@8��{V*֣���7����=Ra�c���@�!�Z��E��O�_wK��\�p��[����g���e����cĕ����������M��q��q{�����KG띯��sU��r��g����)DW�������������l__���:33s�����B��6Wummmuuu}}}]uM-�jF���2�)7�!� fr�9-=9�3:�t`������Dwj���N�,X.L�}�B��p�*<}�z��\^���MnIe�4��&B� U�@�͜c6=Eo�-�[�S;M�s�aS7�[��6�hҘK�9�l� 3��IW�~��A�$������'���F�KlG�^o�O���={��nѥ��c��Th�p~��˿d�������]j�5�ţ�B/n_�*A߹�5�G����I��&���N��@+i��Q5��|��En��A��E�Q���6oD��.6 D
��^�+�,��4�"�+�G�zH��[e_LE��?]�9|� s����^!HKr��i��/Z+�=w������E�n8�yU�����u��c�	L8V��Z������ļ��&����iX�L��I�F���� �����(�oWzV���~�����~N ��/�� q����V2bW��Ep���?�����2�Uj�)��}����2G����a��)���(^���T^AF�YnQ�����7�Ñ�<J����L��9���:m�Mښ�7>��<(L�����/�{������g��7�g���V{��mwɇewǉ�w�cf��r~[i�n>>w�}d��]�兛�ؒ�����q�+������#+�,B�?	�����J�*��NOO���Gn~pp���\QQ��>���`��x�)((��-(���)f̝����;��F���C{�U�
��ڸ��O��Z�j��j���33�0ڴF$@eP
�b
���.R|je�l@6��ڶ���!Ɂ�s��)�c(g9�p3�q(���,�r�/�� �^ʃ�q��M��n,f�ڮ�vjl�E����G]��0*� ��8;)܈���Yvt���{���Q��Vy^�HQ�w��TK����0�^�m�e_"�[^��㩒�����!	ȽX�YyK>����2�|"�X(m��}k� f����6(��{%��	v���Œ�X�|�D�S)w:�H�F�@H^A��{ԶM�P;��4=~�DX����o�OHy�W/�{��wEm��7=��׍�%ʴT���fRx��.[�b����U�7z�xy���G~�mAoSzNS�@���B �ݿ���̮·*�t'�+8	����̣��tI�\q'h�䈟� 1�=�~b��;���s�q09.���P\�2�}���z�&�7�{t��(����JʈQ2F�AiPR�  09�c#��RR"()�4���=�<����ι����l��z�����}���C�mq�u�*�A�6\��_ii��"�6V�~���^��"��P.����k���O�����Y��'�DV*���EW�����<EI�l�j.��� �@FBJoM��U~h�gAe��=�x���ɮX�#25rM�
��#X��f���m��GQr"q�Wh��8��ZH������p&j2vv�E�Y&Z�?1���<�En"*܎��AP�]=!9�����\����'#�'��]����Q(�)�a802�k"R����ez[5���[�F�����z$��l4��~b��SH��sϮf�d�y��ϹR;ZN�^1&P�#GH��@�O�Q��|SR�p  �f�lK��S!C���0�i-�R���	0���p�Il���T�BO�PO�dJh�Fr����E��D
��;T(��)��� �!��"}��h7�,ËG�r��#�,n���ʹ���������QT��E��y
�UO��u�J��0�Ϋә���UL���|�o����������R��/*w�3�P2`��a6tttL2>޾>�,6�­i���<"g�;�hV\ܾ{:o{8���2��0o8q���۳�;�o9��x�sC���!$�,�ӜA�u��5�Ҝ���ϳh.,&ߒr3�)@���d������*P���܂�۟��*���Ӊi2Ih҅�t���>r
Qp��$�	G
�h�HS�j�L?6�U�߰3�>��T�a~ux�j`�<�7�_<Y��ŦK�=���o�z��BN�q������xa�ye�;1��e��(�C�Tr��8�h6W��C"m�=N���_w �u�P�%Y!�J���iK`�:��|@mJ��[SF�ۧ9R�0���m��:�47�̓��Y#�Ћ|�3�p�j�\�X^��ѣ� SM��v���_�+O��'!!�.�����X$���6�9��*�΁��T�E��l��\
s�Vl!�X�,�80^������V\��O�c�OI:�3�ۮ�.���O����<�G}|D)`Z/#!�Q��<`��9�(I�� �m �5᧘��::\#��gZ,g��$�I-�K�@�|�ӷ��i���]�|����*���!,�f} y�Z~�-r�]N�^��]��U��믞���mS4!G�dTq	D!	=�Dn���-٬m8{�I}��� 2���WB-�������k�za&
��5���L㷅�f�C��Ȁ� `�aX�O}"��Lm�������z�{|4�U>�C�B�9E�c�X�!U{UN]+ � /}��ӟ�ܮ�o"T�ן�_8c��,�y���֮t��F�����^�M���4^3���p��!�/�`	u�aMU^������
NEbvEz�h� �l�$]�g�7�W�0��2�������"Q(J`%�[P6��}���0 ���\�&��_�F�L�H3;]�9?�����=6���z��Eţ�
�@�F��IBX��e�5o�	��r�k�M� �`����Vj�v�:�zF��i\���O���ߚ��ýsD��he��XӾX��m�ˍ/�V��7{�t��k'�0:Ga׫a7<��R����\��9QQ��*�yy����p��tZ��pf����R�X{��̔���bm� �Z�C�#x�I@�A<���Ǳ�ZZ�bI�laPv_X����� ��y�������d���~��~�C`Ao�KP�M���&��/��_��ni V	P�����TEo?�-|	���ś�@����5�$r6�p�. �@-RV���'>k�����q��0�GS�>ވ�$�/\���cd��&�$6����n�+��;E����g �ow�X*�ՅJ���q���h6��@�8�X��_�&)o9�f�'I�5�ɓPp+2�&Y��.	��՜$B\OkC�&<~c��7��]��+��`��p���2��s�,����X�ɜ�C[%��^#pT�SK�[�<J����?ָ7�?�go��}��J,��L���;��#�kj( ��-������J=o�}�Z�P�a-���/>	�Vc-��u��s4��s�I��r�KjG�ɂp��=&)\���6�����1=s,�_�/X�8w����fc�ج�˘>s��|F�h*���Cｈ�rI�i�b*���ҫ��/���`X��*��X3K&\b�((��;
�p}"Y�$��d�E�CZ�o�#TL��K�ٍDN�rߛ�I�jkII♤�9sl1��䤞-vR�D8��wg'�!���F͎�Q���}�S�tFSuF��Q�N�ֽ�X����"�Kɪ���((�I�,�N&���<iX�H�A�zI�
 y�V��I@Q�m�d�����m� E�S"�E]���B��c*/G*/G�:Gj^Zϥ���"Y�$��H�%��U����L��c���xW�����R����֑r}����:~����2��{N�y�h�������.� cC�
��?���]�`΅��Tt��S(u�S�$P���^������NO>1����. �;+���А�.�-q�nA%$�$��Z
�c"JR���?���e�U��GV��5etrN�/����&������Bu��Q��PO��9t���sA��1/>���H�r><�z�g��4
+\��\$
cui��oUR�g��4?)�rWn�cԠn�$�\K2�wAP 2qo��we�Ia�z X���[/�Sz����1v|mÐK�B��cn�(���v�±��7��4Z�|�:\�qԓ�!uf�GS����NnA�HR�<*��)�Y�osZ�Fa���>�t�R#wu
3��-��<� &�����B&9}�>�'ix�6�0\���|=y���B�N���v��+c
��1$��3��3xS�����]�n_W���?�g��
�-({�O�z���.�gS�cN*�\��J���Nu�Bz�7��S� @�fM9�;F�+����(���5���CJv����Y���L�w��`���LDp���T�r�oD��l�m�}ABs�{����_Wn�*�o3�'�/����6$�t~ �c;�9�~4�i��JSB�+W��[{��+U�Eܠ���ݻ<&�e���'0@sк̨��&xX}�e� bW���v��рrH���ʓ�8�L!���N�Y7���Ȁ^6�n?K�D~>���s��A�c-}�!:f�V3�x-�D�O/��V#���$s�?�:����r�u�v�r������5^5Gx����5F��rF+����e��������;5qD��P��3�N��6c�M�_�%�]/Oڪ��yV�j�6��b�h,}���C���Z�*A�o��CEӲ����us+F�F9�8��e[~�z�c�o����5���t��p�Ӝ_n0��sL�_����!�t��>3�y���M��lֹ�ு���j6�G��"��.��ȼn�Q��]g[����1x�-lC���R��<^@� M�iɛ��~i����_�Ӹ9C��U�P�[8N;:��1���Ipe�Lwb5B#�>j�8%<��UH7�g�"{�X���-�R�����y=�Π�7��.QK5���ˁ^|<��A�F������r���~�A�awlK�M��V�}�Y�s��y��	�i��r+�S�C���n}��s��p���e�껤ɲ����Ì�7'���v�V�J&����z	+�2G��	ѹ� P���0��$=�)w;1N'+���o�ҧ��+ :&�.�/ �;G�7�n�j��-%������B��'�3�'��]d��ˍ�\F���1�/������_�╂d�	$�\��/r���>y��^q.M1�&yzP�#߃3|�2	�t�^�o���n2�*1/�!�7`��Vm��qΛ09�{��-��7l=)
5Ң1�$3-h��8@3�mEE�I�2c��i�	��w�K:h�;�e@�.[32���C��\`��|:����ii��MLN���xMu�WY~�n����M$O�
~����B?_{��|�N�$���p!�x:���ن���e���o)�O�/|7B�Ů.,�.��®��/wm�O���w]�[�\����ﺞ�9��
�9�9]�;�jS	�����������[�nơbY0	��S��0డ�\�N�TtU�d����*�+.(���D�x�!�8�B$Ç1��ޞ�^#��&r�1��o�]]k��{�����R�����Տ��;�(p�����~��m�-� )�U�'� &��!4�Kx�7H��)�+�hÖ�Y�%a�4���A:�*&:�,����I|�y|�t�@a2��/c�%�EA�f�L��V�=�CD=���q���Ԉ� ��ܴL*Z�V+$��;5��sʟ�R��8�-jV��m�#N�[�������L�L~�?8��a˙9�����˂�L�W���<q�:�I������E�3&_}�X��	�O.O�h���/�(����\͒��s�*O���2�k!k��8�Ӧ�_\F.B��?0������*��6�1�Q ����!S�w�q �?@��"c2�5S�KP���B��p��� ̺z�w�r.R$�����j2�U5X������z�]�-����
I��+��Ц[��H�I�x>�����<��h"�p]Qu�nD~����'���ciЮ�+P����(5�fA����L7�<;��>[֧g�&��}`.�4��'����dն�����̯�`�����&8��t�n����4�hd,�MtJMk*x�H\����u��C��)�77�Ñ~�2�3*
6u=ޅyG[&ceG,�Af������g����ήǺ.�����<���a�{}=�s�˦���wI�͂��xX�vuX���7���ʤ��ޣ� �W��]3}_'D}���|��?n�K�.�JJi�Î/|[��6>0���Ic_��W"��ބz3۠a/C�a���$��d-�()��mv�}kj0:�/э�_�34ugy��f�$(lD�ɉu%�����_:j��Jxȱ׍��f^�1Ts��'N�)M�cŵ�Xr�7�wuh��v.WSNA��$��q�I�����]i1��Ϋ�Tr��O�^���RLX|ͻIvY�G�*�[�Р�_i��d��'�2�(���Ē,����%u�,��C�1|��.ߟʙ������Hdkjc+_��=�Ob"��l�&�P2P*uBm;t�|:W�-��WA��ňD9��r�Gw-�ϗ���j�N�+u
�:��Y���2�3j��R46�4���H���eFPR�]O9Wwz�+2��)1J�>R1�=�'�e(ۿ	���2��������4��y�$��i��7z��M��!C�;�<�hq�3��S��l3#Ŷh-�Ĺ���P�PMS��;d�����L#�̺����#c	�x�C����\��'�9�S(Wq4��Z����H	0J�L�q��4���X�ͭ���z�ҋ���q���NS���w$d�'�܊[� �M�SZ���*ZP�i���[���kyN��V"�-N]Z����e$�[v����$I�0}���i"����vHw4b,��Kn�@
������o�TLk2��	OĮB<����&��⫩����O�[���"���oazz��o�v�.������ṹ\���\V��պ91K��6���n�w�>��<[�d{:�0ӁB$a~��8����:�Ĵ�UfGĬ:�q""(�dc '.�l�#NhFFF�^I�|F6�t&23����m)��l��l�~��Jm��hX��Xw;៵��X�m ��ʥK�5j��R�ui�u�d�ڡ�4JGّ�.�4L�Y�:��IYkL6�7)��z��\���?�����~�k���Şm��{�Q�U3�[�V��pz+�����ҥ�⶞ϑ�
�Y��T�2�vs�{h�S�c)���L�����f
�'c?2%%�X��d�.��7�ϳǲ�IF)���ͽ�R�������Iw����o�#��{>z$��l۝��"N0h�˙��C���|o�C��^nb"'��c}�F��bʬ�"�=É�`hx��$$�4���d���4���ßn0ܕ���&72 �u��)k����Q�v�a
���P��jw�H�K6-ۯ6ƻ�b*O���Z`W��y�cQ�o\?�@b�#��2��I�]��<5SX�����&C�/�¹������hA�'w������Ђ���X���h��&�rY�L���FU^�+c�Qs�ib��/g�kH�\A�4ց&ǔ�ի��i5���LgT��ʾ�V��J�ŘMa%(��`+D��"5or����̭�����^P��v�����q�M�����*g����7(L�����{�� ��
?*
m4��k|�?���[=�x>9+�|9?$��uv�Yvפ|>�uY��]���+�;OX��&��#�}�.߉?{�+�&�=�P��������3؅/�o}���vÏ���Ź����������=�&�Q3�
�P>'53׋zN�����=]w[[WO[Wwww7wg��w�O�-W��������[�y��y@��B��J�sm'�Ϯ��cG�I���l��pn���!-I!j[�G���loz�+Ii�ѼJ=l�f�:����v�y�'��ީ�)��'�q�P.���P���I���9V|���UOXq����PY�?���D2��E@�i�dU�D������{$.���P�X��;l��H�||�
�x���o�7�OjU�F�r��L��E���=)#Q��8���d^P�J��Y`�tn��o1H�]�X�A�g�V9�Mrk_�����簃+3�
�?f*s�Z�@�lq
+��7��4'dD����U�=�zUp��Z��>�2��e���\��FBA�m���/�zp1���!:�����d�;T�d���%�w����$�9�\u�Q���=qݑDO` #�[\a�l���s)�ץ��i�M�wñ�mD{oř��j2�ܵ(Y�#$�*L��1��dt+�L�Q�y�
����b�����=�F5�F��EThʘ�H�$+�7�rqD�����!;�#0�G�T,��VL_��"�N>�4jC;M�&�$���w%%fz[���j�V��|�	#�b��W������#�]�e��M" ����D��j�rbb����XN�1�4�'9R3�x
_��)i����=�h��G���?@���E�ZiO�	~��0X���p�:�af� ������̖�>uYeH�f#,�GW��>oQ�\D���<����?ߧl
-mx|]Mbg��[k�7[�I��Y(��+)M6�[5��|�;��[����rǑA�����Buر���~W�Y�͟�c��Þ?*/�y��@���r�����l���G�?S�������P���xޗ�,�d��z�"K~a�YII~na�+e2iu{�%$;AuD���ӥ�lc��dstFN�ͳ��g[-���I��Z�b[�[������|u `L�L���1~1���E	�L�G�����ET+�¸�}�eN_�"�t�z�S� qb�.#�G ���8�|_\5m��^���]%Ȗ��ѭ׵��2�ȇ�ϚkӪ0ߤN�&����[s0Bԇb�@�L��ܷ����=�Jx��x�JEDث����:u9*��f�fӸ�z-��
���$JB[�pf�[j�ü��?o��@���x��߱:(�}IS��\iv�t����ye�D�<�.ш1�9�����ژ���Z��;�|�Icp��ق�96:ջ��1;���@J�5ri�F��/�N	ZL.����:�
�z˶�,ɿ����Z6mU+���>�{��k�������F�ZDx��i�34uҧ���s�o�7��E���]������4��^:���zT����jN����+�=�i���ӝ���2����޶��J�{�=�x8��QbԻ�)��~|�Y[2��KB/��k=l�D,Y!bM��g�]']���7kd�<�#ǳ�ؾY��CT���!7]*�1�W�?/>V7}L@�v\P���*��4�0ϳ�e�;��24����FUGN�������p����G�wgw��q1uU#�dݼ������%�yp`~�犉�,xxZ�֪\�!���z�(�m���G!c��T�"5ώ�5��HR�B�1�h7�-����[=�d |G He�6�&����IzE�p[8�$ؖ�x5-���r��2���.�'�4"!���2Q��'�Y-.�}��׃,�[�?�,Ѣ���ήyK�oD�y�S:��
cJ�w�Z�b�VF���(.m�.��d��|�� "<5Uu�����[�^�&qߒt���%h�[���d�_\D��t�����r����)�Bx�����7W�agu�7�!*7�_Rlr.N0������3�4����q%d�������k$��=�O����ʒ쨤�����$�vo P�WǞQ:)6�=���_d�  �%;М�}.���x�q�`A��Ӝ�d�6�l)�>��")ض����/F�vo gp�����wB����S�Ҁ�R?�&�7G����8��_E��
+'M�k���pVk�ֈ�\�9l1�A'z��i�*�ly���Ϊ�	��73{�Wރ@ꙏ2���!�V}�$�Х<�k�c�ݭ��� 6�}m�h�^�sr�]� O|8�J��9A��7�$H zj��kc��(��-r��Hq�9�������,�+�O�nΐ�F�5Y�Qo$� TETV��V$!�U��Y�DÆ��螽��o:���sG�zAjjT�u�^|N�6�4Z��ZH���&�%���B�9{Yk��q4C�s�v�;���G�)&�b�N���M㯱u���I��tLmjѦ:�������.��4pT�TFAF"hv	G�v�~/�看d�ɐ��&sN(�\��z�5����bL���~q��i����8)�W�A5N��� ��n|��d���H
Є��(EO�s[�GR�������\Ԡ�LW�?�∲U��G�`, ���SҠz��[ ��[�4P��W����Z=w�Tc�$2esk�â�rE�Q s�7,��97�|�\f�����˶�K�{�1~l��TI4%��^ۮ�%�Й��w@͙h��)�_����9Q٣���沠����G��F���՛�U3��)z��Hތ��|��Y���F +&�'f��ۣk�W8
�?Q��Ќ�1[o�췤��J���l��)Y��jJ�u�J��A�����g�����j�ο��X�.�������ڿ�-�H�Y�s���`X�Ź��s�s�:��]��ۍ�G�546�ڃb-�W�zq�����DDD�$�w�F
�k޴fGD��c)��}�%#OH@`
j&�J*h�+�s7F�싢�k�]����^���\)iw=�i������#c6EU�@���s��Z��ԛ��/��S����A�rь
R�e5��Y��>+��I(E��H$���${����j+���8�gS�?"_r*�p�p��M+��G��}�Uڜ�X^%�4��t<F2K�0�1	1�kE�"�~L�-,��v�H�.���b/r&-�ńt�&�HC*��)���ԃ5�$�̧¿ k�gr����o��c�GdWh�i���MG����*z���4�
�l�2�9�7�
3��*�V�
ڞ5t��R9�S9�.
I(;l|8��5ľ�V�NDC�؜/ܣ|�}Y��+�"�
��
�ХY�n��ʬ�խ����`���!z���?8���&|W*V�������i4k�&�|���T�Z=&�|���&�u5�����Ӑ�)%�����vwi]�+��W��¯�!:��B1TJ�
�� :& ��e�)8ʌ�u�0 :�� �?�]����%���wP#_IW;y����H�D&ǂ@�}i	u{�	I�)) ��$e����-��]|���bfq���ط� ��1pT�����ڄ]A{����ޓd@@��'�Jæ�^=�-r���S�Iݚ����r����?���ܿi=(I˭Q�=�(�̸��hʹ�_O:B?�����������ƒ��tSc��f�2�|*0�</$�p����'��vq��y�5:��Q���J�ړ�#E�8�O8$qI���ReTWG��(͇:��;�F�/��px�-�u��1%1�� �Ќ��5��DE����f�0J��w d?��f��&r���T��vS�s��t��D�zd���S��W�W�jNu�8�7�_�5I��-��X.���eG^���fY>��kL�1�I���b�D$l�V�����#��ʹ���L�^���*�YQϬ��O�H��n�T�o�$����Lj���
Ř��(�IZZ�z{0�ܛE��}��*�SAb]3�nr��}��ZU���}�BU-ʔa�U?=�u�אQC��QD�Jj���Ei��@�3�M�JR݊�3A�"����� ��reY����
y��.x$�G~oV�O�ͮ[���0�[�[��f�Kd�}��Z���gg�\q�7WS����B�nm�4z���20gcbE�!��k�2+��(��^np�0��,��E�������}?1C�5�K��;�����������Sְ�G���m�	_g���R%�tc�n�?:��aq
���P�_��J�&���b�l��_�PW�)����w�{SZ���Ld6�`��Hż'ϒ����z���9*՝j�igI<X_�K�P�ruM&��c$.� D�%��m�#��
�R����W�X�b�|���t���B���mLW1X��-b��BN5�<Q�W�
��0���@��J�U�N�ղ�H^����DJ�	N���a&�K�J\"j�D�"�m�,�F�M8�R�����Q��F3�$���G�4�o��������8����v�6�ŵZ��h�:�+�������<�_6tV�%u���U���̐��8Z�\OGa�j���O�z)�Љ�*�M��gqX�Ju�ܜ����0��b�����xA@�,^W��U�]U�;�;c�P5oPo�D~npC����T͡ O�e�+"�3�%_��K�G ��?�(D�N� xT���$*IY��X�R�yo�G/��PS�������^%��1���VZ�Ѓ3Tm�O�
����%��[����b���j�6n�b4wt����s�!C�EHg^0Qy�ZG+ ��~�Y���\���%���6�!�F ��+pkw�iI��b&�+��И��SG��ڐ�����%�i�S�=������������D������$c�����T/�U ��6Q	�߰��Us_��7�D�F���=��X���1Z�����������sv�y�Q��xF�.� e��Ҁ�,�Xd��ۛ��2R ����o.3�N���[������;�Q�c�Kcv��N�5W[/�A����g8Ǩj7��@¥��Ȉ ��%}�+ZM�قX.���^T�6�b��hb� ��S�z/F��@)nj���r�m�
G��e����<�c�qѯ�x�X|�wC������2=T�r{��i�,A�X�G(��m�e�+	��#�����.S3���`���W�n����SEmP��𮔣���<��Y����3<�s�\";K�r��n���-��e�$�f`�2�j'QYuR�Ű��gTycm�~FHz?�U9ʭȮ��t{%$���Z�c�!F�Ѿc�,V����b���"B"��0�Z`��S��#����z�q���jI�g����_�r}��d�wd�s�+��Ջé}����<w�O�3����ӷ4Wևږyy��9j­=�mա�m����K�Ct���m��}}����T�d�����������#�P���~Փ_�}�_���[w�����R��)n���}��m�v�X"��nG��tw.PIڞ�M�N	�"��jV?$����ݰ�b@�#�@��@��e���L�E d�bbE�������^Ϧ�s���O6��~��
T�������V��$o��`A��Ϥbt�v2�#JŽZ�¨W�#cU-	T����	ΰ[*�
��Y�-W�L�B%��'H�G�R��`��>i(|����o��V���Eu�F�� ��8�VNɴ���5����eL��5��Ԓ��U�V	�w~�� ^�?����b-ʂΓz�߂}����ic��� �XlL��5e�L��1��j���<D���� �dM��E�*<�ʟ0)���O�,�'#$��E^��j���LiJ���e�-rdzI�;�zW�2_�ƛ'�q+z�Pث�o�l��K:�F��v�f��bC���s!Q�?�L��}PV�4g����"��EV���C(�	�H�+@ض\c�lE���Xx�6��<�%�|Ň^��>pr������=<�ˠ�}�<�b���G��i���]hܞ�'Gxz@\\Ľf�}4�ֿ
����}���� ��m�W�#�Ȍl��R �Y81�܂�.ܚ�_-��,� �:�p/����^����3W_RX�m,�T�=6!io�:[S�:���+�m�36	�Ïm��M� B�َ��h�O;BM�3���^"1ug����'�<�(��Z���W��㽩&��n�.Sݤ� �ʂo#c�)���� &J��q�d�O�i������+x�G�\������w*��Gs��8�����iG)����)}��4�o:;���2??!�5�{��T[>���S}�Lٕ���Zu:��޴�-qU�����zu������ڋ�	&�)�iX1���������Ͳ�>�*���Ź���/�Al��wp�`��?Ⱥ�g�L��CzpauK����r3޹�	z��7���n�ԓ�������������s���`r9վs�K���sv�)I�d
�����C(!�ߢ�� ���MN�W��S��RҔ	
��_� ����/3:][Z���₀���Q{����Ϧ
f'(������G��^|�s�G��;�a�zi�m�g!<;J��n�G�F���c���
�qzp��LwA���������=-Ԧ�g^�2�YX�V3�Fj�����ptc_�7��ӣ)xI����Vp;��;Sg#�2�F�����X~��Ny���VS��H̬L�Od�[i.�, ����w�ӈ2hz��4n	HI 1{9	c�"����'d�r����N�WGs����Ќ�l��T�w�C����X��Ug�SX�ڲ��v.B}�Q��\���`$5�ffP�Caͤ�W�oalU�,;�-���λf�,q%�)1��e[+m�|�
I^;���ʑ'lΓ��Sne�v�y�5�������m��"n�w�/!,l+����Hv���\�nM��n��[������ZL��0߭�`rVM�у����=��i���&�5�C �{�g���"�k'˘�`����r3]5S�c��/��u]�O/�C�'���;g�����i���j���+����:O��(�����0t�i4ÉRe�ɠn�U����=���/R���#���څ_�K;��P��`������x��26�v�IHX��>MB��SsUS�|�e�`���K<CE�E�\�6�S���{��z��j�ʁp$v�ZД�yw2����6�Mx�$����u�O�3Ⱦ�
Ir:Yr���ԫfy���l�Jƞe���j�Ӧ�מ٥~!E(סg�������Y��g_Xp���xK�o�z��������i��m�>liv^������ogRQmoWR\��m�Vfїљ��؁Ql����h�ٱ��#}3���q�X�	~R'�Y���`����[C���W�;z���C�ns(]���swrr��\��P����a�����^s��&��|������#����?{Q��,��sAZ��"��R�d�
�{���$gY]��u�<�!���+o4�~T��	FAOS�!��G
��0����'����^8��}ҤVS�9-|���/.�DD���D�t�.bo�wȆڔ�D�Ѧ��XU���"�&�(FZ�RM�����߰_�qE𔰡v���¿������H��}���!4EZ\��~9������:������;��M�cFY���K�%��h�o��<���2���(|݊Mh��eA�&d�V����)�jRsP@���T�*�Ԍ$meD�"��|&����T������P��ÌqҢ(�*��i�V��%��h�#_��噤����������:�jȀ�L2�B`�Z�e�*�p�՟������]��s�]�͖�Xt��B<�ܖl\����e�6U��f�(a:ǿ�:�T)^<��9�X8��t����&0��&5�Y��lĴ\�>gr)g���ݤ��\���f��� �J?>�M4�������j�,��q}��ݕ� WW'�ZȊ-�"�E��yNn��)��h�u�ZC�I\h�? �z�&�-��Up����Vx�?*4� �|���e�b�
�
�`A3,�4�O������ʈ�Y�o9�P'����7��`�6���'�I5G�"W�J���Z>������Fn�������v`
���k��z��7lkt������_:^<� .�P�{cֻ]�i]�o;�ҥ�nIeM3IZ1�[�:������Dc�챓�1�2�ici�L�X�1U��GY������~͊AeB��"L= ^Ƥ�u��g�z������E;b9�~�����i���f��;d�P+�� ��.{0#�Uˋ�/�ٕT�$���2�t	���#T0�J�m�܄���6�@�Axy��'�YzbV:�=g����鏭�#��I*�&�
����9�޽l�>c��G���o���VYzJI�ڧ���";5��te߸�wk�n�oކ�
s�a��NOX���I��.�#ϟ��p�]�^�ue<�[��X��s]:���	!�Y'��z��؎n�Im`�ma�P��[5C��&��!��+<�����Mђ4�?k�%iy|��I"_�y�|t�����3����몌�=S5�L'-������3��Y�(iJ�lvv6vJib���]|A�G�W{��%O�l\`38Š�4�Nj���D1�D��$��.3�8���V@ <��KjQ*X�%����N�D�-�C*���Z~��A��*�.[o�/��I�-��͙���(��*�h~eP0-y�f�`�|�<{���1x���tq�t�;ؕ=Z����^�`4�����;�22�vC���L���>Mϲ��`�z��J����s�~o�"�Ҙ
0�#�[~���y9��W�;�Y9k�C%�N%���.����[�˧I�k)���'����T�+��P
D�1P�i`ܻ=Z�:я�V#칵���PE��S�*�T�R��0�z	�*z����Ã�������l��:3������da���s�z��a���%1��kA��2��rf�il��WƀK0�a���,���4�nsyɤMX�̷�(�M��3:�bΕޏ��~J��(�46�U�ƌ�f��}=�*��������q��Y�����9�F��yJ�2����FV<���&y�Y�	b��a�<hNĪ	��wx�ƨy�����Lj	��\p���H.O�:@S�V7�DY![!C��Xz*"�B]`Ҭ��٧�)r3f��-Q��s���f�sZ���~	kT��wA�F3��R"G�F���T�d�@M,2+i����z£"f>	�<jȕ}ѡ�)�I��J���O?3<2K����=����g�!��E�|�B�&��瓁�|�J��+P�}��T��Nn�䧌�W K�	6OO�bd�'���1��Þ��B�^�>˿�5qU5pW6qU4��~��R�T)[�XtG}������}WOB�� ��_)J�����ݎ�@ƩD�hݜ_/a�{&V�w]�	hs��3���ڕ3���>�K�5���8i��<�����Mf��l��%OR�3}&��q��ޠ7sw% ���!�}(��{�- ��}6r��SՌŋ�0V��<[�O����S��5��o#�5;�/OmƖ��~yt�=9��8��ڽ�(�P	u���4S	u�%/�����E�z5U�uy��������J%�.�K��Z�E���6Ŭ:\��<����C�ʖl�vE��M>I��jj���--� �[�ʚ�"j�)i"����/��v���Ų�R�M�_�U[�4[���#��$;��V�'>g~��B�dm7�՜\S�i��I�2+[�˒��`�-�^����^4�ZTŒCҌ�bdV��x����NH��Zk�����{�,7��Z�BH\�OKi�&���}~	F;=��w�'W`
E�i�D�?A�:���!v�s�7W���
98po��ve�LZ Z�$��Nu2�g.`���x��lq�����,Db����L� �x��ٲ�+Z̞�S9%97���}w���QYܰ�Ȱ���̷i)�,�kj?=�I4'�'�dw�)���,1y2�W{NK9��w��8M���eO���Z����ы�{(f��0�g��<��0��L4)�RW�]7�ુ���u2����{B��W�VMk@��<�������j�{�5�V�`Z(�][�H��[��`�ݭx)ł�݂����K/���{&���K2g�Y�Yg���=�i�Q��_a�X5o�j˿zT(�rD{p*��\�)�U����^���\�\�Әz:�:��-e�/��O���5�������*���g���n����*���oQ�ʳ��3�����Ӡc��8ؑV��[�}1�$
@���纑yH��|���i�`fB�_��;�#֋_H'��2~ Cx!9�A �u��.�((���0[+7" ?��a�g��GI�w���0?n5������@,�r�T���AS�e-��ɧ)��������W��
����v��þ����^�+��ܔQ�W�h�].GX��$�ed�S�ԥ�5$ե��#jBP��!�Dg�(�}J;��e��z�`t���������af���0B�a�VAO��`/$�Sep��>��>���RT����T��u�N#wpK���~��n�m��\�e8�\��?G�fHjs��b�����s�B�=��q)�s�P�&���1aw��$��f�[]p�ʞ��F�0}�����VJ��$��m�@��g�ުI�Z.������'�T��qp���A"%U�������{�ۑ���wڗ�͟R������6c�;[��2)��p�S�P��+J��Z�c>O�,J�q�^1��2j�O��-;R�=�A� ҭ��>�{ኤ1ea�H��R�щru áO|���)8��#��_�κo�bWk�V�����o�
[�r��$=�F�9@��"���!5S^Vw�c'���nA綶Cfz��c��6*����n�9���>[�p,��[��+]����Ll�nl��*Zk�<ˏ���N�Zo���$<e7++�/̈q����9/�1��7�Px=����Bg
��� ���uNK��|�#�B[�&�4ӏ4��~-	 ���:�Rp�,5����ߜ�I5��ArC2�(�9�=�n�Z3�l �}� ��e���KX`��1�@�?��
	�#4����A&=��) t�ͽ��9��5P�_�v� �5�h�:&"I�Yhl!	�;����˪��WB
��e���d)h��V{1cX�%^0���W��8�M=bRrI��¿��9���F�%i�,o��+q��QpQ����f�"����Ed�d����d6��i��K�Im�,JɋO�m�U���[��la����ut\��^��CBб���/�O�O��}ޱ��mƪ���=��g�2��<؟.�ǵO�;�^W���yN���s#o���9e<B�U�<U�|��m��>b�{�4�D��Oz޿t�?|�a�����,��"Ϙ��X�t^�`���iW���9��n� ��y)���s;}0�P��V��ԟv)ש&�[��7��~H�	�#a
!9��d���ي�:Zp��_UeA�D�yR�!q���*��k`���1x��8C�F�_~��ݟ�2�-���L���c����SAd��;�6�H�s�V�\�UjX\����3����%S��s�C̛Y� >8g��br����I�?4�822\ͱ\E��9�?p}ت�I��1_���%�����e�I��`A����|��C9���h�Y6�v��y岹U�a��+�d�(�]3�z_ې�&��"��!i$���@� �0ݶ�|�~�
�Q �E��$�b�Ш�>��|�F�]���ǛDK�/�L�����
�Ȼ�KIq<?�#�y̭���R� ͆����>�&����r��j��y��(C�w�?���a���jn� ~|�PO$?�@X,0L�k�&�`X�9�]�	�S�����U��Q�M�t<��~4�bDU�A�{H&��-�q��~~|�Fd��ޙ�4.A�JՅ�K�u �<��m�9��5ɑ��ƈ�.!7�ms/΍��Sǡ�������,ҫ��� G^q1�4��JE8Ϊjm!Ffo��w���T8�$�e�gx�����W��P��.�ҹ�^������t�?oƅ$Y�1�ac���/�>��a��q�\��>v�k̨tft�S��)�6��-�:�hy���z��p��}X4��u�dY�{�:��k9=�֦H��'�m�eN"��$���pez���4��a��a[�Ъ���䵩���r����|\Oڕ���E橇?��L�غ�/�4��i J4�FqZ�n����X�M|�6��>j:m���AK�+7!��k��dL^]�r���t���P���Y�8]���.:�5�ͭ痔���@M݋�AHa�f���GӘ�g_��ը�OJ��ј�&�2ׂO�)Y)ý�ф������ãS/(9�h9�(^@y��?!o)��2�QSu2st���U���g<�g�����&몪<�E�u�@�*5㘗�G�?��r*�g�0J ���	}\'޶��u��n�a{��߷,�yGZp,T3���FVGZ�����������E���w���u�ĚEOV��#c�/J��x���!�Q��pl�q����Iy�e��u�u�����+	;m~ծ�b#���>� ���6��&��{A����I�
���jϝ��s��ay$G?P#՜>`B�v֔dU�nZ�r!��+��������ix�����m����~<���ɏ�f6��^�zY���!w'6�yd$UX����Y?��\��7m,Y���g�[3� /5	�=BCa���c@�;�K	��Ԏ�3�+�.5U�A�f�!?m���.��q9�Xc�7r���ɔ�y��8�Mq�����R�����;�vPF�	@n��6sD_&o!����`|M�����*�F�ɨM)ic�hE�#�9��%�R�fB����U��Cl)��}�KX,��̋�9�
��;��b�T謉��@�gZ�5��
E.��P����co���G8�y� :)��12�F�xT	�ZL`�64x��������[r��\�e=�%���[!@���!������~e������Q�t��y�G+8����db�6�*�
��|i�5��?+���%[��ᦽ�F�v�,s�7��~�2����h��2�9���� ,������
��Oao�Y�G�k�p��g��x���-0WF�c��?��{��⁹���!�8���/��r�u��|��?ø~�,��߫��~H�;w2��t=F3�)���nBzHG-�AޓaA.m$#7#��A��3����E߅T�䬆4d�d���b-|_�R��pi����x�6J`��rr�а��g��*�fzZ�O0���9��g�s&[�6[�wC�F8�'*����{���k�[ji������c�MB�R�y�6Vp��\�g�$8�S,	�������BD�oi�,#���U�V7I��6�/�`��fw7u�-O2��`/�;-�ք�g1�q<��Xq<�qi��
�� ,���h2-q28����.Қ��2�A��35Z,���Y}��u}��Q��Q��\����
KQ	Z�d<t_��R��)��6ɞ2�Eҟ1n��\c�����3�u�i�yZ�(�-?�&T?�YMb^�Y�bEc�������ǭ�#���EcW g_߻ a��2�uw���"����ʏ�?
і���j5�y��4������,����N@$����G�ԇ�I��|L��B��V��:nN*������[�w
d�Y�C��@J��Zj��������ݓ��}�|8�Y��Ǳ�lE�9Hm|W�����}�Y}���5�73߷��7w\?��u��E��u�_H�M�[����o�=x�{tI�>����x��Z���|BA���>y���N�����dL���+Q^k���<�3[����4�Pw����DBq׃X���﷿���읲2��.�k���a��|y]�su_qn72o�=)?Z%�.m;����[� �q��x#�`�i"_��x��,�L�,������z���w�O�(+>(�,)�ୠ�G�+5�kN�o�n�{D&B1Q��u����Q�/µ�~�@}���������˚��u��if.]9��+*����56��	�_��l�*UQ/�4��L��DgF^U��M66K��c����P�NN7��| s���ct_o��={Uw�]�:I�X��Ľ��ͼ*u/����=M��
�l��)'�����	%�Ij,�������ȁKI��(�d(HaJ�����fx/��s3 ڦ�f	ǦJ��JJ呫��v3e���0��*2���t>�4u��t_z-Tx5-S�x9��Z~_�N�(��_uLwoz��Վ�8�f��nA���`��+,�Bb5��������YcюV��d����kN��/��-������G�N�Q��G�KZ�K�����������NR�=	a N1M�->�;��4�U��Җ��R�K�"gc��,J�u����!�����򦬿뙿ʡc��p��QM�Bf��f���������'���>����f�^U:�NF�Q������ɓ����t5���jʅV��.N�OCtu$<�Ζ�N�)l;��Ȥf���F�qT���i�a�̊�<�����hG��G�z�Cl�w8���Y�as%����D���ȳ���@��'��lE��
0�i:0ʔ��JL�Q�ۥX̾�ɲB�E�XX-d�%[�Mzń-1�!�lb	�u�a�a�����,��|�T���EK�bkǍ>��~/�۳��bI�lN�b~j�/����2N�Gɥ������V��C�ֺ�r䗤�L��d�ի�Χ�_���M�1gw=��s+�`^7}yʹ}�W-)�^?Xnt^a&��ؖ���(ɡ��<KE�)7�^�`�e�5� >��Z.-�Xߗ������ͪ��˦$�����������J�_�nd,jL%J)�0_3����ƻQxQ^/� ==5=-5�б���.�M7K��~/�:K�_
�^������$bxa	>��4
�OL.M�--v�\F�Ft�|l�T��1�����r�5ƥL��3��H��F)8�q4hxkDU)lp��1������Mo�&�w2�+ppT�v�!+ż�i�e1�.�����.����E��F��EǮ��}��*��RƇB�|�l�	~���Y/�)u��YD���C�(�	M�a�F;��VEI�:��M[Urus����A[u������A���W~�Y�nA2��,N2��c�']H3߿Z۪���A�$��A��p�K�*��<��5��9��a-�YC/���K�Kz�$�Q*�tU��U��`	V؟	���3rS�5|t�x�=D_RB_lH�c{̕��ٌO�R��+�P��lOoP��x�ޟ���?+��`������3UM��g���w����G�JZ/�v��z���]�Ӄ���$wR_��5���N���Z� Z)�ֳ!����ID�$���'�׏,�݀��%�����V�7F7���Ex�bA�ȵɑ�����`����2����~j=6��G���F��j�5ָ�F�t��jڹ?�(������W�9ĭR饃̬H4�W+DմAV�3��N�L�G��<�����I�@=4��4ԇ&�M�_/��|q������<ri�6g)��;�_��飌�R���^,�`%��t��"b��y_�{	6���s5*�#���n��&���E�A��/�~��xq�|)�l����>P���y�>�kk]�[N^Π7 :�9��7w�t:�,�%aˎo˞�.��i�]C���1�8�����&v�������?�~6�S2��	1���O��ɜ�l�;%�O@x���x��˫M�����ErdݟK�b���NYc}���WI�Y��G���g8�m�r೐��}��R���wT���.�g�ʖ���"��2"R2Xc��-�! ʭDȺ炈�'�tA)�g�ӿ��Mש�DqD�����
X6N1#���k�o Rr0:!�ͭ$�s�/rHԫ�}cQpZ�՚u�R�ˉ��L6�K�௨����uh�|h�����g�r��/�_������+�}����0�Eŧk�SVY���-V���Nǖg�-#�°���y�+�Gu��q3�*��m�u���U�9-��C<�!���Ά~{�֏j�����0{����
�m�T�o�?��^PTĨ݅cx�{�Ȅ\͐�'[%�[�oC���Su\�&��[z� ��D�\#ʪrr}}}j&�?��j`�^�j^�*2�3�:F�S��'�_�c��l��%sy�j^57�5od�/�i��L=ii{��\�s��k3��&��]�j�kw����O;��73K>�s�O�ϲ$7��v�	�,d����N0U�ڵA�=6}D<�/��??Hi�J��}��b��ȭ����6��%q�ۋ4<��2B��>" �YY��y��b*s�����
a�eV �y����6�`Vϝ��0h633W�2����ӵ����'���Q�P��2��R�Dr���n��\u��.\�{�]�Ei����@>l�Mzʨ��9��w�N���38Q�1W�)ΣAhɻ�Q��u������-�
���ų��'G��6�����8]A�q����^8������]S%|��^zu�t(2�G/4����y�iW�o���y��d��>m�ܓEI}����W�A�&m9R��d�?l8�ˣ~<�P�o�2(��f��b����T�:���?>s�)�J���S;pڨ&�C��^.E�� x�w��;��*aCzB���@б���(�W��(:���9F�Ͼ��y����ε<^0�V��N�/Ǧ�c��'����O���f��ġ�����N|*���B����7d�Xypǩ�/Q}�e:�ߪ8e������Y\���?(>j�FsM���J����W��0�I��9�����E�1�z�.�]�c �^�t�ld�}0r�|�,�Rt-�����J���(l����4k@r����j�8�Q9����R���	���;6R�zw�9��e��p��t�5�a�4�t
����y,��s��bb?�����b��>���C;�g���jN�%���ټ�8�1��v���_�<gqb��`C.U�ϷX'����MN-�
��)�/ZR���y�=%ѷ����}�io�w6��d�D���4���-\&��8�+���J���%�7p#�����l��`6�]@� �\�|w���CC�N��T ����8r0p�W�\��gjitVqU�WJv��B�إ��;��276E0���Qܺ_8�ʺ�,�����y��L�V���[���B@�����^�ּZifXs���	U��n�;-�Ť�7���욜��55
��[?�$;�$-oMJ�2�[Q�Q�G�E�w��N�F�C��pq�'VV���ȉǄ ��\l�pq�<����;��-׻T���[�oyR�_����>1܃^�O�LNv�Gf�������nH�A�GOy�oy�>Q��~k��B���a�U��/j��]�%��˧?��O�B&&w}C���.z�+;�/�������J�1�+��u8��60N��M���OBC�x%P�4�Y��t"�f��̛�-1�����}���Fyr^��y��"���S��?o�eڽO j[!�m��^�l�t*f�)���9ܞٍ��=���8:{h���W�&Ԯ�*Ct4.�z֝L7Shp�����,w/�jx-���6���{�s/�]D ��;3��A �����u�!�qr�ۿ"V����X6�էI[BB���g�mY��珺��~W��~7w0�b�`;�
W��7��Rض�.QX�lĳ�	}d%�W3�cAt���7�����(M�d�����e��,�9���<�v9U����\�Jc����p�2�H��H�� 3J�����%ѣ[(P� �7���*tC3�	�z�������sG�Ӥg�㭧�(�Iw�b[�C,���놧C$�n�>/V�^?�܎v׵cR/6��S�c�]����E4R]@�\�4��������� ���  P�k��%� �<E�ٿ�Ν_Igv����QF檱-�-5��Ib2�G�qJ�2�[��c3��W d�F��lV�-�H{�_M����uR�s@P9Q���0�`؈��o�;��騥#՗�y�Z)��M�����bW`�v�!��:)��F�*�|x4v�U�X��c�n�\�OMڵ�GM�m��ѿZz.[X�xy.[;Ә^�n���gq�|:�U�Y�G�þ�
��Ra�g��LI��&Mh�]�M]�$�r~�sL6}���[�h�ӭf��mݑ����73"�0��1�N�{��)�|���u��@s3�-a���
R���9]�C�;3K���q:n����tBkWN�� Pt ���-e��������b��3W�F��0�Kȷ�5��p�t/ಆ�:U��*���}�}�]��Z�~6�eJ"%���o�1��?d�X�dL�}	<e]�癨bC.ƕ��C�(y�r���5�PV"��V:!K����\U�� p��=T�n���<k)��jl��������3�3`ΟΉN+�#�b�k��	����R��'H&d
�i�&&��'f����1"��n�V��2I��;�٤��\2�V��4�?vNz���
Q�7
+�ً=*��i��}�	YqY����{�c�v��N�
A��`�*~�Z^�z��kWީk�%.8>� d[rx� *b=;ؗ!�喖��F�]ز9����Fl�=�8Ѝ^��� Ae�##�çEC)\��O�5���ڑ�n�Q��"M& ����������������&����E��5_A�ǯ�N�-N�^����9�߳����bs�,=o��Bü,Z����R������_�p6����~Z�]�:[5�Zy;��/C�߬������z�R;�����pۉ89~<]n��r<����1���,���3����X��.��~������ۀD��Y(GENK92��JxtȰ��˱B�̔z��ؐ/7������Bҿ��Ƌ0i��s�~ v������V����eo���0U�q FX#�<��f�����P[>���	1�ڻY�U�6DR��HB��@���������-5���jgf��6�3ԦF���^�F�f��럷V��5�s���N%�܈�p�\Ӈ]H����$]rΒ���Y%�iE�����p5=J�̾�;�k��zL��䶪4���6�#����]�?�jL�����Y�J���LL�Յ��}��.�uo�;�}iv�a�C������:�"�G�4��?	�Ur��b��4��1��n����?`w�9��G�``d�����!�6EQ�KT�7�� '� 9�(n�J�ʈ���<�("ð��¶��ϱL�C��pi��9���K��:)E��^P��vN	'�'���:�����Z����y�<\���}��[J4�:��5�A|��SIO��pc`�3T��N�}!�o�Y1� K[1�D�臲!�˥̒�����(��H�d�d���D]o�4��M�Y�8�Yw�X��G��c��r��\�qo��װ?�E�Io��x\����������Oȴ�zw�pT�����/õؔ��E!��eM�8��� SBM>�R�H�5�;�1W�W@LƩם��-y��5K�5�� �"ܜ8�.ʮ�]D`���c࿓�N���5��4F��$ϫb>����s$��Jڰ��'4�5�zՑIf��"t�z}rܔ���x�iK�S��h{n���;�1W�� � �:��:tQ�Ci32���L�>ń��%�o�1!�V��V���}#�T.���v�]�v�A�Y8$\��.�K�8�J=�?�^�O"��T��MCsm`����/՜���ג^ i��c���e�@+�BW���+>����2�P_��cp����gE<���aN�Ѱ�v�<2��j��}xg9�K�.��%�;��>��V���*pڑ��GP�������x� ��-6�����=��;�������M�RSÂ}�Z�)���hHyQ	�%g�zi-���R�B�ᴆݝ�:�F<ݐS���DH���1k����rE�W��9�3��9��:f���8��e��[y�׮�7e����M�]�m��[�x�.���q��Ş��9�Ș'����u��j�m�'���Ei�Ȟ�</���y�[3lQ%ؘ�t�]�W�gq&_͐Ɣ�E&����E�T�x�!�������3�����z��������sw�����D#��:} �p~~�PSW_U_�q��4�iN5�����!��k��N������j���ɁQ:p}�[U�KC�%�Ἲ�O��k��h:�HZh#D�WH���>M�ʬi�Fk�����4�r��pkZ���hNL2~�'�O�L~����6
k�J��ѕ����Z:^b�t\?�w�/c���=ΰ):�7��4�pI�xn��5�@G�.W�[:f�4�5�W!��|t�Z�h�Cq�/I��HH�#?�UcS7%UC&� /M&q���z��+_<";RoZ��������bzi1�U�Y(���Fdwu��D�Ao��"�oB{&^4��c�H����M��>0�3�򧺣�!�5Ő�CiĹ�����Ɉ6������[������zb|��2>9t�Ni�SP�a¢Ga��9�5�t�v��^��@��`����ߜ�۸����>u�B����CT�q���	A;����Kײ,��Z�Q��k�ᣭX檗�͕ԉ���H�	�j#_j��1J��շ�.��ъ"�9Wg��Ύ�ܲ܎da�)Z@H/�8���^���o��.E_P
�� ��e|?EѮ�P���\7q�Mm�5�f�
�9,��	���v3�c���EZ�ԭ5NN)!.e�N��[]z�T��`�j�T;N:clI2�s��x�y���2J�U$�@��&���2�c����ߧc��P������ε�Ҝ�h���(u!}��3*$�_<տ��E�w�g+K%������.��	�ͮOG�.C����r޶U�5h��k].�k�$P���PƗݠӗ�fL��β�w��'b]���;R�+|)��1�O�N�qp��/Θ�m-�;�?PDM���#B$!sٲh\�೛�eZ4��s�2�#M[�����Y4E0�v�>�!��f�O�6ַ�8:�ğ�*�P��]u0� Fp�� �ID']U%�Ƶ"� �3���JP`��*��*;z���;K�*����[��ܯˬ�}�δL��7��j'�^N��0�pO|������7��l�K�M_�����<%3	P���<=:.�>�]��s��t?��CL��� �m3�QB�]s��M7;��\�c���J�����)%=$
�#p�p���v��M+Q���G�c���*?���7c��oG%OÇSv���F��f5+t�bg��g�G�{T�������xYy>�]��l"Ҙ������F�� |W��!^�&eYYn���\��]��g�q�f{Tt:�)��.-�W�#~:��g��1�؂#M���Fl���A~����ş��,��к�(�У�䴛dǏC�&��F7u� y_;m=Z+��G�W
ԓ����x&������8�����K^�C���Ǖ?*�T��m���م.�o�j9��J@{m'E{?eC� U[SE�/��.2��J���p5<�yGG!]y1������h��$��¤��v��M���hA ��{�)Q�|���WU9�z��=�un�K0��Yڽ�ܝ�?�b�Hw�0��>����oɡH�$/�
,U��rB1��Z�
����j�����݊���O�D�E��?���e��S�u<�]�r�?t��u���vF&[_����zʹP/*Q����c��`:��Q��W���w�H������v�^7��uL���yI�$��#J2��2����fIۗ���G�4�L1uf�5�y����s�3�e��
^`5nLm�W6�g�@����PbbgG�O�'6r$�s��ߑ�L�/~��5m�}��j��6]qX�`� *���U��G���9�d.Qr5vh=z���;V�����_��2�6J�h�-ǒ���� ��-�w���������Wuɹ5h�'ӫ$����׬�]_k��k�.<蝆F����L{0G�F\P��	F8�U-?�?ҭ�M���m�D..�����_f����K_w�kt䁰�B�m��iȃ��ɜ^1�-��ƺQ_�R�������3�5��s��gv��U��G!��w-6��yqx�Ee�
�T����?������k�a|-�^}�k����$��W�f�����($��非���[}:zLz��,�kq�U̰��ʧ�x�6���&n���j�H�n5�)�Y�H��W1�#�;����'��,"`x�EX�{����,%�������f�̀G���Đ���~�rA���q?�	��5+xz���}�|��v-h��̒)�m�o��2��f�k��N��`�B��b���F��?�ͩ I.}�ό¯F@��	�*I�qZ鈨wln�z	W�ٸ�H�Q�Ds8	o>]��)E��Վ�B�q�B��Q��%�H�a�aӾB�g���(�D�a�qb�,���|Agzaw�*�,��)����\L�L9��/DQ\	d�y� w��QMze� ���L	o�����dj�L�2�l��D�6k{��w�qH��`�0����!N�Zp;tML��mQ\3����t���q���y�?�kyW����Vx�V=����� W�B���:�uN��Q-��FTިp#�j](��Ū3�����N���s�a�xP"n���7̋b_#M��m�lG���7�L���I��}�d���6-Ts���:d"�ﴩY��ڻ@=M>u�$T?����(ս��h_�7���1��/q �S8���c_c���]�5����fJ�*�~
XC�nm|&�o	8Ա�bx����o5WG������6�X�D���DE�Lf~��u}I��1�c�O-\a"$nd�#G�)�-⫵*��=���B�o�45�O��65��:����c��霚_ P�MJ�1��ٶ��ڲ89���;����½R����Ѭ�k�a�>�f83�2�8��:�s[Z��ߒEa=K�1֎��N�v��,_��ꝟ�Z����~�.��Ut+M[8�9c �x���!������	l�������Խ�ҭ�̣Z�Q�)S,�_ �wj��ޫ[��L��;�Ϡ�;�U��nMdG�b�y���&4BZ)"�	����Z��b�l�9M��F��󶳐����䰄�柩��ɳO�C�j�╮~�=�1R?��?�[&�Yno{�y�^i����L�,=k�k���;u%{��.b� ��\^S^��X�-�%~Dĩ�����)�2�Q!�㈜����� �9����E4eZ���By��_����>Î�{��!��H��3�ė�Q�v5	:Z�����W����H�66����Q�e%hذ��\V�8hX%���Y���βKl3욂��Z�!ܱ�g��D�*�gq?2���cV�O1�%%�GU��ۗ/M���1ˑ�0ܗP��7��r�>M�� �\��>/ok\��]�b38���DWCWG[e3p}�O�z��=�Lܫz����g�zWG��<!�.|�i~�2���-���;�u�B�?��vb�{�}�u�D!��bC6��s|�~�+G)4^0Q�b@C�ҙJn��m��㬭�6����%������7w�;���z��Fx����Q�_DAȮ;���kK�O5iNkܪ�uz�Y�����G�	�PZPO��GZrlfDѕk2_Z���HRZ4֕��XP���ϡ� [k\�G�No*֝tH����f��i�P<�	�a9�è �j�0 6��G�:�|v?�>0������à曠����o�#;�������[E60'$��Q5� VS@\�Y�/-���36�ifΆ���oNf;�'[E%����s.�y���m��E�GL5�N��?��m�;�c�ktm��sP�5�FS�N�%&��~ ;�y;v܋��F��KI#�� �0�(=Q�d�\>���b��Df�.-�U�����I���������U';�o�XK�po�ra�w�WΫ�wWՏJ�6v^`�;3Y���_p�J� ۰���JW֐� �uÈ/�^�W�r�uwB&�\a�L֠���z�r'8*�(@�H��,](�K]�ˎ�zEFw�ô��kxݪ��?�~Da���-ϱ>���{Sn=���R�߀�ا���1r9�ih�
6�������)�.#���M�{Yu��&E_d�ŷ�b)C�0��������(�e��&�zg4��g�M2���sc
�Vld�Y)\R��쵮z�6́3Ӓ ۯ�c�3S�K��`�.Rco��Ꞿ��:��M�|Z�H����)wf�u�m&�iI���`�!{�E�콤��� <� |��~��^����i�y\"[�p���O��K��^��Rӑb������R�k���țV���]/}s?mk�ɀ�q3���EuS]���tQ1uTn�E�i`vj��{z�w`�ktr��ȴ-�l5�k�;��@���Kϊ�����8#c9�X<#Cܘ�Iw��#@�6,=ir�qn�1�jr�f�w`���yREm��*����<�Ld��>��2L����|���ԃ����vK�.3�n.�����p�"��(F�\��C�-e���u�ߨ��'��D�sH���ݿ_�(�+2��~ҦZRS���Z1�L�W�~�}4�Sɰ��,��������ώ�X'm�Y������#=ʁ��]��X��4(i��XZt�w��^�|W�w�?���Q���_������\�gi��U���<u.r��1Wr{��M����{��}��c�y=E�#����Cʋ��%���h�0���/_�8����n���8;�d�=dF%PG�$�Ïj�9�T"�)�\�Arz�L4:��3�Z�W�o0�&����	kP�_Lת=Mg�{�ǵ�	�z�y������Y���m�O���b�ŖrI��u���%C@��΍�����Ǽ�(yKy�r��c�~=P�Z�:H"љek�H�����a/.�8�^��\��ƈ�DS�2`�(]�6q�-�� �9��k��<�k~���Ѡ�d�����K���/��|�(�uFS�~xದƱo&|�9�fr��=H�����M�� gQ-�_��D�F�'k#����5Ip����
�-�#7��"��
3���n�<��ݯ���p�җ�U��lj6�8�����k�:� �)	��'ѿ0k"�i���Q.@�#+;Ҥd�ε�U���R֚'��R��
E5�@4����H�L��M�؈�	�k�xz��&�Pv�������e%���f�Ћ�;ߒn�OЩ�!���i�v���X);���$��wv��I�ôK9~�`����`ۛ���+nw*n�gv<�L*�$��y͑�'W/��nT3��������}��x�Bf1M�*�-V��[.��1��(u���`�G��ۨ��Qʇl�mT�4;��0\�Fb�������J�?~�F�Gp�~AAI[Uz�U�͙��i��%F�I�Q:�f�ˑ0t4a�.���-<1��S�#� ���;��<~)O9����&�,F"�1�md���"W�;^�=e3���h[/z9�d&�������:�n�^`(���B�u��♻�+@1:I�[�B=(S��x�u�5�(��E�;��Zlj=H��D��$����U5U��#k��@��MZ��72��CG�{�=ĭ�n��zӳ���-{�7zV�#��b�I��8X;���B��V1|��)HߥN���Ƀ^G0����Y�O�����ro�����L�`��J�a�r&��;#���<Ye��T��dH`54_�#�����ͳ��5?�׎h�r�s>I����{�)�1�!����=�=ʱ�
A}}���v___xx8FxR���2������m��{?כ���̶�h����������Óm�5P�k�f�Z�Ah3$�)]�ˠ�΀S����&خ�
:o��#��+X�3�,��X��Nx��΂�����؅=fi�i@����̵����fp�m6��`̕�2N�h�KKҚ�h��<��3�_0�*�Y�����Gi|�g�#�l�6��7ٔ�n�[��U!^���!�{�2\�k�ze�aMW7#���8��,	ӀP���iP��(bm����3�Ȇ�D��sgѼ1�V$ïV����B(�{�K��Qj�x�w8�����S#�u��ӊ K3�Qֆ��C`�����kT�^�%��3*�},E�_d�~��7�h�1��fL��_��Υ�lQt�L�TAY-�R��kM�����l�/��m�_\m�����_����Sp��{���0u�Am}Q�F�[[���R�h� ŝR<8�����-�	���%hp����/���w�~?ΜY���o�5{�Lܪ�~�k0u �D+J[9��ȇ,ʁ7VL#"�̆��*��4��$��5�s6�34��}�����q��@������G�#�:��^�l�ᑨ`1��_`�E���&:��Hr�Q�nT��'St�n6�e��v̲�	X@��<>�g��B=�����ϒԚ�8_��Jo�Eu\S�JW�0V��v**�>Eiu�'��y�H���h ?�F�(]r�RX�EY^��{
�V�-y�-eY��.�G��5D=3)�R�
�2�e΂ub�YJ����0�W�3vt�o�M��)9���.��W�ץ �ĺ�f+JV�l	�E/?�i���1kh��E�t|�Y%��D�%�)��q�/�F9�'E��Ʃ��"U�"[��E=�E��1O���%�3`2�_���Zi�iF�rJ���<��>��"��jz[ދ����"�Qv�U�Ε2���M���MS����}�%�Ld]�s�tq�t��߱��w��Y��$R�x2ղ��d�3��[;�)z��G�d��ە��ژ��U|e��c,}��L��������W- ��76!� @����$F��DQ3��2�Tp,�aF��s�D����=}�kC�ס~��W;?�����fo�<�G���6d[�ɏv�R��_���X���b��9T�����eo˭�s��#�W��0���Dffc:�y���PfsK�� �����P��,��[��D��Z�|��AV�$����n��_��QG��Ӡ� ���	���"�w'j��rhʳw]�����k?6>#�nfn֓=�Ŭ�p�qjM_��-0���m��9�F7N��N�����N� `_Y��R{��ry挅��&%L�#MK'an���f')��խ.�&*
?�t���KSB"Y:�Կ����qw�������ݳ������wnnNSS3���������Y\\���kljj�l��r0�<�//NO�/�R��c_ګ��1.�.1�/�t�䴌p)�k���HC��_R�!�⥁Mf���r��~'�w�2�Oϟ^���;WQ�ۙ���]�4Z]K����B�y�.����v`_^�ɟ��U
o�k�+�a� ӟ������:q<���^5_�;@�u�w�d]��`C]o�����U�瀽XPc�F}ʀ�|qE�,߫ڎ�X(�o�|ܕ�<�� ���2� ��� ��@'�h����K����x�O��[����O�c�������ez�ΰO������9�-ࢗ&��f�g���!�5g��j-<Vk�º�S�j��#�9"�u�������ƙ���x�]�/���Z����I1)Qx�Bl�8,������� )H7=0W�u��5:[�����o�n����j"=�Jd� 6�(.���1N;��zb������$��wޙ��̝#��R&�O����Q��d�χ��]��~��w���@A�ͯ�M��;KK;;���Y�����������e��u;� 5x����71�wۈL�?���F�2�K"7F�Y�R�K�oC�y�Cd��NA��Kñ8J���G�
 :"�UҠ@�\*s���]Y��_��>�w+��$o�|�9��	�ľ��.��+]��|�R^?�}�Dx_��u�Ϛ��zׇ�����Q].V�T���۝���i(�����w�@5�S�!X�pz�4Bi�y���%>Sl�Aq��Oz�^Jm��}jR�4�o:�w���	������c��Vt��n�%�^P�2g����'+IZ��E{��5พ4 �.!+��sɎ���g�� �Z��a*֬�f\�a?�L����>B'��i�:��iH0��� �;��<X�:Hk|��=�}�l,۹I�&*�/N
5ކ��/Z1�W��ܟ��(۪Ne��޷���SM�XNkE�x�I��-8K�4���1��wsx�x��9�igJ������X�(y�^�}n��^Ըw��Ro�$���j9a�[K���!w���	̫C��w��I�3^*���t'^U���d�|��U
r���g�Y[����G���yHZu��֨M�r,0>�������rG���C���Ww4r��t��3�q<���N�V�{���Cdq���L��z�N�R1>������ɍ�;[�q�y��M�t��f�(������k7��pc&�|;���B;~!�q�YC���Z�M��~���;��Y׻N�Se�ӴL��K������w�:����O��Kc��Zᾋӧ�W\OWH%�Xnmi�VPb�$�M��5�QT�0��RѴ8ofꙿ%Q��l������蔦5����թ���[�	Ň�Z��F��fNu���pxq�P�Faa]_(�]3��A]IM]i-;+�'�4x��:4�5 w���w����˃������C}K�($�޽KKO�~���߿�lcSlg[{��[�����y6�57�y�2	
.�����;�[�9��y�T�f2����Ճ��ؑm��*n�j�j �c��6(���4���}=�B=�"ʂ�_ξ]��Mb[��ˍ�Q��'ٱܣ�z=��O��:����a�Q��x�#QW
x�ؐb���*�$J�����)��ov)������'��K��͋Y]A%l���nuL6m��
����d�3
������ͷy�㳨x?����cZ	ڋb�c�
�x�
�r�d�� ��A��f2�q����_��e`���ڶ�����N+Γ6�F�i5"���dr�tr�Tb� D=��w�_o���lܜ#��d;޵;���%�X��3iE9Y�^���~�{��R>͉�z�e,���5��\�C����_�)������N�:O���'��mdUӄ�ƕ~�=4ؤ9a��������	��1�Rn�X���c5z��f�N>I0��ݴ�:j�����y�`����z�/�[���	��@k������1	J�%�z���*�/iW�9�bbBS�rF��n/&/?��t([������R=8xR���~�����oQ��7r����xƧI��Y:HC*, Ar��d��E���~Z�|�]�
�\����N��@�8�L"'�1DS��Nƈ�n���<�+
�nטC�̅--���m`L���h�</}d�c�5_x��C&!�[��������n()aT[1RQ��H�o�c�u^d]@�ƻR�ƾ�w�)7��~ؔ@5?A��Q�$H¡d��	0�r�!dn�����ˎG��<ө�=aB�vW]N�V�w"����~^����UX�7-4�'��|l��s�*�Ju�Ń�����/Koæ���p��,���2C0y?�V����Vӑ��n�9#c\��v�p��e�dw%����+�X�F����8q�Dl�B�%>���E�C���Cͽ�z�q�9�p�j}>���C)�.u����M�w|�B�����`����Gl�W���Tg*��"T��R!�u���؉(���R����ky��Y�6�5x��|�?��w�b��/,�wfT��M��u��E��>����օnK͑�5���v&���J|1a��Mk��ѝNx<�ݼ^��e�4��#�Ÿ�p�U�0+�Gxl�+��d ������<��޵�2E*o�i��O�����;+N^٨���ě�3�\	���>w'G�V�i+����D*V^=V^�O+ I���◂~���d�}ĐI討*�P�^%����%o!�n���a��Db@�Mel��çA)�C����`��411��9������ ������M^��\�?�3C�p^��of�Y�;g�O���,���]Ʃ���>܅hQ� T}"={H���Մg��1��U������U��v��oZJ�Fy�Ȋq)��pJ�W��;]�A�~9̽�f�^�]B}S{:��6W�8�+z5�(/Vϸ��2�ڏM�3Q����y�@�(�U�	���Gɘ#���5,��D]��_��}����?Wwo�����
��C�l3144;���?~�&�� *7&:ZN&���d~aan�������wNX@���k|aAW[ۛ���J��W�(K �w{w�)a�����RQQ���MCCCZZ�����	��ʍ�\�[�$&���H0��ްP���c�[���ܤ渊и�B��$�_ak{��_j��2���@�yI�]�L���<b�Z�FQ����.�#���Ek]K]Z���K��$b���e{}�%�3����Kߏ�w���|o���xnxv/8Q^�S�����i@���Fk^�+)� �$��]A�-aگO*-���vRs˘u��f�S��v4�N�W������?F��8�QO>���/�7m�"����+WR�0o�>������#�[�hbŌ���,�]�'kTƄ����[t�?ȸ+�W�gk��6 �@��dT��Rx7�"6x]�����;�E���MZ�(U?%_uS���g��Y�����@�n��NٕY|i���&r���C��Ki�P���t���Z�2�W�ך ����b�Jc9���)�w��)�B��H:�]k����̢�|Fd$R��'5�&��j��D�k"����=�U�-m��n�OQ�>�����Q�[�h�u{#fN7Y������E��xT�w����鏪��i�@㪆�:����������y�\�6�8�EP�X%�_��e�5����Ӛr�;M#���L�u<�+�iK�nfe�C��BZv��ةŲ:%���24�A'`�i�k�N���L����	�����z�E?77���
�9׵p�|�,TU(k��d���\Qvl�gtVb�I�>d?�i+���"�ǂ&� �ÀF�j�|��KP����/ϥ�8���M���	C�Yc���)���w<� ��	Q��"��2"^�f���4(��H G��yb[Ϋ�8H�b'~�h#��>Hjk�DRN��:l�IJ����J}<V�a0�wDn��a ��BP��0���W�ܤ�]�
�!�;����j�`��E{}�u7�ӱv����'�8�VR���n]t�\����kl�v�*2)��p��<����L	�(�j���z�����t��������l�u�R���M����#|E���5�����ʾ�M��)�ކKhE���[~v�Ds�*7\Y����hh��P�
�b�wG�w�n'�.I�ɦ3��-�1�%�S�
��%�.,N, �~C���{t� ��4������dӄd�d�X����y)� #��g��X�ϧ� �d�����N���Q��c�����Qͯ��y���q����$I�H�3YG�b�Ë�'����oN���Ǉ�u%5?���n�?�|$纜���[���s-_mI"i�?l��/]�=������hE}��|�#���?K��Z�kx7�`��d0"���h|�%�.�w���/D1��z���P5��X�h�!Ъ��$SšE$��٥���i���{�F֗�51��DZj�Y��ǟѴE�n0���g����� 4�����'�w�4���4d"̱��ҋ}Z�(���v���R��8w�4Q6e��[$W�af�Tv�"���;���`��^q�!D�X�((�$5HQN^vj���0��C��7G��d6�$���Nu�}l�햍�KW9&�dX�4�0�In�gL���A�i[���Y�}#F��������zj�==el;<��k�mf�� �W"�#�3��cl�]�`�H�f8Nu�y�S��I�����=�yM�y86ߒJ�l���9��ӧ⒒���ٙ��6����T;[[[Vf���hWW׾�3{^\. W�F�6K�p�
L ��gZ]�����6|l�'�w��;�y�a=�:�L6��@�C��T��A�-���4�'u����0��ϤJ�6,�W���^CG/IB8i�Q�%���C�09h�� �R��`�t��Gr��AQ?�A����n���<i��Z���~���=�Zl�6�m�݁��#Kw��4 ��	h�}eC����4Uz�8�g~�~+�;$��s�*��II��Z3�FH�m�l�#�reI�S ���
���#aWb2�z�����R�w#R� >x�?c�a��K�s�A86�>3�������݃��7�۫��y��]��\h����~
�Vk�'n/�Z�U��B+��kvP� ꔭ�5�/���~	Q�&�x�>R��vR�8g�sP��$) H���B��!*�4�,�z����g��7뢝���zO�~���xȫ�/�*ǀ���n�z䷂�o�
ל@-��߄HT[�Կ7�5pR>���/.R�:�9�<��E1��j���T�V����<_�K`���"���	5����da��~#���0�x�c0��D�J��^CO��"�?]Nܬb��� ���y�z@�1��	e:F��jqe�F�@xPૻ�*���x��(k�.���gv�	w�S�E?����1}���en7֦W�"j	�]sA �I���.g�U�A�u�n4��唃_���9�B���+�����Z��a�;ϗ����vBsm���C����WB+���\o-��;��s��HN����=��4(�wS��� �0�)��:��G�`��i��#��jQ��VU��\�� ���`�+r1S2�]h�P�Z�|,*��"w$$��`!�
���'����YJ@�S��.Z�g�@h�S�d�-B��@� p�j`��B2�c�9�I����cC��,w��ӺD�iSw˔t���7�UO��b�O�徣���<ҡ���>qQ&Iz#�;��0�ͣ�_WK�}l�*��+;�u��l��^�6.F�0n�����XeXBȪ���Ic�#���3���S~3�}wT�z}q4���l�^��r�ZU��jU!�:{���6�ڡt8�ݘ��=��zi��6�IQ�Ĺ����L"Шy4�	9��X��� :��-xؚ�,u{M��粴:8�v5t`,���!��I�y�����ѡ.�E#�$k������z`�V�הл���/֙-���5iR��K�U�Ep���n�H6�-P�)��X<��C�u�i��V+���$�TS��!Q(�q��k*3����(|.;�D�_R�	S����E>�'��<���n��/(X`���sD�p�8�p��z4��i�r�f��B6~�g݈XR\|�������߿���(r�����W�ӷ��mmm��K�Ξ=�ƺz�30$��!�����R��mT������֘]=�b\�@���E��g� �^�CpăPa"J�D����T������X���yp_B����RZ�X�-@����]a��x��a��uO��{��b����׮��l%ɵ�����w�����A__�:��-�sv�J˝��]�Va�1��q �~�^X;H�L��$26LglVkB w��{�W�)�L���G�s߉��>X���)�� �i�u�G2f#!�ʞ<�<�p��6��}�S;���eė0�@�d�����	0WV{BT��'�����({�����'�#}.fN�(�O���	?/����6L�Q��\7�N��0��Y|�b\�_�s	Rf�����w^(DEղ+s�0L�a̴�cv�g���q��x�������{�?jI��\8}���o�T�+��~6��Џ�~��9��ӣG��羙�գ�I�1h	,3����)���_�2#���zN�~�n-/�W��xA���������,#la�xd3^Q΢�<q/��)�ѭ�����*�>�.;��e�`f ����;��c�Gg���t�|8���J~뗈L�MK(��#
"���#'F�LB�K��nn���C�r�/	�I��P�H��4Gك
�����'�����ߝV� ���Z�O'T�Ʌ?��@��l�����*��ޑ��)���®���~t:�y��Ζ`e��G��]~��5���feu׽a��>w�􆍵��E#&���P<�����3K�@~kE��3=(Sx����.�M���`�A��8��g/�
���J2D|ݲ��ؠ�������M :���Z��p�؛֒E�(�7y���#)�P�4Q�6Efފ�h��U6 �J������/�0~�mv?[��{0�p;{���ح@o���/�4�:��uh�����%laڼg�dgj�nY��������"a���S��y�(��	f-
$ĝ�h'�C&����3k�\ �f9&�ĺ�����
�����wy�(4� � �hz���."�-k��OF	�Ԧ�7`�K6_�%m8���CF�N��?V��J�Z�D1��i*0���|��we�N�n���9�Ǒ��9ӣT��.��~��A��}=a= Z�blEwJ8�v��.��� S+���#�B�k\�7��,����Q��da�
��zU-d�+��jgJ/���|���9��S�	�y����tcf��1�+Z�פz`�9F�\6d1 ���Ȓ�Xy�u���c���J���?I�dp\\����<���ɖ	�-�Z�|�2��O�����Y5>Z��g��..-��齧�8�߇�ٝ���мz�o�mU�%�
�v+D)v_�:dY��ʙ}�VU�n[��BU�Sb�D2<)�!`U�3�$87�q�U���DXx]W����W$�e�8.X(�6�zb&�6�Nq"r2N���P�mI�0Ӻ�/�t9Ų����L�mŊ�S_n�]۟�G�
���$���Mٸf��8���ouGs�D2J�����q@�]|Z�[���XS�+�yzۊ��Oi3��Nǽ
�W�j���Lډ�_>�����3v��[�!X�p�<���zp��a�$d��B*Y��j!�
r�����@���n-��.�����;���l�9���z�LJ,��n�IG�X��(ʶ�d�"v�VD�G�e^V��bY����N2��]�����(�e�y���b�p��1��E7�a���bq��T�ɟ�2�z����:/���)��������KT�[�j��`;����Z�e���|�J�I��3Ǎ�t����?<�7$��껒��Az�e�W�����X��s�|]\.��H�ei/�C���/9��3�"��Rd�g�>h$Y22l�[��e�\����v��R��}���dIj	�4�k��DmH�;�������p�^[5]��N5�қ��:= ��9�r���voc�;�-DV������󃕝����R�g�uȉ����W#xwY�}��L*���	��� /���zѹ��	b���6��9
�FO��(�`�!�i� ���4$�s�h�G�=�b"�-;��K?h�f�,q��f9�j��Ҕ8B����7d���3w�Q��.�U��lP�3kVq*�X��OBV��ZC/V���{+V��\ڌ�aMm�f�
���q�\o�X�4i��f�_�9�%ޠ��[�~)"�f4�d�R�bhC�s�K�5`Si'��X�3^Һձ-��8O��{��6;¥�^X�M��#;���.(�`;��[>D��N����-J�+�չ^���V��1�t2�{��Gt�7��e��s���'����*{�X��eа�X�d�C���V!�my���""/������AC� f�xΨ}\u�W�����x?��n�v`\����Ԍ���+ۆ�(���nl�h<����2�Ȟ�I��xLٞ��K~>�D����!'��� r����z�- �	��Q��+L۩ń\v��7H�v���j��������Z���|�A����wlo�A\\ή����4q�����嬚�vv1��z�99(�/�3��T(�Fm#~(��)Uj���:E���՛��K خ�	��^��5��V����
��\(E˪�&@ ]�������=.//��*��_����y4��d B����ρ��<c?j�U�d��_h���Pk~�������Z�F��R�&��a�.�i�2�.p���d�j+�%�ֿ��񀔿9�`���g�;� X��\3���b�3���t��Z����_0���r�̱Dz ~-�o	�4���H�;c7�(��	->ay?�u�Q*<6�=�E�z��mdB*��h�������c��G�.%���ڔHK#4�!x|��
eT�/9����1�cqv�Q��ć~d�6�D�A��~J��u�~���*v��a��kw��}�����l��$��Ӵe����|S����xgU\�rͲa�̥�Nڟp.�Ӻ=�3�ʆt�+t�[[��9�۫���'��b�X�i/3K��V_�ye6r*��i檺I��4ma�����i�O�[�r��t�Hw�?ڷ�r���t|�|s#`D�Ar�YS�np�|$���F���|�M��Ӓ�|E�~��)�5�F����5�'y��~�0��t����V������u"��D��|RV/�i�� zQ=@.`��,2���3;/w�ST��9l�@���C���\8��W0�dO[Vй�¶DE~�Ň�.���@)~�{�!i�r�0Xp�C����q�{qL\bg����[=C"i�7�����Q��:�:�%��Y8fǊ`�Kr�m���u��P�ͱ�29��~3��J�Y�>���VUI+y��;f��nv�c��U�\Q��sRԝ�b���R��1�6NԲ]?�T�+g"�L�_���,�BƤ<���� �@\4:�����͹�
ػ为��On�ٻ֎�o�]���<"�gT��4»H|;��'޸sݞJ-1W|a2a�QM���̘�l����
���Dn���#����ʵ=K\!�r�0��>�1���X���i��������R�����X`��������� a�y��4�j`=k
!`�Ec
��|���*� NsF��@�"革�:���K�#,~�����*O���9B �b�ժ��0E'���ɤg���JS�z�<Ou�����>#�獐��I�Y_L��!W���AO�*v���?��q����������B��jlGG�'�걮��plY��WX��dQR��뎍�����?{��������475-,,|Fu����[����ϡr���U�'"~������z�D����L�v�ɚټhn�GJյ%�+0��P3�z׵��n�h�%T&?�ٺ*Di��Mr��`K�iCWs�l�7�5�A�U@ۥ�,�D@@}�׉�^�ܣ�����N�U~�I�������B�U�Ek <ڳy�fM��#q+��G�*L��EM�d�*;��	F/���!j�ڮ蜽ܲ �h�;gw;���4��=T���ǂ��鴜�t��@�n6�B�Lu���U%��{Jw� O��]b�����S�ջ���;��x���q���q���ĥ�H����i����V�z}I/�I���:���zG�i�0�FY�7T�����֗C�<���B��-�� V0v�$[P�ّ\�k۲}v���@��|*�a�=��6��e-@�B#˟�'?��y϶:Oزkv�m�C��{@�$\l_5��nKߢx@h����˼��j��'��ۄ��㮰�,�\њ1�υ!�)Х.��n��U��*R!�vL� ���`q�� 2Nc�0�� @��=&������S��� �O���%��[��i.%d�?y|�����R��ӣ�����G�x�>;��F��G�M".��(���w��9�$�l���q!叓��6���#�YW)ֲ+]�����57��c�Q�^�e�c0�pҗ�<�$M ����Jՙ���]�;r��0@����7m �i���*uR�����t�\ XA����K"�J��X�\�B'F��B� �B�1�%Ʉ�?3kF	N��RL�*�!K�F�����B�=��J�8�[I=ܫ�����wtlYi��֔�� ��i�q��
n�������h�,��}��A�#���@> |�^qQ�I�/�6��Z��-$0���+��2J%����ϯ���Ƕ>?�V������}=���5l�K��_�m�4~0`�Q� ��������k��e�(�*��-�?C���e(����4���0sÒ`�:�p��������Q1��%�s�'X�S����a���#���B&9��l�����1�z���S2��[VU�k�'��up�׆���}:�>�ͣ�U������������lO�;����<��؞���5���=���k����]�F�-CĐ�T1��r�itG��܇����n������e�'�ݯUG绖�Z���8=n�${=�)T)1 ,����k���[6��2��fff�^������b��,kii)+r���m�4���u����,d�h�Z[C,N, P��+�u���k% ��K �ʟW)��3��%�NLO+LLd�=�.}���%�����/H./�����R���^���ۭ�]<��������4�ۯ��v�UW�l'�/.xr"OCn��hXW��\6��9ԕ�c��6��~�P����k�U kI�oN�Bͽ?�ת�\�:�Y_7�K-�JS��n&��<l������n���_2
�* ?l{yy�����x�+H��x�_WѸ�3�q���Y`U�]/ϕw`�>J��,xm��h�!��dtw��@xeWW��*w�^������2y�5�k�W�� ��-���H/Xl�TjoB�x3(M��00.��^�4�k-�#)T6�C�A��u��٤ŹX̿j��U��@y,M[~�~�ɶ"�1dj{ͥ	���7S_��N�\�0,7�K���.ؿ��V9s������mE����$϶�o/!w7!{�.��o��q@7�A誶��bw١¯��F�#p@����S�[��Fu��&3�DΙ���MA|8�%KV5Y��xdx#��� �d�~df����:��:�XW�����\n8��腜��\�V�{�[�M��N��=e8��&�͓9�Dޒl��_F��<-n^�/bڟ�)�����ݯmw�G��i$jە9/}3�YZ��J����	��r���ăͯ}�0��q��J���|w�5���=8��H5 ��Ίy7NدPb����1����U�� \-��׍W���
&x>���;�/�,�QFVTƖ�H�O�|�3:�̛�U秲�,uM��drX{�[�����J7\�l�����*��h����آ��������8K=�0k��f<>���.G�,�T�͸>�ǌ�j� Xy|��'�Q��7�����c5z�5c��cq��;�?.s��)���̽�G��m�5��˛���2�Y3W��Mb��ڼx3*�8����;��Lo_��M��~ߔ0ݜ��Ы)�ND��6�����3���`=�\)'ߗl�̺�QA�����3�c���JR+��u�	���{ $#�S���ޭTr0���Ö;�{oIn��V�1�X����~1��*N���}�6�0|qz�<[̖,��RW��G���8Q�}s
�'���h{(�������@~��C������	����A	�R���u�Y���*�&%��f�~����������bh�}x8��,�#���f{���4���'֡�x��[�()cv�H)cy���u�1w�ğ��㻻���Đ@����{�`z'yRU0�=r��L�߇�)2�.F���\]�")����t�;x�e���2��3++�UMv!6��j93,�VRÉ��������`>!/�#�_@g4"�Rʠ���Q'�jt!����P�7�H�-~Y���=	 ~S�~u��CY�su��t{�S>v��iIJ!���A@�l��eG���E��"��:�u��qE�Ʈ�i�����g��2�~t:c薎4��.p�z!G�S[-��,$C�'vp�`��X���M)�켹l8�\�;3TDn#�J���%L����!����+����+t�[����נ�u|�.��Q�znJ��3n D`�y�;�� ��T���bPOݎ%\��8!��f�@��r�,S��3�y<I1�t^���+��Z�����Z=�Z���H��������o�h�{e49��P���� ݽ�P�G=C�G��G�?�%o����;�O�u{ݼ�9��ӂ�G�gͪ��rЖ�o���D�����9a]���G���ha�1�}�HSHd��i�������m��*("΋ͧ�+��G䰣�z�߇ OM��Y:��ƠA�a�S1r7-�[�Vq�7|�t��klp�r���B���͉��?oŴ��T������Zy�B�mo��f57+f������K���	��Ͳ�\x�4�K����Г2��Y�9L�%\A]�}�%����]A[x+��2>��,R��Rݸ<<g�~���˓��Aw�%���t�5�sΔ�%2�6+ȥ2��Hy��p.����������a/&�2aأT�4�K�Ie�nҪ���rCA��D�Ca�С6�� ��!��.+zmb�������@�����aJ.�F�h������ ��&"3���ӌФ��\g���x��$w��1��Z�dsk��׽���|�i�f������������QlQw�q�	��žmɨ�n%�0ɮ��Y��)�V����E}�['q��@�zQ��������y��ˤk�o/X���<��K�����1XD�\M5��M~��4n�S\TZ18$(n@�h��V͙��P�t� f���O6���9�`�_Ex>QV��8�?��U�"����#�d*<�!�Qܝw�g�V[�v�.Ѯ���P8�!�\+�'Yˈ��'��2{-�r\"�M�R�a��{�/)��hV�fS�.���1)`�gl�O��ձ���45t>��o߷�Z��	�N�Ȣ����8	���=����oz��::�ci�{�]���*SX�w��l�T;[?z�*�͟d���!��IB�ރT�{�g�5�Pk$_�$��1��8E��#��ඊ��&�����a��W.Z�y4l'�y*�5Og�bY����ݐ/iTEXX<Q��� ���4�Ӧ�]=���=so����tYS�!<"� x���ږ�#�κp�". h�K���UNMI]IsYY+����߭ut=���f9w\��6�c��4��*�X�q$)>C�|�AV��޴����y�_|�6p�N	.��?��'�ݲ���HPY�u�(�l��jO���	�{����%�d\�jF��������~?3Z�V{k��]�L\�&�A���F�igZ#�f~��z����G�^��Vi,���Q��X�qwvU])�ߴ�n#�k��ܔx�P�L�X
"_,~��z�4�V���"Ϗ ����J�̤R*�u��uM#�[�t����Ϝ�6Q�s�S��L�j]���+�O�t�Qֆ�.��N��i����>?F�O�K�N�B� 
�Q��k�������J-F�0l��X-0�]����r�{�)�J���=�=/$?P9��א�Q>�>f�_ɻ޹|����� �ZQ���;�����R��1��:�> W����@�8Ws�$���_��4�Tp�tۏ��Y�p;v3P��X���g�8��?z0�V�ݺ.����1.N��uY��Uo��%����dz���¯p�����z�?��d����^p�������Y�~st���4�V�T���7�p��B��=���Vq��k$��O��ΟCQ��:N��r���
)�ˁ_�1�47/�l�J�^LEӟ���h|�z�]L=��{{����/P��Wr)Hڰֈ��p��P�:� �ŷѿ�o�q:�ނvm���sߺ����o�Z�����ʹ������	v+ ��^p3o*g��`�Z���;�u��`�Ԡ+�45ѩ
��}�d�R>��ެz=��Ϳoi���P��qݬ�|_�S('?�	/�N=�>��u�֭M���?/��2<�`�8Av:�R�;S\H���/�
+��n}nMyN�{0�_[:26/� D5u7[<��d2FA�=S�9��e'��:��c@��4==Rh���l�opv
Tqt|���Rд+�^y'�cl^*'����\�99'��wa�b~���G�P�|��˹��vWZn�⛐w���Q���npo�[����4�i�B��bۓ���t�0�����E�"�@i��(4�T9��Y�ڤy�V �9[�N�#G�0������j�zXy��ԑ�2H�#<o7�%�,S���Ua�gPx��U����O���n�r�0�7�)�yo1�r-�6��R	�@����E-�CA�"G�o6�}/,)���O�3H��5CV�a���C�6#x��GK�*
��k���-B+�kp�R�eU���R^��T���e�7N9����="��C��Ӝ+ع/��"�$p��	��Qxd|��N�����u�����p�QQ�a�69���J7RCw�54HH!]�
H =04������ %�]������y�z>�O3k��8��u����Bi�WC\��;:X$�`)��0{n���UWA�p��H��R�,�����dn�M´'p��f.��k��k��p��1�fOg���_��E������D̬���n,��++��u�yW�{��kZ8���'�ѭC��ҧ��_��]��<�026�Hq�{"m|�\�_������h��l��o6��@dT��Tm�OFL��O�ۘG��Aۂ���rSY��s�;$���c4��r�ڕ�t֩z)�9��C�.��\�Ռ~	q9��~ϐ���FGp]�/a����ڙ�=��|U�]�v.0�#7��į��?Qnw�ñD�h��|4��=&"�����\�i���G��$��Vd�㵞8����������@�1���� ���R�#������iuڸ��
g���S�T[��b!i"�W�n.�����4�t���K�FT��P.�	�����s�p������;TC��d�U=�1�gب��|��O���|��8a$��͵���r��Dʰ&�rrե�8�����/��-�8js����W��q/�O-A��Q���{�ˬ�h����*������?_��R���I��h�~�Q@�	i6�q���N0��0��}��ۥ|���P4S�.�KlJ|���#�1>��'r�?�F)�7�k�:�\�]g��O,*B��rm����I26���$�v�����1Qz-�~�߯�D'�@�d3)�Y	쵲t���t]F͌{�q"v�����'��Ѕ�P�g�&�&ǟ�@�Շi&��#X�"`���,d{�e��aE<��3��|�x1�ߍWa��W��w'�����N}�[���'�\��j�����/=_|�'�J�ɺ&���|�z[`�:R�rL�OJ��ݎ�̿+ű�Y)���������&&�0�}�6g�y]�
�P,҈-y�-�(�JY���A����������]�7��cw�F��:�����I@�>%`���!�w#O�؞if�����]�M4N�{ץ =X+w=�y$�le/V�m��s��9~�?��yt�ǚ��h������{�ef��!oN��03eVN�#bَ��e��ώ0�����e���e�'YQ6�{����	��Zޣ���n�tO,m}P
�q�d
V��
��N���C;�`�駬F���-a���7+H����/A�/����@Ez�Ϻ�'oR�j�-�
+%��!��_9�QY���G?i}�H*_��r��+9��/-��j�&��+�N��x��	��?�}7yc����B�o�?�۷�S��6���WH(;����b��U1q�>�>�����b3f��!������ԨlsC3����1��t�7���<>�|N���M�d�>7[m 7M [�h�4cǲ��y<`�Rh�+U*��k�=�w��@nҌ͢�t�SS1��Ɔ�-�şS�+��ⶢ��F�����2#���e��<"i�YzS�gS�y)�Z�S��2K�sU%o�ڙ:�8!E<	4�X�b��Ld�����T��@�T佁iVPb�>ԃM�<�|K�YkPB6�]{����~K�W���j�k^�
�^�45�IvJ��n�ؚ�ƈ��iva�Ȫ�o0|֘u��3�o����}� v�9��".���2-Ko�١��?����
���N���Hl�P�Zh�]i�wa��.�+2�g%+F�"c�c�WQ���/`��ޢ�+Mw?i�Ѫ햩})	=���I�'&fn�/��g��|qSu��q3��J���-� G���~�l�UknA�4Z���B�&*�y|�3툯鈿�����"�{�c܈��ٹ��i�����; \ra�=��k��k郿/��r-*NN��F�dc�ێ`�X�V��l�ڒ���[X�Ә��&�_�
�|iF�q��hY3$H�<��7��kAp�<�o`T�*C�mdt- �����z�4*������$ȇ�9��28�h}�'"�:�*9|�`k�	��K�E�C<����Y���M�O�����L�µ��%�\'x��2��w�Su�c����/���o�:�s�;����"���`qe8���t3��aM���Ϡ�@7GW������+%�����J*$����+_韰טsx����ʧ���1{���J���c�D���Z;-n�=k�o��7���n)��\D:�H��L����Xo4��%i������8���+!%� J���3� �DI�^����c�T�L'OeD��_ڸ/��U���>v3a�Yb��g}��4���AJ=�~���U_X:=˃Ш�t�(+)o�ҧ��	)�?�s��C��u����R� ˷�c0Y�קP�t>EB?DA�/�]I�3:��2��1jS;��A"n��!%4[���e���[bm[`G7\�k��%q���E��?��w�c(ҩ��=V,�W�F��(�$��~꒧���7�ϔ���I��V�'�Ш��N����h�)c�ـ��,��D�sAɍ�rB�&;�mǥ�j�w^�_�]T��G���%On�?H��&UAf�����핻t��ϫ״l��n;J�N�((M��Ƀk�lN|���'����:�9,�?�(~�zib�[Om�ShJk������$�M��Ъ8--M<��ІWےe��Q�TR�����- :Lw�|J�䔏a5�#��"��n& K�Fi׼yS��k���gj%
,[3�^�7?�v�K얦a����="�tc�NEI�Rٙ�H`iP���đ�\��$�%V�dYWN�T�������

�zF�V�٦���4ԭYL4����ٍ�ɝ�iJ�����
^�}�r?sn}'��C'������>�|6f%)s�e�H����T#,������`�,8Y`\$��&���4F���-'�#���2� Ѕhs*�����g�Hr��.�g?=6J�˗
�1�xh�:�c��?�r)�ܸ$���r5b��0��:�µ�L���2j�w��[�3pA��`��W�%L�M��k\Ɍ��X�R{0�T�F��H-�[85��c'�����р�jT�OM��Û"ד�$�I�m-0s~��X�<
eL�}%��Z�g蜶�:"�(X�%��k�Q���q<�,5-���(��n,��p��,)dp�8֭�ʛO��{�	2M@�0�M;[OB�I��t2��A�A+���KE�]|t$�s���]�jM�$#Q�!���>M"�������7o��+���A/�b��4A��C1��?�V��C~�vT���~�;���`B�h׉�X�H���W��h�b��K���lO�c�[w���W6�h�rsG����+�@窭����L�g��n��ϸ,t��
h%�4�Z����'Z��G�(�vn\U0�{7�cNWk��
�Ej�hnS��u�c� :�<줺��d���A��'��z�0��`ѿ���.�#�d���ԓF(@��e���&�cs"��J��Q�%���_DZf��c ��8^�Q"�b,y^��L���DS��h�ѧ���UM��ƭ�z�t)ɯSU�DIH����u���>�V.��RL|���m����q�m"�&=w���U����O�iٍ}5Gt嬟U�?O�3ں�l�Efs�����&Qg��o�$կM����I�
�5�K��.�<#b�֏)C�������%����Ԣ�$I��2�����S��R��tn�D��r�՘��I�Y�Z���ш�j�Н�wv���r�>wv��s�;��G�/�Ď�B�G��Z�\��5�����|���\�y�н0t��u�D[�4���7r���U�٠B!T�1�b��f��I��d��y�>�n�O��w���G2$����������hk�P�a���8�>���8�����)3CCC(Զ~n߯mr'J����.z_�	;�,a0��y��8!<n0c`24�կ&�@}V%�7��7f�2��5e,�kn�P0��E��d
���P���(�n�Z��,<'��3S<Q��E"Q�eC{~i%o�8)/4"�xV��ZM�>{�5��j3��ߧ�����~$��n|��U^5��N�هJ%cy51�z�)*�^��,�`ge$%�� C�m|D���ױ���#Q�k͔'�7!]���4�"��dA0	$R�6}κ����☨�ޱ�&K�2^e�1�����9cf���R�ܸ��1��REC�c���}�=�勜�'���ŶלLK����v�޹��Ӳ�q�üĕ��~�#'���SVOf�	j�w{m�0��~oh��7Q5��|J�u�V\������~�-0۱����N��9��	�����Qsn�.�� <m�/(h���g�4��v��u�;]��?>�L윳n�4jEi:Ħq�����ay�z��핚�}0����Az�z!ʆs�-3&ì<,`m��O}t��N����~K`��̦���4�����p|�4_I;�IK�������<V�S���Vߨ��{���:x ��u�尐��~�#��Os����\e���Л�����J�y���ڦŋ�L��4�ټ�V*#y#P}v�'�гqޖx����?��D=z�O#m_Eg��l!��C�[|�#��~��������MO���da�h%/�n�uVk�k��b��%4!h'��u�PM~؍N�N�2+Ot�.0L�1U��͗�̓y�Z7��5�[����Mk"8k���*��P�n��U5+��ď�R+�+W�P�XA�?a�*��K��!R�sP�eM��y0$�� ����{	�v��c~w��?�~5�-U#�H��h�W?O���F/䠋��r����ݛ�'��5��Tr���Jh�X73��
dٽQ�	.Jer!S�$�'���wn�-��qD����ƙ2*I�r�]t�'D:��@��	�I�%ע�/�Rӝ�E}��TR93���-���b��W<V_[}��amLNv�tҾ��Md�mޟ���Vhq��y<bS��R;จ�<�2ǚ�wO�ԍZ�ax����f�� nl�in�Y�5L��\��$�~�,Ϟ����[&"P��pg��##��?ݴ�3��|���ͨ�VP.)��	�N76��{ETNҡ�?k�Ss�>nQ$��l4s��3�pᮤd��y�\�hQ��$R���M�h詍*���Y��y�G�}{?�"WY+)XK�}��D�k�`wٱ=�h�߀z�kAv��MbkN�W�9G'�{�
�ߚg��nH��X�ԎW�T�л{%�Բ]�J8��/+ڂ�1QW^Y��^��Vo�+�(N���~6B�_n52/���%)�UD>2���r�q��uUm8hi���Zs��i»B�pf����V�UW�n�Y1 =��lBbف�ΧOH����@�����{*����6��_V��-~�%[��������g�o@��Z`T���q��]�d�3��/?�@�I:2�b�Gy���o��Z��j��o­�xP.����ϔ�0��-4w��s�|�d�0�5�2qкD�m�^nQ��S�ʒ䠿��hv����6p�ԕ+߽G =[\�D'������z(oE^Sa-O�'	(�. ��y:y���ƀe쀈!6JCqج�rg��N�F�z?��L�?��o�	эQ�k�hVr��{����"��?�^���Y����e_o6������8�rg`*���4����#h=�p���U�ȁ�Qo��/R�>�g�}s�#�D�w�I؅X��A_S��4��W������c"�~\�3�ҳ���%�gOK�$��vkH�u�:I;�)����	�x�6���}Ct��U��i	�{�a��OD6�ɲG�o�t�9iЕ���� �틯*��b���m��kG�M%L��[A�c�·x��'��dǤ}�!��_�`��:��i~��;�������ٔ<|c3J�HS��*����xH+��1N�;AG|���ť%�Y+]���l�
�_�i���&�G�?�G랡|�2�P��J��(�@��țLR�3�-P��@^X�U��D�$)��IeJ�iA��C�ǭK9��2���nl�p$��%����CY�L&β�p�\�>����p̤`Y�����Hx�R	�r�_礩�H�q���pf��8ܿf$��b��sc�=d��@�?��ٹ����&T�cw�w��2[�'?�[*5.���^�qA�'?2͉�v�W���)t�S�ԁ�m�R3S}~>�8��O�����5�O�D����4�����dB�4�c�DhI �bU�?�&D�S���2��O�����$��uV�Ѐ%�5+��`�E�d�cJ��bՔ�/ߜ��$��*Ew(�>�WPl��~�P����zNhD���H儈�ʮE�B�tE�:H��2!��;8���k@��fMI2rQ�9�k4aL�J/%���+�*�����-�Э�Mz�����U[��%x�����E�I��F�<���>�;�M���Ɋ}���7�?f���XW�I4q̛7ɵ����9t"��'!����u�S/�ˇ>�u�m�O�I)_Ov7�6���J�9�M�lA8������,�+8���"W�Y`���l�Ε]��"
�w	y?�~j��s�o��u%��6.k�
k���^@���߇�f�1%d"�W[\�δ&T��q��2*�tF�o}�m�C���Y�{�;{��WOe�9�@Ĝj�K2|�lQ��\u2��S��rA�}Xֲp�^/z��Tr6�1�[�~B�E���=��^PO�߬F� X��}¡zxə��C��G�t�J��N���AW�$T���˷Q�.��CuH|����GۗQ���JF~��:�"пo�B+<���J�ca��':ܶ>â�YO�%p���C^��^�e�B=<^����4�2���(�O.�q��oJl�b`����o��m3��.E�;����冃�#Y��K㰋?E�<mJ3�1~魌H- ����o�L����pE$3K(�5��6����8�<�E���u�8!��q��
por`z~�XH�|��x%)�'��v��L�	�f���L������e�kAD������9̆͵�О��q� �QMM3xL����{����ɴ�d����:w��s�/�p�x$���w�_��u���S��撙�'p`�Yt'a��g�v{s�1^�t3
j��?�Q&�T>�n�)�
*oX����{;e�?��\�P5��k`GA��,���i���M
E<	2}�i}	p$� ��f��	`~�7D��UZ�嬫=Ã,j~:�!YG3��G$Uw͘W=�Ma�.���IƇH�/�� =��$��G.`^饑�ƞ�mQ�X*���=E �᧮	�K�L,Hx���f}��~��xj{����皷�����D�9�H�-��m��Ï蝟:C}�e"�ك���W��)�F��B�]�m��{�x��_�:��Y���{-�g>���w�r=��h���Hv���N��l?�{e�K�y�ĆRi�yVh�8�< fPr�ч��0��Pۺ��E�թ���U�x8ӽN��%�ԗ�8�rꙢ�y�K�K��*(��OsR�UjhУ�\pkdߩ�W��([W̹V�Ւi98��]~i����+&7kU�ų�r��[W�O9Qze��e����y�y��)nk76o�6lWS���Tl���-W�:ſ��M�ѳ�i�}�&b�]�r���I�"x�-e���q��ר�Y��<P�Rr�`fNx��[�
�Dq��i贉ܤ}r͋�ٟ��#_�F�h�s5��,��3\�)�z�3G�{uCi@�x�����͘C�p�C[����;�B�J܆��Q�0��z�\8e�{侬�{$���؝bi>'��(�*t�x����=��<w��^RͳGA:�+nט���>N�cfZ����wm������op�+q���d�^j��*�P��M�1z��*0�>T��5+������f������S���V�W���R�;MU浓��HX�� ���A�/��k(�/�	pˋu*�6��Ň�q���u�A��Dn�T0'�D?�Z)��y�#	RN��Z
����f� t�6k!Ԃ_��R���'X<D�>�%x�&jjUG��=C���	�F)��<]a��!�K����Z(������sx���_"i�P�^�6��>�~}A�n��H�(%��c��G&`�1ܴH[4��ݼX�EE��T�ʴ�K��WW��U-.�O�����Y��|v��(���P��X��aB{`��pEQ��["f��ƭ���gX�ɟ��]Aݑ!jJ,������?�Q�Mk��mG/�-|b6I��0��1���ŏ-`s`~l� � ��)���5����w����E0��Y#.괨�X��C��R��_p_��n��@�-��if�MD��)����
_&�L�t+?��l;�Ƹ����c���a}��g- �����Dm*��c�r��q30;���h��U��o�N�Ȳ�'bE�4$୥:���Βsv2<}��\��N�:�|���:�a�#{j�4���s����X��U.������K�;��㼟w��H�x.���1W2^r'BK�}��]הKjG~�Eh��,����(C1͢;�$�7��]�B�ȯ��b��B��q�F�q�ޤd�%]��0{����W�=?	��b�G���`!�*We�]��P@��
���3�J�&�t~G�ӣTV�P���`�~q������$�Aq(�R�s��:�nÄ S{��HA�I�iT��Q*��/��|����""�~�Wc�N�ǃI�1�A�`�_�<$�����,b��f��;�J&��˻�z��k}2٫#.:�ʹ��-3s*v��H:p��GeK����b��?R�a�?eV^Y���rY�q~]-gg8xfE�V���+�˫%�Oud�Ծ��l��͗ý�-�λ�X�ʉ�Pˤ�ǵ�&%���֖�&�q^�w[nߝ�A�ѕ��x��NYU$��X�2>�N	123⥦��^b�%_A��6a��*a�2�TL`T+���1��8�95�>۶RW`��(Ʃ�z�8�HE�3�GQ4XV��XT����5�$z�ToT$$r�XX*���v�44�?��2��Q4��+8�{'�P5r�B|���/*U<D�罫�>��F��.�N�_��`Q��Dm!��Jr��[�Jw�I2[�i��o��<�>�� bıO�A-������J�����i����F1�9S�:��'�li�a>��Ndi9�AF��Q�[H����ƌ���r.���>�A^��L��l�p��Ǌ�=e�-���/׍�4��9}PZ
�]��v}C64��.v=V+��dI`릔L����$�ǈ��f�T-��M\X���{����v�cr�����mh%�Um[=��s�^�3n�+bN��P1���<��hbPYAP���/��>6�N��kxk����x���M�z؆^J�V�]6wH�/��Bk���.z1�la�W͛{��rT��BmYPZb�[�{bq�'�T�7g�W{)�J�+���4�^�D��.����LCEWV���<xr���'p����Sp[��D�k~��uw� 4������7�.��%������a���%q��&Ӧӏ���$��՚��i�:�n�(6w'�"rQ(;�Xb�-�C�/���ɵߊ*��(<���$�-��k%Q:�	»��֍ynJS�:6N�ܫ1s�v���Ԓ.e�0S�~�d~qh'$�ۜԨ�y;{����,��J�����;Uk���6� z
�8�]ɔ�S�dDi�h	�ø��󱶾�6QF˼�W|G/�[eC�\.O{�J>����K=8&��{>Ә�C��i��E}�៾��K��˺�KFF�{����~b�XuF1��)�k�a��.������3��6�����/�r�����u�h%��`g��`_Ͷ٤la�u�~�䙨��G�$n��B�޻p[9,�VDA��؂lʖ x��S+��)�W�"�pf ��qO���D6L�vÉʙ<�oiW��8T�yST��x�r��2!<�ػ��B�c鹕����U���I,�J,'�����.!E@��"J�	V�"�v!���eӮ����Ԑ�s�f��<�̐~����N�l�wB+�)���*�vte�X��M�d� �w�I�n����R��~�ŸЦ�av����/mopG7����Z���/rR<��?�5��ƒ�s��u�l��7�V(�7<ͳ��u��K��F��I��oǰ�b����7��);�73[D�rk�={?�`�gs���Fߏ|(�/[N^��߫ۺ'.k =kZ~P�9 jDu���Ē���SYf3�����O�y�J΄Z���54Xv�u�V���$��훕 x�͊/��ʫX7�a��I�9@��`���Kؼ�u5- +���$�$�_�W')��b1��%��ԂT�[�Wޝl<	���Y;.�:�Z�[�sz����4:9�;�_�m��u<�#��ԋS�]��G঎Z����g|4.����8�������Y�Ȅsp���fl�7[I��'��|e6~÷���q7���U]bb{4`�8Z�?��MT��ݢ�g�)��8u�Z��D*IC[g�F�n��o����!�-*%*-������b�x��S���={�C"�Cꍛg�-5���!�o�5#%"�x^���M�Jy��T�����5/DA/L�C� Aa��Zn�R�2�����_��8� ����鰗;EN����-�����u����%��#Bk��+hN���k�f�h�&ْ�Pf�ç͊�NdoR����q�D��&�hW`�?��slM����:ӣI�s��(�7]Zf۫���J��{��<^��F1�L����ѝt�����ε����e��O��1��L��2�m��r��H��h(̛����_��S3��_�Z�1{���ê
�J��ޕ1�z����]�I�X�i �XY�ݏ�y�'��
��������O��	A'��N��E ��vz?!P:0�W7�}���Arg��@+��J0��=6���<	�G��<*h�.�1�.�|ύJ�S����(q��V�G��}*JbL��^h���N \K~[�1��Е�DT^ѝse�r��S�*l���&��۬a��X���x�1�G��s ؑn���z7k�!FX��>���4o"��Mo�Q6cEj�H$�nl�ߒ����ą 5G�Y�$�y�W���d��g�,c�S��)�����eA�����߾����ui�yV��r���^�t~�.R?yg]�e$�7��I@�6��.��������Y��yp����Ϡ�ٜ6+^�~F��j��2�HV�(� �kt � �bkyEr��������ڰ��p��>I�DgX-N�O[��)N8Ӂ��s��/J�Mq����T�p%{�n%W��c%@����������M�cQL@���]��p�n�5�ԨI��x!M��	ǆ����� ��Qq��l�;y�0�a�y�0|þt�.�R�\7.B-��r^�t�+^1d)�.��2�x��QF��]���ZZD��P�#�:��(De�ƪ��G ����.�bǹ	J=�(o���j����L��މ�;/��<Qް����#HS����%���7`�&N�ڂ��c�|۟(/%�vk�K� ��6������t.�l~�r�����Wo�<`?A��@a_9�_��}�+/�FY<Z-+H�-��iG%�`��鏙R��X�s�ҡQ�t�/+�.7~u�l�WUF�3�_e'/�^Y��=�za�vз�z��a[�W?[]BZ�̫��FC�a��rt�-�r@��:-��Y���d��� �;d����`��t|���g��q�%=�.�7����o
]m<?��Z�aj���,���`��ޠ8�l	��
%�${��,��,� ߄([Y�c����XcCT7|�+:$ݓK*�TT�$*-�[���/¦���ю:[����_�-�V�2��t�Ne_��6y�������*BңE<]l
?n=D��^�$-�����N�ޢ4���g�=	/>#na�˝g;C8�
�/�iE���R
n"�{]�Fn"6�6։.����*L�`�k�/���'��|K�E��hp� S2x4Z��l���H���"f�h��*�a��D"`sܠ���U ]P�ḅ�d�X~�4�<��a�����iA#C�A�:{:#P]�능��1k��1�M'��7�u}�\�β]�c>=�ˍm�}�X��?�7��J�U�(�Q���\���R6�[�#��e�o���.K�u�N�(�ş�}�$���og@,SDͪ�`j%?�AU���Z1���YgW�ձ�&A�)��ņ�v�$A�$C���;��8�4�6��@���^�b��6��?r�=��I�'t��Ђ_hyp*���:Pq�C0�M`�-B�1�0���9�г�D��N��IPS� X�����%�0���5<���p����vnfz�����l3����� ށ�ߦ��a�����k��߫.
bں�5�#��d/]�I2�7�,:id!�1{��]�0R1��3q�Y(�i�3t�{o�ƿ�:��0y�e�_��*�];���v�'�G��d�&䉊rT��0��,�����2>��}a�����!��6�EM���^�@
]d�dw�FX=!mH�l u���:���Q'��o�^���."��c׆���,mx��2A��m���'�`PxK��7S�F)f�ع!�V�{�	Zi� �%�ˤ��dg� R3N&�"|�f��T��� ��k0n�[��$,��;� ������l�0��|��L �$d�};�jEv ������� k���]�v�ʟ��	��H�\�ܟ;����,N0�
��/�('NR����fq�*!��,�e �i�/?Ib*�E������E��ҡ�@L���d�鮯����;�.��}(~����F��w,���d��_�,pƺV�s�Q=�l����j�pO��v�����O����c���#�࿹.���=���<a�Gi����}B�����!�E2w�Hv=,�!
��,�Nz'ݤ`m|V)T�b#�j�g��N�����N����x����,�j��yZ�y���Y�{�*�)�x��i�	�gQk355�%{�Nx]������k�v︹G�� �������53�����t��%�3����E^`Z�E�_�q�'[yR�W��h�
͔�Y6�U�zΨ4��]��Dr��c��8��(/�UBl<Ô��<���{>��?�Q5��7>�{YZ)�*�����隩�}|�����O�b����Ы֍Hƛ2+	�$�D��-h�#��.�A���x�޽(r N*x4��n��6b�\B?͎D.���f�Ub�yS�F������b�>��+b�L�Em�"���i��JH��2��S��ϱ�^�oϴA��K�i�@?�����|Z�Ay�߰bihA�Ռ_��wS���
��+�^1��#�����A&�Y�>��Z&�\�VIhH�p+i��'��O�*@���qý�Ru��^p���)�����aMf�5��ҞI�	�+��)���٤|���kVO�3�]@g���p�m���� h��@��\�&��]��ْ]�	 t�o8���a�W^0�<\t�KR�(����T�˕)��z�pI
�ڹZ���66��G�1G>����b�k�gf�$���;>&7�,.x �#��p��Uz&�ftgU:�ӎ���S��c���`)��U�I�_�����Wa;~�ݽZ\hm������l���Z�Ʉ�yE���Yu`�;t�}��zd\x��W�m��{;qha�[���63�$x�� ��� )v��#�᭕f	�6{RCv-��D���&Z^��f&�W>�z������J;'P�7B����n��Z��ev��#��_;I�Tq�{�v䴍 ��ޖu�W��xS"����z�m&��L���6}��t�7c;k=1�M��ω 3y�9�{T�^*֏��;���E���|t��{� �D�����]�1b㾹H�0� �p��]���D��a��C�:��
IE8d���(C����4=��F�����^��b���g6d��s��D�X6�d_|�{����-xjd���N�s�R���\A�X��L���w/�/o�GeZQ(�6V,�������؅�Q2B�W�_}BE� v͘���4Hv���5dje�ڐR���G��<�)�w��V�W������{o�岽�2���߃ݞ:Lr��?s��t4��S���;ܝύ���h��)��џ7��Q�׮���eF�W��Z�h���5?۫�M�((P=����3XE�Y�D������x�i����zs�bsS����/�Z��W�����k̖������d&����e�|l��ꞡ��T�OO˲?j��Jz��x��<�Y�E}�����ވcCI�Aܨ~
z;�r-����MP'������slvk{!��/
�}�iX��S��~��`kƦP�_�l��v+�k��ꊝ�2��vO�*��hdd���k�ꬺ-�"�9P�JEEZ�ȋ��r��cm�\nEo�=�;	�����c�􆥿a�@�0P�}&�]po
�� 7�L;�L;�H#�@�	߰Xx�iH����4m�BU�ݢ`�^��V�����N��q�as)3�[yR��Y��g��A�D�Fp����B��j����.�i�V\��{�iJ�]����5|�]>h�dx��D���|�8r6�&�S�k]K:��v�Ͳc6���&<�SB_���8w����3h��W�8�k���q�v'�xܨW��n�e��D:�[�Q�D��3�
Цk��?z4�B9�@܉�\	r3z]|��o�r�+!�_;�ˊ�E⼞X7��#�VR��G[%� ����Y�%l��%^�|�[���Ni�8&v}R>����I��A:��������.�8y�[��H)������{�v7���w:27;[Xl����jyI���~H����s���_s:�M�k�z-`�r6��-�~�'����׎���2}���ߗ�]�@��+�Ù�����]!�z�� ���1�q�/�}4�gN�����J�/>�أ�(_���m��h��ѥ�[dC�d������%?�Ą���ZU���DFqq=�� ;���-���>&�I��[���;ſX%�fUЎ3.�	
2�b��u�,}0L� ��% �U 2���]j��XPr�z�Ft�����7�i]A}���L�K�/��"��I�}�����P#k����n	��{�Ȋ��".����q��j2M߃W]�����ٔ��Of'�G��~ø^>�������5��3�"+�ڒnsn(�-���=�$�ȖF��"����X\,��������C27��r��<,����Ե���T̽�$�b�q� ��C#�EI��n��m���[Dw�,��񷺻�8��s���������۩����l�n	>�;Zӟ[�{��.�*YVqIhA�>�ٌ�( ̼Q�?�h��f�7�ʆ`o`%��Jh�4��e�z�*�Y��y`�,Dp/-�X;o@�u�S�ҧMO���Ieg���,[��Q*.���ge�ۉe�8@�͙k��sd��� Ϗ�|�x���߅8ڗs߄9�u�?�n����o�x��}Urc�Nͩ���'�;͡���\��^.�}��k�
���}��-X⬏D>��^}R1�D�vF?��V��H����ӂ�z�ݍ�{����E�'��9�l�EG�D�̂���N�T�J��BT��U��4:
J�_{5Ի;ػw�"�z� u{=LS�t�G��b�����dp�����֙�R�Nj ��6�}��� ���@��L���,���Nq���v2�f�D�h�Ug��S�G�,س��[��U�G�c��Td֫d��-�T�];D�ץ�dw(~���b�UicG�K0E=���ÇD<M���f��� �cvtq0��cO~+�!E6�˷;��S�\���V�U��U��^��~`��<�.�1L�&&'h����ޣ��|\���U�1�P��Ł|�����0�~AI���b� ���Pj�a��$�_��Z�0N���mV�O(9.���y(o��i\/�����������bB_���dV
�G����"�ҠB�1��;�'/a�}��^�2�
Ҫ@�[�����dC�ݒ�@>�ef��&a�Z�Շ6��t���xr�s��ׯ�~���տ�Ö����2?w&o�[��a������H����\=�f�q_9�>0Xі�/&�'�&��q;_�ff�����v|��D���Xɱ�h����#^"��РN0���;�H�.�K�Z(\�l����m�y8%���F�v�M/"��	v�B��U��682+����,Ú~��O�d��h�Vztw�pHw3���(����h�I��-���I�?|�������c��u��}_�y]]t��ϧ�xk�},y�Rtf���O�̙�!͒�����cD�婳t�y�~����#H�O�;�uG��)�|� X��;��y��'&�"�+d���y�G`揼��%��������t�#Ԝ���j?$7�P=�����K5 ����о�k�����g*�6�LD1��<w>��f8C���:�ٷ��ݸy'�)զw��U�Ytc��:��F�(!\�Q��/�w���D�-+~�ߦu?RY2���>>�P�� �_D!�	����/�8����_�p	�(02*��]9*u�s�^�%�bjN_DQ�P���A��>
��ʪ�͊�Ww�(���rI�5]I�k���֛�5�����ź�F�����]X�JF؟��&e�QF�ot����Y�Fv vQk�)WjF�کS/�R_�&���o��
ʩ�������c��+pۖ��qӛ��b�zF�hbr��轣�~j�.T_�P}3��W4����[4q%h�4�����3�0�Qj/��ξ!���np��t��!�H�F�|yP�ք��Fp?k�O�����e��%�/r��r��P`J���5����*7��D0[îdW��D�s�6)]���T_݌a��>�����-\�����rl����fz?�_.6�����i�%r�����n����W=���oMh�uHX_ذ���*�6��N�WT�d��Ԁ�:T� �!#(Dg	ὐ^���gN�pR���Ls2�ڬ��S
���+����i��<A3>���clX�AM��Od�>����9d��F����pG��l/fƦK�ڝ1g�
����zz��:O�h-R�f�D�li����~��V�.��W����E��-/aC���x���V�*=�8�B~�#L
m'R�<����t���Y�dV�Z�GTo�fwvZJal�E��ٓ��Dũ��`Q�4G���|�G�_)�QT܄Jw��!}�&�R<T^ǇQ�}g�p�帎�S�]�(��wPfBڹC���� !�����D3��{����T(&�K|���j��,M�)~�Ɏ�}���|���<£���v������+�l�J�w8N��Ǘ-*ϝ��e�?|-`�NC�FY�i��F��3�,6MHC�����e�����>X��eq�k�0���B�O3�N�B�Ш��gp]�
����C+h�q�<�f����}:ҵ�9g�h�"�{gۏ{~�B ~
o�q��3Yö6�0� �e1_��:�OP��(��Y��5ܹ�QE"��K�����D�X䟸���L�8wd4��8�-�3�tЪ���+�^�c��4Ӭ8�p��i�h_���&���u�9%3з��j�PY�2��vFrV��Vb���г�Ce�ߌ����5��5 ����1�BA����}Էٜ"�Wh�u$�s���7X;L]\�kd1x��Z�:�׷�ute�Nkhޚ[1��w�(^;���Ǿ�t��8��2�tYK�j/��y^-G2:3I�?��q�p�90g���D�QV�vJ����-4j@�8ږuo�;�KVap���M6���G��l�i�����C�֛߆�����N	����[n�OU7��0��_���
{r0/*�-�����n�5��S�C1Me���Bvl��c�/U!�5*�oU��>������ү��	j�7�t�eݿr�:��]_O')��K��rF�Ͱ�d��]��idp*i�\�izl8μ�~ɑ��7,L����e�� 4'(Dgm��W�B�OM���&��s���������լ�&[���'ԭ��ʹpB��M6�3ݢr���Bfޔ#'d��{�O��/��־~Y�q$�;p�n��y��\�����w���ܒ��?�x൝��a����-�b'!������.���k�*iՀu��� ��3�D<�]����b��Ԃ��RߩR��!JQb �٠, �'G-iE��EJ�2(�*��Y�P�@o��N�p���@`B�_����W�[3p�P���^n0|%��acN#]s�v)2�'ؐ���$�N4^�[�U��{Է�ƴ��:.�����4_����mB��Fq��t^��6`�}�t �ڂG�V*�]O6B�x����C��n�	�#9i_�c>M�����m�ۜQ����*¡$����ك ��Pf ��,uJ�$��/0����?_�|vl�U�����3!�� ш�O(�ˢ�9��I��{P��聝��i�_L���羦�Hdgeu�"?�d�?(�-��a��CG��oH�,�����f��j��RjC2���l����_4�kqs�;�8?T�������D}
NT)����p�h7�j7ػ�h�/-<ًUO/��;�9�C\�|?���Z�������s�:�B�*,9A�t�]�Ϭ�:��'��~�¹ �N,b��/4)ʏ�yx_V��*�w�i;F���2��o�rU󽳧k�ŵ�R��3'6����D؁��E��q�J��X��	D�M�������;7ҟW5����PK�[�0y%�M?�i���ۻ/�L�D���ÙyO���0��hfL�{_Jz y���JP&���C�+K�0�+H�;g[�c�*^����˙���J��saCf7VN��5�2��0B��|����L)��7�SR�l�T�ɦr���=Ċ�tt���$M�=:�s���i�>�(��ኖ�53��iӒ��_�˜��s���2?�w���d��LK�=m��W�C��u� �d�),����'p�G�y��`҂Ir���̱�S���tN�h����=��C׫��8i~'��w�#f�<*S�^���ߣ��1>�"���kHn��;6�F����]j��5���h�]����6��0_h�9W�.@ׂr�Y��U�&G�%�U̯��1��<�[h?oV����Un���g:�}zW2c�A_+Jg�z}XK{S�z�-ys��zߥ{�rs���z�s>{��QmЮE�T�&l�)�����7�~��A��mI�a ��p�"S,�T�S�oi �jf���כXO���0}����W�P��Q�����~����
�G�J^�J��g���������z�Wބa�zC����|�r9c3�	�h������>{F��`&�ob܄�I�Kпb�}���yqi�iK*o����PE��:��Q��e:�R�ӆcPG䠏��V�[CI�ITX��6_�<�m�Vn���}HYHE�΢���n���fgY��{;��������_���iy�﹃�~�[���|�����+]�M��\�`��kdohϖ�Y���?n�5+^msQ�Aذs"���gb�Rٳ��vo��
mz�x̌D�f��r�X�vu05�|aej:��C?�`0% �5��94��$?�G.X
]����+�N'D�9�P�z����W��	�ӼB�z�E�����%�Ȋk��3���'���X'^3^�t�$���"�%;o�ͮdC@��7��~�ը��.�������Tp����0�3��DO��b5�śz>K"���#m-Eq*��
��,��"􄔶��]*~&>��t�)��� �A|A��]K�V��N�!��B��|����>��k������EN�m�,-��Y��ҠO-â@ߒ,N3�@�u����zf��%�%_İ�o�ʲh��A�x�Bw�M��#g���G��c��� %�w��q4;��D���z1�1�YW9b�5PU���f�k/��v�M��]��An��j���$�q���q��tD�2���V��[x?~�iɘ=}�@Zs�< � ]�1��-/��F�4."W��h�`X���d|��Y�(�C��H��[��?\ЬUP�tZ(���xw��CQXQ��%��9�@\t|1C��+"��|�[8�Z�0?�{�zn��g
�פ��$'� �3���w�0����]�Qsy�o������[]��,3�ڏ◜ͶZ�Ph1�½�0�����w���$!��$���a�UQ+��b�0���b���U��X��c'��i�!6���!/5�pDI���L�c����r��d�8s���C�o3W�ZU�n"i��P�P�6TyG@�3���<�*2Yݡ�ݻp�I��Gw8pZ�a�=���+;�������uR[����!D�
���&*4z������_�q��"���j8�� Pm��Mn@����:��]1��Nd�gY���U�DO����ך��b}A�̯��d�?��!�g�b���'����D�� E�e�(�l�ʃ͍�Z���IG2�q���%��+OM��:P����x��V�/�euG�~�>3�F�"����T'\��^��?f�%����T�m{v�o �)5���C��M��T@�Q]��w��kX�W�l�1�
�B�+������_���r�7{4�ڐ��]��j�_䢺��'�6�nO�~�_��y��Uy�]����^V�������n5�d�s��/φ��E��i�~ꦬ�Y�� 7P	Yw�;��':��hHR	N
��yӻd�2R��<�op���S�1��!Y����������5����)�Y����B��AD�~��M$\�>ȭ�U�Vq�g�3m�3ʐO�	V�~G��V>������^�˘1���O��W;��$a*�����?~Iqb�q��u���1�j��-�i\9����`����Q��X��t��<�D<䵃m���3���H>�B�y\/5P8��%
˂_j�㦆��ç��×��t����-Ak��A����7�}�6�$��@�p��6#�X�y�E����A1����-;R��?a`On�Ae�l��l�U<fr\�w�P����bl>��,�H���e,J�$�c�9o�l#Mt#��2�7�N���W�����v������ِ�u�����Y�����&����*��PK|K���XG���|6´ft0SK�{��!���-øU��Yi~m��vL@����_��M��e��^�ԪT�
�\hiCdiCϱ�e�s
���j�)G�Gsh%�v7��X��Dytս��ZFk�}�����C�D�Q#΀�VC� ��fx�������_[��*aI ��Ս��:$����Bii��|�N���c�����af�OT�*d��ЎQ$�X��0`.h�� p5�-�GI���0j�	�2G�<������>�&΋U��c��]ܷ f��`����]���@�m�t��9�ˢ�T�'�{a��E���l�9����}��mlru�?b���ÜM=�������2�{�Qbz^��f��s�I��ق�����3ۊ�#�(���l�ц���
 �I�N=��g>O�^M7�#j�w�����BLBp�
�%r�# _�ж�b1'Ěb�o���|&��U�N���;���*g*?#��N)	�� ����$5����ƨ�)8��m�~�|�K	��dd�x��Q�Yd���B����"��#?%L�O�sUe	� ��^Kz�-�(�}�o�������<?�6�9{!��?t�*"�0S������0a��hȱ��ԀY�᰷��Gs<'����{� y��9h��>��e�y��~4W|�G�����s�R�Gc�:�ւ%,�� >i���~�,`_��t����eS���nm}if�,�s��M+iO�j�ǝj����~Xxx24���=7�&��ٌf��e	�)ž�
������J[/S��˃����93�\��r5���qW����2"�F>^=6��/��4n�$�\���b]���t����y�/��8����TW�M=��ߺ�u�
�m��a��D�Y�F�]�F��U�d��:�U���*�+9��qsPu�D���������D��7���j�u>������NK���Ɖ=�F�F���n"��Ɂ��q+������0��H�A+�I[�)�jؗ�vi�E9
��C�3�����54���0Gi���J�
�G�,f��<z�N^8i��%g�5�{�7�\oW����f�\&����6m:��k9\�l=��e�v3TZy����>%%����C��Xݤ����^����
��3!��Q���*�{xi�������c�/�E��+G(�ur��mI��7�h/=łEH��w�a,bb��S7`&�ʽ�����Π�y��Tѣ�w2������e+	�� ����~XG�@�\&]�oU�ģ�]'�O�d'�J�魶<8�t�Z ���I�g����)F�g��e�	B����
+|E�iW �k9(�&�VrE+�z����c>���F�w֏����|��z���m�`���F��xe�~#�:r?�=3��R�ij�EL�j����i�儤>�A\ WS���E�%�=C��}��9b�P�2�*���J�&/"e�Ý��
�9E�`˳+{3���'~v��=�H��'j�sS	���a��z$3��6zʜ������$bN�4c?���c2��^������P�1�43�N��꾚�*��7`�MT�����S��č�vwm�"{�O��zE���Nc�Py6�� o���ɞ[���fx5��f/�	�
7Z�:�nn�Z��r��SF�2}� ��#c�ݖL�Ms��"A�<��e>c�/s�_��R��<jg{���R���P�����k��b��8�����s��h��q$Y�t�t�����>�v��Jfڧ!�\��h�d�r�Lp�#��G�F����q�r�'�v_h�zM�=J;d��/����߯��a�5v4�3�P�Q
L�G��#��I�����D~�`�4�����v�Q_)@�!{,g'�M�!޵~K����>Y����W,�j��^u��^�us/�8�T�&���΁ќ�1M�M�2x*/5�_����߳XѦU�r+[7o��N�bt
�i#O�%�bgv�1Xh?I� ,j��j���ʱ��o���:���d�������	%���wzld29|t|!l~�&{��U9��@w��6�,�	��e�Ɓ�s�RD	p��O�>0�[曗�[��"��� dc��i����d��]��>^�;jt	�,MsY029�����ϵ�ՒO⠩k�O��l�p�-L��C��������Cu�H����=�Z�N�xMG��"Y��Ơ����Z�5�A�t��ѕȸ=zP�+k�Ag�,�煶-�wu%S�w���Y.��0��u�.�Ub�9����a�c�`.݁�)\Bִ��!��������5sX#�'��"���2~&;L�����)���Ҫ�5��߯y)�s��D�V���yP" xs���:(mH�0��-*�ar�R��*��P;����hZDw���zM`z}I`z?C���xߝQk��{�>۬:nw��қ���!���1)���f����?�@-7���6>uԯ����t��T7��J*���|���q��i W�QL���O|��e�_�&J�5K��l�q��6jY�Q�D�\�ބW�A�}^�~��(-:�Ƴi��LC|Hs�N�[��ό�xY��̗��?l��l5g���/�����VC�I�}`�<?N�k{~VjdWtXl��u3�L�d�s;�w����Dq�G	�85�M��[y3�AO��!r��O�(*!k����q�A|'G��!�SLUz5%1j��N�l�޻���^2�����xp���,RX���K~�J<��5yJ-ka�I�2"7�Q���Sp� eR�t/~�?��A�+�y��N�L�&k��̵���6"�%�+�Eڰ�(�o<՗ݱ$)�8�D3���̙��E2�O�&��3�ߛU�U��Aë������il�j	"���kb`Cٹ�D:��֛���%���|lݑ��̀�cT����@�QB�8d_:4��f����@\hփ��(�
���s7�8,�F��f�gBeS�>I�hY\����])�jCgF������K�>{`����N6�;�0��U�;_�Ǜ��u��Ἆ%Mxd[0���,P�[�C�\-�6�Y/FGN\u��TҎ�i��&���k��SԊsE���LZy������v>�Y�vvc.ݘ�n�̦�^%����RA�F����/<QO�%�Gw�/�M�ٹ����lp�޿�1��>���Tƍ��Q�,��<n�����4 ����L3�^�B�]Z��-�L�
q�o�*�/8�D����faP��	N�v�N��z��_�]PF���7�/U���,�[0�.~�6��Ea��x��lN����,6�n�<�4�6�2�6��.����ҁ��<��0��yb��v����	��|����q0ɼ$�����!�v��y�Xa�ˊ_����1�.���M&����e㉩Jb*��m���ڄ�Wg��EΓd]�ͰH|
����r��~II�!me�A��6V�(޴��_�<�Z	��J���ϥ�<�&�Uɛ��rm�Ӟ�!�#XF~�Lvx�?�G�A�pٍ���gr%If*B� ����I��+?8���%Y�j7�а!���fdDop�o���0����L]��q��v7�}8~��V�5�_��������z���e����K�v�Uc��dCe��0�@7����zB+hd�����X��d�xs����9��l@]|��IG6��tJ�8飹(��ċ�=����{�m�IO��i�>iv �#ڨ����5	$6h�ɓ(�$�Q��f܊�|y(��X^m( �	F�-��>���Ϝ=z_��sBti?��[�G�������'/�'��(� �=���{��J2;���9� �#;_IO�c-T�zOK@��<N��w4 �Y�)�o�p�\��5m�������ؓ�U��7�ع��5'�-J��>e�cz��N�i.7�;XH�����sLh�a���C��N�Y��/�ѩ������YtJ0�lC� ����(����U�	=5���21U�y����`<����PYK@��l��l�֕�p��Ѣ�
Ա�,:S���S���E� ���1�O%�{@���:��a�}�����<*�=����W՛ �ϕPFz#Es����O��g}|<�
L5��4\ow��O��!6]\ԍM�[����B�,J��o���DQ�����j!�h �H��ж��߿QME�Y��D�	�[DF��.܀5z`
!���|�4�uV~�څn��{\ę��ꡕ���.��H*@�.�jr�6���6޲�+������N���N'�fdd�嵠2:kc��L,�N"��S�
m�0�<�3X�)�5�{#��� �~0�pO~��|?k1l�Z��bi�I&ZZ8ݿ��S�U�7�i	�ߺ[����N/�(]��fL���:�g�\kh:���c��+)��?4!o�����l�*~���O\K��u���&�6O�Ibs+�xt^�M�G�p�=�RJ+�L��
mzMԀ4%���i:ΗU ܊�R��%����^"?ˋ�|�ҎҐ2���z��kO"˲���r��B��=܋v�~dj��h� R�֡�R�ٻ��~���g�~�%�j�<�hd1��д�,��Yb�q������I���E�{$N
�r�=���ƪ�
�2[�C����!d9�SQ��ot���^��>,��VL,r�\8G�������øb5��Z7U�i}�N(]��J�|��P0�7#�|ۋ[����gJ�Q�����/���#0��Y��>�i��e�7t���^�i�?)�mS��?��{�W������P̔_�`��Ba��)&~�g+�Y:b�Τe���{'���ڌ4
�^r������݌�_�ޞ�^�s����u�lΕ��j�r�j�A�-���I��=_��_j{q]��+��_q��F��"� �HUpc��J�y��^�)��i�d�ITG+>��ѡڹ���e��6��O�V����P�N'7N.�:z�B�0~a�����;d�����O-[ȏߠ�c9X_DQ�+���(��L�O�_P�m�D����������>��������(h�i-�
a�'�&k��۞���떖G�ȿ�+hg����c�x�t	`���k�*Z	w��?�	�x��ּ\qt��'� �!|�r�����k	|�����9O�r�H6	�z��uv����	Ҿ�L�3�Tf{0��<��!� 0�	Ŵ$��\^�x|���q,懑}s�c8`.he,A� �Ąw<4���#����`Az�_Jа���J�_,�Rd{�W�-W�̚_�%���M��sG��7�:�w	�VM� v�V���|PM%jV����3�(0e`��!���T�t$.�	��<��|��e�x���oWEY��8�W
����9cpF�v����ȯ�&�l$J�����I]�pЩ���cìj��|�7|mH���͓��e�L��?f�K�R�0�.�!��N`+�2�8w��\�_G��=�-�r{~����\�\���
��c�,j�)䄱��K�&�LѓxP�e}f�/����0��S��x����)�nsLE|���0/�u��W���<
/<���*��!�쏙��X~h��mƍ��xU�o�<-�ԇ�2��g���!�����.&og��o��ɖ�D�'��s�~4C�oE�����%9�P�B�s�.����mM�ɿ�5��N�&�R�4:A۳ӢޛtƩ�i�K��Gki�S�
� ����n��\X��Y���?��j��v�� [^�����`9B19����&Ͳ��QM� ��&�'��tWfx�?y�����|ły�dѧ�v�<1�$5S)��}&B̉ȜG-���)=���p����Rл�]I߿S����������=K>'ɢs͞��Z&��=���?g��V��:�2����>��.^��A��)�/�ûHL�H:�������������SN�ʴ6u{�!��"��K��v#b�U��I3��V�W�J_�r���y�o]o�[�>������<e ���\{�dƥ��u!�@6�H�g${��e��.��i䃚�dGo��_�N�ʗ&a���`Pw��8�R���A�5�4��!�nՊa��a]���>� �ó��ߗM�Ƌ@X��%c,��֒�k�����l�wa�=�b��^��-]˽��\|��@��^��U�ݩw�]nm���������ee'�����D�.����i����j��Aέ�㛯)?�Fe�P�ojtE�����0��)f�@�BK~����X��f��D=	o���8LvK�TD������'n�+�J�&
�Vq��Wܛ{H����bI-����jP/l���h�4���pf��KX�a�)]���u��� ]+K�J��:	���}�G�@ar;�F�5Ţ��_e����`�å��e��"kCZ`����KUѡ-�M��v0#�5{��xZq���c<���W�f����t1��I��i���9�9?E^t�_�鉓%iL�0⚉��5���45ċ��ԅ��Pm��sG�ӵ�^1W��e8ö>���-]<(f$ϓ��M��c0�UC�4�ME���W=-�_ڃ�͵I�*8�2���J���,n�/�P��.��d���%&���k�?����Z���|�(��ً��@� �E#�:��*��WI�M]L�p�R�9�鈧���	l���]�g�jM����`����F'���$��B�Q��~��c�I����!��[�M�2#����Ā�qU{P�c��X��|���=�f0CXJ��Ձ�m��$�m�w*.#Cƺ���N�%p�P��s׫2W�}�rV�8��%~��t��!��b�b̟)4�賜}���S�� �W�d%�/�ò�HO�+ ���*�+��(���v7,\;��?�^��4�¢������	�u�j��ufa4,���O�N]�!N����9��2W��m� ϒ��yՄ��n��(��M��S�?Fj�tD�����E��2c������Xź��ܩ�S�2�'�e�o����7s�������]�k$B�TTWN�0%�ͤxw�P������SV�5��B��5V&���Z�A+%zj���1�E�vMu�e�kk냦�r
����k��y���/��w����;wЫH����������̭���s_�������)�I ���[�?�:	?Dw��YyH�ԇ��۱��������yp���\j=�7�K�<w���ט�;�
�
"A'=5�t����Ga��By����j^��T$ �<s�$V�rC�Ji�|)	��TGB��g�/��Ś�u;Ǉi{���{���t%�GK����參no�_��c]�l�.Vi�VE]�VL42���K{�?���Ff�.��Q��;�&Q��A��,����{�VP�C�6�Z�S~�ƊY�9��2)����y��ûb���1)_䔶�Ԇn�{�Q5ٌ���uR&� �?����\�Oo�FH6�������Ĭ���J�3�3�DAԝ>���!��T7.S�®^���I pѳ�{]� ��.�g�Ã����i�S1�j��U®b�&G�XDz����ٜ��tᯟ F����)dH*b����:��Iㇹ	Y�X�Z��j�ų;]�����ӥ�C��c]��	��֛�����K]�����y��W��o�~�St�����@0�+#����ű$d�Lej�u[)B���Qn��M�y�%�SebK9ӥ��<m��yم��<*�m���ن�ApH/(��)�wzQF�]�M��ϽU���'3|�lh�ކ�&\��/�m׌�E���Y�i�)So�wc��kL2��i��N��;����9w=�c�uH�?��>L��_�%!?x����5����(Y3Vֶ��vM!P�uf���7Hq��ád#*�Ã9����96L�>���'�|�c(��poU|��蔞�Ȁ�|OGB'9z`�E�p7��E�(�]�s����NgD|�N'G���Db0���}Zj!@V�I��8��3b'^3�\����/����'~#ڐ�Ծ����}�w%�_A���p�ly�e*��$���� ��I�������91~l�����;���[/Э ���/V}%�7���y Z�:Y�^0�jP�{��8�lBq�� �d�T����L�;�#�|$sl����2������Ԧ�O���F���;��c��s�ۋ���?��>쾪15t��^t.�m��	/����� ����)*ZM����425��D>亸ݟ�ǹ�M[��7�..�J;s�����w�!C�]��������N��3�;}��<�Xe�Fi�K���j6� dq�ؕ�Х�1wq�ل�O�Q,�d��q���cW��d��,�1Y=֑]����J�F	�_�dZ�����
	�@�-��Eo[MΣ���,��Um֒ď���6PA\+^>B׍�(��ꐛ��<�D�F�u
�u�}V㽫�e��߷�M�S��^6�[͑9,�>���Y����n�*�j�2���s*n����X�<��>h:�]���pG�|��)}UU.�g�㵔T���z>�l�./|�%���|�}�e*��d�z�9�#�s�xŖ�7U�)�#awXR/:�����ypi2�H�p�Nx�[��m���GK���#D�C%�n�t�۞�"��VRO#/�c�Bٱ:6j'��ʱ��{���zygq.�s�i����/r(9g=����&����	G�33�k ��4�U�X��9��w�R�B�^8/i�v�8�P~({j�e���y'��i0ft��Fz5�"S�DZx3��Q3�g^W���֕��s-E}�x�k�����T�Ԩ���堫�Z�/��w-c����.I��4%���?�L F��Ӄ�o����u(ƨ��\�k�Z�U��A�H�^��BxH�wm~|�+�w��} �P�(�>θs��%�����![z��U�oں����}�7̭e��C�Wj\=��UX�!,�\��x��f�x˶a��h�d��w����L!�x#~��O��?/�U��&s?�ح9��{v'��8M��^��_or���.���\^O�wu�d���7����,�2^�Hn�t�+��U�<Н����7t~'|�����. ��J'R�M3���Z��(:?E�F[s�'�����xcCs��J����$�W�~t=
YFJ)]Uc��&Jګ�Ɛ~���)*�EA���3a[��Pq��<�Irހ}�Y�ڧ��|+t�[��e2 c�m��ߓ>��43��j�iU���W
��Vj������?��~&yES�2�+��:�Y�z��\���u
�d�\o�.�����Q�����~_d���e$U
A�8��Z�ΕʈRZ�H���߾&v�}�؎��Q��lFzO`��ik_͢�.^l���0}f:���*B#~�C���x�@Z������Ɲ�_�E�vݐ����X`�D���9+��G�՟a������`Z��ݡk��s����U��y+�oV�h�+Y�
�+378${��n�e�}u���Ͻ��&B�Y�5�Z��Fvf�^����D�j��o��΁3�^�B��!�/"��n~�7��*ihx�zƠ�X�iE��][EdX�����C��C�ӆ�]�A�*��]H���h�Y?y}}����t:c�:�	B�������TǛ��x��������sJ5���s_f����_z����h��]�a�y�T�^	�6��@F`ތ��Z��z
Zq��V�����O��g>���w�Va$MQ���l������p�������k)tۯ��
Q3�}س�7n��	,��!��c�M�\�ϒ]3���_���t��3<������{Y�'n��8���	��$%���x	��(��[���j��'��'�h��sD�L�ed9٩�t��(�[V�"=�_�� ��]�cA�bE���`�n��#ib�"}�A�IpHJ��b���hߓk����:u�z��������*_�y��\�딐��QoҩVn�s�gʔG�MkM���wO�{�����k|��A�˫��dJm�B_	�Mzvo&�o5Z��M������W5�<���T�,_�_��tw}E��FM�S@�*nG�P8��Y@sHzve�:Z#]�H��T�wW�	�l�UZ�9p�_:�R��!�zN�c٥�W�H���*�7���_l�(wE�î�d��9��m!�+�%�Z�}�qTv�J�$�,�%ꝵ��2��9U80|��-@BO���:Z�k��1�������-��*b�i��U[44�ñ����n�ʛ�v���'R���D��\�m\��O�?c���;mD��ZC���S�~��N__�/n
�7x-��ʎ8ӵo$�ǆ;7���+�B&*J{�kG3�-���{-��-�����V9{_�ď��Š����:Z�c#'�� �b�KC��%��qO�:5�h�|5�O�lJ��Ɣf׉�W5�����'!������`G���a�`?c(@�4/��
�P�ѱ��ΰWlT��e�d��������m�(�H��[��LW�#dw�������7��ЪMw"����z��g$��:�_5�}��!����*�s-��>?q�B"U�;XzFd$_�V��-q�:5ph��K˺j@jb(�s��a �����'��A*dh����S����oS�n�X��'��$�Nz�%��66vJ���Ek���޷r?�f܋��b3�����jOa0�Q�R��
ͽdF:�5�4���q��3k�p���q� .��6{����X����7J��{v;[Ϫ���+]�g��.H\�Z�$�������?�s�SОl"�r��	i�ԢP�&�k�P�
Y��'S���Z����<$����_R�� ��`�}@AA�#ϳ���و!�ķ[�,`���� ���l�/�F>��I6^�n��/��/�^���m�Z>.$/3r]A���^��}����Q��?�a���d�9+�5�f!-�rPقo���0�į��� k �bb�rV��
�T�@W@Uu+�3I�>���S���1���Uj�"U�b�
�$ �+�]����Ɲ�^�da#x�xR|<t|�R�CVS�|���7`|EHJ8��Uz���u�������2�	��.�u��.6n"�d܌��Бд��%LsE�|_�84ޙ��TK�����
��n�߆Ⱥ��Tqu�b�!���є�����3oX�'�c��uH�>}�R� �u��-�t9	Ƕu�0���\�3��ⅭN��_k�d_�(|�7�9_G-c���z/���`"]�$��N�]4I���[(��8�� ��	k��;z�������U$��	���0�c4g%�Pf����ଈ�J�(j�)F�����z�pO9$J3J�f#�AA�:R�a���C�R@`��`��t�42��K	�;��w��g�s��<��}�s�BЦDv����0��j��CM�l*����0d,ed%�JY �q�M��$���2є��/���ʾ�@�:d�('_�b�l����Z��\:��Ǳ�������q��R���.�6`^���Y�Xn��x:u�u�TW���KϬN~��aR��H������볢��e�L��&cUBz�	HВc��n9r�
>�"�ɶi���G�ߛۆ@�ʹ���_����P ^(Y�I�9a��Wj�������ty�W���i 6T	5��a4�!s��l_�M���)�-@.T���E���x��.����Mg[�����K�D�6 ّ�|�a���|:�8��et�T���~		�԰����Z�ۊqVMu9Z�~���a�tb���3�)N&S�~�Ք�?/{q>�=���I�N��d�	g�c6��O��G��Lّ���b0���:����3��Pc:y����ve�gEC�W1߷1b�<���-U¾���xmΌe�H�A�`��En[g������$��|�V�p�� vz��vޘ��� m:%5��D�o�h"�><�ȵ.�0������6��a��qh3O�p����P&j� ����/wY�AKg���bm�+��m�y�R}�i��K�|��N��VX�Pb� ��s�P��q�}4�.ܬ�h���D%�x{0�c�ҵ�����������6񬹫˕����zo���5%,��+:�?�L<"��￉
��[��[��[��gS@|�6h4�`�{��r��B"��be� ��ͮN޾�,��K� ��
go|eZ��Ȑ#2�G�:����T��}zp8Oާ�#[Ci:����l��z1��lt�0O�e�5��Z���'r!����љ�.Ӳ��CZ�5$����{`�����I���N�� ��_����%s�3~�d��� �2�j�ڬTz��A9~�n^��q�_�QLW :�85h��T`�P3�\e�ố0���	�Ȧ�����Ե���A�oʟg7i��'2:Da�?!�#�$8	Z؃K�خ��D��`uÙ����`2'iR�_�ߗ���_�#�"ݏ$t��9�� ���Ef����~�̀�dv������h:������P�F��~D"�� �M��{_(
���]�J�?�Ij!6u �>�j�s�Q-�������Zg��p���{�����X%m\t��bm�7sKq�^�aa�!�]w�,��X@kޘ�S��	u�	P��.� �!M%)�����Cbg�w,�������e3 B?��xr}Ơ|;��̬�%��X"gd�ǵ��5	�r`f��K�Z	���vȈv�,��7��P"Y緙���������X�M$:�ZFH$G�q�"�O�Q�nL����Q��e�l�#|$4[o�����/� `�R�j.�˴F��g\�F�cI�Z37m�89�w�0=́��U@����;H��6@��ol�
���c�7�:7�<�߼�E�G8R�z65�'_�{�D!�Ϥ�F�G1�����2럠b��qމ�]З��vt�����,��\�~7k���'v���?I����-MA}�*�2r�1y%f�;����:���N�X?^���ǿ��z���w-^O�f7�˛�O�u�����Gd���\?�%LU#�W�{V��|�tE�|h�����k/�����eoi��~Q��b�$�W���|ps%8�����2��䑶"E*L�lE[���ec��>N�#�xL�(����I7(]W��i�i�x�cZ��uĎ@�a�{�ә�����+�,c�Y)��q-���b��{���<��6 �06Ơ�%<��l�!Y���H�o6�l�ۆ���C҇���>��B�(����c�����F|�?���Li�8 '�\x�mŦ',�K^�,)"܏a7W�6<��	��"`�c����l���z�/˿坿7[Wq͗ge�-�7�����/6�ߴ��J�-;�H>�?����1z?�MIhNL��Fv�a���Яr���_��>L-Y8I��#ix�G«���jQi�e�X>�(.��.�����Wl�/&�?��R2��6���#��)�^T����gTE�%vVtfnI�mo$~W�d�չ��'����I]_����
ʵ\ܠ�tc[\�b,���I'I� M�O�k�y�u3�P��Ch���/�8�?A6!&��8�H �d��,��E?�Ј�a�U=�4j����
�\��ռ��WZ�x'�al�\��#�K�+*�(���5��H�e�M�c�&�i( �����z?��S�i��_v�׿N�d���VZ�k�������X�wD�zPR� _��/�vFl;���J���ԋ9Q;oz<�/d�p!�m� $r�d<�p8�D%�B<Y���\��5���ڬ�m���8�G?s��`�q!��b�7i��\/��ve�8���os`޵�VC�ؘ������G����ш���$g���޷��j���W�y^�\T j-��+�T&FpZ��cj�JmsK��v$����
v(�=��ߗ_��xp�<��Y�$$*hCkh�i�:M��
�|���5���qkg�������o`[̮��Ց��v%I��x�.²�J��7z7P�z�4	����C��#�Zh�Uo?���聏82nm���iv�LE4r���B�ۋ��۳JNZ�?F�R�Ơ��H�>��Yٓ�
���0dd�r�xO����N₁��&oLՀZ�zRcQ��w�V>%�i���_�`�+����E�k� ����пm`8�=���3_�?0h�`��**�O"2�R�x]I'u�dZa�J�!�%�u�j�5��F�?��<���bQ�@�Y^�!Bo���{,E��Ng���NL��WzT���.-l	f5�[;WVT��P� �э���HAZC	^�nߧ�� �xQ�2{��Q��֏�#��ɱ+�N�����}�ʜ4�7 w�߆�䩮�Ъ�7��N���3�X��U�A� @o������}�i��#��I͝l�{s�\����6��?AF�zʱ (��۶ ���t�f���3�yK�H=	�ɟ�mj��E����8.F@VeZ@d���~Ƀqq�,�e������`ʙ�BZ��<0���+Q#b��cEOz]~�7V�Vzh[��V�%�o=�P�)�����
C�П�FY���7��j
�ϩu�|�ܯ�j{>n[-*'�6�XЄ��ؼ�j��ӡ��I.�N��9ɪ*���d�r��ȁ#��ޒy��F�;M
��䰱��WI|��@����\�����`�*%�"^H��|-��߃u��Ӹ�K~�H�հv��j��[ݑy;6_X����.R�n�&�e���;���,�x_��!�m�N���-s�V_XxG��g��Ǌ����^�($�Z��� I�\��?�sҖG!x�QĔ��}$?^7F�>c^�C���⋇�Y���W�� "[�eD*#�x� �� ��V�Sr�oI?��H���JEk<9EG`H���8ˈ�T���_V�(�?�Ku?�4!����7�'_��\��@���@��_��=�+٦9}�@�$=��#M�K���G��q� v�����ͨj4q�6��WB��	,0����������㘯�EzZ��������ŀ��"�dCI�����+���q�P0:�����{u���6�!Fx~]�[�+�<���[�F�Jz�埽���s���?jSޠƒ�^�:�w3n�v�ҝ0�A=A������ >y$j�K�������*�/=,	���;_R�����7�G:ђY��Oȅ���A8c'�_�Z?:h:�"���R�P�1J��(�Gv������* �Z�[�
�S��#�?�-~A琫�����\�wd��[u�ڢ�V���)�����8�C�E�
���ڞ;�/���h�x�`�P<c�ENUm��ǵá��ht���M��E�T��n��pűnZ���x�]��#e(��^�P���=� ��m��{��� �J���i��Y�/��y�A�R�7�J�~��_Jm�1�׈:Htq1�+ŧ Y#\F�[��k��O�qU�d�%XYL(�����o^��qj�����P�9���\X�L����G�&��\�|�9��m��$_����,���})��g�3J���H�G:�b��=�����-P��Q�.��N�XI�b��h������Jk�kD������M��jB�<�j��j�Yo,ot	Ol� �{'�"ZT H�?��.6�U4	�v����dۭ���L�Xp� R#)���mm��r��ŭˇ�q��������	ʑ\���~��_R�LU �I!���nW�
ɽ6���bld��Tb��Q�4�U?I���&1̔��z�t���(u������K�S��a���٦�F��c�O�7��Y�A�'�T7�s*�A<&q�3���N�*/���W.{�n��/`_k�Tl2�x��T�����2=^�1ܧM��s���ѧR���X���<���ޭ�x�`Æطo�hD�Q]<��D�������l�s%��$��F{$��H|�ڐ�z{�������6��M�5���I��`^�n�����N�Pٟ,�?m#d�̺9�r�Q�(�$u�h�3�)���T�NzI�º����T�Rlv�cL��w��� (�D3�A|���ը,ŪE�}
��/�лf`,���	x-ᠢH�w���;B���H�]|�Zy���nF3�q�X��T�}��Փe��W�W���65��u#��׹�Ʉd�U�����E�����vm���f�88�'/�)hŪ��V�Y̎=*|�@%p�Fhe��Q7[yN҈_�����Ȣ�Ƞ���<c�V��|��w�w�I��k����'���/c�?^��ԍ��Q�s��\����U�U?�?�3R,�@��:�Sf��	��LɪH#A�:�8*��� �[��!�s5`�r�l����u���%u���8{��9����{��W�[N�8
%�}�rȎ:����iճ�>/������,��d �T
�>&+}v ���LT�u	KK�]�X�J���'x7l�"^��U��rj*����b�er��F�j�/��h
�����s�+�\ܾ1��9����f�(����0~�mM��:������1KI����B�j��L��D���mE%ߥ�i�B�?;����	��e������ȿ�[��"ޒ��H��|��&	�9��Y����u��ܭ	6�0�`)ְ{Y�l���{Re/@�z�__f���t��~.�*>�MoE�'��Y��zFMJ���V�B����X���l�K~�zeE�t����[���b0�6�������\��;`e�-RYI��ԤH��(�C���[�CK�?%����(Q2G��W�DH���)Ǌ[h�u�w�.#6ZL���g�җ����P�Lô����a�f���[���g��g��UuG'.��d�=�]�Q\Uw]�<V�0�O;nsq�n: �2{
�%�:�E�����ב���V�<����.�H dPKfK�*�?��}x�xV@A,Oƾy@�c��b;�y)*�~i	��Ƀ�8��w�Q�C��m'�Bz�_��+�A�XYz��ԁ)6=��I�d�X6�"�苑G/����jJ������l`���J��I��J��U��O�����������[�f]R��:�c=%��%�����D5DM�!f��T_���o�2��-(W����؝&�;7/�`�2��>{�>~��;K`��h ��I�Õ ���6LHb�TƩ�}3S���`�'��~�7�8tT�'�X�ѓ��{ҫ���#�h��J���������Ź��1����'��2���G��*e�r.}���gL�N{���n��o��|�����@ؓS���YG� ��	���������bM�v^���d�E�$C*)��v�?ũ��y��� {�[|���F��0���򜬌	���Uxf��v^����Vs���|���|)?(o����_��䝓����olRS��r���{ܝ[��,6Ȣ�礼\*��|�F1�%�k୰��s1�oʴ$��OAq"!�p��_+C1_%w+S����h;!0�9�;{6"U���>�MZ��$�u��{����_`���iܢ��Y�N\)����b�j��3c�i<f��C�͒��Y���o�^0�qj�O���L]
%9�yŸh�ܷޤ�
CZg��9���g���y�R�韽�<�/L���V��G��3@^�JN�8���oo��	��C�Vf���\�~M��(Ę�@Dp�a��iɒ�ycc�B|�Vx��T�ى�!봿�ع����,�¿�A��#�CZ>~D�m'������{�S�\0��M͊@N�����ʜ���V).�G��	1��B�����Ʋ��ߟ�H̕�-��bà���rP^�^hf�6�дc��{�A�^P~�K�9d���Y��+৘0D�Wu���������&!�0�������t�m|l˥� �h�������7y��LG08�i���K�0��-z�w^�h����U�%]������t�!Y������x������(��/s�P�G��)�NfU�,�ǗN�b ��uLs��ЕSqu���´E����?��[�w�֪�I7�mN6���Ⱥqjz<�t�*]��z���P�úJ*�Y=;t��m�_y���[�8s�i^�r����-�(}�H����2�`R�D���r-aC�E��Sw;�M(�dA(P��2:����7]�xrXS3WhPR։Y�n��Y�@�;T��䐀�c��m/_!��4��,�o�ѻ��`!�kC�N��	-��w?P��*�4U���Q�<�2f��[�J�z5�M�h�>S���T�gY����vw�űM�@�\����*�-�ZH�D��@�Ǥ�m�;x	�b/'���9�ぃT��F���
�xU����e�v���7Ң۱Du�
w���T����
gяq�R�c�����v�����?o�%_Q4�B8ׯ�3/&[n�[n�ooj�[.O�X�n�#���ޭ������om�����������_���'���C��$�IeN��GG��Cp-�&���_�"6��7@`��߇2�c�5���B[2奠� �h%T�t dEJ\�}r"v/#�
�/3
_���?�O�8����8Z欍vUa	�s+�KI�L�%���v��S��wbN&c�f/�0�*���w�+�!#,��>e��f|�4�_�0��� �q��z��C�����y_lA��\���/��8{����������y7_o^��FdJ�����H���X��wa	N�����z(ØՇ=�.�ԯ�%ww���K6��{����לX"g	d;�<9��<�<�R�mr��#���ͷNˇ�,D�v�����jHN�/01�>�W����������Dvn[��,}�B��&��}�D炔G���������z� �	����H~�y��5����| !H�mヒ(��JɅ��UN��F5� �O��W�}ј�����u}��1̔6-5��>�Ƣ��5�.����Zg���)�V�I�M�}B��pE4��nm曟�������� ž�����H�ƥ��$'���?'w�Pn���*t�J1V�s��0���#Ag�~dB�\��ꆿ��:���ڞ�V�^��'�3VՇ�dT8: ��>9���J㤄��=��Ѭ�iS�
���Q� ؔC%�w���x�u���`@e��Є�'X=>����X��N���X���X�y��hJA�t������
U�k#��C0��\�@ف��,,�W�H�r�>���AM���e݅p���4�3�.`���E�.f�����M֢������&Yo�ʲn���1����}]���|ΞЗ.�"�/��I��<��
٤]��>� Ka�6�/m!t�1�(��bw�T�.)C�s�p�IyI��e1\�L������^���|A�)=���:o��;_����<-����}��� �Pn�Z�U5�G��T�����R��&�v�Wč�&5�e0�ХB�ʝ�%,�.q��G�]ֈ����\/��,M9���j�?��E"��T��~>����XtȞp~>��������17�{j�Wj���})Y�GK*�1f�9��ȚZ*e̖�z��u��Zt����"���=ڼ��ykz��C+X,(��{�v��Y���b�}�;��6v�/E*���%�Jy���h�p��SF��G.Za��j] �,���a}��U���������]���{�uޕX�/�n�(�����+����Z��/�6�>s1�x�i_P�-H������
�*��K~��h���/��.�<�����v���Y�KKq@l�%�^�Q}����m��%�y�i@ea���Σ��F-����SX��|��ǭ����\���M���q��YZYf�ߓ�����N�Uu�/�(�g���LhX�!9�I����D�'���}F!����l���<�1�;Ό_�y��������a p�����DG��NuLJS�q�w���Aٶlr��ϛ�~%4ݍ&�s�Ǖ�
i?�P]�]����ˑ
�t�	_ւn�i���}��8;"�c��װ��|B��$�H�3y=,Eģ6�:��f?�}3��=Kek3�I����V��;%\�U6�ia�3S���𪛒#�9;��ŔK"P�Gq�Yif�#���:������]�X_Q$|���n>W���
.�f�ª|��:�\{]u>E��c�N%2����?��TT���j�E壘ȥ>ؽ����W<�40IŹG͡���$�m�����nZœz�tT��0�|nf����Zb-s�O�؀+�R�e&��h,s���L|5���!K�ڻE��G�,}���ЁBh��ϫ����h�p��C�KM9S�=�Xq�F�G�!��"6�ı%�U�l�<��4�;����li�{��2(���^T�7rx���he�zAw�| �Ai�)w�rL�P�E}�8/���E2/~�F�1�ύiZxm<xp��_�ˊ;���. �@��1��ZXS-���i�&�)�c>u��pjO:��	�1�3x�T��؜�o��IQ,�V{��/�Z��`f��z�贯w|������
��ϣϦ/7���x�)Wq4[�z���#\00���O�+�A�^��<��0�ń���!)2 v섞��/ӤUR���oC7p;@�5I�H����G&�Ib�s4�JmG�iձ���aU����.��2t�5B�5����:%�1C�C���چ���GQ�S�VK��]��ᠾ3@]��2b�'e)��DOQ�}�ݧ%��g��:ׄ�VUkA�$ѳ�S���pʹm�2c�
ςᶏ��Z���bs��,���ehZ����������^�������AҊU��^�f1ķ(�����c�f���w(�=�=��L�`�)�����/�O����ka��D��o��hL��uά��� +U�5���K=�T��OE�>��'j�f40��7bT�[�ϐ��Wm��'p�O1�'�cLՀ6g���O�`��Kl�U�'�����7�M�e���F;5`>ݽY9�Sݲv<�rj�eh�i�� 51�v�IR���X��o2^���U���}�8ꔟ�%D��K�f<ݏ��f7X�ݱ�ܕ�;̘*�k����7hrb5��ȓ��Bb+��莞���c�>~kNQ�Y(:q94CO�S!��r�U�����#-��$@۶��5}ݶ)1K9i�'��a��%��P �Jyʒ���G0d���ڛڷ�c��D�w�*b�N +���wȝ���^E�^��\ޜ6�n�\��]�?��o���~�`�4oP)�v���$�x�4��g<�.�w���+@�������8���bw��J���T .A-x�K��D���� ��bt���1r��J�gJLP�Ul.���e'�H�0~��-�5S�r�B���P�~�y��N�������E�w��*>1�{wz~�UͽԽ�{;s��XO���
�C���������e|'Ph�PT��T\�7� �ݡ� 7F��ч\��Q�EQl�3�U�n7K��k7;�gǣ��Y��v�Ǌ"�2ӛk�|l����Ki�N:Ѹ�}����@�;Y�I��2B9展���+}��C���u�^���N�߹���䡶p.?`V�Tv/��:�`�����ʧl*+�2�Hu�m���쑂�k��}H����Z*MjLv�(^�'�� J���@(Ţs*���M� �+��^�-�������J��,��j����(rb���7�҂pPq�>��t����Q g#�s��tj瑳h_��E������E!�~��}���[uf?M����As���H�=��ދ�<��� 9g����+��+� S-��( �������}	Ur��m/4�����(X�����P��p�P���S-Y�����E�\��`Y���ݣ���v�3�HRˋ��d)6�~��C�����WF
H�-͑��'U%�x�'�P;Y���}Ea:g)��.��Q�Ƨ��Ȝ���0�lr3w����d��w�/x�u�wӯ��~9)׆<�S���g���݂9�Q���3�JQllК	B�t�g���]�ՠ�㷿ۦ��p��T�+���ֵ>0E�4�g�Wz�3��&�6��s:>���iQt�EY���jf��O�1�Yh>����=��;�����E�[O�C���m�^�%�Ng=`����h\y���k1����k�/�!��Թ_��wh�d��^Pͩ�2%�_y�`���WS2���W��3_��V��t��������� ����*�����(�������ʔL��E�&���#)���
��ו߬N�q�K7~�^;i�Y.���g�ɐ�uT��xT�+Ĥ��H��ͳŢf���ĩ @����_V-~N;~�]��^���S�X��ؽP�}D���!��$bǥ)@��*�-��-
�D����C��J�c�N�����l�o��LvF���ר5�n[���Fν��UaeC�����
y���ɲ�Ӷ
��^&p���-��,���l^�N�����
�^�6|꺹�J+NSƘ�̟l85��:�	6��x�m��5���0_�װ��;=3�w��J��<�p��-G�?*�a�磺���Cs8^�;p���(_�%�Ʌ�&�7��j�T�)���/�P�����V�����.��E2�e�=hyVfK���N����qg�������tZZ���u�����&?�z��~I��&װ38�i[B�N�~�s�l	�*�é�V�/���n@��6S�~3xh��&�+n�/��<�vF��^�:p���z1�������nw�l�u��Xf�x���N���q�n�rS�_+�5�n���Y�P�����C�1M����5IK��Fcdg�,=���?�X
1o�B��a4��i��xQ73�6�3p§�:�#�B�b�69�_�ܓX����4��������)�=���F�}!�`���_����K��sm�#N��P�Ù�%�2"��&-��W5�r�O!;c۔��c��~e/���+�|$�QV��ߧ�����A!��<�^��7aJj�7�F>�gi�tq3�f�U���5�K���p�ɘi
)+�)�d�#:�Z�1�a:R"�0���b>^�"6l��vb���2 � ��^C��s�%m+ h���r�y�}t��/�,��=�k����G��eK+�Jx{�� ��t�����1�8��j[�D*�]ّ"=�G:�5���pz��pusj���pk�1�o��39kQ"��p��WӅ���I�o,��i֠�������v�ϫ̟B߽���OaTPjs�K(�N|���?!���/6i��r42ʔ����	�J��?¬/窠l����Ҥ�8b��<?���L}|v֨g���q�K�P�O�* ��E�r9�fA��������M&>��4	e��{=�>zC�%A,ws�ʸ�o��{D�V�y��/&! �G�M�,�(e��v�h��n��2g�̾o�d*��'��A"к�+�I����ۇ�����vN�+	�M�4�x�<��V�\��r7|��pK٪�<�C���7C��b�!vX;IY:���|��Z_S���~B^��' �V�7�P�"Aqb�E��!���'�O��DAH\༉�|�0���\�j���|>�i�:Bt6�oM�Ǩ�����ؖ�ۓ��Y��ٖ������Æ����ŀ��7���Ι��7��N�u���4���/͛/�|8�2�d�,����V����_yA��Q�ib�C�
�H²)ߌ�~��2l��ua4�ۂ����<}�`)����z	�E{�b�f����F��n�	�eP�|u��Ҥn�С9"oN�9���ϩ��K�&�����l���E�_w�d��֪.N6�:�n��u0Q�n�Υ���m<�尲��t�E]s�>�C�?8({Z��:���۲-��}[�]O��3ĝ�9�l"���;��5����e]A�@7��&���̆�n�Z	��ǵ�\��ݵ;��ޣF�P�x��������`�Ne�l�8vaLA��G�)��/��J�����{g��Cc�w�"���c�W�؋E�h3�j��{ӝ�f��I0N�.��=�����گ��
��`��������vʵ�ZeK��S;A�gOQ�ݮ����PrmlL�r��`��T�r�	�TL��qk$�,���܅��=>��A�8�2]������ƤN�cr�Ș�H�yU����5/����=9
�r��Ŭ�qr��6t�i��KR4��S��2�DOe7U�5Ǐ�K�ܲ�\�ٹ+j��8�_r'~����Z}�3�f�sK<K�/ٺ� ?h,w�..?� [:ֱ7I&�5��\�h�����]���,���%6��m��*f���ܳW{!����"A�ͯӌ���wς#�%��&�<	�i�i�D� �]����&�U��"�l��%g�S��N��^��$�.���/@o���Bea+��'Z/��Od��B�8��֎�ue�\�|ܘ̚��8�>��k����jلo�']��0��>P�N1��)���H�kF ƅ�>Q�뷲S=w����p�(&���	%a�fe(}��%��r��G����u�5�C�Hxà�V�ړp�y�6Ҏ����.ɣ�<Q���<$�<$��4{Ŧ\��D�Ia{R���.��b�������[Ƙ��[m>ec�Ǘ�Ou�,(Ρ��d��G�Ґ�}��E+�Zxh0y����:1j�u���"W"��O�zCj����=c���*���w�;S�i8��w}R)E�� yu>�ŰAn$[�c��}�mT��7����>b�7o>��Z$s��&V��C��M�ɋ�B��n����υC�)�������{�y��)b�ib�(�$�}�@�juT�++�o���߷4���:h0��Fú^T+@C�HH��L���	R}U�rĜ�+z�Ku�Oc=�T���U�kĪTa�_Ÿ���jW��-��X��T#���b��Z�������j�@��������&w�O����܇�?-F0B��~(�-��5�c!�M������7��)}���^��TMP�![ȷ���HP�ev��J�1�ltH�_Ș��H-��BC�C*Z#�٘�y�Q�
 ]��A](��MT����_	��#)I�����c_�t�fW���7��zEy%�e�Ɇ��E�`4����ʹT��r?2ّf��BT�0�R"N�^�!�R�'k��J�"Q�/���0���?�P��o�����~\.�&��?}�q27����1W���U�V�щ ��&P7����mʜ
$�SA_�^�+\m[>�\���
A��+Im;dk8�_OO��2��zG�q��VՒ����[�!,Z�#�"^,��-&A����Y�B۽���Ę�M[�w�d�;i�h���'��t4���+����P�â�8��ɴ�����D��aOS��a�Hd���Ƣ��	6��v��5U��� qZ��X�` Ibp��}6ֈFK
��I��U:ȶ�q_�j����/�oo^Ly ��e~TgP���Cv V�:�q �	�6�����h�B^2�����Ӿҵș�n9w��mW��Oݻ�UBe�*��2�)�đv�����m^|��
,�7��������!ӦH����dk��|�8T��E�����˭��bS>RX'�������'D��|���,���������')���ru�t8}ݹe��k���d~.;��eg�Gl�|}No�r��3������-և��㭡��_e��bh�w`[���+��_�Qw#\l��
;^��N����(+T>ih��_���ѫ�9����Ro52g�]V7��T�uuf|_Q���|k�5����}&D����=�nݨս��!#Q!����y� �L��s�I�C���e�j����әTf�� D�H�0�,S	x:B9`�_M��?\7�h�#Oo����H6�͖kw��
�ė�a&0�	LU����⭚Ȇbn&���y��&DE6��|�!e��İ%����p�y^�xs�FK�(�tVjC�6t6q�;`�G��v^��_)��C��<$�uψ�S>���*cz22em`Bi9�3)�e��z2F�2���a�c�uU�>�3(pIc,L�����C�B 81��%L0��t��X�ÿ0$6���=��٫z�>�h^	�z<s"��y�Z�Lq��`�/�_�����j1�������z�b��hr�����omi�_�m�$���������!�
���)���So�&龒��]Bz#��n����4�+���-�`N�R�l�5�a�/&4a� ���I�_����8���R���[Z��Y�/��D/��+�U�P�e%8���+o���@�	���F����	�%,dah�1�^�Hj���(Q�w�o{����%�_[Kh1\K�̞\;��u0'5���������h<���r��n]�Nc���>V4`�#�i�f1�>X�K��w��v�@�/�Z_?������v�˩��ܷZˎ�2�O��t�+ol��Fٔ���9��ו���J��4��5��&w\s�Kj�C0Ui���Q���T9��wbR�5@��u@�dǥ�jd��`m��@l1�nLb��l������딤�A΅W��/�^�7��L���$Y�=�6	��~�C���~�˭���(���z���Mk��my6�ɷʬ�/�6���Y>j@��)Hg9�����[l	�k�ՙW��x���I1����h^�	K����*���G���*�����E��}��7f�7k�f�] �n�
+ ��$Һ���Zӫ�P��Nlw�Pg�H�#^Y|eg�QK�(-_G0�C�z+��2�&xBk��^�XE���-9!����@�8�.�g,��A0�rKk/�
L:Ń�笈�y���N�
b�Y�<b��H�U+��4a���Xv	�}7��u=p�<��n�WաL2��0��"��qJJA%)�65�0����<�X�|y>��������b��c�I�������R�Uޫl����htrD�����,ë��ʺi����O?�2��8�]S~��;��f�n��㈘���B��ǡ�SԐ�ۆo� cKH�f[��v���*L�����[�d��J�{�:�'�����7�a�ĞĞ_�^g@3����(~{�6�9RH�0�A?��k����Ӣԗ�U;�M6�+ �([����Rʁ�k�Շ�3=~�D�kj1��>�{,���ݼힿᄿ��f���ᜊ�mn������?,kԏ��}Su�|L�N�����ɲ�����uP�G��c�f|�pRc�х�G����˹���2LC<F��r�8T"�1�0s��=��V_.����X�VP"2o(;׫X<���`ح��UY�������0��8���88���
���WP@F��dZ�"��I/bHg1�����4� 2�]tɗDe�D5eؘ��w�&{���Nm�Hj�E̙̠U�N���M\��m� ��1�E���?�^>�g�c�NW����Kퟮ-J�i|{d�9��K�h�@J���<�����*_�B+�dփ)������I�`�BN.�̭��xAbw�Q�<M	��N��� �ti����G��?V���&Q��|��a��z�R���Fy"�����ˎ]eGE}���'zL��Ub�M$�����rMn;s}3�����6��hc/���I|8�,���7�/�>�`����������&s���x��6���l��wJ�$���VV�*w�Y椮Y��x���3�7Z�j�Ֆګb�V��6��A콕*��;�b����+�����5.�߽���[�;�3����0�\�m�Nŝ�<xj�\8HJ'i�ؘ�+�,�e��4N�Օ��,�H�B5'�`�W��f�Ma���xG�h�'���/$�����nX����'x��Ɩ���
.�h�Sߊ>.����*1�	����$1®���p�B*��{?N�埞
�;�Cѻ,tt�=~I���OB��(��"v���aX��BW)��)(��-���ȉƏ�)����}y�>w7��@����,Ӧ��IfJ�`��c���[�7�F���`�v�����z<&A��c��d�M+�h�E��{Dj������,�1�n+��aK,�MdĜ�j*�qr<�k%�
�A�l��+�΁�'�અ��XN]�o]�]���@��0���MQ�!�9���Q�Vk �(qq!����x�ĥN�Ӫ�ݱ�����ґ��׀���a٫ҟ5�oD�%+�D&��~���v�6�5Ē`g�~��u�7��G�S�)�[�VF�B�h�D5	����|���n a�
�R��7�2Ӥe���LP�JۈcV���m>�y�׉:H��S2���_c��w�&�U���l��j^��#v&��p�yP�� �Ìt�c�w�wi��?/6#��$/�"�μ?ns��ws<̞�O���}�.o+~'�f: %X�#��<U�cv
��������F��)�i��v�4T*�k;&M�j�t:�������Z�6����X�Ьg�/�(4����'�t�cT�H�ÞZɀ����:#j_` ��J�Z�e�Z]�q���i8P���B�b�F٤����y,�,��cRt��@;M�P��s?ı��	��)��Y�����U�y���Y�Z݅�op*���|�@N�y��2?�������D`��Z��3$���0��O�>����Id���?���~x��O�)c$��vj��I��V|w�-��z�.O]<��F�����<�{��e��T|3������o��G����&���+�`�Lz`4��D��������({�g`���y�Y�N$G�2��`k�h�9��y�&��C�馿e�P�U��=�BC����ɩ�MZ�
��]w��#�`�@���|�ZxWɶ��*��C�!�sH�tB�ej0_9I:�Ll#,:z���w�&k��tg��x��h���'���W�Lˍ''[�R�7��f��G�d.�K� ��z���}��������Ϊ/��yo��&g��_<�?��ʁ��&�%��ƬhEӰ)�;A"]��nT�d�R����`�u	K�%�|M��f�m9�lY�,h��W����v)"�J�K���.�	/gra���ȖMΕI�������)���sO���e|�Q�K��*��5{{�,o~�жqtW#:Um���GQ�'yU"q��Bs�q�̞���j�f�(g,%�<�=
��Z@�a}S�
���[(K��u�~yrGg�l�8��U05���F�6:�-�逥�rfO�#Ŋ(d Rt�bQ��TF�,n��8A��/J�.��8��"Bi�0��&��I|H���j�aS4�D�^��"�7dD��xC8˞e��wy�;ܓe�r�i��O�����Z�æ�	�(dI�J���?�
Ɖ��������o`0ѕ�h:�~5 z*B9��Y�{ڪs��^�#6;�IIH��rL�#���O�9,�g-�����6s$9�������ā@���u�9�2��H��Y������w��7�xǚ�o�8�I����ۿ]1���"��iE���+>��m㮾@S�3�F߳�
Q{v�Cfݦ�;wK2���=�
+x8��/����;�������Ow��Q�]-�a@4/��؉)�D\��V�b73�[�����-�*@�� ��8ڔ�Bf�����6�����}aq-� �&��K:�I`�h�Q��M�K��!:��H�Ω�L���t��^�	;~a��V�������i�!�1�s��N�D=X�۪�4��#�^Љnnz����A�����n��&9�L���N�-+K�W��O���ǜ`��.`�k��'�l>a�%I�kΣ��FU4r����y�hρ�%��^	�@��������E�}S��L����(x�K��R��=R>$�)b	��������uޟ_d�:-�)qϟ����_��Գ,.�EGe�?W�kz���]��}��r�r}<ϒ�9��ӟ+]jWQ����ɏ��}�mw�G�Y��^��9���?�?(]����OS���P�������U���-��az�NQ�E�_JQNO�,i�\ї&�@:��'h�ZJ�kG2'L��~w����xj������3���w���-��k>�/u	o�����Al�(@T%�*�R���4#�Q�֥��IT���-<BE��E�T�g	��Oh]R�=R6��6[�i�xԓ�K�>	�<+��+*f��(��(R��GI�~+���|6��xm�0��W�H�6�c�[:������B~�7c�\�1e��d1頔���a���u�xgA�[�=� �g�]�6��"�1xWȶ�|sJJq^��#��钚p+�CP���w���� |i���}�J[�JWL��I��B�-��\Bڀv+�.�vBZ��Ԋ�����Fꚡ��*	sG����t�?�'m��t�,���3 `� �绎���Xώ��2��Y��XV#mm>�����j:U�>�V h��÷4qt�-5�i�������r�m�`�0~�BO���C6���*���V:�eXW�{����|�"���&Cx�*���X5R����
��D��ά��H�Z�2u�BWY�])�QS�v��B�Xju��=d��f�*;
B�K��L���o�Tm5?ї1H�̝����C$�
���䴖�=���lN8K��z��i2�[�&��3>![F���@��ڦI�8rAśq��"1��j#�h8Nk�f]$|G,_�N�xEo�j�:�"��i���LuDǞ�Mw����00�������@ "g�ܱN^p�o�(!��qPG�z����!���
��y��Σ��HZy��h|D�R{����H�9��i�����rlN��a�&����*��.�(��� �@G���,��8���pu�����\Ie^.�(ORX`a��@rԞ 56.F�´��?�^���+�4�3�ӧ-�nW�WSY_�&j���)�om�5"��)w�[2O�F�&�s1/کDo���sw�������!�S��d��D*c�,IO���W��W]�7a$��n��c�Z<.w7oS��߭?v���cQ������ ��A!?5������!�G+R��#�}l�8��6`��v:b\�d�)2����_tH2EK�<���n�ؖ��aeܷ��-��Gg�?��o�Y��'*X�B��C:F��;}g�C�f�JZ�<������4��S=-�VJ�i0)t^L����i���t,�C����GZ^Ƅi��QnH�K�C(�"!֜��36[��.^�a� 3}�x%��E�u��եo$u�����g�)T��i�Ȕ ��]'�w�ͣ�T���֨�R�r�DWr2�50���QK��U������v��kl���?���.���>�ۓ��혝P���b�Ү�	�
�D�4�@�f��#��Z�ù��,�[��@;P����F�a�&�JѲݼ�U����_*�����w��k�6H4�i�w��r��5��4�܅��L���Q+AS����$;e-�j���3?������1K{�¶'���B)��s�����$�hɅ(����mM�� �%�ʩO�]Y�/%W2�#W��f�H��~Y�y?�m��9~>0+�?�=0�w�Q�9��"��@*K �^�<kN%*����gFA�����e5"��w�{1�Hq�3Ő�Ad���9fn���+���K5�њV
OCA#�_5��oV���ח��$}|���\|���t�~:���X,�)�)��׌[�#�߂�����<�����WE��EDBJ)�Nj��C����N,��	�:z�a1�T�)��WM�.����s��)Q)���܋T���t.WֲJg(��,��p�,�A@�%�͈~��<W���sM�Ń�Cc�JC�IJX{�/A?��/gY�4��>��ᡔ=�6qf~a��]��^_u�%�s�^,�:�'��h* OA��4�����]Ȳ-ş9��ys�v��w6�X�͆&�y�n�<h����t�bZy��4D�c)���������l���`�r��,!(�Jz9�7�]��'��Y)�q��$��_��^���esZfF��M�l
Y�4#��u�E�.�L��s&X���3�J��H��3��|��]�y���\��D/7���ٔێ&����~.�ʧ��F��D�m!��1��%�>��Z!�&�����9]S?χnԁ���r����+o��Զ�������(��x�/%���D�����Y��{t���ؙ���7���:��;���j$ʫ��d̞��B'ԋ~v0d�\ø��j����X���F����vN6W�`�EՊɯC��ѹ_>T�^��٦s�2f��/��]�1������wӑ�__���y�akUaW�pİ����*K.�u}�aɯa��1�����	��A�Jn��d�}� b9�0��_�M
N�q����u5�k �)1n-OhR#�P@1$�u��*��������J�$���88������p֯�y:������OcI�4���F��f�PX <����3�P�r}W�k�=X������Է3��I>i�uO��B?!���=3�a'��|P	u���N/�f4���>K���;l�kh��6��Y6f��P�':�G�ֵ�C��>�r�JۙC�i� �>7�-1�]�)���g�[k�����n�6[ۻ���u�omH���^�Q��W�i���\[޸�s���2�^G�`�����^7矨��@�"m�j�
>�)��t��i4'L�A��X	o&��_�
l�	��j�{�_�@�m�t��U�Y��g]I���J�����P>�L��`��I�k!�_��a�4؏�yU�VV����2eL���_�L	3�{�����ͭ�ѧ��挱�e�r6�~%t�DHru<�IK��I��������.i�}�F��M��kw$�%AYbaD^a�\��~���f��n��D-K{e���'����8K����ܩ-4Y����������+�L��A�"SaY������'w����0s�S�����f/�]�<j^��@��Æ��jh4=�������Ra�@���t�6��4@�B]N�H8��Mu���:��r�8�y�$��l;���1�BB8:eǖӈ ��R��v��5��P��Vu=6��γFQ��JF+(4�zA�ʏ)-+	�?�����Ϙ��S�*��2ԃ�ya�lP����3����;�b�`d���/��i8,�5���b�g�a���uAb0FC��ʝ�x>��h�TϿ�/��]��ka^y/�͇Z�=�~[m�^���d-�^���J�ܟ�z:�8��/W;�&�L4�8��v���`������Wp���p�(8{�H�K��17x�4F<	U~v�V��pҹקǇo!z|.��'w��Q8���)�yc��4O�B"��B���T��0VP��Zr�O��l-ϺVC������/]�=dd �/U2^h(�̊������(Wp��.�MU'�x��f
�F�Lbf����W���zw���[��h"m)r��v�����%�L���#���<���a[CY���h�R���4�]3�2�5%�F��ʏsy�'�4#���1��6V���U�B-����;�G�G����(�H`�lZ�_b��8I��C�3�)��������ъ�������뛎9\�h�V����M������[/U�C��)�x�1��O�bGW:��a�D����<M���8x
�Cўy ~��f��T�E���{nq�Z9����|�����<���i�Pͫ:��;���}iAT�(GMْ&���a������Ъ���H�	SL��ߙ����8d��o��܏��]�]����ty�����w�jC���������M�wcK�
�.�+T����Q��[I�b�xI�YF�NN�ݤ|�m��sx�5 d�H1�%Ng:0�) ԃᡐ��N6��O�쬚1� G>�,���ejlІ���D����f�XL��~;��l�)Sg_ǅ�M:�=�"Qq����ˉ&��k��gT��hݺI6p��o�EF�1쌀h�a�~�IV��,��f?��ϛ������������_"^�)20�Ŗ� X�NUUv���`���E8�b�j~���.�P�m�\��o<��f��r�,���>��DYWo-�ל��t����gI]�|�{z��w��=�j&F��g��0����=-�F�h+\�d���2z����.�@�[��������8�� �2���Uҫ�	f<O'��J5K�@��_s�������{���<��Ģ��^^ѽ�xak6 �g|oF�hI�:�,؝�X�3��L��H?#��a���N��X�P�>�1A�n�	%J�
�b� �R��`ԝ]��q��I��zۃ_X|�4�f��ۃ�1�0ǈJ����n0]�����ҩ1��L�4E��煝ܨA���s��5���ɜ.�-oq����>��+��yp:�E�ݷo	.�����o�e�5s��b�(�^u����}\P$/�5[��}E/bf�K��Br:�DIWa�4�m�'~l��a�&�^ҩ�#�x�2��Y�$�z�	 �����F��W�ԁ��M	�j ����Ɋ��%t�SCb�����L����^oVG����aYK@���� ��N�Q�'=���cv/�A(?�J�����5r<�!��q
c���C���.�9`���?%2�E
������g0�U14*e��f��AQ�?���:y/�Z�/�zZ�%�./^շ^܅���_��мw\ns^�
��ria��e�7u�t�pw�1�O3<��p�}2.��1��4�Ҡ>���P;Xl;fB��9 
�q��j3b2W�Ǜ�����ٜv�qB4��%�Ԍ����q�p�zo5��s���q9Ζ6��!<�JC#I�*����ĵ�ɠ	_D]�ⳕ��'=���F/�������I �m�:�ڄ��(t���ޏV���jP!{�P���[��s�>�eJ�)������<8��ψDcI�r���pܙCE�^m����}ab0�N��cn/��������3�Z�;��������ٴ�6e��տ7O�@��8��e3�=IP�僺Mm:�$����;���}�*��1�"`��T���omt���J��P����IѲM.H��ł�M ��C*�r&#��l�]���|5�����É��n�~=!]�Z��=��g�Y0Q���"�ϵqJ2�p|�]*ST��?�0���N�*OZ���]fWa�ޚּ�R2۠�}����b��w�ځT���]���_���዗��W��-��W#)��������>n��9�w���h��t��`d(=l��o��DA��M�D�.)�;�,Ia�#�bP)F`��k9��Q�0�\z�)w�S�&�t.޾ş�βl>�7�pW-db9�}��7��O#U%�W����OV���S^
؏0�Ǔ=u w�DtV�\i�ې���1K��?-�"J����ٮ���Ds]=-����=����FX)2���~^#a�a�Oj�x�$��:�0�o��%��<�͞VIr���m��ȨIN+�#]��j����v�1�9�3?�Vk�3�s�g�N�}M��o�X9xe��"N���0�szu����]����?.���t�So����hk2�/�����I���|��w�h��Ro��0[�?�
�+5%���נ�1����O��'	���o��������	=��=�p�������5���=��ap1�I�t�'iۈdbcc��ߗ	�GS3���t�SLy���"��^��V�iv9��)񫍷�6Y~�k6˭,o7Ӫ�7�LV�6�zr8��/��D�f��}jD��s�i+�9�l�LP�W��=������˳�NpȰ1D�A��Wd0�r���s�&a�9�5�o@��k�u�߬����+��� �A�E�`9�s�����;o3财��4�bMm�  ������i��i���������>d;����D����w�W4N���O���*њU8b͖FĂ %k��:BN�^����׶Fk����"}g�Hz\pǸ(n-�#�¦�C�qU��@�,DU,D��B���t�-u��8=I�"e3��Ka��'^jL���t���ŀ�n���H`��z�\ZG^��vK4�,m��t?R3&��{���F���}�8΂��Z��p2��.9X��XV5J+��!.昏�H
i"]�gVG�U����k5�x��P��|��Q/��=Ɇ�w�I����������rc����iz\I�zy<�ZI�{.�S��0U`�e���NE���AW|��g/{��"�5�^�R؎D��
My';�W�q�ޞ����ڂ��Q	� `H�HM#_�NG�Ϯ�H�ɼ�[e*Q�*Jsdӱ��,~İ�Osޞ@�_�F9�p�i�/������A��|ʬ�q�l�Ec�=�'����-��-��o6�,<ޕ���%�ME��hT��%��0����g�
(�{�w�G�=������|!�ø,"Q+��i}|ҙ��\�z�TJ��^?�y�,�Ghd�;�b��b�(�MW�Ѵ���]<��)!.���G3�Vs���2�8�U�HQVn���D��h}jĨ��8���lu�)�H� m��Q?kN�B��ך�7�$�e���kK�Fs��5o�h��bR��Z�,Y{��w����q���V<���$����r�V\xt���z=<��qퟙXYOm�yu�� ��̩hq1B)��B����<��|)��f����F�nѬ�+=�4��k��,�]z��1�	��7~�l�i�d�^�	n
��f*[X�#�Ȇ��\Љ�M�Uo	%ݳT�D۱�����མT�
����2:'��^���ƀl�ȿڹ���B=�L�����g~�B���~)_�����7�����9ÎD}6�j��o�,1��\!yb'_�@⥒�L�M�si��ڴ!!�Fk�ր�$(6Y�3as(�����`½^:�b�+��0A��ӿ�.G�O'c���p�������z@�#�ɞ�a���V�]�W}�\��- `�mY�碣�9����D=џ~ܤ�:�x����xl�FrKzmm���
o]w�?_����n���d��]���4����>�-R%���n(`μ�n�'�K����J���E����ϟ�"rs�	�����ኙ*�?����p�����r�c��H[F��cC���[�ǚ�l�K!^���ݛ�܅4��P\ju�G��xP���fA�%+��y��j̹�����g��("��`?�U��z��dUԕ�y5�=!z�8y��6��-�� 1�w@A3א���7��--꺘x�A$�d5Y���=�ʣ�A����m�G�\3�
kr�ϕ\��[���4�����SPM"[��'�Z�ŏ+��blJ KI��Q%��n� �IT�4�k��L(�
"Z�/,��.�u�M���7c1��aq��]Gq��� �e.���C�O��s�G%��Og�h�$�[�=%��Vo�^�C8��Suk)����(w-��"^�b�ƿI��Xg�(Ni�Z����o����EY�v]���Zc/�@��`�t悹�e�~i��Ė��þJ�]�#I��c��;�i39�֪���(k�	�]#�R��2t0�gʂz�5A�K�솴�E7����t���~�w������ϥr�K-&�t� /ًJMY���C�w�m�t��*Of�q؆M��`���~��5oQrxV��.�(�?y��/Q3��~(�G���t�ѷl%
�����3�`v��m.�P胶����Gӛ���I�A�-�]�(�Z���
>j�<�q��$�h��R��/��7� {s^��:�5�ܝ��E3�d��� P��"0�(�V>��$�x �-��\q`�<�{M�='�̙O�91��Ab�G��_��j�qg������BI]�Rمg���B��\23-�(�MmG�����x�F5Y���ԡa�%4դ����z-�y�I�lju�/g��W�~d;��_i8�Y�2�ts2��|��w���残����'��ѩ���ܠQAO�����B�^x��FJ�̽�)ۈq-N!6j��ԢB�['O"_�q~�F���4��=�z��u���ح{�j��Yn��4@�
�-��< � �A��N����A�D�/��RL�kF]N	��_
>�_�L���B2��a�̆k(Mֲέ�UaB�?����?�g�F�~��V����:Xht����/�_�	���^jp9�N�ߞ�JVL��������Q�;��D?�g���F0����E�B������� ����y%�fa5`�뿰�U�A_aaI_��ȿ��W��'�L�f�/�:QKvn�+�12ѕ�W�ԋV�Feo��,ȿB��>���[_a�C~j�C�0W�HjPlto\��.�?��Q|Y{\6AO&�F���;A]������g�f���"�}Y����>�|�$��1�s4��}�� ˖E.z��\P�gY���h:ח2 ������B(�%H�u去>�fe(S�4��P`c�����TG2������,���VY-�ZU
�WDG4�K{�lF��,F�|�V�ޫ|�M�CLQM�SUb+��lcW/�J�nﶙ[�|��c��.%�λ��g@�+~�V�����]�J٨����P��a��nT%p��U_���V�"zI�i�Z��z����o�[J~��:������i�z*L�f_���!�xJ��e�v��F�B��s經�q:��Ӄ��8]�1�V�l���d��ςG��S�~p]T����E!Y��U?��h�k�;-C������&V'{��M�B-?�D�Gq��DyTS�[�"���\G��%>�&A߼�{�R�ӎ�G�sX�%��r���k���q{��5~�BE�?@黎8��C�:s�
�,�y���JAf��8���y�	�t�٠�{G�c��2��E��_�$b��i�?���0�7O����a,-#�Sf�`.���T�~a��bD���s��殅O����]�����S��#A9��r1M��A��qrM�r�g��*g..��g5������� U��)��YX��$rJ�J��Úc�u7^K+iCyfZ!a���5�D(䀺�,H��:�I��h1Ih���"�g�<�a8�!��g��ޒ�{W�舣bz �v�ǔ��(C�/��]��c�1`���l�a����O�hW�X�f���$�/���aK���%��p�Mie��Z�$]�h��A�&���b�����p���$eiY����%��7�B��"�H�Y�uK7���6������'co){�"�~��&�:?Q�?�2��#�����/��Ϟ�_�1>�#v��A�X#r��/h??$�s~m?��-�YFwco3$�P
�tk�_X�=x_��6]����:��"�T����̘^Z��+�Q��Ƚ�����+]&�~���>�e��I��>a8��|B���u�7k����w,k1�zg��I2���Y�n4�{�!��3eM�Z�A��\��b��<����0E���\J�D1�����'VT]?��`+#�J�NwRa���3�.q��Ar���u�OeyQ�q��Ib�#Y�Kzp�O��b'ޅ�r���8�Yl3k�#m,�1�%d,¿�&ӑB��~��u� ���OZEљ`@}��n!fP ����u6� ��Y�����7�D�����R�}������c������ҝ�8��II}>����$�~~�{fE�kr�D�rK����ࡓP�U��M��R�&���Wc�^n�Cc�7]L��G���3�]��_���bPuɛ>�υ��QxF�vaA7��u��Bk��t��4��JkӋ��G�?���z�������#;�>@Ճ�U9�xJ��q[b�/�t���{������[�`���O�H���6 �$4k1kVw�'}���<���E�	+:	��?����L���hㅬ��|�g�V1�>6&�i|B���ӂ��^sɳ�-�Hu��#A+�L�$��L�&v��_M�F�?:;�r����e�8���;�A��
*�
���'��M��3�!�������[��=0�u��9�L��ln��R\��*�WyO��/7I�ua�t�Ω�1�E�+�ǭ��W�D�	���-
a>�'24]a��0 ��5ɳ��έ��� #w	�e���P�D+���l�t��e&"���Y�����n�ߗr%�ˁC�3D ܯ���hP��4�F���&�z\�2���qa�X,���K�9Y���4�ׇZ윺o�7C���Ŋ�G��/��x%�/;"�Sx�~��nXy���ܺ�E����L���4H���̛.0��&������P��`�q�!N	<�Q� ��ȅ���a���ض�&]��y����DD�Y�s�L���~n��<���٧.\�v���4��_��/�|��=
��	�<{�+�B;6�;,9�{�VbZ����6<�5D�]��帧�0�C���_9���m���*a���n@K�]��0�E)���c�P,$�������V��O�gJYG&�>9U�KD<���l��_}b�^"shp�qP��:N�<����ٲ(ͷ��tCԑұ��0lb���[�&n6��z�P$R`(?M�.�	I��i��3?�L)q�L����ik�4�
[�u��kY?��MN�b ���3�F{�C
�����t��������U�5k�+�շ~��'N�jϤ��e�Fs��4!����Qt�|�j_$����,Ȁ���qP�y�Y`�� ��C�TV�S=Nd'�u�[p��g5��q�����'���px�h�J��G1�j�%:�MZ��oc�R�K������x�{I�����Y����#�R��=	�)B3�G�a;E@jm��}wo��A%l�j��j��F�\��?���m�9�'�񊂜/������5-"YG��޹�C�H�9[Cg��N��̏@Z���P@�lL�Z�۸ЍR����&����y+��meADE�0�+�;P�B=#Sb���֘�U٫�H5�7�o� '_/䇄!ˣ�;%S#:�Ԟ���*�Z=�N~�+�\�]��=TQ��X�������ж�5o�85�!���_u�Ҝ�v�n������^38�b�Qb�?K���k����p��h޴���Y�0.����&��;����n����'����}j ]FD��|�A
���Y]�0�U=��nG8
!��Bۤ��eu�*��Xv�rޑ���� ��L�iN�ad��!�A���.�(��(���pΐ�'���� �/b��\�٪9�XAr"
��_0������`t��O�\�=�y9�V����t��L�}�	��MA�����x(-XH]�ڦ�6g�����o��TX�k�4��G�����󡘣�7�M|Gs�k����O�U�٧a��ej�e����ƭ}�7rj��6�p�fwi�5���)�|W���p���W7�)��#A�7r߬D%��i�1l1%�o�@�,j)���$�}ovޫ���n��ʙ>�F���M��9ƶ�وS<���Z�.���j����1a���]o�?��ޘ��Ձ�R5p�ex���r����e�2 !���{�w�n3I�e�'��ui��l.d��r�`i��&\Wͫ��{�:a�į.�1�r���f����_�=fi1	�rq��i���8�|_q����CY�K��ߌ��;�K�
���JO;B�D��t�!��<B_X=���S *�A�~wF�O��'g�ABT���������%=�F�I�~�M�>U�.��*|�s7�FW��N�t]���&e�����=u�l�#7�Mj�x��<�����@m��=�SxD�n��K�
�d�^�Ni J��=���K2`NHQJ����S	dɒ�G�ԄO�r�����{q���quB��d`��5���iW�t�n����A<�!�\r���B��X§o�|�J�y�3���8m�$���m
�^4�(ZRu"
/E$������}�0���l4|����+|��7�7������[ǈQz��2�וC���t#���VU��:�o���Ƈ�� Œ��j��Ӆ&NDI\E���"�߭%[bU��E1�񷫘����L �������yGíŨr�00��]�T�6�z1� OC����M�o�'��/��̈́*2�9�z2����x�<����:�KM!�ZC�M����ƫ$J���p:�*Q���x�&]�C�im}}	˥2�!H�}�md�tfz<o���1��聼T��{^'�[D��E�6�œ!5�烬�:�?�_Xy,���+�{�b9�R���'����IA>�ѕ���y�@�m�B�`�vf�44x(�5[t�3�ף�I�R�,���4��l�IU��v�_rČ�@<�r�<P���i��=w��Ͽj�*�'�{1�Cm	-}�l+���v���V��U�4<iP�8�j����ֺ��s�&�j���_\�s�F׵ޤO�,�㹲��V�ӓ��̀���zc��Z�9G���e�mP6��&�����̟B���$�N�7"�@����2~Q��Z=��J���p�	V�}r�s<Bz�o��5-�|�hu`�2��=~@�ͺ�!��wެ{�����C�)�����t�\чgUmO�J��g��FD�9�2���S�^ܨo���Q�����b+%���#,wl���Iz��(a2�E
���F���A�j,i�_�{x��n�K�s�Lmz��Ψ�˺�r����T�Ы��E���ӹ>O���7�'ӈ�mbC�*	�E�)�v^��8�M�v�l�7O��>jAʺϦ]1�9P�v�:��a:]��!�c��gE��ı4d1~oehs���P�˸��t��������������� ��9s_.ǐƀ���w1��J�;�Fo�J'�*�p>��P����.���w��r�Jtd�j�j���L�â��� U"w}�<�c��9�������INǴ^my��flf�Wz������ݣ&�J�ϻ���t�D�l��R}���{l�Y�<�6�!���������9�Q��O�١o/M�%3�(���r��2��a�0K
m�q������j��A����3�m4;֤נ�ԫ�Kt����'AP�`j� ���� |O�����m$,M�q�%L��Y�z
D#v���I�c�S� ���O�a�F�
����G��8�����XN+��j�
Y�ע�	��%�ѕLX���J_����m������f���ۉ��^O��"� `W(V�^ՠ^'�=)����F�`�(���ģ�|��l����h��f����*�����M��#���}+��IO9l��W�H�y��-6����
�����,�L�X׵f�8F���O;� �t2��s&�5�}����Y���ؒ�-�7��"b�H$��T��z�.'��B�l� NKl�(�%�	%h7�(1�ۭ�y��v�Z,�E#�dt�D#�h}���RI"�b� $�K�3��
q9Ok𳆭N/k\��i�X����,�"�s̰��������q�߻�əQ�f������_f=�]�ta&��Δ��T
'�#%�ͤ�5Q���������y�Ak�MA��}PB�S�ȑ��I����*Q��Q߮�J���293s�N�����[~�jHHL��~��1��(O� W�i>M~��;�H�|:��aú��d:g	�W�ɟu�PX���U��̪{���?�:������=>��Ih��o���~Yso40J�y�NȮ�+{�	l�2i��y�u5 &�.��M����;�#�ۅ�k�֌�Gl
 0Q%z�k��X`�a�\�E�U��X���R_&��w��Ғ�h=�U�tL��/���y��Pv��B��� 'g)����I%d��Y�6���Km�;�`�ah_0޷��uQ�ݘ��7�EmYe�ɫ6��uP��(Y��?�����<W,2�w��s/C ,XV�G�_��_�}��|m�<}�`�X�Ҕ�ޱ���Z)ĭ�^�o�
�����̡q��:�*o0�B��lIJ���+�J��S-�`�BT/�Ig�F�va���+Z��Hq�{������J�]�R���-�ww�}<����ʏdf�}�}͜svڲWfO�,L5��?�D�V�Q0O"l�$-�1�>Ыd]�O����sx���l����4��sw��N����$�0�#������.4L�v(�KA�^�I\�}�X�G�t����10�!�4�O#��d��.�S��@n����ZR���;� -�9�bf�(30���ԧ��ڜ��+��e1�a
٣�Q�����9ړ^1��_�"��:6|.Q�.�u%�0.�pP;d�oWK�?��֛�w�tii~���&��1�'yT� �V�����_����*���s��,o�˞���[�׎�>�8��<<���ػd��U��� �4��>�o�����Pܬ�����5��4����%�@!���aKW;���a�R4���uֹ?m�#�����b�r�����n��wl���� �ۻ�ϩ�H9['O6��VϢ_� ��;��L���;���P4�(C���R�"�x��i>�|dY �?2�F�>y׎�Wy��m&r�)4�B�|�(OUIR	ە�����)Ə�zO�$�Ԫ��P*���7T/C@]W�b*լ*��B�ތ��m<��"�n	�A�AC�
|�J�0���������#�fL�w�
`�!��(�`�J<*�׳���c�8>��@��ٰ� ���
��ת7b�tR���рy�~��+b�Y���n��;շ����?�F/��k)�g���tԩ{P�Ob�Ϧ��|n0t��r�i7�i�j�ҡ��VJyImQ�v !��uH�/�u��-3-�����
���1������S�E�W[�g)�`��[�^� �!H�8<g%�J�j":f��͍ۀ��)���v�_rܑ ��[T"0rb�'ez���咅������O���7
�-$�A_)w�;�Cj�,�͕Z�W�{..�YU~���;�)��Ģ��ǏRdٚRd�����F�"g��Ӧ�����{����q�������ęɨ�7�ˢ�ۓ3�
L��Bw÷ц­~�=#.�B�����9�}�
�lz�
��^�1�ڌRЁ�1��`t�S�#^W�!�ɾ����9�a�N��%���a�F�QF�*�J�li~�U�/ (T�|�q��,K(��2��u��}�%M���V��)�6�B�t�d����L���S{�Ca�R���������?Fؔܚh9g�� �ߧal�{�cv�\�#���$���3:��fS|ڋb���:l|l-�O�g	��,s��>R����G�Фv���L�a5�� ��Dl
����[��tw����胯�ad���!e�:9ȆEjZ�N�x�k��3��cK�WJJ�1��Cz����]"���J����4P�r�2�s��7��b�g�ӈ�5m5`��,uA,3���| ŖW+��zCF_$������������m���ӴqߓE.U��<bR���*���̡K���c���=�'��'���Prz3��J,�(�w�sk��8�9�����E��8(��,�&�_6� _n����d��/���5ڗP�[[� `@ @�5��p�"�\���N�T���@�+�9Kf� ��
��'�5a_Xa��d��7�[ډ?F�4��~�~�MlϤ�8��o�VtJ��}�A�D9��Z�
._����n̹��g�2��gw��K������P*܌r����1��Cw�bi�V�L9#�w����H���3�}�r$fpLII����,_����z`�h��Bz Mg�Q3��pC��-?��E��$���:K��C����^��T-Zn<]5<����*!�k���(U�Y;{�-������2]�44cS�R��w \�܁�F`#�O4��-sMF�6�ߵ�=����T�J�_(��}.��	��|����՚N�^���l��/�~n�*�
8���gv����t��*�bP�LLj7�^fk��Ws��_�:kژ8؈ʝ��;{�{�L�҉���5����[X�x�~�{��}�����ݓ���˻D^�GTë������`̊ն(�'��B��«�U���y7&��pn	3o?�[�zed��\q��d��p���J��9�D鐊T@
�.�88�絙�zgS�j �-v���f:��-Ugi�9��P��}�=��;	sM[�F�27F!Yh��ي�9��]�/	�o(��������jMp��?����)���I�"�}�n5��Oo1ۿ	�/���F��>ib5;� �;c���^J���Y�L��<]9��o��E����*�g`;���2;iE0Z.oQ��R�d�l�~>s*&sHڨ秾91�LLh��&ݹ����/��>My���⫉"��ܟ:�wRJ{�Ч4��@{���o�+�3�L?Jp%�j�t���a�MǛ�Œo"L�k���]Z�Ki/�Y�Lg`�;�A��f��Y�ݚ7����ؒ->������D����]���
���'sr^�AZ��y��H\_1z��f��K�L��^������͐�dW͇�ɹ�
_��?օ��o"�=��@��<�J�I�0뢄Z���mtI�r�����1�ŉ�N����j�''3������X:e�+Ǫ����&�?\�IB:+*��Q�cI�J^k��0`�p!M�+�h-5��և�3�@DI�?FYaҿ>�0@��A3T�qS}qUI�Y��ëI�C<�E�@1^���>S%�����FQ��V��f���G9s����̭bI�jf�N�ب,}H�iE;3��t�y�a!3	rd>m�*��bt��*hl,h�z��uY�"8|~�\%�%<�&̖����s��QtX-��>d��<x#�߳;�8��_�wPl@��Ap(BC��������&�L\�w����.{�����>����m�e�!l�I��$6��!?E|��gC��D���s�������k���E'��a���z
[�x93�?C��Za�W���Ը�<�p�Wq�@��\<�Y7&&�(�]^Q��(�{s����c=(�Gzan:��AP����eK����m���~�E��֟��QtZ♑�_�z�iM"�,�j���:Wk�''���Q��(��k ���D�� |����4�ת=�7��^�8�c�|��oSշ�ry`�lN$�	$H��hVRt`���[��à8W��ʢղ�k*W�V���V��6s{�¹V�O ^�
.>���J\Q���rч���%Nѧ������M�%I��e�PG��E�/lR�}�(�v�L���[�C?��h����K$�E�Y��a&��\n�hBa��%�����:�f|�H� �sU�b�K�\�G��~�T!mg;�՘h	�V����b.�sr~O\�qa�z܌w�$@ة��:�)�V��(l(�MF��Wl�"Z�C� ��z�<m���o�AU >�0Y���2��x������o��8�4����r�6�z�P����U)�?E���xp�h��3�$g�FJI��ܺʛ��Ib�Sv$2$�/�l��`��Uӿ�B@�ϳ��j������v_���F��h�6����w�P�Z�tM���%ɽ��o��M=ʾ���%B�ˉhbAܠo�y�e%��b��P��Ʃ	�G6@��W���"�
�J�J4�Y�غ���Qa�]�oU_=�k���o���k9��"H��-��.�8�M�$B��5���[}�7��4�POa/�E�Y:`d7X�U�RF2v�+�F��*g�]7T_G87���Q~hw�����֜F=������������x�5�DC	'�v�ʰ@�
#���������NR�N��Ϻ�TJ����?q-9YB�mW�}V�+'**�*U�}�}u�9�Yt�Y�ELDELz�U�{����Ц"��xJ�y�؟r��s�;����0����䨼R�:�W4��˔Wt��S��	�RO8��>�ަ����cc�R�%m1�~"u��%�A�9,�����+���,w_�=�[X�N��v�J�ݸE�;�/]�����X� �W�{�\S2
��8�##](�y4��ŶC�{�7�x+�%��[�G׍	:Lĉ9U�`�p��B5��%�?���T�Bg����}��.E�WN���Z�Zh�9��<��u/����d||v\-s�/��r񻸰�v�M�*a�r3>�b3Q��i�lRK3b�w0�{��)�(`�n�P�d��^�*�y3ݧ�q!߳f�u1C)K_�,O���n�tr.Y��`��a���J���~[��`��N�w-��0H+���PG'M%�J�.�!���98�cVL���"�&�������_�0�AM��ɲ��Y�!��p0p�����(�Ŝ��t�4��vDX��V fQ�i3g���!Z��Ʌ�_����V�)d)w~'��F�
˳r��"mOC���5��Rl=$[��k����]Y_*e����1ܷ���Io��Rͤ�㉫�?�Y��ļ�e�b�'��*L��k���+e�eV@����6��1W��ʏj�ͦ�Xk���\t��~jX�y~jk��m�m�����>p��
x��Ľ �dc3Rd��~�2B����A�i��k��C~���X?eDy�1����������˻���.Η�\��G���Ӥ��_0܋?7�Y:>�%"�s�eyy7��ú7�^�I8��H���oߚBXSkC�����e�<J���/� Dܲb�<�">� �8�;�_�Ľ�?hb�U��c\�$	�2p�r)|�j���֪G�h3�V�q��֔ي�QM�R<m"�E���S]�������xgbom����M��h=?H��8�weZ����i];n��TWF�
�T0�x������z��IU>�kf��VpU3��b�������;˖
�	 �*!��D����2�0 �+���@x���zyfz�Ȕ���#O��LG�|P�,��T��bR�>� {����3�wC]�de5���a�6�ȳ������ܩ���At`h0GA���7�T�t�,�:��H���@i�W�aOGO�r_���$��ۖ�&l�H���]��S��x�B��3qHqo��ܦf�aY�����6�H�S�tq4uF�����~�J����~�qɬ����Am����ȩib���q��_�1��\��d�@Ð@L�5�C���J���I�L�H.qjʔ��~�w�w�g5]���V����q�n�XVk��F�U
�y�wf�#E�/��=��R��T����ڼ:I<'�K�X1$ǟ'ܤX�F(wC ʣN�_쩴��ʃ�Uh��a�eg����*ib9��u�{zx��C����VxG/o���1�pu��*a�\'WV�8���ih�ȥD��>���C�7�f�d�`\�ѝ~67�;��I���0d&h��� �m46�]I���NI����� �_hש:��sJz��t cdf0����X�5�v7����i+����Qvq��j<].&|�c���Y����2���wV�A���J�T�nH��%�)��s�AO�J��6nc ��2��tunf��B10m�DGd�?L�B�*�=���-����^�K�?d٥��D0�S�B�orU�w�%�{��ih�&��h�bS?��p~6>�ߛb����;���o�x��"�r�9��Y����H~�����?�u��p�/:��F��T��������2ݓ���u.F ���$Ef���FIrB��z���.O�*�um�U�P7I!�;�Z�rL��P���0FS�x��ҟ��"yr�Aܹ��%"��_-a^J&ն�gY����(E��Z�j<�{6f�`�9��Bs���<S���)�Ƹ�V~�P��j�1���%���yr1(��.��(Cű K�]TW2kM��,KH�y�$�XM�}"�y�i~�>@A���"�5g��=���Q�k��낤���t2�������2aI$�u"��LսI)�.�	l����q��߳0��PR	�ܒ�42�K�����?� ��mR�b��hdH����Y1��)���� 7@�[W	�/��[����~K����>۱����R�&�Ne���Ϫ��D��������oA¿���V��hY��\aF�>xB=����f���h~wM=�wl~?y��s2�ÏO�Bk?�Լ�x��'�tr>��@cZ��Z��\�W� �=�[|۲�� q��|a�qiE�0�`���Ǣ��K&,U��ꀳ��Q����f�9M;B1N?%��UN;h+a+D��K��$��*�1
c�.Fu<��6z�;��OόZ/��/2[�/���w/oݟɍ�~.�e4��R���*��D� ڡ��A#�S誈�J) �K�wmq�͆�p8lCh�ͷJ��hs��� zV�b�i2��'}c��[v����=�kʼ��t2&�4 4(��^{���}�P�z�Zه�?��׵c��J�>/f���9�\��fx-83�=�6��*��/�wH�����L$ɤ$��o�5ҡ8�sW�h�������p-��k���V'����X4&��þG���2���5m*c�C7���W�6�'b}��ě��|1xu��kRs��:��0�@JK�L#BP��<���#��la�4��{7U���Y�"Ȫ�t��p��!E���gQ��d��5	�|F�KC�"�HHϊ�c�ZI$�@��3���07+�����̑0+��*��6�� �I��ש̩��ΥLv�����z{~׵��ę����':&y��r�,���C&����u�*�B���E&� ʅ����}�`p"�Q�Q��)��1�$�� };iy��aM��k���ǰ��9�T����L=�>���Y�a����d�̟_DO�/?�b�t&�{�o?ڪ2e��y+�rV�r��}Z��0����#���r��l�VsW���6��L.{�^>��-�qi�VjR��l�+�Ï�զ	 �w��ʤ5�d`[l~��]�g�K�+�K�$,�9K�4�(	 ��Ú���%��+ĥ��.�0�; ���%'R�Y[�g��y�F�J �2��/��5�Q�*g�X��]I�g��d��O������.�R WD�����Tn�$]Vڸ��*��ף�#>�ّ\������Hmz�ޞ���`��ěmV�ʦ��Ω��c�͕�BXA����hXgm�Y*�8'B�Y~����6��RA	K:�F���	k��W�ى����c9�����s/���c��S��[w�]��2�3���bm���&;�`���Q5��r��{����˹�Ҩ߷hMp�Xr\U�*M�����r�Kj	K5��Z*�e�v����9�*%!Ϩ�m(���M鼳��ihRX+c�����PD+�&X ��W�x�ߢ�{���>��EN"uO��������&2�l>����"�
�g�QT�3̗8I8�q���Ro���>x���VzR�JDɵ��mj�n,�O��$[���V��sR� ���)��0{`p^����!	�׋=ɡ.���@^�#�0"a?�3=\h��Z@��q�9p �S�B~��Ou�=~	�q{��oq�R������Ӝ袾�W��yko�)������?w���-�2>Q1�}��6J�QJbj�V0�#��P��M�LJ
JD$�U�YD��K�������"�Y����5H��b�~�b�R�v�6��66@�R��ӿ�o6��v��=9X7V���A믑��gDOcgG}A@�M3�5w�`�V�eS2Ρ�f����"=K�qB�}Z�1���`)��ȼ����hg�J�g�To�6�R��J`��e��d��_T* �����(���%�AT�g{�9���>�fI�9<rN-n%K!�V�3���Ù��..$ه��܀*�r��WTψ�$#:kGhv�AC��뾁HIHͨ��
-�����Z����d3^yj6IUG�Y��7���͂[�n��8�t�F@��t���3���l>M�Ğ�س�ǧ�zн���7����uwݑ�A�PQ�Kou��P��&��"��W�ѐnTd�g.�+������*iq�K4�6HA@�fpEcҒ�/�K�îS��G��{j<�&���{l?m[UmR��"��������%�uj�˪ihJة�m� ���2��'�4@�?85��#9Bh����B�[V���[�y���RTz[дP�mf��2��wXD:ȸ�m{����ȉK����M���'<�ӛ�>������������76I��W�tQH�w�8�+�0JJ88�ۼ}�r&��+y>ĝ|�7P�Z�/k�#���0��UH�xNС����M�oz�آ�����͢�$5I�g���.���"�!���rH�#���e��{uf�~�I�kC��䈃�����`?�6z�r'(%�q6��;�m�0��ppPX��DV�`g�˂"����t�ד������'��ZGT�ճ"Շ��o s��l�?�O�'r5��	�2҈.��h�?�\.����}�}��8��n��Z?.��{�[z�^�Oմ�Li��W�+�TzB�8eO��	Cq����a��w�CI"E?�|�KQ 9�Z���H��T�k(��O�zj�����/������o��W�D��.?�^������~gEK��$���Z�"�A���9->��;��p�[b��� 2=g�B���i�6�������m�a;�(�=rb�^�g�{=GO;xS:g�Sҙ:E�d�KZ��8Ƣj���yHqT����7S7�l�t
����f�kQ�g*Ϟ1��$�b4,�����|xG$h)��Ǆ�^��T����f��J�z�Y#`Z�j�"�>3
�=�3��M�|�Q��Re���:��S�B]�΁u�qR�hJ���D@;�#��S�N��h��g���[k,h���9���n&���֫v�Y&����(�ӝ{�f��{���Z���s��n���?�ө��}>���>��g.̳%ֻ*˳i��'�	ؠyk�
�̂-!�J��a�����A����n�ۧ�1��_�ZE) �"u���<ԗ�^��i0Z��/na<`Ɏ��q#�?Z#�w��صw5Ġч4��V������5C��y�������o�;V�)^5{�]l�-%Vg�9
�&QF�'�&B�7I���K&u�w���=��v�=NΛH��e�J�y[j��>�e*���U�#��L�n��w�3���:���'���Ve�
]8��絝rm���vB�6qE��5ƚt�O���p)�)C[�OtZUM��e�w�]>	|��HZݔk:@jBdg�ə��6蓃�־`�]9���A[ٌ��3\xl�L�Ƴ�*�9�����������"=�%OH^m-g(O�`���� ���2�Cj�A=�qF
u����J�)��h��~�uy�H[��~o�h������Ǳ��.�"<B�F�v�l-)�+s訒�/(��+ѥO���L��/����e&6I����vgj����\C�*�Z�cN�MÐ��s��5S��wK�1wƤL�Ւ��c�?+f�w��Q%��K�肻�����2���>^�P�R��(�q�Z����Yf,Xb��8�3�զ�S����.ؙ�P �������
| �$���`I�������ď�z�m�:�x�C��?��Z;��[��qe��;��������V�k��n�.��I��*�;.3z(��Ĳ��[��b���3C����Y���s��	<�Tuajy�dQ^v�?����f/ү%�Ժ�Bp2��D��N��VpX�՘)~y�1y�γ��Wj�D��xs�E�޳Tb���?u���AT���
�xP�ߨ0�ګ�c��n�(��l
h�̒H�U�=��?Q��@	Y�ۮ����M4�$n��,>`:r]�zR�|����	�2�礦�Ȋa�h�b�����-�Z��р*���A�L�bl����t�% &�п�I����E����`��Hz�_+{f�W��x���2�ؖ=��<�_�Gth �Ж$��D��o�����نY�:�n�c�}2�����G��"�3������^�G���'T�6G��ԫ��+��KK�����������f'����]�)>0>�ΪʌP�j�eΕ\���d5�Q��>�z�����'S���F;��C�.H�Y����n��7 }��{Z?�N��<!���Hnr�_L)�E�wb�ṥ����B�Ɇ��lז�̪۫s�7�����,��ɬ���!����l��F�\V��-�M���	-��;�>8V�o��t�U���D�t�[0�Pi�b��Ke5UJ �!�u��Ǟ�l�7t6\�!�p<3��eg�����K��]u���ߧ�l���q���N�l!��&7�#'/���(Kg�پ��3/!�������i,��8�%hf�,а�C�X���QKi�*���P�?=�.�o�&U��Î�����q���Z��~�呺�9o<������Ղ�fW�\|�a%A �f���YƷ�6�h������v����ђ@` �v5d ���s�@�:IC�v+�َ�XK�8��բJ� 9b�d]�.]_r*��ܸ\B&���j;�%�&�s�f[H�BWn�%�� ���!���M����SE	�J�Y����pL ��Ibb�����v&��a>�᡿]Q�X_�c�jb
j�~�#DV�G����c�J%�O���~�}�����YVٟ�6l�=����)x�Dt�d=��^P�����̠h��o�3�ޔ��jI�'��-�"L|���\�����~�������I3>�8O�A��7���RǿO�y$�__�m;nR���ݏ��3�n��x�.׋��6��LU�S�ۦ;;g����U���g��ѳ��c�+i�7F�k��/2��Զ�ji�Ň�L�n���8�p���S����2��k?�����^��T�CX�����Dx^��U��`g�	ϣ�!K����?� �v�y�}�w�j1�΀p�ewe�A�AR$(�d�Cgk�Za�*`�ai9�q9�
9e�v'�؂)�n���S8����ҍ뷰�M -ed�/�FW�����\%h�9Ѕ�9;��V2�+u��aK���"�:��N�TR�NiK�:/�!����7׳E��Zг0Z��_@�>^��|��<HK\���d(8]g���c�tw6��'n
��c������Mc��(�ٿr�0����G5Ք�0RY�z�ī���߼j}�ډ+s�h�O�R[V�u�T�&�S���6��Ў������oB(�����T�������	��������͓��{Z��О֙�>%?�[\FDz�t��#F6�T8, �rƮΉ�NL#a=���sR�_8;$�~�����%gv�:��*ݾNv�4N�^�n�?Ulk�\�+6��t�?z6X�g���R�\��-YjG�+�Q|�Î�k��*�	l��EҸI5WкlP�R���4q[�K�n�p�&����Y�v�Ee`�S�Dl�#��o��y���m ����p�w�,�Xf\Шp��Mkz�����a=����X��K"Yb�w�	�\�N*�X�[� �xj_��k��5y�f^'db��G��;P��Z׈B��#XaY�tN�@q����z'��v͜��Еl/$';��	A�0��!��1��)1��72�V�%S�;��^����:�� �9C֊R6��/��e�f�T���e�i��rvS����k��3��./�M�أ���b���lw{��� *��`T�������P����iį�~�9�)K����p���� �M�-L�ۺ�[��bj�F��_��kCaJ:y���;���@��ᓪ��ZMZ�a3�(ͼ/�D�b�_��K�ʒ"���2�c�ҙ���~���/�vy�9:���>f�8Cb\
��������q
S|�>�Q��u�mR��K�}��<�oM�9�:^�e6��:�}��Ҍ���l���g�Ĕ���L|��-��x~�bi����Sя��g$�8q�}{���:E�p��/,☬?ِac��v2�V��ƙ'':��i����7~��~}h��"�%dy�c ��7���5�|u�+.���nnj���<[�-��m.�?ڞ��w~^ș��ٽTztJmcZbo�2?��j����}�s��N��9�����6��"���X��p 0@����t�SK�9K7����i��|��ě��ϩUu�SH�{Ƣ=� 슾��<Ci?*	2�j�����N�W&���7,K���������;\�Z�rs?��k�ہ�S^R��`Z���s�@�x7���1|�EB���9�Y�����J[<{�S���"�j�/A�n����F�������Ǩ��P^��>֕9=9LNF�i�Y�Win*;rN+@�!	UdI01O�P���vWۭh��A��W��r����G��_&��p2n����{�fY�8�;�.r�����DB����ɒ��R��Wh�����) <cd�=Ln��H;�	BK�W�2�?a��ٿ�nz<:A(����1_�����.ƅ�>}�]���T8$�5X}~�(|�{y�Y}:���}��6����[I��x�W>f���ݛ�~��78.��W�FC�.H�3���t���M;�A�<&�@g�sP�L�� U� u�?kL�߻#N쭢�o��-=�� �q��mR��ps�����vbKYv_)8��L~���������y��]�׷	�̧X���~��^o���Tgm�U�mn�(�쩕��-��+�T3��Kv��x��~8&��ٳT�:�5iB�-=_}J��^����R�2�e���^�2zI�Ի�_���डrSsB�ٌ���z�Q�䍎�#�{��_܅>�1[O�srh�ț&g8�"������_����v���cWq��<�3�
�1��]���<�L_�R3�I&����F�C�T�Y�zX6�Xv��l�~�6�|m�o�s�0y<�9j=n�M������j��>9b��t�n~��8�]*.?���"7�f����xB������64w�ܽۚ���׷��D�<߀	=�(Ѳ8B��b,Is���?��$�V� �����W�Hf��Gsa�f��O��
&	8Uh���3��~�7�Έ9�$]�U��<]���l����cu����K�:��=�=�y/�4]!ݺ��C�n݀���=�%���w*f߫	�#�t�0��P�@�=���C�&�'{l2����5��I�]ɧ��AJ�暈G�3�C��.̸K�ol<���+5&~��a�;�I�ץ%pЗ��<��~��O֐����鸮� FNQ��Mީ����To�-RYoH��:�:�VwK<�H���L��G��5����aDs�#+>�T'n���g��Ȍ��t�o�yʌ��7I�o���SaS@K��[z��N���������Ʌ��9��^&�����ZD�/V{�p��><�?cݽ�Ok8�xj�=��0�����n3�J>��uO�p�Z(�R��\��l�G�����Z�i�Q����٬�K�6�H�?��8�	^ٙeZ��Lo�-mD��(���wû3	;O��ǥ��5�~�)����f���
�����jtT��F�vLZ�q����h)���rL�H��U�i~S�jy��C6���^m�N�ګ�W!��l-�ļ��ص@0��7Hڿ��D��l�I�aH�-J�:%����lQh݉�R����^ C�iaUPR#�n�4�h%�5�	.sR���`�l.$���#�$����4���y��}�:�i1�( p�ԤYi�Un�x���S_x+*	�[0��+!�@��13���^>(u=�;=���)X�<k�t����NL�f���w��3�He���ג����_R��/������C�� ���4����rZ9��`�Ϟ	�)'�ʼ�%
�%E��s��mm��(� V�y�zש<8�
-�ZvM��V�O�4�qπ� �?�Bz��<=^��z�ɷ��mΝ(;�������26�Ҹ���5J���ˋgË�7�^�:��{��f����ª���yu�
��Mo��˪V����������p������du�o��*�xg۲���l�a�oq�h�ɦd�� �1@6�i0�����x��yl��1�f�/�_����r���`[q�3@�̈��%�2�#��\�8���&��v�4E�|[�w��\�@<��z_暡"z�B)]Cn���YP��5�ߺ>�oѝD�l2��HQ!j��0��39���ձ����J1�)����è�)����l�d��b�R�v��ª`���f����H�*�OPU� Q���R�x�%�o��z���K�o#T�G�X�����w;�r5�r�9��$��Ϣ�e�>��b:������Nyd�u�O����z�N�T������#Hr��M�}l�-J��p��cKd�b�QZ�픉)t���ra ���z4ʽ�`c�����ϗR��xW8���}�}�}�3����~\��m��9+fZ­+��_�i�ә�{�z�����[�e��G;�3�c\��?�	1��?cv�|����P������^��qaC�*�;�e�<Y ��LI��%���,�m�*V���]W$oV���/l��tfO��ٻ�%W�;4��l-�W��5@�T�&~��Fs7��|�p��*$�c[�Fi	%Lޤ!G�*����i�'�ų)��~���v��`�H������_�Q��4�9g\^�6�w �jQ-�1�Ĵ4@�3Tq���%��ph���~롓�_���6ud1Q�I��D�s�t'w󬩡��ԚBJ%��Au�c��]�]ͼ�K+��ϩi�L��ʗW��,.3O���K����F�D�`�[хߪ�'��	�p���G���%}���+�����-K���`Tv�Wa�UU$�w�� F���o
@�7��)��t7R��M2���̥��.�bw��i>a!��h����^�)ؑ����'h�I�L��v�7m}k�Ȁ��sp���ѦAG�xJ΅��d\Ӎ�#�Ե}7~���H9�(�>����,�p�$m�S2V� \�qb�ay���lE^�W�`���@�X����E^^l7��<�,�͂W�W�[B4���b���DTAG����;B~�A�x��M!J����,�4�^���~~uIN��o��-.����y�,���57G�32oH��f�xyo����^�zؚ���xS��rע��l�c�W�UwA���|�jԘ���Sm9\�9�^RIcD���|'W]Zp���;њ2�9�D��Mm�J�'͵���.�2w��\vU��=r��Y�΃s�v�+�m4s?pXa�!2�}J��32�A���������Gc�_+�mܬ�И���CJ����?^���S�R@�\�?�=$����(����W��1�Bk���.a	,�n-�q'�B��d�%�}뤸tɭq��@�ͻ�Q�K,u�*H��$�����M:r�K�7�𜰚�H�ڡ@aS�L4tGG�y�
������[�NŪ��V�g�Wb��d0��������jV/m���p�����	b�ty�l~簘."0_�RIZrBt˹�����������)�ƣ���/�a��Qc�\�$+�W�r�,,��?R�dJB�i�~��?�Q��-VGi�K*F���T�CA��R��-s;^\6rW�����,���S����@$�9�2�Ü �7��J�TE�j! �S�|#�'0�`�勲���� ۔Wu�N�������8X�"\~>��"�(�:��CE�#O���"o��j�kk�n>,���O����.��� Q��c�jq�pvw>싪e02qv��>�=����%�p�QRQ���
�LʲC��c�6j�m�ʥ(�Һ�%;д�����Vhw[��0�� A���/z��o�Nq�q�覼���K�ybg�f��1bDW �Y���d�5�t`�i����a	8��=�ts��6�)�@������iJ��ē)�@ÌTC}0��5[�2�Zf51�e�]$׻Fo\fmH�R��|S���X� ޮ����/iN� ���sL/���/�/7���Ͻ�����/������*����oݓ�Ʈ��{����N���#w�`E���8PAEZ^ ��S�����3��:��hK��N��\Z9
�$��BSV;uc�����6�nm૿��m���m�]a�o�s��������&���b̏�V�z�,��s�����*&DD�#��1	�p��Ȟn��#���x�`�kT{��+lp�6���	�/�OC{�xհo��q�/�	Ì��,���Pbg��CD� �)���M��ęg& K%�m��kS]���MMf	~�����R��1��{h�,�Tc���t�QM�P` ��"ҽ����(�5�Si�QC`0��fH�n�������9�g��l{�x=���z�{���Ԃ��,����N�Jj�|4�iV&Hhq���e� ���~6/�>D[�t���؍����T�j��\)�HB{���b��������h�v�`l��h�b�)[��~��;?��B�h�f����!ͽ�z�oѱ�M)����q`�&f�����>�L���T��YK�q���0��L�sX���ݴo��?�l��F�?*J4�WX@�Yl��܈��c�Wm�f�MZ��זּ��i �b�u8�Z���V�X3'ڨG�s{Q��
#@�v�:�ѳ��I�<�=��;MP�d���\��D��I���$�2��o�����0���^x���%���-yƧ��+b�O����/�P�g�ٸ�Չ����~�d)�`ՉV��[��������[�g�X�:�G������O	��x��I����\��xzDj|f��p֟�ַxM�`��_�#ϔG@��Ӹ�D�@��2������X����_��vU�<�%�բ�g��NZ��B�HH�^�����l�:]	JKCMx�!�`��ʷy��ʢK7yg�I
�@>�h��ERp5ꭙ��ynL�2���7���'��4I��⠺Jx�?��/%H����X�F������M�KcQQ�_�.ͯ��k.�k���\�^�x����"�=�-9:���.�NLM�/��9��x�ʯwq���͏g�d����@�r11���W�����mǾ��R�_@�� ��7���_��
Y��~�e��N�Z�8�#�X��2�#LzJj��	A�A����q&�}{�b	+u�M�:	׻�~�/��4�f��	���)�	D��4|��]�󆊡"�rȷ[$1)��^�ɡW���s��1���@tx'�����y�z�CӪ�'O��oל�i5A`�D�2Mj/c�	 F*!ɞ<Uխ�~�?u�	�~,�C��v_K��(�7�M
vM�Y�h�V���
Z��SA��ҸD��V ����V}[|��J Ҝɰ�Y��$�Ɵ['�⭠���f.x��V�K��{K�;�/#FQ�t(ݩ,���ω %�O�6.w��4֊M�iY>W����^��=C3�ޠUZ��£�D��;E���vi�؊JM��W�����d�|��+�ka��(%��t$L����%�&�=^9���W�Ez�a�{&�&潄��M`�Cǰ3Ϣe��5�,���F�&�6C��2�
�ʡ; �(��� P����e��5��9�E����R28�r�	L9G}��G�8b�Z؃�b��'<���/ݷ{ކ",3��̿����J��S�G��@�������O��1W�-�vM5yÊ����&93�W�+ew������~������W�>����������2�v"�ꄅo�G�ͯ'�y]��O.D��<:�n�r��@L�7���}����:��>jm�d�������έ)������*������Sĥ�h�I�2Z|1�������X8� ��xS˅��߻������E���s��g����`.�Ly/8@R,x"�}�*��;g���Ą�@�z�G�.Z���]�2t H�� ��1)n!*�>w���oEiZU'�E=��"7���أ�&�Z(c)"��^#�4z~��z�%�nx�� 9�ڃO��$�S�"釃J�FFGP	`�m���X
����@(��OE��nB������ǂ����H?���H^-g`~*�ɉ��pFޭzQ_�M3h�����)�%���Z�gS���B�/[j܎�7�J�\����T*�_�S�O�����Y�tK�
�w�/7��"�jD/F���9v��>�^W����ҽ؞�۸Ԝ)�������R����5�<�֘�NV~7K�=�ns��Z�Q�K� G�X
�R��v1K�]�_'=au������	넫�������u��mǯ����2�4D��q�}���*�h������|���zc�jS;X;k�f;Y�x�X��e��Onp�����UW��n�;R�M��SȖ��O����X��xOp`��U�%�~��= B7���p���<��Y	�PX���{����ok,|0��4K=�KηA�=\�W��Y�-q��u�|��vz�H,^����t��_F�+��i�,*�߶��/����C3����>�VY�iW��+ �H�17�ECXL�t�.�7�	�,|�f,�J���:k�>F5'>��I���Vw\�︈�v�N�签�������
����#*�C�65TG�f
����y4���{F��'��>�Lǫ�-Ą�s��2 ~^��dN��,M�3)�l�Ub�^�_�T/eu�J�՘I0�SX�"����
�����޸���*�c}T�Эa����}����F%���U��+�t��_Z��PJ-��;���d�*�^��\�3�d=9(y,g��{���H���`s�UW��++`0�Nqږ�i(3#��R�������y��.��R1E���98��Ժ�h����\�m	��ջ$Kݕ��+�q��a%M9|����lS�O�4��e<��)�?euLr[V��d��?�T��"NkE/�u^�u���o�E�]̞BC�k�V������?�b�����A��|ax��g�h-�4p~�h���F��O��0nR��t�ܭt������+!�e���=#�$����c�K�d~�&�c���4��'{ U[V�l��gg>o\	`��.ŹuwXnc��[%��d��r��-�7L��Ս��������n͸S�'��q�XB�S�O�	h:����fVL�M�#�*V���Z�� I��Z^�\A>�t��@���H�8�O~+�XO?N�.?�kd�������G�z4�ikz�0��.�M��=�N#�}[��rd4�	�a�C�"It�a����~�p������[IǢFS��G��k�K3���7����<���~�Abf64���3�����>���3���g6�m���b��uJ�tL��\�9>���Ԇ���[�c��+si�5����8\�Q_Γ�)��k��ትU�͑���'�u8|��,6���r�m���zm�c�z_)�/�^l-��??,����F 3^6,�(70�f5�b������d�!w~pg��J̀�o�S�a'�=�H|L"ȁ��H�:k̎��K7	�N�}^������i���w�s��S�j�4��k_�����l>�pGuAHߚ�hZ=���t����]�镗��{��]3B_>}�l�T���9���rcA_X%�g�����7��EO:���!# ��q�A�)%�S�3[��H��"��hV��ќ����h ���(�<�y|�d�p�D]z�+N�"��-ۛ���P�%�1�_�8��L�7,�V��|�нز�9�=G��Ξ#�
���/�/�v�vgp�ч��,h�j���3���(�l������T�	T����#��J��9`������j�l�a(�j �2�����X)��Jy���V�o_>�㐘��Fσ:"���gG���Z��&{G�$I���_��>�N5��N0���V����9p}C"�'%�ſ=���{�?�}�10�w��0Z��:
�cxg:�ӊU=Ϲs�F}�JC�,�p�%vM�X��z���q[�����Ez���36�/���J�r�������O�_R�&(�&UQ��bH��b�qË�u��7��FX	�]S��|ۦ� �Mʷb��'U�,h1�x�`)�hD��58��tn �_�r�~�B[kD���S��������g��!&����b>���7���+!އ��m6�m����}M�Dm�Шq���b�-[�N�:�;J�\�n����D^0�Ԅ��ø o6̨%]׀��H �a	��4H��Y����1_��J��hC�������t�q�p���]��:�0ޜ6��i��� W���8�<�+�tO#u�χ��k��ޜ	M[)T�c���A��Ń��iŤ�9jZ�4���N����Oc�i���t��m��L�1q��&;��J��u0V���PaXzX=�>��H�1�c�����BR��oY��Fd���0��S��u~����zDI�+��*��{�tݺ�XP���A`z�֎�O�cO����dgx�Z���>F��1s^a:�����o�*Ӈ�����:��6:�)��ip)$ 8��SZ���?sDld\�#.$�_��g
�O4�M=y�1[�7�9}p[�5�)@֏��?@�~;�ڼ�ӱ&�o��}ǵ�v����o�˾(*0�g8ʟ���������aO���<a�~XE����xǘ�+�/�VY���y��@v�W'Diͣ�L��u�FU◷�|B��VJ�4M��Ix�^1pV}�L��R������kdѐ~���^����ӓ��rܤOT�z�@�WR�q�����+��
���y�hm���|R�8E�΂l���j� >E����X9�  �x�_���wkV�4��n��� ���B³'�b��ǥ�]�~z�|��l��u��[#"�pz#^&)�$�Ll�nL�s"���@w"P"��? �"��)	�K\V��"'5�|IX�b.�l �.O�gj,�ǋ�:i�6/��>���?�ڱ�;㺻P�}�۞)��dg5�+K��Vz*��i�+zD_S��:�R���[<�����2�����������'`����m��r~��܌�CdqqLE7ʖ�
^��f��8n�j�4��q�u&+6K}���Ԣs�N�#��=����sK�|��M�?����KV�� ���Ȑ51�Ӓ'C�������HO����w�S��9E|}�&�'�����j�l�9K�i�n�-���g��~%k,x�%c���|X.`8�Ù8H4��	���m\�H��p1�������X�#����J��uT�2��nb��DѮ#P��;ҡ��
p��WN)��8�Od�A��a�]+�E�Kb�-_cS��~��*��|df>5�+AR��9��^��0ҽ�����Y�!�ʢv�MR
�WR���7�h3?�������e�r�+��Gar �p��%�N@z־��l����9��@yVf^�C � ��v;�'8��V�i��[</�<%٩��aP:�V~�V��-:^A9EM��a����`�@\2���!�\��~k�j,n'.��3$�~x>f�q�cU�#W"�3Ū����)ڑG�ܲ�u	Zx���i�^[���ig��L[��"�[
R5�97����2�@@4�,~��p,JJ�n��<�Y�G�p��g���Ob.�_��V�L��+6��2��'[i\���Ey%�UK��`�v49Bv"��K����Y`ty�_��P x���M�T��}��	����O;���n?�<�3�J6ۍ��c;[����=ۥ��Ɩ�Ym�}κÒ����=W��;.T���TE��5��^�r�H��q�`���)(F;3���
<��
JWJ!� ��о��,��&`Bi�_ɟ��Z+�*Ԛ�Ѝ�<c��G�j4�	�p�_Q���`�"[�O6�Ω1��4m��EA�4��4z�'�Dkoo�M~b�x�T �:!�����ٻ3�'c����tx��~���"���G�Z]N}�_R2!��"B�Y`��Ed��[��`-���7�ߓ�ul�[�;a[H<�p|ENkۧ���3�����'%��aDOM��ERq;���%�W��0�51����l����*�X�:h�cS&Ң�c�{�By�(/4')��_P7�Ι<��x���7�,b��Ԉ����:�D���tU���R����X�_�v5|�E�X �U�W���F�����~+����X}C�t磸�߅��|���5��-�@���?�բ��ӹ�b��eS���=vm7#VĆ�R�����㐤�~϶�V��]���0��:C�x%M���
�*��DJm�.��O#���z�.w6~�F$q�1������8���؏�%�<ˁ����O�.����[�!�eL3%?�N&���Igt�q�l+䐗��?��7�,�i��@)ԡ�f���(�_Ԕ������S
����WFt0���?�*�#H��'��wOl��ԛܣezỔ$�����{��1����U�p�̋w�s�f���y%��t�Ru|�AkG��J��#�R�̉�O+�n0\;�J����j���wO�W���n/_�흷^���ԉ_oܭ��.6��O.��}��į�A��l��@9�\�ڎEP����P��\��At��^�yh��-֕� �|q"��r0r�~�ϯ96D���7h�^����o�L��yk�sn!6�q�;g1��L�A��I{�`4�`�՗���[������� IO�7\�뢾�~* �G�үWO�K}�U���ɥ�$ǽ/[яH=�b|�/���e���� �f]�n��X�Kp:'�d��υ�lV��\��	=���-_�1^D�=���I*A��VذU�p���y�Ya���k�΂͎3E�g�D�\+�w�K���uX���W&��*^�r�l%t��j����7�9O?�� Ц]6P����9�|˙(�Q�~P�k��N�B��4��.\q�?��0|O1�����Q����$�J}|��jD�ۇO�?��Ʒ<�妑�?�Q�~���!�(����뛜�]n��"2r��֮T���q�ɧ�
E~=���le��ECЊd�PR�_Xf�ݜ�=�]�ܳ�:^���\�m�8|N�v���l����.����� �G�]S��Î?�A�'�.P�+��WMؖ0�����gP�u��@�o�]]����"�
&Y�\��3�Z)t�21��2�Q4u�сDZU�q��~��_:���
/�3���i,�N�/_i���шw���'�����߾I���s'��P�3ͦEO�[q��O���jߐ��IwW��7ъ{',�-vۍ�Q�{�y��3,�/6P��(�R���Od��(��V�Y�s�/���K�%�����,�������/�hY7�"R�ク^ʊp������0G��-tms;�Q����}6c�g�Kȳ�M_Ҋ�%��|K^�Cj��P�*���M�ۼ:�V�2Tyd�ivcKiX�����^6�{���.!��䊝{��K�"4Y����i`����dX
���O���t0��S�D:
�u9uԃH}�(,��ø�����i�@QhBu�'��PٓJ% ��ʭ$ڿ`��/�(�_��Ȫ�!!q'��s(_���6��x��O��]3�E�B&r��l,ےޫ���,.�T8mb�EX�S@��ؘ�i��j\K��e���B�Z<��h+X�i.i��߻I�zq�*������w�������_�xFZ�Uua)\�1&yHOEY�y\շp����Ƹ1l1���6���z4�ߚ;��"$DS�ГC�;Ƈ�D�@�����S���ɳ��&�˻��*^�?_���Tx�栴�[>f^λ=�g�E�Y_N���Z����q�:��*�?��zbP����E�Z_ߖ�����5v��d��ߦBN�iBA�oH��Kӆ�8~�F%T��+> �8_�6	�1���v
 �Oz�p6@�Af��F↥�UP8�nSN��H��@b�6!L�b�Fa��t9�!��;�+,2Ui�8�>��/�3���x� �y�!W/-�֚�V�we��Y�f}��=��o����MW�O����_�_��'���zf{�&���w� ���О��\&����۷/u�~
]+Ud���	��o���Z��ՑS{4cn֋�i�4���p�qN�����o�fp��,i���3::Z������7�t��(��|a��x8���Q�����:���3_��q�{�R�"���!��yGM	Q{�dx�ښS�@#��n}�ˣ��;m�V�"��}2�a�d�xV��Ѿ ���k>�������(����0{�Z�A�3�(�_�H����7�7���9�lܣ����
RTǱ\ қzJ��e�z�9TU�9�@���th�x=���k�;d�f� T־��d��3�f��=o�{��,P>�fo%���������l�����oc��NU�K�Eyz�_�����$����Z�����ub����R;q�Ru��p��������$�u��$�ʤI��u6Y;��Z��p�Z5�Y�7�5�r?y�"%�� ���8�U���({�����+r9gA[��C�_��Ռ��&�a�q�ڋ�Zs9�׹�{�H��H[��J��k��х��[5��г��� ���q�CV��
}p~K�mf\����c��^�pa���w�Ii9��'�O�ϽN����9ꮔ��[���g�,�:�zYBH�+WVo��<)���T2*���BC({�j������Z����Ӎ�Q_�}�E��.�zd��ۅP;�"���k\�=���en�	�$���f8��;n��}b%�ۤ���B���l%�2��J��'tOx�E9���RԳ���C��^���v��/^�O�`��ꔳ�[X���w��x���堳4�+�S,��IH�x�=�L2�*M�����:W�a����"���zd�Z��Y��5Y�3;}�����z����P��_ ���W.�@�_z.\�.C��Ȕ||:>��Q1����6P� ��+#��!��լTa�؉���-�I��ԟZ+�T_��s!C�lf�ȓ���q��ͽ��X��/y��ȉ-�"Ɯ8%B?gU%��V4i4R�Qh�0�t �&%��tHeլJe����zK��������O�PC�V8q��vJ�S(��T���%#��_�Q�Nk7��<���	J5�7�t�B���� �uګ�ov�c�'��������#O(8\�[C�K���N�$�F�(r�_,��Gi�����aG��-%��b>��w��GU���3��ʼ��u$�(�=�9i��zB��(ٓ>���'��&$��zn��� f�	E5����,3�TG`��GgyY#�*����hzF��I~jv�x���i�5Y�!+҂�3�w� �l�	A��6	���@�$��B�-�;��|ۑڑ�9V'���z�:�l��@ݼ4��b�)�SI��Øw`<1pv��!UG�0-i�G�T���;QQ (l6��qxm	�Ru.�Iy�z��81���5Yˁ��D^> @L��\�|L��B~7/)�l�Np�Ay���q�&C��8jG`�1 ����oʞ���6T]:�Yv��p9(0���&p0/�s������@֗�	&.qx�_��|/��E�C�yx�;��4iE��S�C��Y�&�ҷ8%��s�
=Ғ�K������$�s�΢E;U�j�*�B�q�z[�
mARU��@�4�t�';I��(��iU��Њ!��}���*s# +M}��Tp%�t>=B�����gGΧW��'���0KXpT"s�{���V�+ÿ�o�g4�چ_Tq�O_-H��
<�w
o�d��|19Q�jW���̧RX�g*8,7���Ƅus��C�S��f���Q����G@pW��������_Y>g�-�\S$�zZ��M>V�6 *��t�:-RgV�������Z�߿�#w�a�z1��<��Wd:�Ԏ�R�'��Ǐ/`��A>cb�Z����&��t���u�*��*\����A�Enf�Y~��m�K��ʜ��儘R��ڢ�T�7�,�k�w
����Q�ďe�I������hr��7���
P����C�ٿ_#���8��b؟Gw�d�T��hI.�f��82hD����
�,�=�>߯q��
+H�u�$K-{�Q�ǻ�s�m�E,�5!E��&��T��L��{馆m(��x��h���;YEfX�q���� i�v)�tt��*��![^a�^$�d����� :'���V�xrʛ�HfC��r��8�tr�ՙg�8�d���i�� '<`��I�۸�>+����m��I?l\�#ȣ���+������J��ԨΫۊ Ϋ9͕T\�ʳ��H�C+��э�G���cU���)O�UB��ot��Y7"HL`n�5vz�s)h;��>'`���������|K�`���$n���;Ҁ��x:b����䘡������M����/|��W��&�_nWY���3�	J��~aF����$p++'�7�_.���+�ٯo��־B� &z9쵪�!B!����_RZ8�����tC����#�(�_�,ֿ�̚_Q'	��zͺZ݋���2*)��k!d�4fX�@����� �uDA˂I3��]�r�K	���q��!C�oYK�La<�v���� |-��Z$�L�xƳt��� 
�c�էEV�*�^�z�d�q��ڌ8���]�J��er̓?&�B}J�ņ_�4�0;q�Na�O�Ţ8qt�T�}A��o�~�7�q#6��"�x����&K�%X���~Qx�^��L��*P���q
���D�s'��"p��e�l1�¸`�-�o����Ӡ������"u��ED��(D����\�����o���s�;1�LZȃ���W(��.?��_b�������լ�IW�Nu�[`]�"=��z�S�)��~�YtA8z�6�F��=M�<�`�CY���.���-0r֪���Ė�߿wԡX*�N�?�΢�ּ�����d��r*
jf��|��d������j���ܫН7����o��S�t=��l�@`�b����_�:0��e�#%H�쐭-/U^԰����5S}�
�hL)%5	�j����m
���ά��2�&�m/���0}#���xM��Ȍ@�S��� � �g��+̤���A��QD�~�t��e���Py�KcӨ�d+���
Ɓ=��GP���"�	]�
�V�~�#����_�os@��pq��z�u���	kл%U�!��n���������Pr.3
;�nG��}.	��F�4�(�����s
��(P��c�3h������p���?$��x6�(t?�c"�6/i�!P^	�e۪|���1��jK>������xW�X_�b����B�X�d5s��N�A�(%@�V�f�c�<������Nӿ"�~�^��XP�����'�V��p!7�)����x����^~@g�~��1lr2������rWc'S��4��M��� œ��X?q���)��⁨�4�� �c���$��yŨ�^{����8� �bT�h�[�c;�.|�L�/��3�a}\�����lȄ�����Yl-�}~7��\s�=G�w0�}�� 6"�-�P�`L��
��r?�!��^��̬�/�YW4q3�Ys�| *g�O�.Qz�T=`�]K㼸3X�;nhC:�|���A�\(�w��s3�g|��t�2ŗ�|v�o��|�@J
őPMp��ݏH���s���<��
z+*W��	�l ��*��UắN��nG�����U󟽜���_�^���Ƌ~�瀼��^5�=���z���>��؛]�^>�Y�V2�G��h)"�ޛЯ|��Z�������r};����U&� �魂y�x�H+�D������E�����!��4Aj��~!�_�1.������:������hH�\���jd���P�ɨ�R��n"���7
�n.ʦ���Y�)��9`T`�����糟,I����!��\�  X5E�*Zbsi,$�H"{���z�/øaH2���a��k��h?�ܯ�]�� P�e�oYw	t�Z�_mV�	3��R�S�N�7�Hs��p�3<�w=��ޏ��^�G]~��[���%���=|���@E�1��R�6�)��oW6�pTܽ�U��tP��寂��JU?����,0��!C"����<
�QTR�]�,��H+�j>��g�1M��'L�M��Q�2����%I�{�} z��A��d���W"�����;+�~��M�|�s���W��Ov5l���*x]a'�:+P;�s��d0FZ���)#aA�?���uc�;l�Xf���M:"���^��@����b?�����+G1����TkF(��e]B�-	D��}ޥ�i�����s�93�݊�;(bfw�2��Z��`Q�K����tw?�8h����0�5�D�!���-�lV���oʅo��*&��E*�~����k�b5�X�M{�ȭ��C�2w��/��Vc��v�/F# �W���
��ϭ�>�KKy��l�O=_3���g~��y��zoΧ8O������K�vn#K�Q�G������PY��6y�Y�4-�Qb�\��VFcU�'Ge0������fQ�k��,�2 ��D�`��� Ll�N��N�s#��X���r,fqC߱�;G>�g��f��Ό}KR�`Ť�;E��o�	�{��{�6��������8��z���ɉ�.�I]7���%��S��2T�2�'� ��)$���2�(�>�|[�|���AӐNE������a6�}_J�}�iR
�W���,�l���︖���g�x���FU\_���K%��`Ԙ������_�>h川�+Ц2�;��/xH��2x<%_��9H!^;&�X�m�݋�y�*��v)VAı��h��!��PT��fHY��4���(��;�~�2ȖL�hK�T�*r����&*`��C E>��!��L 0���w.�7�^��8n0�/��h��?D+�%��VH���;�|��uҳ�ui#��Oڼ�w!���A'�����g+"�O4Ȩ}z�����n���`��_��^���$9qWQ���I��1X�[jt��LEy^R� 1��u����:s�E�8i:�X�>鿫x��{ҝ_$>��%�oxCFtŰb��xy��L>���1��(��N0�L�Y�[�N��uH�k*`-F�L�"�A�!BT�� 5�1G�ȍ[B"�B'�)��׌,(����O������J�թA�ܣE�?`���jhDN�5�T`�H�� �g˝��:�2�s��YW��ӰJ}�&R7Q����5^!�c�u�"�3wkm.F��'��VR?�R~�� nzXgo�7[r���)��",?��YL�Ьt9�x�Fz��ؤ�_i:UM�����F@W����k��X]npZ��N��EP�q�Y��p�{�}�e�qgt���Gr.r�7ջZ�%6���'����p�ŗ1뷕�Y�S\�?���Afj$(҃���q4�*��ɢ�Y�~�c�U���Ǖ��?gq�3�MN�h�ߨNk������Y��(��������D�����.�� vG�9O���� ʗJYXk	��3�4��cĚ2�
h.>��^Ǳ�+�֯P������c�fN����}��l*<��o����_��!�~�#��<հx�����h65����`N�r�uwp}�g��S(�=��I�Z���_Ч�q�����<�cz��*��3����:���<dCn�_�=��r�w7в�}�C�r��ʞ��i\8w��=򺻎B�s��������S`���Ts2JHm|��	�� ��;��ɯ��|��������M�&�N��G�$������VM�(�p���s���}�+,Hr���o
�:0��"���� ~�$��0����
FH@�H�Ն���VK�Usք��ȼ"�������5�˂�A�,ݷ���;Fi@L�g܄����ɮ7�Θ����lY_Ë�g�IA�J�2m#>ϑ�F=)��ъ���O�~ztc&��òg�3xJ�Se�6*ҧ��4�u�b��7�8�+����C  v�n��g�C��ASZ|���e�����i�cP�,�`��PHx��H�?^>�C5ba�]��D����H�N,9=|����fG.�G`/��%�W1���g�2s�)�M�ǫx��gTr�[~|���!�SL�
!�f�4f�4������ys�`�J������l�j�|���+��c����B�I�-�Gx�ɼܤz!;��co��^N���$՟�n��t݈@ʎv%��F�4�n�,�a��ͬ?���9e2����<2��b{��S�C6���h7��Z*�mV��jl�A1��率7���
4u�۰��*,���� ����o���g���쾕���!�y:�C��ök���@��Z�}�ǀ� �vu@B��,lC�Ⱥ=��f36��B_G��4"��]�]�tH������HRd2kT�d}�>I���ږ`Hߑy�C��o��+,â��.P��g�ޗ%�<ZyiŷoLXpmj>#>~�h'NX�k����FU�Q~!dأ&����0%�T[��Yl2�xe�3ڶ����ҕ�L��a)$�Rl�ɊgZj
0@�l
�N@e�S�>w?I�m8�(��8sL����@�:��A�>"����j��0��/�=QL���.�W";��8J����li��[s��=��q���IV��G<|�.e����/�L!��aި������k�G�u�ۅ���ET�hPw�.�5��rc�K��ߙAF������λ=;���I��Sq�/V���ee��uuu"Y��jj��+i�eLF@/�\��˱ {r�� ͌���Hd���`���5����hSq�"� ��mh�e2��4`]A� ]�1��bT�c��g��?�+b�-�D���]V�e�:2B�@JBp _^���tP;�}K_�ja��'�Նr��x�o�K��R�z8�.��y�����v��~��@�p7�t釴NAZ�4��7p�����Y\!.���xƆ��'r:�K	��D,/��n��X��%�/[�t�9����ݖ>�i������Q���8�9�l�5]��s+��+�0o�F^�W�ztO��7�~Vgx��wۉu�k�\���	�X��.G����&��e�Z�$��Ӌǯ�O]��ؒ	�>4�&#C�1��"n�pIȖЯx=�6J���ci�((�V�)�H���E�ʌ���@��M��75�V��"/��7�9�1�OU�����NW4��|���zP&��[�����3-���r�����t���%@Ϡƣ�r���f��߱�B��[�d,}�����%8V_��p?���>�W�xE	�r78�%�?���A��{h�OJ��e_�CZ����D������kC2mH�]��涿V���\La?{S�u)�ǳ�C�ީ�=�)Ј?��+ӽT�"W�HKY�0��܆���� ���ޚ�SA���o��l\��f�ǌ5��ڭ�Qv������,R�?�8{��B§��&{-��=��=Y꽈��*ƒ)c�"5����ϻ�p3/�_�vE���{SŊG�����F�ß�0�:�;n��$U�H��E|x�c��/��eF��zj�W�2פ+v���k����d�����)<���ҙ=��������}e���4lD��⧤�s������TJ�����I
�"5�������Li@����{a#  ��4"Q)��Z��ei�?����\�C��Z,u��b�=�<98Hd���M�����i�^�:��%�Y��C�s9<�*C#��v��0�wĩ���1�4n:ʚ�<T��o*\�֏�U�zx-zf�}�TA�7Uہ�`�\3����D=^���,Ջ�E�l<���{h$bG�.�����7\�Ӥ*���(O�T�;�M�o����
Iì��~��s�*�_�Q���&|'�\`����+%��~�W�	�����$�eZ�:��jR�QxU7lp����]�j�k�1�V������?�w=��X�l��[�4 �)D�'c��ڏC�����8>����1�x�Y ��&�ad;���`|��x�%�<���aI ���a��Ĥ#q��� �e��ai?���#��
�|�*�K]}��O�(I�����^��Κ���I�S,y?�F���B:7�fBQ��(���H�G�#U�C�0S����:��n�y7��[ӑm���A�=��V	�ؚ�@�is0�mWM�{6�!; ���JK�M���y_��Nf�}Sq��O4�2x�����6� i
H�I�����)hIG�	����)ڼS�Ց��U�=��P�
�T�jq3�e�&�L�g�3U�/�A]x��%l%?u��{י&�(D��P���f=��ϋ��2�ۓ"�˿&X&0bb���g����'K�����?���+'@TTT�AJla�4���������ױ#�Ξ����=�][�H��g��sn�yY�&��ұ�B����`me6�\ͥWPBqR(�4"�~x��hT;k�YP�4B{����?�����O�E-r珛�T���3��Bڒ�=�u5���ڦ�HJ,c�M ���^��8�J��`�PY%ƀ���K�.Σ�D�4YL������t�Ye-3��"<�dY��G�Y�E�=\��.DXivI�iX�;�Ni�Vz�ZXZ��a�e�.��x����s�g��y���9�Μ�����}���r��da�f-����,ʠ�5�$jH��O,L/�(%��&�G%���DZ0����������p�4����.v��t���p����L�Rx˨�לbyNə�v�/�ږzؓ(fb2�LF��F}\l.�Y��q1��uR��a��b�u7-�G��t�Q��0���T\Wf����� r="|��ÀYɘ'\#�֢y(�(R���C`��rG?���*g����M�՜�<͸���r�A ^HE2~Q�{�Y�O{���`�Ŗ;Sn��� � 逃�s��wRG�����s�����9c��:|��*k&A���x�&�����󈉖b_&�J%�*��iIxG�~�Jlw
V�VO��Ȁ�[G_��9W�O�ŭ�݊Bι�NC�gW۟?)(�ޥ�N��X��D����O�ނmc���!jzހ�zv�~G�,���}�w9�۝����4Zg"�A�A`��*���~�m&��3����� ���D&b�>�H
v_�/4�BM1���fPR�4b��9t��%-��P5EK����٭
�Ζg7�f5��PI�j.Zb-��F8ܛ����	����.�/�k6�4.�¼)�-�Y�c��a�1&�:�8��W}�f�m5.&)B��|�X5���~+|��ؿ�ۉ��I� ��կ	�Bo�i1^�dd;�{��m�"�����T�\���O�^d�p��Pv_FO�h�x�M�.A2CמY���!��촔%�-t��z�%�Y�����E%���M+	��#�S��M���D�b�Vd��;(�����H�6e�U+ۦ�j�V�Ǻ��ė��RN9�UB2��H���:y���I�v�-��h���*����dZ�~=���8芈�?9��KH�o�}F�_s>c�@]��6�fx%4[z�����؛[��W;��|�Dy �T�Q+J1cb�5�8��F=u�1��%�{3GV5jk�0��@�R[)Y��x'��W��Ȣ��a����7�$�<���I�K@F�����o#���_J�lA�1�#�y���#fܒ����v����,;���Ɲw����W�g�7&����E�������t�e�8�\e��CMt��.8?}uWX��E��A�����F|+�� ͊�z|mbBB�d���������/v$�*����H ��ש���6��OX#xyC0�3����2�~qN�[?.�x9�@�_|�ݠ=�تM��kh��AL���+�<��� �)R�jh���L'Q�Wm��@���;M4*�`2<�@݁�=��T �����9����M�EC��C�7���مd����t�;���|�=O���l�${q��ڹl�sy��,'�-��:W]zK�HD��/��������h��*�Jq�Al�K{Y�#|��W�Uz��&3�=o����H�W��p��[I�<{��W��F���٢JP�֥�egɖ׷R#��*(o�I�m����Ar�Mxe����l�m�:C-�6n�a[!���dm����ɔ�߬����9H��]4��줅\�ux��ja�'��������t~XL��J���l��%��W%���eѸ�%�6z2�$�؆��Mf�S��%qX0I�)e���YQl�zr]���`��=;}��*ԧR��xJ�y�~-}d@J�`�5�(I�Њ��9@�����u�]�%j���g ^���Q���\���-�4�����ɹ�ݧ2����f��H����&����ɾ揘/��
uI����g|����,�����`(��fο��"�T�����F� �
9ɼ.�8�a'b�#���ڽ���4P4:dl��̇	c��}�<�x�m���7,�ֻ#�tgn�X%���s�7��¥��?��ET�%�; �z���ո.y�'��<Q9��D	q�6d����O�~�����"�,�D��צna�S�_8��mY�A��J�en9ޥY5QP� jݽw�0K���ǖ W�%;�����@5�W��`���;�� 	��M�B��ZUa7d�gP��04 �n�\�]9sH�kg"e� `? ���[�18&9�����(�I���s�(���1�c�o^a� �5S��wG�W�}/J��IT�\����@%
B�e%8�a�K�kW/�g$������~8��?������\�w�;lsp�c꠭� ��<�3�>��jOT�LL�P��l_�ǜ��?5;ˏ��@�*Le�s>N%,n�� W���I�K�D�Nh�y=ګ��[�	j�Ў��x?�{���#J�ݹP%�%#~أ�x>����)}����x���C*V�I�GO�,�f� �Ы�l~���[^� ?$�0�J�BTkK�.�+���t�����0�����G�1~p�{��@���i6�K�=4w�nhiy��y�[ϭ�U�ȗw�]��M3�.�=�azlt'���)j6���x�4|	S��3�C�LHS��	��E{0!���2`��oC�4L�vft0��_i㍫����f�)!�	 Fw�ž9��f2�@>"�ݢg��@Ͽ�c/'�V>�Q�����`'�G��&��升]��V��~V�%�h�&�s?2~}�:�'��\^\�
�U%N���b)��!uj��/Bk��^C+�{{��yF���O~��M-�A�������e�;�SvJɗ����L��6�4���E�H�a����d��'���r���)`$a��W�%�t'��P�˞l���OlI� x`<,�!�����ʹat:�9��?Z�IՄ}᜸[�_3;?�/�Ƈ��M���.빐w��>���]�ws7&�����/�l����(P�L�A�^Э��mp��Mߑ*��0*"�mE���¾	���D���H�D'�w��4�|w;��v��@5� �K,�ci* o���ş�?s��*��rJ���i�O*���kd��&M3��%�eXH}]o=(
\�"P�D�ah�6̉�Y+S�-�
H�Af�`��b�����q�J��� 2�`���n������5�b�����(���C��!.�N�����ՙ����P���@�_?4�	�2yf|B��W:dIL~��~�Sۭ֧�>�3���LA�0JƇo�� ���9�t��W�"g+��6$Z���im�g������?����%�벳�w�� � ��N�IQ �[#!�	tzrm"��j��W.���C��S|�d���FF�1��s�L����j�GO^T�K�?������-��V�k�i���tl���/O�;2��&�L�g����|1�S�dc{7d���ט*�dL̜���vH��D�S����]�$qr�ه�H`�L�Ɯ=�R��2O�
�yn�f`ϭ#�O"��S�����9��=�5;GA�X����y4���O2��U:��1mV�<?/���,�[,�/��W/Z�l��K��GB7)$�S�ͬ����=Yy;�z��7V����}�Tg�Ol���y?�U�S�X+�%_vihM����X	�P�ʅK�g���7�a��^���Z�4ZTͷ6z�ZV.�@�c.�̾�Y�y+�ax��/�X�}����,Ќ��(�3���x�%�8
�U��x3~#TܬjM ��\�_�[z(,��;��@��Q�%�Wy(S{�ߝ�R����g���5ƀOa� `2^?�Y��2m���!�RGm��F%og�������;��\C�<Օ�q�J]S[���5P1��"�������z��&�x��J�n�����y%���Wre����8#��۴����4S��kZDa����;M|��Z���B���6D��#��U8�#�Uу�b��]�m>��CΖ&��"��U�ӚU��D稾5�����4�f-�/~CkɎ0���[JrJ���ہ���=IV�{����b�U܉�Џ�qt��f��:��]	�^��R}W�M@�1B�
�����{�p^kh ��r������O��(�i�A��cv�A��a��j��$}z^ЗII���V��"b�ȯ����c��S�93���F֗�,Y���
����1��>�u2'��]�}A`�Rv8t�%��Ĩ��V<�z�Y��#��B�:�_�c�<h���#�2T�3�
�������[8�t���y��w�����A��R+9`���V+��4�f�˺�V+�2=J�N���=�T�����Z-��é4ߟ9)l��X�F��+';F�M��a��gU�c�����,��~`�"[xBU-����ٍ�U�]o����Z5�+�&�a�A�����N������@S}G��W��+��x��>O�a���5E�st���6��B����E^�v����z#J��u�����9U���p^�D���ۛn~�}כ��>|t��������0n�͠�'����cһ������HQ|]o�+6���/�`�����ϳB3&
���@�C��`&��,�����x�;�~	hGBF#!%L�PlW���@N����&�r'�b@b�Oc�
���ڷF�7����aY�Đ�@���n��7���n��{S�D�$�9�u�?[�Q��_�;�:��,~�����|[�vu<�-N���v.�G|3���s��L��(3��*"bM��#�0����A��z��P2e"���w!L&�X3�v��
/�M^�R�/b%MI�n
@N��8�LdS�ʽB�km�G�L�&��e�����z낏C<�$���/�?��צ���{�#4hMߘ��f݈�E2?b���J<��KN,t�=��:ܠT)�\4�G1�P�R|���brl�6��!��+yI���C=���P��w��ѐ�c��C�]��$\㷭/��t�������w��)O�kAF���(E�D]y�\[��D:�=�H2(TÒ�$G)Z�mZ^Fsאؠ�vS �Ii����V/�U��� �e�)j�������[����G|,��Q�<E�_S��G�h@I�(�I��v������K����<O��X��d�7Ƕ�!<�F��t�P�l���j�Il��Ѳ�^sF�Y‘���-y��T^V����v�M��Q|U��DQ_/��vs�z��"��eo��߅��ƌI����D��3����D=q��������������ˤ�mg� �qx8z����n~��:H�?-x�[��s�5r�,��D�����DAX�Z���Q��Dx�_��xA�����6���:R�𩏷�Å"�9��	һL�(g4NTG_��� !w�G�1F>s �V�t��ե��˭�h����Ђ�[-8$=6	�\�D�#F�JV���|�:��~H���f�L�tRĔE�>(�����rݝR�3R� ��?ͱ���r5�Z
D��Բ۪nN���BZ���Kw�9�?s���>�ud�V�V�t�V�8�}~Q��A�׬7^�PeͬV��e_i���o�E�oh�R���`΁���}�O^� 7�����#aFp��wB1��;��z�5mv)mϒ15y*�*hfz);;��L��$�l#e;�D�W���.�ʗy�㋛��?�?sF����6!8��$:��=�n�������+E'�L���?tP_���(=y��Гq˻KM1e�c'(j\��bI�r3*D�>U0��nR��̏�π�#h��-v/L�ELѲ]����V
�.��#K<���]r��9t�t�"��&=�����x��u���z�?{��V��ၼ5	_����"Z���+Ј�L��5��(`��u���)~O#sY��r ����I\=�x�R�h�{�&�A_0����i�8���V��=��ʘϕݙ���Ƙޞ}bu���~������#�(n�5)�Y���S\h͵~	.Kcc%��O��~�a�m���4;�u9c�����'o]����p#n[����ԧ�&5�Z�{�"A��ji9":&��[QO�T�]��]L5Dz?QHZ��}�������$%������!�7�f�]��ͼ����y���.jʠ��.���J|�P.���,�Xހ���쾷�ĥC���h�5�v7	7�>VSU���w����I�P�V��3�����_�o��J�
x���RE6�F�3Ww�߶o/crN�"c����ǥ�����%�����R+}�*��HU��ƺ'�M FV�]���T�|�E�?|$���ehZ�|G���E�*�.�������
�X��ƟK��9�?W�.�[s���9[�|�����TA�>�Z,�9x'��|�H�Ũ5��:��7vM��'����W|��wf�x���Q��
�Ȣ���>���[���Lg~4θ�P��ƹ̯��d���R{��9�#1e>�]�Un�P��ڢ�g��O����d/�
~�(-���]���Mz�,�h~f)��0��7˄,�䥉�/C]�i.�]����("��>!�)-߳������^MC^�aҸf������}T�jn�Inɗ!p���9Ņm� ��D���F	A����޷�2�ud�y9_+v1.[
��}v�S�&�9�} ������Emp�-=�H�1�*LJ�c���PS-ߖ�\���Ѩ���~+D�0���|�ɭ|.u�u�җ�y`�[�x>��*`�O��jx��T6�e]9�q�_:�8;=�tj��w��M�l;`�㣽��~����'�~-���;ݙ�x����yqG�v�,��M��i��F�vڈ��=�CpUo�� ��"�y���3z:$�^0^H*\�$��B�]�1�Ո���U���Y��hN�y>gŧΆ7���s�X0�K�"�ax���� ��Yn�Կ�%R��'��̞z�Y�{Ž���Q��z�H����!f�	�I�:���#�q�Bc�YnbE6w�~�������S��ˍ�������G���?/uy�r٬5�mgj-=��M�ʎ�:i�ͨi*2Y�a|5��k�a@���V�=D��8ܛ��PS�C")�T�Zjͳ�?�X\��\�٩�ާii�V�)L�eM�o�ȥ����1���X�ZTH���5���}]9W��V�/�g�8y�Ls1���w��ݜH'7*f�aQ�{�_$T���jF��B�W�rڶ]i�~\n���w��l]�>d�'�F��9��5Fkȵ&���]c7v���#;m��F*���>��GD��h�4?B�Nl^�;*{y�XU�>8����H���vj�V9���1 �����L�?�xޢ�%���@�es�Z�spg��^�\�,�˼O�3% \sh+2�C� x9R�l��H�.+k� XhnXy�g�&\�����a��W\	*�ȱ�^��#;�����-��ۘ�"*4���k@Qn�B�w��l��Xxq��"��]�c��N�{�O��G�JX2>b>���_��[��_�о|�?Q���;W_��i�
H�׷w�.�=..�bcc��Mڿ��y�,me}�mn���1�vsQo��dz+�N���/��R�gCMMCS���B���κ������ᡓ��c�����MN<-Q���#��j�?x�6|j��6C%��\�)�3�_��O�5N��j����NZb:)��y�3�`X�����kC���ی��T�^я���l���%��W|�Kj���螧�M��d�]*	�~#�zq�AA�-˟�}�u5��:�����mv�����3�5�C����$^P�݊m-�+����ErF@���{�;'t�����@��K�N���{{`�\P��7���c�ն��/�����<BaO�4uǺ�2��w�������bN�͖C��H�����"��Z#T��ڇܾ��u�"�\d�bR����vso�N�ӣ~$�x#�����0�Ph�JsHk�0���!a]*���>Hj՚��%E��)�W�b'p����n��G?Y�Z�9�lGLjË��i&�U䙫+ӡC��M���*��NZQ���4sAoC�s��һ�q�"�a5��*�)b��O�_y�¦�h5���q��2������q�$��AP{��}Xp�A�S����L�q��Ɋ�-��I96W�`�o�����H؉W�w�Q�z�rK��*�^$Z���L�e��������HXxx�E�M Uخ�-�F�]>�������Tdcx�)D��p�=Q_E�����<Qj��J�2���WL��2��S�^�����Hڊ\�K�t����������)�}��;��^�24�)	�Jn&ِ=&
���'<��h՟�����6���ד��֔JP���y�RyY.��u��f34�F���'ɥO����d�ľ2s���k�+S�)wP zbl�	a�&(PT��wb§�l�\�0��<��Oz���{gΧ1'ۃO��9�{�>�~&3@5ԡZ���b�U�85e�}�'e�2-Pm�sn�15���.��u�`��vٷm	�{�|@������L����ݘ��sP��Y����f:/:����궜�8�Zb2�2�z��L%���]������}���E��m�q&�aS�رm�ՉʻS�f]^��/�K*��Q����]���j'�ϝ��T�]E\�[���2�2&-��U�Y��10�ц%��:��f�gt���{���v@Y�����5�6�t��	�ܳ��>��_��kʩ�	=kQ۸>c�`�"\�Q���B�٬!�Bx!kn�.����h���������~7�lP%G�<��n��t���{���M�(�i����gŌm-.�{[�b�/Ӫɗ3E����0����.V��qC���h�e�aF�7S$��7�|�(�Gc��YN���CV~��7Ic�r��B�7d�S�-}�-a�n_���[h
��m.%��ݺ�����y����B���`^�:�EY ��(�r�ͨ�jf�s�+�Z>Ԝ��bM�����$ŕ_y
;��
v�L�ⱉ�� |���K�s���6X��7����g[.�r.������8@ ��A0*��oS����\_�������/�
bG]�%m��g皣�-��WΛt�v�|_���|E���|���mp��[�8�=>*�A�ciW�"^��%�W���ę�(.M|�n����M_	]�&��US�ǎ�������'����gv��/�9���������2d]����sZ�5u���6g��G&����n�<����q����ƛg�J4�Ц1�9��G��s�&dj�F��P���*U����5�Fl���I����_���^�ZZy����/�o��O���MҷG�)燢ç�ﮛ�HR��@@W��w�mz[c�CLI�g����6T� �cǃ43l!�u���9ó�=3���n�%[��/5`��)6,.�UG��K���ڨ�f��vk��̙�)<ۄ�1��J�0a���|���,R��NsE$�0J�*��Ǹ����a�J��DA������80R��oa0K�"���M�j=�;�-7�M�?Wa�u�K��yP��l3�Ip���>^j.0�xɑ�旟�n�˞L��+���Mq��_t��w��I�C��#�Oܨ��o��������c���j,�ϛ�ĒEW\��bPϸ�B�%$A�x>F\i�	�ry3v�����3�Z��!9�D#�T�~�<��{#���As�u�G�a_H���km�CK����Ls�'�*Vű_<�࿔]<�Th}:Ǔæ�a[)Bd����76�~8,,p�T̳o��{�'��~����N�����K#6������Fk�vS^3LH|��¸���zUձ���������2�������wY~����m|^�z5��p~6&�5��m6���t{{����Nr������Q�Y񸠈���`��F�g������׀e"�;��E�䙝�fQ��y�ߩ	�Zy�-��������_>YU<9������uۮAC�oc4��aRh�z�~�_���Dw`6�Dö-��2������鉎��y��;eGd��S���w�%���.D������+�M<�:$�����Ʀ8e��ъ�I�����y��b]���'���`&���6)��(���3z��uEy?*��K��n�1 ��PM�RN�ﻋ�j.�m/��Щe��W0����U�pPd�o�	��E�Y�z��P5iz��&���ͤ_�9@�Q��2�=�|�5��V�蝕�����n��N�S�5�����E1jUs���l��ҏI?����9U�}��[�>�jO�Nޑx)��O��r���]հ��O�9�(���T+ϕGP��[Ŝ���EVw��p�d�۵�_�2ЭbM&�)Hd��:+��n� K�n�bcYЯz��^�����`Xq��cbjė>�|��������ɮ�0S�/��M���_�=g�12q����z���Z�<���T��F�8�A�/Jw�hY+��h%��#V�1g)А�ȟ�.�#oT�E*�X�,�4ҩf[@�S�%7���P@p:����֟�)����ag(������6���{�$j���uBA��c���Hֈ�/�Xy�l�4���p���A��=R�~����3h���&���Q�	�Tq��.��p���0��d%pְmX�(��&�,s��H�}-��Վ��õ1�z���:�F�kRx(S��ɛ_�n�%�6Zg�&ɭI�+��jSO�۫[���do���ɜ�[H�c�7$�23�	���vS��e8SmO��i�6���������gW�T�JpN��~��q���=��<�=�^=�Ɗ=lN_������5�9����?�`�2�sH[���96/��9�0�d�i�>�v��.3�o{���	�B>0��Ȣ��1%V9a�.s��nP���*՞H���!"]�4�����|���RJ���VY7�?�o�g��hl?|�b�TA�J�
EFv�7X��,���ۇ5��5Ňoɯ��p$w���U/'Y��Vŵ�h���.;<�x-}(��:���j��X+�as��%^Ѫ�k�v9�n���lU����"�M��¿�x�pz�� �H�?[��?�Ϻ����i��o�r.�aM���6����G��w�{��[�?����.Ƅ<cS��R_9��U���9��Vp�Fp&����5�ő=��FR"�N(9�׷K厨)��W4�����N����c�H���ڲ{����%��HY�$���q$R�	�R
�A}���z��<Q	�~;���!'|dFzRI+6�Ͻ�I�`����gy����M�N�$��W>Yt���ƚM�&|�X�(;�F���p,Ś�$��TV���:q�&m-*���8^-fk�s��ҸҜ����9H�8&.���)��Z ���%����#5W#�6������x�?���2�����.u��*�K�U<����Vfp^�$'�t~Ѫ������������,�p[�h�2�;��M2̞��&��?�=�S,A4a����<U|VK��Q���65�,ip:�;=d��|�Vn��vR?���L��Fw��P��q;+�%�6�u����ߜ��SY}�k�gLko��������[M����?!�ك����I`a* �#� �2���"�R�K'x��L��!���x8c�T�TY��]%.���T�:A���4�D����%�VĽA%��;�|��t��6�j~M�I�B�3卢��#I���K�T��qJ 2w�9o�!��g1P�5��@2�ȷ�KK�׶@ ���
e��c��j&W.�Hr�%E�����y�Sl�
�R�pM��Bɀl��A��c�f��ДZ"�i�";Ș߸�g&X'��l��cϰ�v�w_�48߂^�=Ѿb���W������R����M�T����
�1���z�^��������hݜĒh��^��):�~��;���9�ggg/..b�n�oζL��_�%�廻-��u����}�
�V���'�����0io������u�/�@tww��;w�����BO4�F���@�6��r*Y��}����@������H�\W���="W?6�W��k2�2��~Fw�BHdSQ֡m۫�*��F[Df��1a�,}B���}��6����G[Z� ���3�òg��0���/U"�����_*m�J����&G��>x�+��޿�HT"��«Z5�w����5���/�X��������t���k�Y*��l��.K�bd��j.�@vEß��ڜB��-���l�}��P������O	���]J�J?k�6���i��=��x���r��
�Y����O�"ilԳٛ����d�C�j6�<���n����W�o>sZP�����ݟ->�`��<�^"�� �/�tk�O���q^n|$��F�?s]Ylh�tq�1�n�:�?�պ_j�!Cԥ0E�Rq�q�<�v�*"SvJҼgB[]��ZF� بպ���ސX���i����n�Z� �(��Z���8��������A�0�X�~�X-,�i��~�ީd�QF����!B�������mo�u}Cot�t�ύ��ds�2�J=v��]a3�6���/4l�z���� f����n+�f*?�-�˒h���8�=�1�{���=��+ � 5�*Ժuͤ-�s����Y�p	%��Lp5�y�Ȅax�*�q����S̾Q@?ľ}�K8�l���Cs���"z�Pϕ���l��E8^��iO���S�->����O�ō[J�!�rK�����/L�~.<f�Hy�fE֩��,,���`��w��4=��4֑�$��F���}
����ʶ�ـ1�-���BT������ꀼqd��B��
=P ��!x���x�Z&��&5P��L<~��F˵�4x]���nD�b����	��4/P��"tw������Q+�}������q~�9X~t��k��r���0B��U �8:�<���ls�w;�����rp5�o���Q�9pOԫq�D8�����` �}/#��~�6��б兽�R�	�����Q���)`@�۽T�Yc�G��[�d���"W�a�ޕ"·�/�Á�Zc"����Wz.f8.�s��{�8�s�YQ���yL���Gkk$'x��2_�&116�у���g���xĘ��>)yC�9x^�Q��<e��Fb�u����Į�=o�o}Kf��i�H��]��5�.A��)������w�oK[��]��G�9q]��	�uǛ}��CO��b��f8�B�P��� 0�V�ǘ�w��~�/����Q*T5d;)�5��~��i>�v��Am�^%�m-��2f@vPq*�.Q>6#�k0 ���_ER� �����<R��_�bA��&���o��<��*mJ=M7��Nk�.����Iv+j�G_e���e�b�6�/�u��ףe�e��;������ �u	�9`�J[K���i��3[S:�wg��'�Ӭc�Y�-�_k�#W!% r�)�t��tX��ͪ�����q�2�u�ԏ2H�4���m�P�V��K�6��͡P��=�e�v�E�Rѱ*|7�V��^e�h����^i8u��:l��d�9��	D�`�Cw4z�vC������I�'��O�V���*���(uY�h�ټ��R�
�����?;��h"˭��� ����x�5�ܖA�dc�J"�cz�� ��0��Lro�9D&@q���z`kƼ*���:�Dbee_��Dƽ��o�ȐP���2�i�@�^}��K��Ŧx3��7��Y&�_q�ZR�<�����䂤0��S�
1��`@@PF�5M��-7���U��2i��ϰ`�ق
��l3��P��ʅ��P�i��NĊ[,���෍�~٘�V�DEj6�����������Ӵ�w�ldg��������Ԓ����7���?�<s罣��� �j�Z�s�Y-M�Zl�*�|�h�`���[�<��I#�6��	 Ch����Y�����d?�4x����Ȇ��e=�X�l8r�Xzc	�Z�G@���󀘼��{�l�)𤻙����Y#K��<4��Q�re��H�R�4�Vp�Wa���
� ��������`�߿cY���6�lMZ}.���f998889.5y���ڿ~����s%abbbpppuu���omm�������b��i|S$�>���R-��X�L{�ڌI�_���M�e8r�'���f��k�~�T ���M$2��9�nR��4�]�DkC6���o�n.������ ݴ	0y{�,���ȎZ�e�_C��B&�)��1HxK(��<'*�"ͅ�8�Ѥ�vE�d�T�%�Y��ǳ@��ޤ]�>�Fc��~�?��@-9R�x�l������jlK���(��
l�e����/�u��_N�V���%������s>�Y����L�����R�n��H��W(f�`�Ą�[�b�(�](d�7��+���f��ۦ�RYH�؂Xko�/O;$�}����XU��M�t+�Я�,������g��V��g�Al�a�rǋ� �A�="�m��3�t��	��	��QOܱ����t�Χ��P�������%A�I6�#���~�C�$kf�Uv�/s����^H>�WcI+
��k��ޚ��Z)��<�ؼ}?sX�V�0s:��j4�=u�`�r�Q�|6��1	�j���1�z�x���ƥjRʘ�#���-�_ٔ�	+�rx�U�)z=Lt�� ��nB�0W�j�5�Gܔ�W'�1��i��~6���NG�� ��D���1Q�"d8F�5��������6�%{���F�V>�4�p�	��K?c���3|#��-)�Q39;�D���Z��P��z���J��i�i�JgM&М���f��D�<wV��a1��~m�f��s�:+#�h���-%��E��{���[\��8��Kc��F�%�ՍQ�������}�7�������ߵ��G1e��� �9�Q�>C@a:�9@�:�,��&Ƽ0����?��{U�����c6uR������0l�Ǫ�^ݘ`P}>����u *�5"�.�Քl��Z�iӨ�݄�?�įO��f.���n���8O;�:�v����p�����{��!��?ྑ�����}K�̎^��IM�������Q���ђ=W>�L;.�z�*u��b�	�2u!��@g\y�r�!��E��R��k|	z���&!n�q+ �����a�N�-�,�XA$��(�Wx�0��+���U�?v�ֆq�)���$�����������v?��'�2���.w~�b���@Z�3���˙������?� ��Ԥ��4/Z�"+�{��67��I�o��2�4�h��+�i�P4E�G����IZ�3&��C>�U�ݖ����z1PD+�p���\��,�I�U���ȩy�X�Ҭ�� �wSs=rژ�^l���8m=�ZA���([��wZY6�q�@Y�jOtz--Y�]^������<����A�JtÌ�aq��S��������b���F"��NG����mv��i97)wZ%x�|"��V�aU�E;f��d��u&��E%�m�ޘ�!?7lz쟽�Ԟ�����A!-h�=��l�9��Q��^���������W�����M|�n�.zb�qĕ�5x�}��㥽Hd!�Tg�J�Ҋ�O-P��s{F̬؟?���(O*�c���Y&Ҋ���}���ɲ)��q?-�SP�0Y���UZ�5w�/E����oJ%���tr7|��6���s%
'I\�+Q~D�heXUi��jf��bt��H^0w��()�d�Q�����\zi��8�'��q`�� ��stp����IK��q$J|�M��N�Nߕwm<p��^�w�X��qxR�'��	����@�T?�a�ڛ���/�CQw��)�K���eh���CH�u:lμi���PD��e�a����2���q N�3��B��#�V�	/86�l��|�dCOC������j�8>G���rC��@Q^�/�Қ�T���4�ّ��!��|���� m�H�t�,o�n��A�`"�z.��A%�x�L2')1QK__��@���������tw��f,S�ı����p��s���&("�D}vvv)&!N�������EEE��R���A['�!���j��,��I��˜���x�-��!�>�k�� ���&*+�v���'�*M�?gU��+#�-ꪁCЬ3�<}��+p���8��D�=@C�挆虿N� ���5E�%D��V�O#��51o#?�}66
&	"",
��@��x{_��c�Z�2����s}�/1Ԯ�v�����3x{�%��`�a���X8˸����3 C���3t���--9    �R"=t�!��!1����%���<o�9/�眽��]�\�h�+�;z���G4� t�z8U>/�j�+j&td�_k�	/wr�VN8B�U��qlN�ۙwl�a��\(�M?)�)��|6���]���X�2I)D���Q�����R�o=�O+��|�Tbt2�*:�����l(������.�é���D��.ۣ�l�]����QZi|���@V��H���%�V�u��Wg��C�kp�_@gWWqٗ���*��o)�MwW���nݣTÎ�f7��W�# �Yg�\����fq��"f�o���N� ���ڮ�s�C#V5"\i��{�%!Ul"�a�Nn|�k��Rӭ<��D�I0h����w��^۰�E!rk���E�x�0�hr��u�����x�ja�8�g��*�g�,NF25\��Т��Uv�,4VJ���z���4|�'R^���O�2!Q&#G���th���#��^�����M�*�Eh�O�!ڞ��x��]�H��X؈�pmI�U�R䏂���p��]qX���F$<mGb���6��U'�ę�%D�ӎ,� r�|�9,PҌx�Ԅ~��r�y�O�Y��?֌D��._�f��¤�`Fn������>�����k�	�q�����2�h�{�H��?=Ď5���rxx�u���`	`�ᄘ�7��䐢���C�>l��P+4����'�m\ �M���kffe��q�L�T83�4��YZYs��1�># 9��O��`b�����-���Kaf�WF�Q���=Kou��m�9r����l+���#*���	2��������m �b"�Ue��8���*,+�L� �}>���H,)F&5�z�$�XՁ�o�Coߢ9�&A5 9߈xv�������Xq��1
t� k�Q<K�v��E6y���c�}�yo�������+�M �Zx=WJp��9$Oh$}2�y4�H�	�>�˔��Q�}�����uk���#&��&ÌR:ѽ��Z� �k����b4S��V.��q�C ��4v�C����H �-�D|��+r.0�*�ѱ)��FM�"�6ΏX�74Mu�㾞k�h�z��N��^)o�X����MI��~�M���*[!%S%!Qz[���v�K��c@Z�/�	}��o�߮���}ֳ�C�I�3��Z��N�nL�"��*ϻV�tܢU��L�=�J��5}�^��N�ܴ��N��ي��T`��!R��}�ʨd�٧��h�z�&̈́���I�n\�W�TZ���,U�[�gWv9�������m�����U��҃���+��͗��We��չ�G���B��w�G����6��}�jS&1���,Kz�����>^+�0	Ead�EPk����w!R�uE󐠮�l��GVv.�Fa(��s䭝>�'E��R��/L��_�}*��z��C������l�Qf˦@����Ne�\�
�Á5���'1
@����⑪
FV��b?��הy�g���N��D�T����z���Ly�I80��:�[�B$5�4(���A���K'Y��X�*����9��4v��zͪ5��K�j���̄���n�Y�F�֦0�#IZ�8���^>�>�z�K�.��yd�:R�kkD)0W���N�(0����u�U�	��+}{�e�͖�T��	L���Z(˜Ϙ���-�U��9����*W��W�r*)qb�x�~�)�Xs!�',x�Ld���86��?��X����"�����f��Q^r�W����%�H5Zss!����oc 	����ݩ���lſ�a�:rˮY�J����񕕕���'���*��K��Ӯ���G�������Φ&��dGQ�7.^_��I�V���	,��Wc��X�i�kY;ʯȚ̩D�i�bs�v��ƚBr�g�v$!Y�UOO4rB�i�Z2P΍K�� �@�J�^|Q� �;�:a��9����L�0r���6�4|J�i���9U:%Z'���䙚Vr�9�F�$�;T�a-G���~��a0ޤ���SW&R��Fa��A]BWɈ����҄����u��fev�eT���-3��њ�\p�n�<�w�ǫц{VӠ�qK�V�.}��
lTeW��o�/zԫG�FR��7"�Ǖ�M���2YL�mj�^Yo�e}`:��X���r�3�I@��988�P���/,9���,K���#�,���H9n�Bi��=�^�Ók	_��:i�@�`)�w"A����&������z�����\�S>�wk�����+ߋRz�ze8�����2c^��� -�+�$�0e��R|�����Nzn����}{b�u�ʫ5=2FSf7�8��}B����9Z�,QK#懎̟��'���D��/)��+�M+�+����Ӡ�UY|r��:�����XGyc�i��ص��r3����F�� �>E�Ijz<�k�`�Ӏk��~=~�K.�>���=�9�Ƣv]����X.wh/��Z4��T<|D�sV��C
�XP��6�P�%����Wj<A8sW+�����u:�4X^>��A ��jR,�m��4�̀��v�d;f��P͠�K�IQ��L�����L8�|�g����=�#�r�K^w���F�6b�x%���z7u�;�=��g��d-CF+��s7+F��!�xFП<��#��82�&u@k!�6�� �f ��kj�����������^�ܖ�<�LٽYh1�c̞}2.����&�� �A�[Xs<�I������z�{�1��~\��{��.��p�l`�r��B�Wt�c����Y��@8���P	����j����J�(�J�gw�>�!� �8N��<dB��]{���bEñ�(c������.�	��k���a���s� ��C���$�{��\��=*��,�D�)�����
Xm���>!�+����UbqI7 I�PR7XA���ZܷB�~�gLk҂,.�%7�k��Z��63h1�w宖g�����A�f��j^#8�Umo��!�D�n���ߵ��X>
*�}��"��y�RȇO�2^��uI�Ն�S�1��G��� ?)̌9��c�*��LN^e��%�HJ�[t��ܫ#ROlM9M���Ġ��2[�]�V�-
���9g�BccA2J{Q�������AƆ�&��J�;�?�=N}�� }����gr���u�<`��F-���P���qPr��MNq}�'����y��>�tB!-3��z���k%'�{P�����FN�I6��$�/KM��/�F:�7���zq�0��e�R3���%,��t�����f�:G�#\�d�J�R�����u>���i�	��L|�����	I��(�81�%ln���>tT����H��Yz���������_��3���g.��M���[�ܡ�#����Ɏ��a�EQ��l�D'$%�Mew�Hj}D�V�^єv��E�&�.	'cC�x�)�J9�3&T-�m���	q������{�9�Z��Y#��i��
Z[0"#X�����x�aQ��U��z�L3lA/�[�$@���bm��f1�+`VLS�YV9t&�2뵋 @�֠����0N�I��g@A��(dj�	���W�)�ct�ꠧڴ��9�_�;����|굿��:�����ƈ�Ų�	�U7G�~:U"	�a�-��2g1�y���$�j'4��)el{&)[�e��odD�>c�~:e��RH���,A�v��;B�
��o�N���>��:�������4����F�[dz#����b3#�Y�7H m�~��z(r�:���j��ƩE|]K��9��3�� ��9���D `D9+���I~ ��嚛����t>{��}��� ���P���N��E���,�DJc�=�_�W�em�Y5A��}���t-M�^X�����ه�?��Ф"�Ȫ)�`�Dط��ICZM����e�ax�J
�&��,��LiY��0O�Ͽ���q��j�ԉ	��HpHٰ׌��)��GY�[�����h��c�S��Y43a�c��s�6$ >J�@A���j��e��/(�{2AIɲ#���)T���>�%�b:�C,ŀN�@���*��6�S1��SE7�<�'��,���v��p>�B��]�+�3TNw]?���N�}�"u��
A�%.[���g�x}�ե�I�~X�k�F�j/��ZlX�r4F�O����@�Ap���W^;�BMI�&o�qˮ�٨}��S�B��9R��߿�o�M�9s��|iin�Y)�p�f�G�w�S�-6&��n�x-�v�de��$�$_���=|�~��-�xx�%J�X����m�+���z�ۂw�A��(�6��.�n�W|�q���O��_+f�K�#V��&Y��y|�T߳��%�S�e>�.�O�tU���5���|�=���범�>��q��{�+z��N�8ϥ͝`f�-h=�Щ���������}:��UHqn{��K�0�	�vBDZ�����	�v�ٱn9�C@�Ff��a�/�����c��	A��{�˨Y��`��Bv�G
�����&-,�<���d	�\e�6s0&�	�n'A��Tv�qr�-�]�g�Y�2�|��h��(��썘)�����x�*���#]�.��q,r�j bĎ�����&Z�󽐟�Gd,�(�֊��)݄
P�eyU�K����;ۮ�$��R�#��H �˷�M	da�=4�;jN�[��B�L��1z�fۓOX-���8��*�22Kf͟��pP��~�+̈́�}B��rX}1jY|4��[�'��'!a>-���A��\g�:C��(�X���#R��s�`k�=m�v:.z|(�2���P����
�/�ׄ>����A��T�^�x�_;1�?�#b�*��B1Ę�^X�#�X��8�S>�ៜ�Gi������{���F�&��E��o���R��e�]��S<bF\�+�v�� T�A�E@LN�b�&?�M��RҜ���yKB�C�d���A�x3�gmiS'�+�CܽC�6L�;̥���I�9�]���!��4�$�.^1dA˞B���ȺVHJ�����&�Y��r��a�������sYUZ
6P\�5��&�ÃAo�4»����é��kc���P'[g�s�q*�.j�Q����KF���a��+H()��_���$�+����c�R�n���m�J���{o!}��u-�)���61�˴bi���U�q���L�Cb�����H�k����?��hB[����6��q8U�IW��*�W;K)�ٽ��G��t��j�'Ja.�����*,�Ө����UC߸��wnw�0�PtQ×Ȳ,�qN��i,��v�-ףi�e��5�y��J��)��R��8����2gBhs�}�z������B��!s'$p����#��w�7l`����/�l��w�BHF�Y�J��"�{C��Nug�U����\��J�U�H�u�����%���}�_��0�����d��|l����e��M�gaJ�z;h��m7T5y�4Y�S�Z�ġ#�3Sި@:�9Q�JWUMh��|d�\�M����L1t_m{h,����tĠ�qe^��o5FJRzP�I�1��׈r���i#�_�C�]p!ǆ���������W��HWL�:5�����\��n�«_$��]}�7[ܨ�L�S�&�ȓ�K�Nn���nZ�22�Q��\���qߖ��I�䣠j��V#4+5�f?�T���MR�i�!�pq����}cac{�b�(9�����~�T
�F�龥�e�lWW���䱎d���k E�����Ss�~�L�"� ��;=MP�zIx�=Z�N�+�װ���OTC�m�qqv���S�:' :A����<�j���S�wb?���n.C�45�GG�*5-���rwwи�C�f��O��� m�n�|
P��p����e7e���Yܕ/���X� #e|�Q|�>E���_&w�T(�+��jL��=�-��7�]�!6Mצ�x��4�p���翵p���3�A<\�O~{Q�kx�����AT�}-�ߟl2~
�&Ɛ�̀��aA/ǃ�V�T�N�1I
�z�@_z�P��Gj�t�rrF�"*�O
	��I@�O�)�Ͻ�:TL�
 �<�h^U�e����`�?,خ���A3�j��,?p��!tE�>���B]��F�g����*-K���Fq_��fN��L:�!���~���2�p���>#x�@=�C��ћ�R���m�?��U�M9��9��������e��3g~��]%$؍k;V��U��-d`<��nm�m�i������ L���*�7�|��a��
R*�:��8x���wûoFs}�`z%���[r9��*M��zy���5�P�Ձ����^�0Ʒ�GǍ�<y���'l CQBA�'����]�GkN������p/���;�zV�z�@/���P(M��i V�$nU�6N>J�k�x7s'�+���5�HA3�/ʷ)��b�a��`��;�$�h��D�X۳�ar2�8�hv���{�r���.�:x��Z�4�']?��mi;����ٱ�0E`QM�)�E��S�0q�8J�ـ5<y7Q=���@���0o�+���|N2�1�[9�
S9�x��AAN_� .�~(H�O�X$3�J�P��$5���ՏȣH�?-@AА�� �6��2'�D�Bu�9�]��,ީ����gjl����C�>�#tB��A`���@4�$^ݜՓ�������vg��p(���J���s�w�A��0c�
7$4�r.��^ﴭ�����4�$����6��ڵcx�ר���>9��_Wk�����|\Z-GZm��\�a�HIxn�9� ço-���3\
���^g+ti����!g��W|M M��� ��g�����v��*4U�	ִ 2Qk�&�u������
��@~�Am���U��Jlv�[�C�\V�T���[�c9P%��3��L��3xcY%HM����}T�}ۊ�l��鲢m����L����� �x@�֟�� �{iකЦx��������²&�3����G�Q��9
�:YH�I��/Ȓ����{O9��s�4ڧQՑ$�	>=t��o#���R���~�B'kJ�����V��l��8���)�!���v��+���Yjc�6Sظwp$��p<���K����o1V"��m	�駸U��_�۵0�^�|�|��{߫ݍXP:D%/5E���C�B���i�M����./ �cB���IX�}�P��6\�~��ވ�?��hVTLq�e*�����ª�Oѩ����E٦.T�c�{��_��*Ѽ�O ]�?n��~��!Ԡ�ː�{`,���\Z�~��+4º�`���#�:C~(��|����Q�����<��/�o�l���L�[x��e9q������x]~io��q��!O�@w��NpQ�p�����F�U�^:�7KPc\�(���ۛ�����]���Vj!9����Ac�0��QuՃU����ͤ�ۛ�A;��������y���3[�Vg�µoH���N�+˻�������q��o��yk��r��+s��FHon�X�m�η�9�r|ҕ2�CwԽ]�ݲsE���<�!���\��Yϸ2��� ���\{�0XK�^;��ـ�k2#'��S��@����N��|De�>~F�o:Y3���f���KZ��Tή�O[�Σ�a%.<w0�"N����uC!Y}/r<�����%<����܊�	3]����5�5sN�{�RX���Av��29Z��׼�5��:鑅�����2��S������D;�>�7����J�;�to�ǯ��Wh��*�kS���K$zN9*�D�rz˂�v<�)���Ҡ�@,>����Oh��?~����kkk��̬4��l��l���������㹾\I٣Ӯ�h}�P`Bq��D�ɱ�|S�O���(Z/h��I�o�n�����������MLI����CC�;�\�����OI9��6*
��4~1;��:�6��nKp,դ�
Ftօ���t��"H�����"sq"̬���a@���s�It(�=F�X/�̔~.�m��H��n�+�2�E%7��s����7�qÕ�J5�6��>���R�d�:�Yd���)*��ͩ�.�$��� ���Vet��������`%��D��� �gMo��!���@$�$D����)�,z�v\Y
�DH%�%��Ɇ_ʩ�ep(I��:�c���Bt55��8t����BzY��a41��Z�n��.�a.���.:<��rN���D����!=|/�L35�JcR|Ǳޛ�oM;�T��^rP���N�[��:F�����P�E"�k��ߧ�̾��&��~y�������7
u�����MZ�s�f��D'��YSi,��~���������ę����͡�*u����JT����`<�W}H(j�����(�Ȝ����i�2 �,�ǔ���3�0��Z�}NC	��D��	��/<�٬�"_��P�<2,h?���7v'�����Є��si�BQÓ+'��D�J6��b��J�)���OQ�x����ӄ�;�,�ìt������;��?�_r�sC���=����8�ū�<�/��7��n���s�s��7���ǮFn������yϑ4�yO�p8qqWM�W�Wp�(�`^�������wx.+f�E�4+��)�?v�=�SEG�Ҟ5K	~y E��F�0-*�i�u[��	W��,Qb����4�={��O�z�+Ah���ah?��hInnk��<I�����K2 .�O H)4.�<�F�F)���?/�Lk�es��}�hT:4-�f0%��5�u�BGۋP|��1A�c���>�|w.���j!�'�*��c�Zs��Þ�aŶd>����3���kSf:m�}�4w�J�R��0�v]W�#�n��Ӥq��N}S��g����N�f7�$"Ŧ���%�y�*��2��{�
���� D8K	�=����Pc��D���m/��f�Ig�wi?_w��ߠ�+X�C�޽/�P�f��4���ڟV�Y�r��Ft�ɚ
V���:uB��I �'.R48�BJi+�Z4�@��0�P�����z��#C����S=��t&ϰ���~�0F{`b�D���d������4//��D x�J�޵�Tߣ61r�ݾ+$9vS:�>��*�.���N*�,}�����r��^1��sxm����w)��e[�,�v�])����7Ń��<�i<:�qn�@�B�i�/!��0���7�^�M(�I#�_��,��_.M���zsOM��bs9�X�}�Ӝ�i	����кS�5'�uˀs`��<�hA<��9n^!�o��cG#G���N�{��!�{��?U����n����E*���Z%pPp�s��^�v:��z�u��x��w�J��ؾdZs��0q ��a�kq��K�70&;����������}���+�M���c~�,�,)�|x!�a�j&E��¤������#.3�����b�V�Ɵ�\zl����� [�>fl�E��{.$�����j��b�%��� p2 SO����I�"�4W����l�'�
�E�-�s|�<�Ebuu�Tһ����������1���bVGg'��$��$������i�d�!�%'s����Rm��������Ul�gk��y��`������;��_��貗7�]�^��[�֮��w>������0��|^O�/�% j��io8������̱�d.W�!b��
X=Y2o��3wKє�X��WCRω�g-��D�J��K��jR����NS�|�vW���)��µ������������u�����o�xv�@�tT��4aU�د[Λkm����_:m��K��ӊ�W_S]��1^�Nl�����kK ���e��
b������1�d�,_*Q(�qmJ�ɨ�� v
�g�ʈ��lû���H$�<{��#!G�L���Yy��Jofjm{�P�n����s�}�Ħ]���E������_��2� 3~���n&F��@�@j�F�5��y�K�����5�c�u9:ܿӮ[�].�۽D\�FҠ���DN�u�9�c���>���̓2�
�iX����"I�m��>PPBc�T֋H�q�sC\�D�W�"Wʙ?�0�<��HII�����@���|?�������2j,�fnΦ������)�P�8r�亱m?*3>o��-��Xv��m�rg���������#�J#&�1�#<r&<1P�����K|R��	+�3L%��Ah扐�4AzeOӧ�F�¿cN�+�vh�1��t�����s����m��S��ķx��������佮�p����C�;��k�<�|[?��L��l�,�um �7��'��B�U�%F�T��fF���a׸��P(�4bG�a&��\L���-� �����!0���1ϒ{�)�7V� J~:��mrN��ۋE�4%)_HTҝ�jlc��%9�+m~�����笭v!i�v���p���ީϱ0;��F8�%��,����/MP�!�JC��>F����]�3K9b���F���� G@^��s=V��3�VGL�'�4>J�m��	�i)ͪ����;���h��y�/E����O�����a@A&��0.d���a	E��ХH��A���1E��)� P,��)OJ��/���p�Cۓv�x��(l��m�}O_��0��e��AӤ��cucG���gA����K-�ݮã��9�����;�]O��+N�u���z�ͪ�R:4Tz���}BAB���_ә�w��z���/`M���Dk��g�W����܉��Exr��p�97�'h`�|`�}�˰Q&�wy�N5Z��s�%�	�V��M1����G,jK�۸�cC ��%�QÞ?�k:\Aif�����p(��6ɪ0_ Z�b^-��D'�]R�1Ә;���(إ���]j�Meλ����=[�N�ɨ܌W�fk4��5.�h ܧ�Ce;�ors."Eۋ�x>���%��.�I	`y�iX�?���O�*\^l�G2�/��fa�gs����Vi�S�W�����'�B�{UwWǉVƉ��b҅�z��|���.�:G^�X�C=���|(0Gy-5��|D:N%�0�`���-�/^����1 Q��
AL���gO��M=�\��F�+�����^�7�!v�c̙��*�^8&�Kh�E�Ig�g��zC��:G��n�X8���hyߐ��(�R�!��k�yn���x?����O��	&3&B�xZ$3$V��V�pD��"�!�&������W{��!`�(�Ts�H:[2��$G4'���YR���V�z^�W�z��u�.�.����o��}>]�T�쭇5ۢp2��Z��õbt�c-�|��Ņ���a��~lkt20D���x�yq'��@�K���]Ve�9?
}n�XfED|L�H�X�ʷ]��1ö�y��5���02�Ag8�����
��xN�d���s�?��a������&�Jeʒ-u��2��#���uf�l�l>�1���M�n�|*���_{�H�����&����(�=�36��͆_�)�#��Gn~l��ܹ	5�Q�:'��5�s�YfHݦ6����� �#4�l���q'��u��A�%����Cõ��o :�d�,?o���]��m4��&Uҭ��[b1U4��?[���a�`������Y��.���t�:Vt�w�B��+D\��m���l��iκ�;��7�ɗ��ɇۑj��V �ѵ���'����p%;�{�OW��߿�;���[:��<ܿ��T	��&������k�l�d篺���ޮ�j���������e:�l����_��vܾ�w�����������1]�(��[Y�ϯ��s�ɗ0Q�:� ��+�+/qۍX�b�r��A��c!;-��щ�XO�t��/}!{��o��.`ui5,�q�{��ޙ��m�ٝU���>M��g��x���[���j���wO����W�>�{]u�{���X��K���X���X�x�1ȌS-�y��"��F������T����ܘ汚/fԔ��zk�R/�A$�)�/(�N_f�d�xͣ�����pr��lu��_�7��ُB�����r(��)��{CUݪ	.�l��������S�# ���@�����`�.�<hSa�����1z�����ӣKM]�yБ� �a֨q����yl4f�m��>.]j�zp$X
��ǊkA��|�90f̟��(1cc�_�r��q��6&�g�b���-�Q�QT��i[G�"����n�Á�S����cƊ���|J*�p�ر�1��f�"]�m[@ZL\��6���Շ�����V�~w�T%)DK$��D���|Y�vHΛ_���Z��g���~�M'cGl\�TԼvƼ��F ��y��]5�0�����w�K�����8�Q~,���\���o�o��4��o�].XY=�?�|i�It����6~m[���I���9�Ǝ���8�ض���\�<b��6�����'�R DX���I�K�^_�G�!��DC���N�BH�I���0U
Xֱ��f����m�YH��.hܳC\l�/H7�.�=bG�rdﴸQ����Я�k�������*<Kĩ��(��1eO��{q���`CA(p�K)��S|�5�dϠ�������ih��l0�7��`����+uϓ��P��tɞޙA�"��	�zGa�O�c{h�wY�������G[X��0��YK�%I9�]�Rn}����Dɾk��i%d�M�c\ K�FV���F���D	���/�=��r������0�����]˝��.yHgB>�9I�nB��^�Z��Ե�Y�^�V��ue�tK>�}��%y7���@�7]Z.m=C�OY.�ű� ,�N㳵��i��̀���v�s?�F#~~|��I���ci������ע���v��c3\x���`�4m�mb�/�ub` ���f�'T�	���H��h��W���7/�H�6�O���4G�x
U� �0.w��	�D�!����{���0��JVl���+�+�B\�{�8H�zS���R���q �5+�����}[��uQD����ۺ�	HT�\�� Ԣg*y��k0Y����u�����O�h��dc�#��AI_�rE�fj2��������m��'��AP�h��߶��m�A������)Kx�G�X�}&�4Y����C��{�Z��b��;>.�[A\��V9k%�?�2�C��J�iM�1$tf���Q�K{ܯǚbSO7̤��n�Ǿ��d/\�8r��ô?l"�&F"��@��S�d�l�sLe�l�����ǈ�%�Qs��LZ�H�>|�w����"�ǐ[�Ck��_�I�6��$�^}���=9��_�`cq��@���מg�sӺ)B�%Hvܰ�N���1~��C�ߛ�'w;_i�Nc�o�	��#�����/���j�&�G{$�����_�[����Y-�z��|�4�-x�Mwh��0������%9Έ�tl(�W;���Lz�/�4���L6�a[b��F[��H�~�
�,6�j~�V1�Wz_�����ٶ��:];��x�M�!�4�&����"���B/L�C8I{�5VUj#�[��$��0���M�	x뻓s����C��mQ����	���d�,)3���x��D��	.D�S��� �a�a;*�G�,�s��kI�θs�,\��Ia��B�Gd����$�
��,*7)E�#�ҩ�f���5��6���ᯗxu]z�I�eLNá2 �1�H�-�����\��U g���5,N��hx
�*����Cqyqt���FJ%p��4#dګl��aM$���,8}����y�������>~���U�7�����=�� ��}��mEg�w���; �w�UW���C��,�Ag�����]�C�U�]tڿ������1��Q�υ]��⾻����щl�����ů�#��@a�t9�����.}�TR[X��oJ���x��E��ED�I+�F\���H_�����!}%����S�����!��R��r��7x���7]P���7'.r}���q�A)ڏ�������x�~(k�z��j�#7�t�$+�c�7�On�O����͑���������/Ά���_�9S����Z��H?^�&�s�R�	U���Y���b^���fp�.��l��B�������� �Q��_�IxѼ���_������-�l���_:t0��t|v�%η�_�ɹ�i�Z��8�	ҳ?p��Nc��t�[�l��N̚1��мk�2���T&� �̓��N}'	\tm�/�u����ʀH��6���opC~�Bm�`j��J�ߴ��\�=dqO?���y�1����<��⋵�b��5:�K���r��R���L���,.��1�dآ�r�:o�G&8P/Pa�P`�`�w���y^�mQ_Zߕb##��Z,�W�A�/$� �`��'�ƫ��Ǣ=�'��[�N N�!��जtD���1��O� ����|[�5ѥ����$zJF����ն�L��;��?�߂��V�^��w�u��x��Lqtߪ>��*�j��J#��=
0e�n���k��F�W�U���t��,H�aK���8*Js��O��}�{�b#�V����K ��c��za��M�ؼ�f��mlu0�hf�Յ� c_eQ_s����!'
n�ţ�Q�7M������/�J�� �Y�(���:3��/�l����x�W��DR��#9m8e\+{��~��>��P��Cu#8�7^C�Q���<Z��阂b��Y���N��ж~�5Nvg�Y~�p���-�dZ�j��REQ�殧ġ+Up�6A�_}�v�F�b(4 �^�*فd�XT]�JEcg�9�Qx��L�Q�ye�8�7�v	8#a�ʳ�v��2�v����ot�H|��ې-F7�Uqz?�����V��B`*��2ui1uiu��N=�Z#;k����֮����Sd����]np�8���M�N���i$�P0g�Q2SН��z�<)�o6NfS��8�U�P���x>�}��������KǠ��FΦ��eB�B�V��F����8`�Ҳ�"{���6����0�3���+��c�P��&��Ƨ�����x-�L�fFj�)e�t�?u�7�~���� ��}l6�s�;�x�R���C���!������~dмa�?�%uCQ�kň/��轊����5貃�mm�3�d}��]|;,C�7)a�1�*�檌��Z�K~��i�J�}x�D�GL��'��7ݸm���S4����Ǥ������-'������_x���?@\Q&2,��qAq,Z��#�c�쿠�	�xM.���<Z\9�FPP	V��s'XA�!Pj�B4�Ϭ@:�jnzT���+��g���م�$�!�6아O�P$ז�}2v�'�NU�}�f0߂F��<��(�޻�!y�����K ��$�!*�ui��d���1̨�0L<x#�d ��0����i�%��~w�T}{��AC��3�+L�)Y�=��+��Y�W�ԯ:ACߺ%l���U�X&?�� #�E����2�;j(�)쑧�\�C��ɃB�ޥ &^���;n�D�����^�nϥ��e��d����k����r%H�aZ.�o���~5�z?g�hVܥڣ[�cQ������.��Uv'o��X�!�A�?a�7r<~,2��+n<^�^v)]˳<꾸��%�v<[|�u�k'�x� e��3O�l�cB���p�77 =���u�ͳ�V?�5�;��� Z�Y'!�=�e0����lz���O��M���qm�fP6>����Hg���b
�t�*W5D����M� �~!�Ot;�XQm��z����CW\8A\����
`�
'����(}��2Kb֤�-Fg�@Z,����+R3������$2e
Q�H�P&��(n=R��-����d]��T����^}����(jEx~2�u���xvrQ<�ˎ�D0t�Z�t����ȫ6˩6�DZ�]L�ܖL�t����<�94��g�oZ1s�i\��kX�@^X;� =N̦7L.�&ZR�[3��|`�n��[񿆟w�J�JJ�6��,�J��N�5�41bX���H[,9�HT��&��&+�fh(�ō�I"h�[}gkd=�V����hC��o%._]>��:D�d� w'�쓱C�����j;Z�����^1<����?���2�[>X�
̆�H\		�cs9�i���)��wxe_����tVQq,��4���'�����2� 8����2�{pww��;\ο�k���]߮�U�,���K�����ˇp(Q���*����#���������5r��o�@Ir�p	�t��q��n��4X���`v�;����a}��� <�]��G�tjs�X��$��G�'Ed�ه�A�̲f*+q(6(���:#)v����R�`[��n��+�d�+ׁ�GL�ש�a��h�Q��~�2S�}4�/E3����5o'k�z�ǲ�%�Ï�`�K`׽��^�A|u;�B�)�{*l;�\RT����/,�[�����,dE������A[b�*����D�Ƙ(�N���5�Z���\���M���4�cZ�3�
���=v��BH�3�,�t+.��rC5N��}�#�W���g��/�O�F?|.�����Y�wM;�~b��J�LQ� Cԩ�d/&�������s\F~��
����9�V�N|��-I�ұ/d�������˪*}oܟ!eȩf�PY�pxe"�ϱ�4N�%ݦ5�D�_#$L9үUM�T�gH0�Fw�����9	�&>"�M�0@Ԑ�6$��I�>���~&��QD�/C%����K��xE�yA�|@b����K\� ��%�*�����_H����o��Z���`����A������62�2�l���y�fE�8d*�Q���L���=�k8�P�K������aO��)��n@��f=���m��1=aH�=O��)qM��V%�����<t?��v�Zo[5�r�Iv�-`k�M�F�!��Z�j�0��_�'q��T�����W�0���:	��ωx�����2���P�Y ��񜣫T�Pd��|孷�r�ӣ�n�z�.h�Gl�P�{���bY����a]��.��g��>��.��g�y��+,���)��:�@���[���I�� �'�\�ՆC�˻�.u+�z�e�dU$�,[|��k`<])_���8d��2��3T���^h�B4-`5��7�՛B6��K�?�6�����ȱ��,�e"F����S�?�%�4gE�+�;�s
Z?YQD��5��k��рo(o�] �`*���rD����q��FM��|�S��֨�3A`��>�!gT���V���Q�V��� 7-Y!u�_��>|H�L��.��S��X�k:�G3t�c8����K9?��$��T�)���H|d��T�sl����k,���=�YCT���7�gC����PT����m�l:�&�m���(X�;����o��Kޙ$`�yl/�Ձ��`��u^I.�	����F��"�����l���<���P`�Ò\˷��h,����.��8eXE��w�SH��ڱ�4|`ˇ�s�?�|�]}Ҋ�#��;�������wx9�ST���-��vRT��+�h�9BL(��~*�s]�ŭ� ���Ң���+� ����xFQ��2���6���gŁuũS=~<�J���7b���j�$c��G���=\N�w1 :���������V.�:�`�����p"�.)��V����6��O�+���)XM� ������s��� ���j��&ڝ��z��6��A`~å��f�:���3��h��������V��Fݛ��r7J��t��8��}g�=��mh���ȁ�i?B>}폑�MK:g�M|�؇�U��F��PK̆(��𡧔~4��a3�=`m�&�u�bȹ��n��#q)� AIm飝�DNL*<
Y�=�7ۡ0�a����Q&4�E���"Y������-���p��WfL���q�N�EN��"��L�3[���B�����p��3]h�UJ{�#��E�"U
i�m�htQ�T�F�.��/�k9��O����r)9��kK�M��m.�>��dD-|K�Z]��3 ed�;U}�
}�Y�
 u%dn�U� ��I�;fV4��;E�S����u={��,b���,#�I��I2R�t��w�2[�:o_Ɗ�q}��ե��?�e�������� $�&��R "�b,$��{�a������O���[W���lH�yJ�����)z'g��c�L۸�/^ڏ��\����na��3�7��sCߗN��gVx�����3�uK�v����׭�7�HZ�i��(lO����������m��ӻ�O���8ȟ�+ۀ��ܜ}pZ��q,*��]����E�a׈}M&����	�-/�_Rބ"�
o-]3�����5��>W$o�E�Y����E�	���9
��ܧοt���j���d��Zp������s�S"���U�B֭Q�? )�G"���I��A��+��.!����>r��rdt1i�`�Ч(���������i/֟��{�9'Y��l����ƴ�^N�	
p��h��7p���r�JS��R���Pc~�x�n ���ꄹR)�ݷM� �eV��`�e�p�[����|:�U�4o٠�]�[�������ӄ@F҇��Ҵ�H�A�,�-��6"���?6;__�fT�O�6�{��8�$fa�*�=�E�0��N!��D�F��n[+=�)(JZ'ױ��MJ)u��C����~/���~��Jd�#{���#x|)al��N%�#æ:%���A����
2rQ�  qq�3�8 ^wn" ]!��}/������A�"�/{ �wr8\Mq�>�ml6՚�nמ��t֠rl��1�9�1l��9n �Ż>Qs�b�h�Ԇ�p6~�-���"����'	`��xAP��]�]���'��2�SEN��
�ೋr(,Z؟?K����n�N��C؈U�˩O���?���E��f��Aׅ���ukI�\���S$�t.yL��6��m�J��yl�˯1<�?s`L,�` ��1|KN������C~��*�L!ڊ̓��SO�D�y*O�4S,�/�B�n��(�L�����ɟ�� �>�����XK��Ԫ��f�v�7���X@��4N�_�W;��]�����}��Z�]�5�BB&��N�Ɏ�H�IV;�/�������ׅl�^sO�Uw�ɸ ;����`��v�"s�V�;������(E�Yt�ǲ��򥗌#���:��\��ʪ��M!����3Sx��1��F��!b�"�0��ܼ9꫹:9e9�8�:'��4N�t$�3R�UK�����fjf�y;�������6�4��j?j����ʹ��o[x�vְ��!~�1�Ln��k�$r��4�6ӔH��څ62Ь�c*�S�+b��U/6�.%��FL@�gQ��g%6��@΁y�'}	����Q���_�?�J�}��D�Ȏ�5�m/��~j���ߘ[�q9]l�$i�WzMѫ��[���,s8M���0�lI(2(��s�Lf�d�������9�^8�����sT����)Ί�>Q�1����Zʔ�Z����1���Q]Ɏ����
���2��q����mH���������@вa3��L8Et�кZZ��Y��^�b(��Յ3	�Ԭ�(�}1�I��~jy>\�K8j�7[��?�?�3�RL0�-g17����ΚVy�M����?ٔ�U�eu�e�gp��	�Z뷥�68�����3�F�+h����xUfaD���ڼ�^v�+v�wc��wn2���Z��X
�A-=��"$�n�<{��рu��H���$: nq|�2��O(�x���ȊrY#��(����v�zI�lI�`8;�m�<�w��Q�u�E�rz,���w,�m
�����D�˚�!��q=3�2��&�i���r��5z>/1�<�K]�UxU���ڮ՟͕r�<0����'��to	@��b�礽f^
��$��id$H��9�Yq\��gl��c}$��q�%L�M��k�aW0�2E�tAh�Y\�6���8�ŊP���oO��V��X���4�}�;�={:�x�/쭟lZ>8�7&U�[��XO�2���T���\]Jǻ��(8-Y��MP~j�EŐ*��r�9��m ���*�)���j��
��;c`�q�o����D`�BE"XձP4$D#�� xP���H����f�Y�"���PIں!m�"9�5�]h�洤 IT�I�\�JU#IM���������'O��)�e�WkzF͔��[M�3��5�?Z A�V6�:�:U�p6�Y��9����_|c)KY󪡦�Wvs}����߄�|1����D�F�BP����CU�c9�սw�c��賀��g���N�����za�״�KX�@����č�^pD���Y��QH��f���f���R����l{�L�M���bG�~��O?u�
��0�>;��=�
�{��r*h;Yiv�5U-ɩ��|8 �k��I3i�3_�&.�`�N���P�xU!�P
>X�	�� "RO�Ai��<�����"Ms=\f�Y�T�����T�"��`K��d!�˙�@kG3I���>�[G�o�z6URFX���W�p��c�aHaa�a�`a,5�0�K.���a����Hd�D8'�[&����@;���"Y�=գ��q]%���4h�P�)G�j0a�~��:����1�[��ٗ�"d
���H!~��i��yY�l��X�=њ^7�n%L&$��W��v�列��٧Ə�6��F^�f��߽�� [y��v�Go�������~8sǮŲ��}oթ��k��������uo&�V7h����Aˀ!�2/��%~?-�x����|����F�N/N��<M<4�V��'bA��O��2�9nNo�[�P;��A�f�}��B���{��qJv����Ө5����c���8��=f,������
����
�цN�!	(R��L��[F��rWh���E�:4.��&ʖ͗�e~Ihӭ�6�	�T*Z>���q�b�@1�k"�����U���"A�	k. &V��O������m�w�k|�<�0��#qmS̋���jG+��U�ȖܨPtN��?�I�L���ځ�'[7�����B&�� ��F�����Ε�����g�P�5W��^e� s�׀V*�p�\'D��l100�q�qB>T�^���,�v4�@B��j����(�`nfv5�������pS���q��4��.7T�E�J%��5��AX���oL^��E��:� j G;��u�h�������ڛw&'���������l����8z{�P$ΙR����[KO�0��un���ݖƌF�:7�����������kY+��(�<]1\>9���:�����8�����/�{y/�>�ޅ	~��l��r�%z����{��I�n��ld����@9;M!gP���tH��n<8<zI6@�<��ㅞ^2��4�ѱ^Q��Y�8�f6L>��B��@�ZO#�&|4�)5 �-�m���r�e@�_^=l+�BN��<�S�N0���A�F�ɡS�ɬ��4De�;��p����c×%��G�N��h���#�ΩJ���;��f`F�ٞ��;����K��C�#1��I�'H�P����/���#3��M��`�A#��}�01��Oo�����>�=BV�0��F5�{�!�!]=0du5��<N�a��v���$�TU�l��*#�G��D}�=��io#O�%�d��JS;�w�}x�Ȩ;,G���Nm��?�K�?�
T��%�b�Ι�3��n.�E.b���(��Bi�	�"'���U��Y���=xE�}7�M.������k�D���h?.���@:�l�:��l��x���."��(�f��c�	�|S9��E���V�k)�3߉��8��?�)Bt�h	���*��#
���ӏ\Dfqox�v"��Ss�h�Jn��\ =���( �^|@�vE��Z��i2j�z������;��}w1~�xݮ(��ٻC\X|.&Y���}迥�Q(-�9���*�g6݇�uֆ�z"�ec"��g��V�8g'gx.�K�
թnY�L���F��$ �WҎ�g�t_���l(ǻ"�{�/�� �Q����{Lk�w���+��9�!�spPF.z'� W�<J��Ȃ`X�U���6E�F�)�c�EE,�\���.E�1�"t���e����W�[`�4�E���Q��F�
�z	�Y�e��<S�a�ԍfу��K�lO�J����=�"\�G M�V,���E����6Y����@�<�@�2�@��~εU8<�ؗU"���T��L�C�4������U��oA�I�R^�(�"|�m���YǓ'�"=(�{�H��ӳF������oƆV]��e�W�x����R?a���Af�E,.�J�;�)��F��W%�Р
�E�x�����4��5��*��₈�킕Kj2El�	��K����ۑ�qH3a\ ZTDݹ�כ9�D�h@����/@����#�\H�c��U3"�/yu�6�)qͮ��A=l�r��)��isP��*�0~��K�l�]Bm�a�/�- e����	����&R�*����v��Q*O�d����8ݯb���Z��@�!K'�a�o�]�Q�5*�$ ��� 1�ﾭ�����'�[	�ae2�K��F�r���ևD7�vxZ��Al�.N�G���w��o;��/�9oGow'�o6ʤ�Ϙ��-�ZS�]Xyy|.%��sNn�N,ngN(Zh��Zj��ﴷ_w�X�3��$�_&��_!���YLJ+��k�>p�������-%1E�M�Թm`�g:vV��o�	ɸ�"3��	wP��D�L�=���!���i��%�A���4��fٚ�h'�.Yzd�h�[��7㼎f�T&km%�4��,���L��3�� ��	#����C,�~���E)��@�$u���s�!�=�W~�$�mg�)rn��x$��*�ϥO�{�&ǸJ	��-c���|\S|WLS�����e����/;
��*D?����l}Eyp�@r�~�P:6H��1���-���e|g�uwƱ��q�����x��N i�}�؜6��t���s�A�%T�BS��%U��M�T����y:�UҠ��u�6�z���U�RJG��C�e�dDNY��{�2kz�	��r��L^�G�����_A�T�f����u���eT�@V�x��\uM
ߟ>��{�"��I< �a�wZl��� �S6���ж<;`SW�>��Y���XX&�Ɨ�����Rk��;��	�Q
�!�&�e���n�	/z���<9:::<Kںz��g2��']6��n�>nna�������#�һY��L���`Y��Ѭ�GMcO	��TP��W9���B�����(�'��J�������������F�<��U�`o��tCs�T=�����j�;W͈�8ϒדy��gNؠ^vGM%�nr�3��auU�?�2��$�:�C����$�����KZKf�i�;,K'�t�~�I�rN�/����3xRHD<�h�vL��r�C�5G�čL1�QJ~�a��C�b�u�Kw97��������eZ��HX\ɇ��J�Ӱ��6U� *P�S�X�W���>�not
��DN�s4txC\q6�����h��eÂ��C~4+����Q#���)�C:r���z�!}���ꜹY�2�6&��X�e�z���M둛��g��Ѩ4�E!%��z�g⟁+��,H�e����5ڌ^K���U	\��\�3,w��^?,>�tKG�7JǺf�ԡ����h$��M�j����k|���t�<��g<#����l~�S�ٍ`ر���ű����0<@q�}��ӓ�'�/ A>���'A�l4_/��������O����~��V��U	�-Za�l�s�t|��P�ʢ���+	�3Փo?Y�\�A<��j
(�3��倣��Nv���mkh�Cs�R.4W�(�
B#/�\	GS�=�Uxu
�,�cI �Q7
�=�<���`��S�b6�	�n!�8]�C/����]!�]v�l�� ��"T·�t�%�J;!y���I��Y���,^�����bb�	��h4N&Yp�q�E�;�EJ�o��eӞ�7�!�/�K���=�Cy�T!����He؀	T��Lq��6s,CNd��&-�1y5�wr�Ϸ��~�<)�:$;I/;Y���v��t����!�{�Bh��������8�ND��L��t-���8��T-ʯ��֒������oF��3�.J����߻��E�������v���L��^�"���kB	�5"O��Cl*<L���#�"[�A6DX�#0�gm~"�\4!o��+e�YUYe1��GS���/sr-�G'�PX%[���	�B�&�r���J��R����tb�}��ћ�R�-_ ���'����
��0�;�.m"�����Fm�1؈�t�_A�p�����b��!6� ���� P.��tD��r�R�"D/��ꨖ�s��;#Bl������;��:ymlgRAqp�g�$���WjǢT1�Ȭ��5��]�����$��zp:3𧢿�%�28�Oo�.0���e��E��E��5,�Ȑ�ߐ�א^H�>$I7����kSs����	i�X	�(x~��jyJ��0c�l����,����_�7H�z�l����ǟφ~�A�Z�YlC�0nZ�i��N(m"�b�1��y�$��)$����)�Q�B]z}��*q�lBKw�2v�*P�������R����t5!vɋ(̭��U��J������~O��R8���J�rt�m�ð�7��!����!����
C�=g��w�p�Ny`]qS����XY�W��z��d�I��0��#形G�!�V��8lF��aO�t���pY��=�Qv(5�N����Vs[?��3'Cle-t���vY(U5����bUh[*�)���Ƿ�Jm�r�=cƕk�O~ԛO�}g�	�.R�jI[�/"�G{u��d��bD �r��.�t�9�s藑,����j�X2 MQ�s19�L�$�}6'i�*�,I1)�(ЌN�6��P&�V[pؕ�){��"hPL�ь��.i��DrR)��oH�o��A�b}�4�8�h�zq
�S�\?��������EΈ�B�E���5ry
�O�������a�_f^��G��t�=�%�T�jǧscEl��_� ���?�i>�q}�ć�'k�k�*�R��6s�gL�DJRFh�c�<�`Ď���r4GFF��m�iV ~��-#�V�$Z�;8�{,]�F/���k�;����q�T�`��)b�xȹ�`��μ���0�������8�v��R�������f �a�T���[�sԖ,����i!}�Vf1�ڂCju��5�qx�����D�G➘��(��UxT���$�C���t��	(�J���3��.?S� t����T���C�&�\��hn\��I���\ ��ۦ��yaɈ5g�ʎ?2�d��M�1�*��7���П2Ļ��E��G�b[�g�f��2�HD~pP�N�9�4��ש��B6���R����_,uZ���Gj˂"�ʘǙ/�B�H��Cw:�"�>P��#��xp��'ڳ��8\�tD^MU�H�Z�K��%�ر�+U�(ź�1K-����A�v�ҕtF��e�Lj�R?K1^SY�9�5*�AK)}�]ퟙ3���Ҡ>d�>kl�Y�!��o�d�[P$��kd6� D�`�@�=m-d2�6�?��42j>��T���U$7�FCI�4��'I�R�6hѭ�c�ŗ5c�A��d�D�Ƃ��WNL�\�ʴ�C���� Zg9]k!y'���yS�}wF�%>r�:c��v���v��3<At���e�<A��k�c���#A��o��/���BRZ�KP���0������{2L#�F��A5�6����H6�"�\6�ʦ�g"�F�2I1���mV|ʘ�7'�T�m�����q+(�x�G��$����%ޝ4�=̾>�ǭ��J�8s笪�m�]�-*&^����V����ʄg���OEE%,�Y]��Ͽ|vgea!*�-Q޾��k����i}txx�f���33���+��]�Ãzz�f}�2<�'�f#jld���e��]&ղ��Q��#ɣ,��G}LF�NZ �6=E��i�����S2��yꐙ��hF����ҫ�zb����+ �F��)����rn!�RN�2��'�"��T��*%c�GK���8tT'����pv�T	DX����m'�{�Ns:��'~�������덈��u�b�99�L�C�D�A��&5oYrcB�L�7UU�6ɧW�*h�a�JT
'ur��� nƸ��#�}kQxRE�l�������q��.}t��u^3g3��~��8O6���甎ys��Ek������/��?gd+'�]H����6*����g����k_47��q�أ���[3��� 3T��T��u|i�뮹2��A�֥ ���7�Y��0�߾��?C�Jy�X���;/�*(>Q$�-��2aɎ�6�����O��ƿ�?��	�=w0���}��e�
�b�5bXo_�z�~���. �|��Ѹ���s\(�����Yg}���������N�T>����{orc��qt&��c��z�k�@P�K�0�_��z��r���OӬ�oѶy�]����ɥ[�������4��V�%��P�X��)Ot�� �2ؖ�T�X��a1L�X�ڬ��!��X���8�� �KŔZ��/��<�����> ��u�ozt(������@�շ���E��&Sl�oT�ȋRA�rs����B�BTY��@þ	~ ���@��<�p v��3=���0���B��j�o���,O��D;*R�񳧣����\v剎��n
�.�^�}&��i�M���#�t
�$Fڠ�F�{��x�'���mf:IuJC�]I�K�K����4��Mv���έ�t�����)�Ccڞ@ݙT���3	h+�{�*���q��YS�:�F6�/;LC��6q�g�C�~g����ZΊ�U�x��d�MX�Z�\{c~[/��X['����`��yĆ���������4�%?��C�����O ���6�,V�ǘ1����\LM1�q�@8θ<_^���[���4��U�P��Ux�!i�Diq%�;@q-�g}���L  �����6���^t��z��1r��ZQ�j" <�K�a�h��A8�̧2p���؉M���"&Ԭ�����k��Uu!�����w~�J�n���9��0��;�XM�5j����jblko�cv;�����vao`�rPuۖ<����|�����u�����6���Cvf�k-�f�����aS�_��3M+��sn�5��5��5|��X&L@xy:��!=�/�N�	��T���B���½���t�[�Dv���Ft��$u�<��=�4��vnqa�a�MsS��1�E]���@�ݽ�05�I�R�Y��f��oP#zI�˷�X�e��������*s��?�Y,��v��N֑"�������8�Nmi&o"	��m�.�E��ھ����e�^h��Ml�E�vY�%�S?�Ay ��$���N
��ł���?��~���I��$�׻"�k���G�=`��o�Mg�C�=B,����8���iE@��Ay+��qI�����Y�t�K��b�,��li̓d����Й`���o�r�x;Ԅ.�����xq�9�%�2a��`���4,X��_ϥ1,���*F�+��p�!ď�w��rL���	�G��%��f�Uy��t�h�%�[��J��(��B��	��O�spA,Q��O���p�I�Dh"dB-(��r�U#�H�4�qS����Mc�M#a5�d�2�ZJ��3�U��]O����^aq=p^�l;i$�\�ZV���� K-�%e�~�:1'9Yᙎ��/��k�5,��R���t���]��V��tO-F	,ߵ��oG��B�y����п��݅���X(Q���W�s�w�������\'��)���y|"SJ�/cLǵKm;C$'D)�qo�b%e��u�����n������K����N�Z˛��QUc|��llM��]UR�a��AK��d�8�1.��Y0�|d)��	��`M��b�ЛK���/
�����V����|�F-׮�DLp���`���$���&��	���[���E��A��N��x�tb�(�^0�m�7熋�*on ��e�#�V�=��T&�����`hY��km�0���+9_�(A�k��E|�ND�FA3J�Lq� X��B�U�-��\T�'��䡼x�z�����vP�t�/�@��*�8�Ėv����/�5\�yXEh���V*�B��8wcS:���
���g����| n��{�U�1��ܼ������G�� `A�^BQѶ-s9��QnA���6OG/�l� ���u�i����,jݨ��GK�� +ޝ���U��/Q�x.��*[���	!���
�+����}7B�~!5�7�Q��[���YE
���%�%�e�%]�
b��Ζ��Po8���P:��vc�������}|9�|{]v�|����n�1���0�j��W<�����p�v���Kb/�x�g�ݫ7����Y��JX�"AG��Sz��OU��E	�u�5�%�bevbL�����9�~;|Z��P�FF���Ι0vn��Q)T��d_:~x�(@�p
�ӳ��rr��]-�xhgH1&3&˱�UT�[[WUU���\g��IKK�����;)++�C��3{�]�.
b�T�%����}q��~S�w��T;�b1j��b kuZl���%�b~&Ahp�CC(*%�rt�#�ŗ�Gm������cHF.��ل	[���l�ic<��!~M��ڐ�*�������e�^�7F��`�����K��%�mS��x:�����;�TЫW�Em?R�CݤG�;�	��/0���-�q��4 gԼ����jhnQH�6��fB]����N#%�ȭ٢��K�"hX���?�F�eC�>�W��U�1:��S�N8�R�(��[&�՗׺�Vbc�hmQ(���ie�8���;���zYɥ���m��������t��]�3I� �b��ٷɄ�$�۹�m�$��e�G��E���_�&>�t�Jq�H���1��n��
���\	�2��r���u^��k�����L@�xrUR��rj;bY!�h�5��`.����ږ ?+%))-铛��i[��d��,���/Y�ޗ�V��V��ӕҵ�:��W�Ƨ����I�!;������Te�l���N��>ʻ�ϭ����T�Fk^��W��|�溾��\�n~�:�!P�2 n��t���_S:[�ZM�TB�jwG"[�#k�kW�f*X\������&���a{�+q�υ�=O
 ����O'r W&�0��$v�̠���w���WN�i�@Q4f%�M��"��4{�z���<�m���L�}3Y�M�7\9������Q-'�J�P�뾏<�,�A�Y���&���������ur���T�cȮ�9l���N۴�ή[��Ȗ��:8f���.#�	~ʢa�vk�/�'|Y�:R��q��͞� oCy/i
/]�o"t�~��B*�g�M��zpH�/��>��<�Z�{��(8�Ș[��:��=����X��z��p�geX����������XvT��X{����%�Wj��"8��\���6˪�"c9��ɯ	��2���c�~�����	(m�|�$[�SN�8H�����MB���ζ��H�q����P�:8�8�:y��aՖ@�ʢH�tuTY��J:�ϖTDȠ��;��%��� Ƕ�o�[���2��;��'�G�v	����nfd���g<?�
t-����ƌ5���g<��Ħc�,��ZYK��fbv�z[E�Y3���J.
��5L�5{sscI�\ �nh�&&�{q�7��l{��0����vx������ά�ն�h��hSw�=	����iن��(���bqF|�H���|GY~@qPT.k� �ĉ�}��V�  �*���:�(J��?\�}ԐxR���j�P���KW�z)��/�S�E���B�MʃԲi��{�|��n��a����rO;��S\m�ZfON���^����������l�FD����D�H��;և�|����D�qZ�Dxm�}�1V����.b���o;-$q?Dxt��1|��x�7��v_�6�������銲O�O�� �4�'x,{�2�c|[`�V�t:����7����~i���*�*C*i�"��܁h��* N��V�E��9&w���y���]�������V
�#�iĄ@�Mk�z���.t��ϲ$SU ��[*,�N{�s�ОCJT�x;(BKf�+���I&�cX�
Y[�A�Wn�4]�!�7Ȁ���������{��籝o����;V8T⥦^H�u�TN/�{NC��I�(hif��%8X�"d#�.�Hh�df��C�sk��02$���e��k6�n/wF	`��+)�Hb~�l~�������Pk���k[+�P*����o�v�F�$&��"E��/��l�{d�}���bos�Y�q�_�m}�]�x{y{>�O};]q|�	�V\o)�n�Ky��u�U�6�bA�m���G]4�/|�<���Mv�0����j=K4���.��?�i��tD>�/
�tGW,^�v˖�.*zGe�]�EDrL��{��[�9a\5��8FD��X25���U ��l�D��Xp:��/5A���=S��J���Xɏ���r3��T϶K�**�]�`{�dQ��:���i�k�Y��
x�J`mW�a� *g���H22� �^\�9�p��)�UG�s!�`�\�B��8`թ�VLB6{�>�b�E�T�3�1/@��v� M��WC�3.ܵs�-��?E�zux�y�T�Շ�J�|J0��h&��nt���C���V�`���hp�l�$��(>^dVe\��z����{�����92\���\�#4u,A�D�(�DC�2Q�}����e�LaS�y�I1�S�E<�B�e=��P*ZJ�籑����щ�k>c�"�`dJ���1� �o1H,A�����.��2������3���Ljr�\��hv��tnI1+,�F0qF����_e
�d�d=���t����t�4��Fv��_���v	Մ�=�5b�
��6��⥽�TJ�Uܜ�u���MM��yyy7��\�!j���wO�����HHH|||����GGeee� ���`������?������͖���)�&�I�Y9lD���#�8uE�>oq;�ّ��⳴{z����B�����-T�p�
�)�,
�m���E �@ >��CN���8ԣXͳ}ĩ�/����t(~D�|uf��/�b�C3��i]x�62,������%�'_�C�0�>/�C�2D�YS$��pt�_��݄pnc�7�vJ�Q�ꉐ_��`�L]������)�m0ň���;"�	�gU��H�f��y����%��X�@/֠ ��I���b�&0rށ���,f���;�TN!&��� �:8��%IwB�´H����'۲�3f�v�/�)��.�H�4���K��q��qȶ�"�>%�Sa��ϵ��o��t���=��2�'e�G���m�*�^R��,]:��u�%%ke�M���1�0\\TY�����;7�!ģ��mlRo���؆�+�{Z��3h�ht�Yl���ܟ��;�!%���%F�w����|�dv|y�u���̿��W9�L(Z�O��m���o�{��cћӧ)O�Ƴ��[ݳ	�ѣ��u�߃��Q��G?�\��P�hB;j��f�k���������(ؚ���Q$(e6W�P&\�w�ڝ�E�d��҃�cIiĮ�+��Ni9I�?�PG+�$�d����|.`d0�a,�I}���p�6�yɭ��_��5;���<0q��=2��~@��b-NQ�Ub�.O�xQGT`˚�)C�9�Z}V`��KYbNiB�6�r�]&�����@����k�m\k��Tx84oc���\ֱ&��I��"��{�?K*hH�/�,'"L&�K.������a�O�M�ۤM��%'��C�v��e�L��͌��2���t��G� [��$�ʤ9c�
{���F<�d��Q�Lܷ��}qa�(����SHy`���E��ϊKD	�"aڞ���Ff o�:	N���Um��՜��(�ܑ�f���^����������\�0�\���
CJ�}5��&D�$0)�U(�/�χi��u��_��q�l/u�m	�W�PN/e��-^�\�d��7jU9V(�JI���@.�y �Z�c��sD��ߞ���~!;^'n�׷/�\~�!+��BRz!�^��mHK�.���t�QQ=�)�n�\�wi�a������D:�c�ZX��D�$鐖�.����<�s�}1羘3�̝�̜�Խ�3�\_Z6%_�]�9�������pP2$�~BNٽ��g�	S��=��D�g�Gnn�	N07�(�5����^6Q*��I֣����V�|<�X�{��G���wv1��6�UYet�+}�t v�Qw����������-���M�kJ���@��'��N�-	�b��n{��[5��R�ȇM��2m�L���2�mz��\C�)Ya�5`�̡�ǝ�������=�?�5ȯT�h��]��,����w���4:��,w�y0<�.~ȷ{�Ǧk�k�ZN�߯E6 �vaI��Y����E�*cE���j�c�]r^����NHv������f�TAնSH�7z�#�^R`��2����R��`0��P,�"��B;vU2�|�_�g%8r!))� _ՏI�d�ր�H��#<WjZK�8��$�����G�+�Qג����@x����@~�65J�0�T�J����?�<�̵���T����rh��۷nl�����W�-m�w��~�+�z�]����cG��\1n�?eY�H��1Β���h�o�R��&���ۡǣ��[�ǵ�_^�\ޝ}��W:hS����( ����ӕ+Z���0X����w���Pt�����hTșP��;��
�+Z�4:
:>*�BAD1x������v�^�����)��}T�A{��i��F���G�/yX�o�w.lx�5d4{���N���������7uq����^����=��?��y���������a�����7�֊��6�������;��Uo�_��5���b>�*�[��h��&�3�2d�S�ǀ�Q��*�R��Fm4U(�#4�SS��2��ɍ���=-�i�+ ��Lw��d/��vIGCz�6��a`cņ*V�F;����qc���qoۖrH�T���{��mh.B��B��~<�-�%�)5q�!6!���Ŭ��X8	i�R��u���O��K����8$oI1�8H`� �ŐF6� �KH�	��Uq�_�����Q�����K:�Xi�O�i�����Q'#4�{�f�\"�J�
ߗ����ڝH�܈�}�ਜ਼�]�nNE�/����z�wRj��xV�9amX���Gd5��M�]B0��C�R��	�V�Oc��׌���ǚ�#C
̻f�	��PDx�� k�Z��_*(V4f^��Ck�0���Q`ńz��z�E�65�SQ��7��n�0C/?\fA^i6�����,~@·r��L�@� GC *�=�ۣ9�x���B��� =0$*��3�}&~�1��[�4�S��/rs�TmO���k��tڔ�RU{�y]7�
e�����2��ɞB.
�k��S�(p��a��*��:fb������ee\��CC؍�,,�Ӹ��5%%Vff��;P(����������	��D"�������l�K<勋����}���˼_�"�ao\ڱ�Gx�N@����k��BR]rRF�O��o"���$�슺�V�5�>-_@W��t�rs,4�.��@ŖH�>�P�Ww����A �ǀ�D�Z�7��q�s��|E��'~ū*(d�QN-2���E��&��fJMlf��<���(�B|3���
�`N���7� OW���uf���Y���8>��}A^���1�M{R�I��c7GO�����I�7����|8�p4�%��/�^���1|�r��t��Ț�����g�a�����F�3���;xMVR
ެL�goõw����)�����(���E��E��E��.��t�j���r�!J�|�փ|i[�.�Z8�"���+}�#b/+#ؙIr{����L!.ZT\P��=}�����7-�!�Ps"�&^���{
X�����w��|(�^RD��C'Ou[xv���zA4��c����}�����r��>�S� mt�X��u�7ul���Y��&_� X�W���lZ#Y���鹁�"w�s���7�v����5uQcʝ�AKH��J����L8B��P��+�"�-D��W§97�4(6�ft���V��~t2=��[����f�K�|��a��b�kt���ߧ����[gr�)�H���%�+�4Sc9b�>%J�$�������>	��~�Da-м�솜�O,��52sfkAmg��%��O�l�"��6���Jsx����u;J�Z����*��C$�2y��ZL�Y��緢�32��D*&��XFK�dN�w����l�͐���#7o�ai�i~�ۆ�Hb�x"���7�r\7" ��;WԼ?!���V����S�"��(�:�7Z�$����H�gX(�(��]�L�Ⱥ A�4���}�[H�g���r����rH|/�K��~|��Ҵ׎�N��L��:kq��C�H��h{0�=�`aA��8��h�f&ڿ�������6n�����sz&����8d�!O�!O�Nyb�<�S��O�����5��@�À�3?!�qp��7y�N�rb��}:2\��3罡ПZt�Om�NO�������}�÷��o�q���MJh�F>�A��4&?��\���������x��u�5D�"1M�A�)��nL?�	Ǖ���ibOu�|�9��+7-��q�
����ͯqЊU�^N]���I�!�f �Q�u6�#t����Y騄�[�,�L-� ��-r�{b��	xp��	zB���+��[�{�:U�S{�.`�,3 �˫�ު���8�i�O�Յ.�c��˽�{��.>�i�[����\�/�2��2�,�o�P���PկS�T�uX� ���^�z[uы<P�U{E+K��ݎ#�e��Y3`Jw��֝�����E;��k�ee������T��Qsk��2���e���Q�r�&c��:&3�����*��)
��f��K����Ʌ�	��P�B3
����6�sBY�<�詠��Y|�W�YQ�	x��f��i��賬�p�yN%bƗ?ZZ-<�>ތT�>?xj����"�"b���1����>�tr`\֟�p^����c��0l��u�s�>S��։�5ZTX,\f��k��*fxBl����â㔊F}��Q��RҒQё�b��%M�y��p �O��ivؙ�4y/��:J{�띏0~F��):�ԕ��DW^;L&�x�Rp�UBG/���h��-?tS�����]&����ؽe�~{.����{��W�Ot�����%2���P����PK����;��[�k�n�#���~m��a[Vj��U� ��~˓
cJC�O���z���k��D�MVS?lk���K%�Q*��d\��?���h��y	���m����w�<|��}�S�r��'�q�u����3z�}K��c)�kO�4r�xq�b�~#�~\F�ѫGGw**�wc��x��S�w��	��P��)��I��x<�{F*M1.��Wp|��)!�q���4�����V_���N2qig��2S�mgr�j���D#���"d��#���잊I�E�
/���p��S�_���ǻA��
��H���{CD�������	k�"X��' s�TO��&P���
J���2�Jǯ�R~ͨ(�5+TjwXҖ��&�m��uf�0�GI���ֹ�@�����R��/��N��{p4���M����N"'Wt�	�tx�\$Ĳ���p�D>�>�A�{j�Q�ۖ(A�6��K���v�~�i���	=��<>b1^�Z�d�>�L&�����p"��vx&�d,���̅���J�c�m� �k����*5---%e}sQR�/��R�*��`���eee����yk%����_�������P�Y���oy���!�xGƖ�>
�:xO蹋���j��Ժ=�_�]������t��s-@���f���g�� c���4�-;.����LT�)�c�T���짫X�k�r������}z��Y��'�ք��gO�l�����:]�*�X�cX�z���Ծ�`B��2���B��Zd2T)��W�������،D|L?�XK��|��G�hٝ$c��>��q�W�wF�6};�ٸ_�l�$4�AK�g�Q�F���oK��L��ih����Z��+����ʯN�=Od/X�ץ��myaq�TH]���<����?����ͭ�Q�`Dg>�C�����P9V ޛ9�H�E�S�(�d>�V�*L���IVU���%���X���Ռ��J�^�i���[Gj�KȪeO���TbUJr�O&g$�&d�'���_�=]l�-fG�e�{�̋k,���=����Gr�~��):��\��Xx%:���r�fB�h�ss5$�-�т�>��R��TE�v����>�6�)�����m৲N^��(/ο��I߱)}�*V�B 5�ꚑ�ض�O��$b�4?W�'�:�"�'�e��V&e�/�n�(�4���XQ���s�ݴ��vѤ_L%���͉~oGĮ�v�<���(�+3�0L#n�M�_-�ec]P��)Lk��|>v���>�-�kV|X`tJ����E�@�rc�����>���.�2�=�[��-H�M��������2����0h,CՠV)i3��#C���"a�	�h��_Z�G6�Z.���45���Wc�݄��Lq�Y�}p�j�_���yi7cv�'�~[�6[��&D
g�iR]�D�Ag0,����H���'�M�V�L$
RЎ�3���ɄQ�3Z[3%GS"�k�2;���}N5щ�L'p,2�d���6��0A���MT,�
°5[��,ud��!��=b�y�!rhV�O��f.q&��+
И�<<m~�˶Vɹ��O�-%�gN��b:��A{#s�Y�7'6G�RA$���?��\)�N�2@�������m�p���'
��M*�>�����+�t�A����0kFz����F���6S���ߝ\ ��C�ݵ�#|e�T�d~n�ycQA-����v����ӻ-[fQ�3APy�6��H����׀l[��`}� ����yNy|�Ο�$��D��ͺ�q��靚��?������;�&�]�V ]H�r��<��Pf'@����tF�O��􉃯�U�k_�ϋ2���K��^�-����{��P�3�A{�/7*Ϗ8�Y�Q��:w���䋉N?���l�����>�go���6�w���l��$����ZB�|�-/�ܥ	����8�h�:������ɻ	Kc���n�5���QT�������o�C"u�����x����d^D4>>��(��3US�
UM���A>n���e\���-�e՞(X����q�E�������\���������t�����F�c�V�u�NI�SD�s&�1�T�b s����b�df��R$�	V���n}m&b_�U4���G�Q2�c����"<>���Ճ W-�M����'߱x���7o�%~���v���"�)�veqVn���6z��NI{��0K�C�%�_ٔ3\ �Mjv�r�;B28}@���wu+���a���\����������9�;��_���f��K=<�p�>�ˆn�D_ �*ڪ�Vi��(��N4Z���܍s|k�D�x�Zi��e�W�����z�0@!�]$s�J$�5^���A�e9�ofl�6d�P�ҌN�4�P>XkZ=\j�b ��������k���ޖ�	_�5�I���oM�^R;��!�o�=	�?�*v$(��*ː ♹K��7��=^�5�UIFa�F�v׎J���ű)Z`��0P��p�� 	b�>�FsV�XI�T(u{�{1P5�2���"x �_�hp�������
�r�fT��t̅L�*xԥ����[�H����R���2�}�`U5N�:���l�ܢ7<����|��`�9B�nSB�r�;m>���hT���{�s{zp����kEm�ge��el�g���֐��{c�B#�D�������u�C�
_�P'Ţ�P�\�T{p�62E��`�+�-������]*{L���>qe��F˜��n�v�3��S"��Ŀ S��-6RPu$�;%9UWG�Z��l�>�[Yï��<J(t߲[`q�A���B��w�M��\���R�^��`������A���M.�� �ɀg�Q}�����z��t�kḊ��2+��L��� ���**B���L��`0�)ϝ񒨨��RMooojjjK�����H�*�'/�TUU333�;�
��^�`����GG���gR�b���r���[V��v��wzN�FT��j+S>M��^�n����%��?������Ne�� 
8|.l�0\Xlh=b�o(�=�J.��ۘ��
N���>�^F'\_r�dS��?Y�������c]��ԟh�{��o���b�yx��3��~�ֶ'�$��s��;����4&��|Cы��.}_�-D�Ǫ<̠p�y?�X�<����ֺ����]����O%�qjՌ��)���e������rȑ�?���oSt��hv�pl�L�)�$O�ac2��ܥ;���0�p�'�*����+ �֭Ez���(w��.	sz�E��K�s���2��=wUjM�g-b}�"]���|��qkڻ�y��9,L9��/^k�lp��4|8�C��3l�m�I7��JX��~"U�m������Swv�;��sAk�����>���/�+�칝�R?�ٞ���q$hy���P��p�3 li��.5>�>����WRWw�yS�_�Z[)�S��aί:��Giu�DЈ��B놶����A��!T�őW�Q���0�S�d�ͫ��ؗ8eՖh\e����fW��ݶ�����6��'��'����
��He�f�$��+b{M��I����64o'{
B'0{�����4����4o+2]f`���O�:g~�ǭ[�1��k���ܷ��M8}H[�>���Tq���ಯ̪ؒ����Sltz&�1A�c�+���}�]�2�/��ߴ�+��;AU��>B֪�ܿ�R&�?�i�b��/��X�Ҡ���I�Tqʴj�?��ڀD�~�lL*k�(�L/~�Y����9 H.�*�l������3T��s!�/��[E�@ ��k�e3M��K��N-`�`��T\�� D8�T*�tծ#@_��Ɏ:��>���b�2;,9or�� ��\lq�Z�Q���.7_���a�+38��Xb�̹=���-��q^>�r5�������{a+!5�а���1*l�b���>./?1�)���<^����{\閶�g�3�¬��,��Q	����~��"�<��-ON~0�h���L,��a_C{'+�B�	�N��̬k�'z����0��v�`
�o��@	}����tH%�#�A˟`gR�ش�@�A)Wr����G"���k{|��i��=�8ט�õ8|��C'�-Ơ���,�����Ǽd;=ЎM��ˮ���dS�/ذ�y"񸯔����7j��2y�t�@����;2��X6>���*1v#ą�yi��ow��hl�R���_Ï ��U"w��Ǖ�W�ڹB�_���a��r�g��z�����?�����ڶy�fZţn��MB�\����e���SƢ���l���ũp+�]p�H�!�;l�4�Y~�R����v��aK�w��n�%2����+�5<*�ؼ����W�e��jU����򖍢|'L����#÷�M�H�:��!�h�S���Y-�W�W�#��W��VV����S1��4��<֧�WG��Ao#�＃.����^��-��M8�]G�yW]�H��߄l�.n�_
0��ʼ����.���C~g�D�u$dk��$��+���N��W>�^-��tD�<뢽���a��`�x�a�Un*#�"C~J�&�dE��=
%�V�X�%}R&�*�)���s�7I�w�W�<�)�w���5�����wf�n�����?�i��m|�2�ǩۨ�9j���6�̀�� �)h%_:u��Z��ġ��z��Y��+���0j�;��AcC�ɽw���r�m�xc�g%%��?Bbq�+�U��OԵ�?�A��_����3�L�PIT��Z���1���Ց?���E��ĸ�B %uV�tH#*x;��qsΰ��!�m���3p=-��_7�\����zi�ST���b������b����օ��x����*�{��8EN�/XވԠ� c����Y�"����r��.J��t��0Bu��LF,�����T���2[������5(kat�&{����*B>�zc���$jpW���ncO�>.��f��zAs�lm��[>É�c��i2�z��z�Cs[n�>o��!���]�Z����BF�cRAY����r�*R+TᏖ�]f�U�@3 �/���?��z̅g�[�0F^�,?[z�4(�"u�54�֭���4��Ϛ�T�8��YX��`Տ��ϗ�z&~�" �{�( 1Gy���o����,��<n�Q����D��Ҹ���	~f�������Z+��`6o�.�$����S��3�YĿ�8Q���*� �)ڶ�I%<|�������>T�x�>˴� x�d�TTSP��>�L-�>#;[&��.���Ą�@�F隋Ċ��}}�M@�Z�H&x�e[oH�Ug�h�
V7-aq9277geccc��z�XT���ږۂ$�(����� �-�[Q�`���Z���(�\^�-̏'�8~H1�����1/U�/V�/�c��-m�����.�<Qêҭi�g~��?[`�B��rLi�����<��c󺪩 nZ�.&dn��-�!$g�m�
/��#�5��qd�?:��P~��o\T��j�3�36��&ҡ�G���G�*<�6���`O�����3�Ȼ�S1���$T�P��bW"/V<�vh��:1�8ѫ��)�ㄉ�tu���M"hWɾ��u�=������"����*w�d��y��!iS�m�hˊ��c�(p�\��8��$��WƢ�O��ҩ�WOՍ�=�E��S���}��+�h�y�< Yz[b���t ��7oX����kD=l|<,qxX��?.*��9fLH��Q�܈�e�4aNTIuˤKJ�~�a���y�-���גߊ,U�L�m�������j�N�B=����% L�w��̝,��P ���?�����6!�m��+#�+G��`�N��?=����I�&3W�PO��}0C!�4����$�C���A@��6)�
*B���@�rDpOp��U!f�I �:�$�b������(�.�ʓw��v-�1��3�\HDg��&S r������Df���Z������lQ�9>�eE����~m�0@^��|}���z�]r����}$?`��b�:���D����j�M�������C6�o�r�{n@��}���)92���#�Ӣ���(�:������7�[��6&w]��)�dAl�J�"}qp
�Vӽ���.�O��I���:�%'�s|��0ُl�x4\�9�2��{';	o� � _J�� ^(����e�`��4��B�pzϒ�Ya����9]?���|x_���S �)B.�=���w�t�Z���{���Tڍ5%�dXr|n�߅0w"R/"�	B?F��&�5J�	u7=�)(���#�5G rX�N��ˀD���E���E�V�=Qi�^�g%�4�u�g8�="k2m���$ӱIf�$��U|�G�3���X~��,#�5zE H��U�Z�"��=���"�}p�Q]�v��䲏���!N!'N�A.=Y7��|h¡)r�G�3�� ��e#��G-�d�Ԫ�&�a����;�1���@Z�Ȇ��e���ȯ�q��^㞿��ݯy�(��z�(�et8w>�q�Ѽ��P7\\��Tg�YŢ�&����2����laz�5���}F��cV�1s���h)l�ײ!��t�
��Mqȕ�QH����6nKcJa}���]I��t�$e�e�>ƍ��w�݄��Hq�a"�v�~p�Paq�n�`�,S�ҒQD��3����H^�ϧ��#���'���S�V��,�3#tm��W�w��GRCe?B>��h�k��Bn������ۼ�x�";�a)�*�EН�Cgۗ�\�˦Ǯ��oMY_���wwAC�n6�oڃ�6�_���������
o_��(h����c��q�2y�љ!����(3}(�bW歧�7��$�X����.L�))���������zbY]���P�i͘0�,S-���Qk�hU��#�	Ҷ2R^ޏ�ld�� a���$WcWe鉬lBy���/s�K
�S���x>��1&������|������U�uL���z&G�4m���Ξ��[�\�BQ��HҞ|�y/��V���1���m�{y�d����o���dd�q	���]����0��q����!Y���G�%{c�u���+�?�7��)��3�XE��F7F��J�NzP�<O3�˻,�J,g�ZY=�G�
J[2T֯BZ�$�H�z�\��o�<�T4�e��˓FF+ߥmY̅����6���������u��Dp�2'"qXi	Q�{̟�g�ƅiPDB�GZ�9jn�ފ%5bH�a-� �Q*LpU��G��/� X���j�;a�Ҥ��5N����h��dʛI��Zv]�h��|��B��cv����D�y�z��s���	�Z*�uq�a`XU8�:�kK6O���"\$%��S� m�ܙ�R ��c#�P�	U0�0� ��y1|���X1���x���)$��"��o�DGD�;ug�.k�Ph�7nl> ��b[q�ԡ��G�E�@�-Eh+�di�ꢐ��D�W�`�g_�D#q����@��W5�wZC���H��5�V��CV�"��t��Ԃ��y8�-�7�q��n�r	bn/��BOO~aa�m�d�m�T�Z��-So�څ_+��]*�8��B�uC[�LMM1J��/4���_����&�慽昍��oh�,�hL���0=_���I'Ch�	��,�ނ�HY"���=����3B"�٬��忻�/N����maȡu�4�������_CC���Z��%HW9\:ǈ�D��{�t�ߖ\h]�Ҙ��<L?����U���o\�l�W�8��[��+���e����-\��	xf��wSb��*E��^c��2����ѯ� k>	����j[�m=��\� r��nA�2D���`���#�:f����r���i,��݀;C�V�?iM�ĺ����O������@*�$t�����Zm%���s͔��:2����٭�孟��S���K#�ߘ�������1p
5�0�5ʅ[z����L�H@�6�`RÏ�Mձu)����� a)���m��*�Z�~�Xh��_�[�+ ���g���~��Wh����T�$�r �aAE�`�qlFm�PQ������čl��f�*�.��ݯ�Z����	9�M��+��c:ڌ��.��s���
.fm�7�|�-\}*p�J�)a����%X�1!����"-[��sm��Xy!�H�'S\���?��N�2�:r^�'�@�4�-x�������z"n��A�P��@4�O����M����*�jڋ��>����GU�G��z���[@��p᯹�5Qx|���Y�q5���o.�8Bꤪ�C�`Y߅D�"������䟫���Vw�9"�nTz�z�U~b�XL0��n�b�@m�����@�VdEN����L��3������7��M�u��̉�Xe�.� -+uA�i�J]�FV`���4�`�/yQOs���\�� �V��J��Wz�߼zq6$v>yH|��$%�'}G.2F�&�,)�QY�̯����������E!1�3�U�u5C~�M��`� �M�+B�@���4b[ɐo�ab!p/CdGO	u1HJD�=��e
�Bj+�b �
W@b\9SL"�h�1���>�(n]<"��#صcr� �#> �b��mOp�7�������a�}�HI1q��cӎ��N�@q(y�����`������e^���ǚ�?]!յy�^&�NM�F�q��EʤQ��ݷm�4@1��|es��^L��&�B=��;�4�����i�6s��x�Q��z���:��_&M���M�N��+�.6
�2���o�� Wf�Ip'��C(�E��ҿ���-����q5��<��/_Ƿ����@f6��°�W���%�O�'�^c3I_�a��I,��TՁ����qk�E�ZQ0���^v�)��,�Ե+o�qt�ÈV�\խp�T�������?��E�HQﾷ��М��Cƴk1�t�����r�p�s�l�]��;l��z��u:���]���mq�^�꼛:���Az�ᚨ``�#�L?�lŀ�_��\�c]�/�Fc�}-.��͌�f���C!C
����?c�s�s0���(0T�O�H|�A��������}b#6�1�r#=����[�U�єk�զ���@#w�{��ѐD�k�hr��oXH��"SR��7'
8Lɔ6[��}�3+��l��>�������<i���¾�}.~�C'���	7(��#�o��3�n��7�a�y����%F�<C�O����;Xno�F����_ƛ|��<�}~ ��������o4�7�������ծً��"������&��&��A����Y&��4�:�����~,��.-����2�k��{�Hͽ�?���Nr��a�0����Rڗ�`����{��RO��j�S�y�����b����m�(���K�H�[8� N3�"�dq��sP�\c	�}Y��`c��9[)|�"��ɜX��A����%L:>�<�=棷:N\G��Ɨ�WY�w�+�폥����V;���6߄R�O�6�6��.�1b�n Y����6ؒ��UD�U �0����h��s>�?�]��/��7Z^���gqno^��>��"e�cl��G��~O�W��l�a���Gj���ut��<˩��2\��j#�t~A�����96��3-P}��I^�o3��{�å:�n�lLr�����s,* S�~�a'_�-]�ɰ'��a?�V�me({lix��K1P:�(D���@]|D�Q��2vlQ*��w, ���1u���n���x�PF�.Fy%�y��\��Ss^n��$��ɕnzٹy�T6���'Q�֊-�{|�S8~��Vo�Un�Un�֯�4i��ǟF�|�'���N��QM�آ���!�2�S�Z� �q�4��I,T��DH�mzbKA�0��k�I��zz$�q�Ea���,���K�_��7Py�Dv֚�5t��>��&��	t������;>ZM��	�Ƨ�B�0�CU_N��~H+{��AFE��5r0�D�x�1�����K�鎢��wQ0�i���{����j�H)ïĄ��ަ��<�A�gt�� ��ku��֍�=��ڶ�	��/���N����ߖ�p7�p?�p�0�����K�M�H�68����61X��y !a�QXw!7�q٬oz�C,H߳��s'���'�� �P0`btt4�MYIYY3W��r��A�z���$�~�*4y5'��1ua�	�90��Pcp��yʧD��_(T%��.+f��ZDM��� ��E�$���������+89֢Q��ۚ㫡�@��֟&�~}Wf�P ���fXM��(�����N�\I�$t�4������e2u�S5�+%Ԓ��B*r!��e{����"�e��)oN ��t�-l����گ��Zͧ`?�-�����J��������h`�/���N��K,�i��|��ִ�v= +pL���}�OQm��%A�q�ӏ�<ab&�Su�?u�bKLU~;��т��J�y'R9tEwiMw�����(���A�������]6J�u�QJ�<�WN�9��י_o;%�:m%��^*�H�w���ݗ`1���X�V�Y��>��^�,kd��]{i�n�\Յ�ڊ����ߋІ���=��1mgkG������)��G��3Ij�������'�R��S�)D��
j�	��c5Y̺�kV͊������i���#{��(Y:&p�2���/�
Ƙk2J��fm)h	���Z���f�M��3�H�46���'g#�3-�RU*#;�t�ӱ#���雿5�k�L�$���є�rҀO�Z����d�1��^�i��H8�ƌl	�y00�|\�������x�|]{�y���%�=NӪ@5�(ɯ���z�Ui��]-B\�UFϧ�|ù�;CY�o�y�����dR?�?sxELݿ:@��ɕ�}[{�{������Y3+�^��ւ��܂R���r7�ΪAI�R�?r��(Ҿ�VJ-~b��6\'/l��me�i}�5��%�Uqs{�?�~!�ˣ[ϣ��۵|�Tx1x��3��΋���/N��i��U�܉�R�nv���4R�f�v��c�VGd�I�ϗ؞��AP���{4B�k��<[�)�$?���e\;�q����J�^T��{� �W�y�7���,�+��c��BL&^Rw#ζj��j8���)��ס�n�M�/�RYw,�>V����| X�Gp ��!� ��!�bq�f$B2���,Ӕ�������'ǆ-.>�Z�;}zK������&��lC�jdj����8:�P\m�l)�r�8h%,Ύ����߉<gq���i���K�E��1�/9���Bڕ/��C.*I�p��#��O(  ����s	��J�V�M��K�cc�w�^��M�ȥ�����������_�� {Sj�������%�0|G���AFx�_��䟎���5Q6�{����:~�-gS�FO���ze&��������������*�����?ݧ�{u(�ۗ8��G�S��Oɹ���R�r�ZT�j
cƄb�ښ�A�ɍMtK����%��;���5��OAz ���RD)���I�*a�m���!7��d�}��5�H�?9�T0D�%�6\���@C�.�3���	cx�Y�k��hjd��U�>�T"2�(�_��d .�N,{VI�R��1q�J�zW~7���}�vSdm�0.��G�|�e���EB�<!gD4!~y's-n�Կ�H�@� M��/;�J^��&�o)��W�Ms�0���W~�K�ɥ��L�"�{����!�~Z>�DC���3�;C��}�/�#��􏌏N�S��t��2R~�Y�k$���z�h���k��A��ge��k�~q��۩�@�P����d2�E�뵧tP�`OX��9+e�������ށ���0٧^�P��.�Æ��GL�Z��V�o�d<ά�.����F�����wO��ςn�گ_=^��<ܚ�l$/�l�=��έݗ�Q��W~Xr?�\j��Zn�==���|�6��Xﾾdp�njh�/���J7�Te���C��9��[g۟Շ�4�� H��y�K�~z�������*��5Y�l��Ӭ$��NB����S��MBX��h"�U6.v
Q���}�P�l��5a�W��+��������e�Îs�헼�����n�f��E:F�����2?
�4:ʨ�hE�%�ϊ�a�#�-��y�]&x/��$4.��)]K;�9r��G�y�R2Z����}����LmM۞�Q��S��C�4eK.�)�V�_�(qeHLI��7�쓿�Z2Է))�����7�*<);�3���
e;�}#�&4�N�qL�?6!1IT=�2_#��u�R�
E%�r6"	X#�,�82��E�&�h��~�����BV�oي�Q�T���6�t��r7Y��>�!�o�ΰ�펟��yXA�&Om���(��1���9��iX6���Eu0��� �ᑑ�HIIQ1�t�����b�e�a�?��iq���h��L7ɢ:4�$#֕*D!rPv����X���ڹ��OC���7ĩ�쉉'8�T�x*�4l��\AY[뽆�J#���e�뢐�{r�ARq�Ys�ފ��	�훡����X�\M�� �+� ���D�~�O��"�;��-����;?+<ZG�����b���v%yLw!R�!Y����1�3��X4�kN��D�b����ి=V�RA����`?%##;���X6
ΊYi�X9$�R�i�c>�c����{���%PVW�\�I�ITD�2�iJ��l�����5��@G"1F!�8:K��E[qt�����(<�NvE��.Ll���b��Ҥ^�|V�\N��\*��~��Q#���i�s��XG��Kme��g���Y�D+\LO�/7i�g�dW<?Զ�,�9� �@L�j-2�����Ya�r�7x�' ����j\�C�v�H�{I�r��r�5XG�̣����*@�S���)�khj��� 0�*�t����*[ �5���D`�[��x�U��2��<^�k�'�d^�ʥךUj�RkP�Z��o����TOB�71ϗT�K.qz�	._qBr�7�ƓV�L��x����Fkj�%�Ε�;��@fUOvM_Ji{Z�s�����C w����&OV�7�ޛU�M�JH)�K,tys��$�ΥP�2�T�	�r�L+W�$b>�B��&D��h
K�0���&se4���Wxr�X)p9�	.�' r;xv�j�rsV�<���/~��W�Μ9���[��b����J��;83yj�Rameٮ�̲��=5i�Y�x�@+樸"�XaSj�z�ݢ0"��"�F$W�dr�͠�8T��#�F[X��Sh�9�����8A] MM��M�n�����6eSSX�b� l���E�u�2Q��,�.����͋��,�l�b�'��J�$3vޘ�6�$)#
⸒:!��K	�"ܘ 5΋��DM���������K"�垖���~a|f�����}���W�@+�T!�D��L*�T��T������������5�fj�� �i`��s*	��F@M�>��D�|KS��'BS�����aq�����<iE"���,��T�{!�/�'=��xϤB�S��+���J�}����57�R�&^sէ;��8�M{ģ	��������Y�+����M���4/�N_�"��bRŀ�)���Y�ףi:�P�ۙ`�rUP�Қ�f`C9a�f�&<9`j`d�Fʌ/����LM��`0�;��~5�006g#G �PӀy�f6b������x��U���������i-ahj����f�=%J�5G�G���̵g�Y35������(������	 ������g��-t^Zl_����15�f/�"��515����Y�)[�*A�����R����ã���OYlm���Q�{6f<AMs�#���}��9r��r�:)F�
���-�&��u���YX l�=SM6�@Blj�4��ʁ"E�|�\eM �	v����W�eįi�J���d��	�� �H�蚩�q.ֺ��8�W9OW�/T���\+���<��L���U��n��Qܚ�y�A ����UwS#�"^pW8�%���J���Y�7{z-�45�[��d�]��.���' ����y��	8�i��@��	����S
�c�Wݻa�� O��G,�c6����G{ȧ����b�1㖔q]B�\�0����B�y�4�p��;�����	���q��;i�tIN��N{�536�E0�g�*��2��UNا  �j��]jB��ШA���t�?aLM��\�� 
�TH��Y���,Յ�-�+�w��M���>9t�L�s��Wn��q������7ܸ�vy��ĉ��G;�.������~���_��_}���������o^k�x�����竮\���A���5��=����v��7�
W����_:Y�z�����[+�7��V��;Vp|6w��l�/g�>[~���T��J�N&�J9\%|��R�JjRKuJ�^.����p|�;��[�c��`B�Hrl(�VE߆	ݎ��0�v�wnŐI�Z�쓏����_�������o�����U7
�*��}{lX.6�I݉فG��͑Q(�p4"dG�m�C��ٶu�;��x15�~M�}kT�T�NT�,l�S�ɰI�m�'bj^�~ij��B0~���-�a9a�k����*Uq#�	�M��]����Z[O5��t���Q�j-��ʶ�$���9.u�AnV���Db�	,���ұ4��`�d���#��t�u`q��Xoj`X���Phd��/���8<
�FP(<*��D�$ĆR�a,R4��ʹD�������4�2˭δJ
��DCE�)c�(�IW����)4�-6#YZK�meq�rm�Ɉ��Ez1Y����1d\&�R	�����X66��St�D�R���_�T��?���s0���p(
L˱X,���j�¤�[F��T��H�%:�6�D�a0i$2P���F#�.`z��A��M͟4�& ka5��5��P0����Լt4,X���ǫNB��iLS6���MM��c�,<���	����BMxDTXxdxdDLL�aP�,&U.��;��j12���f����d����:11Mͱc�Ν;���[TT��z�N��h���EÛn.����B�C�/~E���Mʆ�°NMl�2&B@C���L���)��W%p��s��4H�4��)�iVӜ!nɒLMG���-7!T��zj���-����FW_��`����؜���PV�H*���rHu��6UW����tCc�iw�uO�����dMe��*I�SG{�-��<�\p�qW�Д��	c�����_�<P��(st�;�+���Jk�c�`�� F�l�hd`�S0P��� ���LeMo)R�&�i���>�/$ܚ%ݗ)���P�&A4M��!IX�T�	J]��8y�Y���B�\��Tb�F�S�MZ�ըu[�^�=��J���t�g'�'��  ��IDAT��%���d֤�ԧ�4$e"�ƔP��/Ը�Fo�;�.�hoVe{ZikJq�/w\;cK��&Wؓ*�+R�=��ޔroj�7����M�f[��֪�ke�X(q�r�j�\)�hT:K�b�C�|ڠ01X��!rL�V�h�.p�'�U'T��7�����k��4$4U;jJ-e���=����������w��Kϟ�ym����ٙ�������~����g���]_^�|��wY[SFm��8ˑ�hLs+=&�CkIJ0ĹL	`'3�j�X)��94*�G��X8�a���|��ɭ� ��4y���N�Դ�����/��w4�W��L�s�" ���Ƌ���9��8]l�)4��
���l�L�b�+>��ϸ����=���ʉ�qqJA;,%��#�aF�=b�1È<>�C�H�w4�g&�GѧN��/L��?�Ⱦ���\#��Z���S	�31�s!�i>�?�0?dѡ�A�ѰM����������i>�����|�����5S��@u��<l�}�_����a=��?��_HEϥ�g���L!<U"<��PjD��U��h�w�;V���z�f9AuƣX�H�D#A�����u%�#k6cӀ�p~��3Y��u�ҙ�����Ж,@e�����'(k����&�f��`XM��@Y��P���`��s�6����F�T��
Z�	vn
<�h�7����f�R���Lԛ_S�2��:��W7�cj�[�e�	���P6G:36550�&PQ�����Z867M4,'_6��n�&X� ���n�9r��ss�KG:����,�[�oY�ۻ4�{i���15W�a���"5/����L����KY	�c����hj )��Iz����m�ZM@� �� V0���^�?�삙u3��S���NV����x�`S �	�5�{�fd��,����ٔu�A�J�:�H6o�u�ھP�<�r�t��t](w]*v\η_ɲ\M3]K6��y�O�O���>�c��׎(�x�#���IsU.Z᱗�%
e�@\���I�p�q�������Fd́��}��%i�9�}�~�����#:�k��Ygj������:_�A}¤ ��_�<1���+aޑ�q[Ƽ)c_��/K����zFB;-���r/�E+nŊG��U_�/&j.&����x���2{�Nq?�5���=*��4��u|�W�&�1�W��2P�$*H
D� 	PZVQ�&�k.��5֖����=:xhq�����\�r����o�^������ׯ�|e便�g�u����������?�?��W_�ߟ�~��׉�?�u�l���U�K�/,�V޽Sy�fك��n��]+����r.��霥�y+��W/�A�����N�-�-_9�jo)�I��5�$�4��'T	%Z�X/e�R�5b�Z.�J�Q��1��Q D�DScB���$T5,�Iݹ��c;�����������?��O���~�뿿��YFN)�)��&��5z�TD814����7���؝a�a���h 2�3b��;�پ����}�o����C�n�ܾ�I�� F��c<Z~�S�m�Yyن��;����)E��e+���	P�U�����45#��Cu��j{w�����^��ݕe��
��L�ҥ�%	��!8<Ga��L<F�4������F&1 2�JaҨ,:���!���-G$a�4RN�!b�x
�����EE�b�B�1!dT(�%�cU�E�q��(�,-pi�}�2��0NZ���hC��1G�;߸������R�l-u�γW��s��>�H/��hhjp�蘨�����H0�EG�?w��ЉD&}�L	���E�P�i<���r���N`�s�9�Ŗ�%z��b0��_bfjZFJjNFfb�Ǭ7�Db�I%�p(4Rj%:&�_�,���ERT�eUZd			A��(�f]����Y'h@G�i`��oS��x�����4��OI"hj�S����Te}���l�ħX�tX�nVxDThxg"�{H$�8����ku`wJ�?�r�H��r�l6�J�Q"�������9rd|||fffnnnrr����555���&�	\��e� 
��ঀ{�������~c��`'���a��؈$t8���	S+
���*��~Y���N��&�E��)e��0�SӒ%�����)�ԝEڀ�A�j*M��j�1�wzj������,MY��0^��F�u	s]�|�,�%��qa��أ*���(A	6` ��'�*����6@C��>�R�e��4�d!��`�v����􍙦=���ǁbgW���ܵ?��Qd�.3�TX���P�e��6V��4V��k,��p�<���4_����D�tj ��G��4-�����-�K�uC���+�IV��%Na�S���[D-���r���#��\��ϑ�x�Ƞ��2�Bf��,R	�Df�+\JU�J�)�2�H�*�"e�\�S�R�L��(1�:��9#�))�&>���orf�mzK�ْj��9�i.g�˙�v��)N{�I�P+�r�B&�J	O�It
�R 1YL2|b��K$�X�Tΐ�DV�9+/��1k�����������±�♱�ũ��������ޜ����+�����~�_��أ��>����~�t�Ν�C��&�����K}0t���g^�����ɫGW�/��p���������M��e��|{Z���P�lz�Co1H�|	�*eb�\��������6n�[P����� ������_�p�$
�RE��tfH{r�y��\妬ˁ-�A��9��饩	 �`�	��-4���fs��Y��4�W<��[X�M�)#sJK?��L�I��D���:%$���CԨ!R�89l��Ȍ:/ĮJ	���ާN�n���;�?6)~�S��Z��R���31�37�i`@͇t$��}暩��������~S���!�#"M����y��?��M�}bj�b�wИ�,�K_�B�b>�r^�HD�I�ϥ�����T�T�c@��J�@%�S��k%����6�-��J��b��G>� ����^ʚWE���5���=��5�u�& �\�����y�hZ��`A�5�^��כ(k	Pпn�ӂ���T�M�S�� �Qp	�0p-�	�x���}���	\�x�4��jf=#UF�i��	$@�*�f����&�h^aj�Zto*k6�����MM�\{�������鮲���c��O-:��ln����2S�ͷ��љ`Y��_������C����n���~ɯi���v-�5��ֽ&��_K�V^�5���R�|U��ռV�|-v& ؄{Nt�Gӑp�=~�@��Y'k ��5��@�7�o��S,k��w��PM�p� ���<�4EH��	���u�+E��MUXf���Վ�jǱJ��r��r���R�m%�r9�t=�x3�p�k|�!�&�x��|�ߏ��s�`@͊��Ġ]$��&��*
5�*�xC |=�i#<�)Ss�VEx#��>����֓�=j�iL�i^%k<���J��5���/!?a��	��y��=2��y a�I�x��ߕso���e�+R抌��`^P1�ڥ7┷u7Sגu+��K>����[���M[E�F٫�u(�TH(��MM�W��U�����2�TI*VQ������g�ey>KINbMeAs۞��3S�'O��:�y����-�n4_��|���7�._i�z�����V�_���w����_��_�՗_���GT?Rq�L�����d/-�_�Zp�J�ˀ�[+��/e]9�~�T�c��Ng-�ɼp*��b��T��t��EO��������Tj���8���es4`z,���1*�F�Ƞ�r�P�EQ�v�"Bpᡸ�(
ň������Q������(�!R�������>��~��_~���_��8��C�E���u;*$�3��]ԛo���N�[[#���-4z{X̎И�!�;vF������o}�{o��g��ͷv��5l�6:�&�8�(�3�D4���4г����P��|'��-p����Z�����($���5T�Bʂ6��}5��*[G������gS��ҫ�w��-J�B���2��cq�԰���2�� f�<������It�BP�k�rh40�%S�2O"�	�@D�`:��cI$���`q�Xll.6
N�3^>�GCK8D���ӓ�\���c,����ynq�WZ�*�f�ru�������=���l[^��c�D$�$DCS��������FEE�cci8�Bd�|>����_���d2X�$0'�����[5ө4!����M:}�˝��������]���`�Q��
E�`
�4��i�K�W�hjv������	���& k�	� �05�oSP�5S�M�[t�Qwu�2�%O4
�r��G�S1DT**�$S6)d��˒I���h4��ۨ�{��p�l6�k`���������333���`=::���^]]���N���f��j��L&�TJ�P�����7��_�&�Ԁ�� w���V�=&|;ƣ�h�x#��+q�J������~�Gq�{?5���+
`XMW�.��Sa�VZ�$�ZwO�����Rhn��W��
�%Yv~���b�'�x>/�,L6��L" �Z��vy�S��V�\*�Ή���k�=��.7l* �ny�K�tJ��ʼU�G]��%ꊓ�%ɆR�OW��W&k�L���9ֽ��}�֦t��,m[�����}�Ț�{R-x�	�	���MMM@��� �k@ �5K��iR����$�L�%�j=��8~��_��Y��2���S�
�Ka�)l�G'�$��gQ,��NR�|2�G�s	8�!�T�@&���"&P4��/֋d&�Ԩ�8L��x_�+!��Lћ=*�K��K�V��"�b�Rj�)lz�ՏY�0HyR>�˦2�t&���3�R>|ܨ$���;m�D;�+1��ڔ���ʬ��:���Z�--��Ό�����쩑�ũ���%��E�#�c��wo���/��������s�������������ϟ��Á�WzW�O���ݛ�~���{�Fo_=t�B�Ջ�7WFo_�����X��侱���]�sk�
j*�K��Z�@��hYh����g��8�6v��W����q��4&� ����$a���45�}y��������e ��3�`S�jf���������J��i��53G��q-uBE9� O�HSⴘpX���s�c��r�)t�y�{����b�ײ��y�E?p��~a�a�̤��N�#��G
	���s��3�c.��i5H&�=��C6�_�w"�O��4������<'�[L�f�� �������
��K�=�˚���"�s� ��<W"��J�X�������u_+�o�߱*n�T�q����	�9�KY���Ԭ��i�q�$�F�%=A��e��k�}�|@`0��kM�?r�^C�?7j]Xt1p��iZ����JYSn��h ��ԀC0�&`j�&�	_F�@S_mS�� eX'h^���4T��Ѐ545�u����h@M��ȚW�ה_�@_�5�L�`Y��
S3ۑ90o�� `jN����?ttv �hXN�k	6���@�[������N�,��?1�rq�����Ks{��Y�Gd��l�kbjV��Wg*.�"c "kfaX͟���:���� }M �&`j6gk]��i8�IOk5	G۽��S���f�B���	���{�#kG�o�=QeyP�`<V����f�T3�2�&�h �,L0���M	�3FK�E�J�����-V;�T9�V�O��ϕ:.ږs,��������3���y��}�'���ɮ����	�;.�-��V�*\b3.R�K�e�*�p���%A�a�=���������ɀ�
����Ѽ��$�B�FM�1���L F�l�5��t��.�汀���5%,�#)����T#~�=P	�����kJΪ���b�r�oǫ�&��'�V<�Kq�sq�.�Q�|�&9l�8�:f��ޡA:v�Ӑ�jH�4�Fa�Ԩ��D��U��T����	�Αҥ�L�$?�Z��,�����>2x`z���ٖ��[�.�~�����7n�y����k7�W�4�>�|��䣧�����S�/�|��|��ر�����)�y;g�J��J����k+y�W�._�Z� ȸp6����3'3/�ͽx>�ܙ�Ǽ�����9O�����Ԏ��,�ͦ�ٵF�T ъdF��,�Xdb�BdR��*�V%���X,3,N�� ŢYX</��h�EDa��(N$�Kc���|��ǟ��o�|���?���~�t�Qim�%E8����HbT5:�Aپ�g�D~ok��[#o���ֈ�����Nțom��￳�{o}���z�ͭ۶�����b������I�zA������먛�~��[�dnjj��0jo��� �Sf�-����W�U[��,���r�Rˁ[[����٘a-O��X�)F�U�WX|����0X���#�����k���iG���HM���q�M������5�l��P pD�(d<�����A��""��N"�	8$ኌ�1�DLM�G3	�2�Gň�����g۔nmQ��0AV� .��}��4yM��6K[�m�]��]�˱��g�Y�R��X>�����Fbj�#cb#b0Q1�A���T��ԨT*0��j��L�1��0��}pA!�)"���
E�����]ZXT�_ �9�iI�n�C�R�<:��i����޿�/�J�,���;��G����>PYX'h�"���mcj�؛f?�ɚ$��&QZ���uʒ"����	1�����DbP�TDd4��AǢ�4�L�׫U��b����@�45�1�L0 GFFF���fff���:;;8p������������_�V�T*e0��P��8��?���k�#x*��O�!��!ĆrɱZ!^�ȱ���E�}+s�����"�Q���Le<�/ayI\@��R5-YRhj���DM�˩�
�@�ڋm{r���2��0N�e�y>7A�q)X6=N�w�y ����
b�I�h�'Y`c@�M�bW%Z��$�,�Y�H���T�2ͥJw��.u��T�`*�K=�
��«���*��j��>E�'Cݒ�i�ѵ ���*������2��Z���u��$�	:�`S��M���m�Z��S�/SMx3��B4�	��t�K�B� ]˲�"B�b�t��!�04*�M#p�D.�F�Qp��G3i$!�(��T��A�0irUF���h:�BĳX1�)aЄ�R��+dF�� i�|���* B��M�)"]*aIe��#��%2��>�ф�XR,�
>�	8x�y�T*�q�t$W���	Tj���*,4��'��[48�3����J��Jɝ����Lf�M,N
��LOO�߽�3���|�o������?Z����?�~���ُ>>�ӟM��|���?������w{n]︶�~u���R��K����=stp���œ���/�힛n�=�ZT[^X��iU<�Y >8�f^��Wa�V���������a5�\�no2PMMG��;K~(G՟�ؔW�A� ��bC �	l���8�����f:_7���H��%Iƽ��8���5l��h������?-&̈���Iv���`��(���iZ�q���tEFyj��
>��>w������`b�����Q�����R!�s��s!��C6�E�4����L$��{{�S����6�Z@�_Ӽ��[S��Ygj�SV5 ��N�!��A�f=�q��O�uj˅H(RH��V�P'}���i� �4�{z�]��Mqա��8�Q��g}�	�x�'<���fֱ��i�����;@m�#e}@450j#�	�(k^�k:^�YVp1e�k�p��GLM���	{��w35��"5 ����@A/� h�b�� 5&@��_S����f�_�f3S�4~l��	65PӼ>�f�15S�����N���녦�������K�^vz�����Y@ �f������ɕ�3cK'�����k;?�|i��4�{W��,4�>�fy�de���dj����@/8- <�L_R 
�x�f����^ MM *����N>х� �\C_,k`L42s�.ث��NO��`45�;�D�i�}�R���`�r�T5M����5��H�45��j�i�f��	�P�jS�%�2Z��	PH��*�b��X��D��l��b�u9˼�j���������{����>��DǃD�=��V��]{լ� �^�1��(IHU�8�m,�&�xK�@S���mM�m<	��|"P ���D�C����<"S���l��������Ɂ�&X�@;�����a]+���5���$=a�8�\�#>��HH(�?1J�����ya�?�˞j%�4���%�����d��׬���^ͪGy�-=k����Z�VɌE4i�8Z��tji�Zj��Ң%��"-�ײ�4�?UL45��S���'#e0�|L�K��h�Jr�ft�쟝ꜛ�<uf��sm�W�n�m�yo�ͻ���G�q���r�s{Ξ�w��/�������<��?�������Μ�[Z��u��ƭܫ�s�]ϸt!��r���K��+�r�.��=�~�dֹ3����;�}�Tڱ�ɋ��3i#i=�]Ҍ4�˥r8�z����X$2K%V�Ģ�������$R�
'�G�#c��x.�"����� �5D�MS��z����ٴ	闟|p��z����|��'�?���!׻�r��$ �����@�b�f��5�v���1o���#���on��[۷|럽���ww���� Ƅ�(o��ZN����� 儍�<�?��Jϵ�45���k� ՜!���e�����]b<Xj�.3t���K����mE��"��<gC��,^�mQ$�e9O)`�iD:M��I��'G�V�f���h"���0�@Ģ6C#�iD*��
"�N& P�42�JBCHD,K��Hi�H�"�\�2�@!`)D����QL �A�f������L��أ)K�yd�nn�WT�����T����YS�m�δ'�lR��̧��q�t$��G����� ����h4�D�2�`�%��\].��0isr0!�5��L��<�Ec�d���ө�޸��ܼ����⒲������̬$��j4)$R�M�҈/0ɇ�kLM�������݁�ט�WTfۘ���O_�(MMM�ďR��̲��\����x445���A�FFń�E�E��M���KLF��n��`P�T�	���9�Je���V�������Ʈ�������ឞ���֖���uttTWWdgg���x<�á�j���R.~E�,�ڀ����:�q�������n��F�吢4|\�����'�����	�*��ޓ��5MhL�m45��uW��oj�ݥ����u�:ڋ��9��ui�,��K3�q+�v)�  �Y5�
��iz�$�X|�J�P� ` �)�N����x�8�$�^�`Ws�K' G`��"(�(�0�3M2��oS:��NE�KZ'���\ts�f_��� ����Wv���t�U����[���H�`X�&�i�M�5SS���	k���xA��Wb�X�I
����C�1�4���Dbcñd4��a�pl�5��P�\����a����$b��b0H"������NdS�LGf3��R�R���B���qh6�ϡ�Y8���8B
OD�i|�#�2�(>2
A��$�DSP1l"^Ȥ+�b��d2Y<._!�Z��$�� G_���!��3i�'yt0{~��̉�g�ラ�G���-��/���/�V,��_^�����'_~������g���OV��������k�_�}�t��F>����g�n\t޿}�ѽ��'>}���?�{}���bˉ�Ǧ�ϟ�t���\��@mgka]yEmYJ�ӡ�t�<����+5q���j'��ūvs�������(�w4�@dͺ4(hjF�������/�N� �f$I<���y����>�!�i(#2;��L	p�|�$=NG�u�QbƩ1ӌأ\�y)���uW���%��)��!��]�#+�+�/L��?V�(��4�	����q��^���k���yN#�`ӿg�-7�"j�������p����Op�'�5Sx������k���� Յ	��I�iTX`���@�} �ݓ��+�@'}��=6ȑ�'���L���4(���Az�$�b����'�����$�X��5��IO��9�� ړ�d]��+M
s���@��	К"�����&���Ț���~YWp0_7�`S5l���/{E�|��C`6�[����5S�j �(t.Э@Y|m0���\cx�!��`�f�\�GM�DGk0��a5Pͼ*��p�{SY�.�f?-v �fӘ���ܩ��`Ss|���L?45а��������& k�����ՋG�+gǗO�/��:7�zazϥ�=+�-�k�fun}�D���`�p��t)45W�+��ofj��.�,M���350���`ꙁ�S�|'z}�{� 08ٗxn0#�,ȅ������e��I=ٝ|�;p�'�Lo��C`�W��G��='f�&^�n^�J�)�#���n9���9�̷x��$L7�gv��7{��K<ښtd��p�}��1����k�9Q�`�`)��7Oҝ-��J���� �&O�W"RV�`j��߄��5F�u�uא��2�|�j��e�3Ŷ���\�J��r���Ps�k���M�<�8x��{	��N�u���Ny��:ˤ�'S����D�-�6�vG�Ԭ�~�^��
�Ss�H�C �%R��d��!���B۔GT�FS�B3P����i �jxf0PӬ35RH�hDV���a5��4X�摀�X�|"b!H���e��%Ou���%熜yU�Z��W՜k�5�l�!�`��O���F��I8m�O�cZ���ѧ�u���Z��֪�4k�MZr���.H��������jbj*�~S� ��)U:f��U�a�KI�\T<+�$AW�hNq�o�)����N�]X�<~�����+Wܸ����=���{o��{�o�lZ^�u����C�^��O���7����}x`ui���ƥ���W��^/�r-�����w�/\̿|�����K��˗WV�Ν˻p1�칌�'S�&/I;r,���#G�G�����uƂ|sF���Uh�]%�DB�TdS�mJ�I��I9
)�u�g�"��RB��H�4����Q<[φ��$�X���N�����W~������|v�_^~��W���=dN*R�����L��B�k�2Td���FR%;1�wc��D�F�G��	�ykG��|��mo��c�����(tt:l;��d,"�G�N�2R5�<3�@�3Q��`L�&��zw�xO��� u _�^��(�u�;���E��B�B]k�q_�e_�cw��.�V�`ȴ(}z)x��"�F��04���Qp�_Ӭ�=}S��,&�F������l�:SC%��D��E�������`������	D*���F�jDp�ɠ�4"��c��T����`c���K��Ņ^SY�����p

麪LCy��,Uƕ��T}q�%٦4H|*���"�"0���aH�ZD��"�bbI�L�3�"�P,K��P(s~���0451�
�0}	���<[�P�������+JJˊ�a5.�!=�X0		�!��D0�G� �F^*&*::2
 �z�a!;v�n���+S�VlS~Y󺘚ʚ@X�5�VF��Y��b��Ά�:��nve<�*�W��� ���o��ͬ�g ��5���	h�j��D9�*I�f��)�&E��sH��~��OH��ذ�H�c�+0�թ���aCT�2#���-��x��h4pa�'�Ñ��VUU�����������ݽo߾={�ttt����߿���:333ɿ�\.� �D�'���5�р�,����tHDbj�1!lb���d?�:IE� y��uj��U> �.�ĭO�@S�
�͔@G�V�U��)3�UٺJ�]%��b[{����֔a(�*���	�C��I�z!C�"
)>�E� 8d�F��rS)`k%|�F��E\�G�g)�)�,�R�<�R@W��Z	|��e\��gT�MJ ��~pT%�L����q��M4E��2��(NU�Q֤h�Ҵ����Y��|Ӂ"kK�/�,�"��
so��`��`��P�я��\?Pa�i@MG�
������`ܒ!F���5>N�����15�� ABVScX�!Ԩpz��A��Fo��G��$
���1Y6��ax !M§��$�*��%B�L�����#�б&��t,M�W$:|k��貨�*�Z�s�\����9x&��b2WB�I�!�-�29
�!G�Rcci4�ᐈb6�cQ�b1�b�L�Q:�o�&#�US������ln�g;���������#����c�����ɉܩ���G��?|�o���������g~�����?y����]W�w?~6���mw�V]8�����;��\�Ұ�T�r���rӕ����u�O6�8Ҳ8�q�H��cmӓ-�C�������ʳ�=�NC�[[�R��EN�CT��U�eM���w� ��=��}I���k=z��`��/[y���y�P�v�@�G05kQ3/M`�_B�p�a�H?Q�/���NSL&JF�.=jf��C*ʸ�6*!��<�a~���d"�4#��qb�%�u^@��`>�^��_�_8e���]�;��6���_�D?�����P�d<!�i���`�2H�`?Ϩ$X?j��T�s�)�MP��=�#��)��H<&������|�i��j��X�M��@�K��g0�X��|�}!ﾈ�@&z��>�ȟ���
���\�H&�/�`X�]��Ar�,�b�/�)/zTg|�>�\�i���LD�N�*�#y��$ށD.`�����['h�K�
Й�U�'(k#�
S��*��&Ve�:;�	$@A;ǁ�?jj����@�X��kM�i#���C%��b]o� `ԀK�+���XCS^pS�5t4�o�K5���
=�4���L�z����wz����LM����=�u�:��䅎�bg*45����A�{��:
&:K��95�{|���t�酉�G�����񹯙����>�z����Cu�'����ZY؇��ݫs� +�kuj�gkV�jW�W� �+W�VgK�̗_]���Pvy�du���|��rhj�( \������x6��X���L����sCi~ϒ c���H��H���,�š���������u��O%�IBN��zj(��`�����g����?ݟ{�7�dO��CKc�#�'�2��O=ӓ�2R~y���|3��|��٦����e�>�3�?e�a�3������
�3{��z�+�g:R'Z}���Sm��u��*�`��G뜓M�A��
#���}I���p����2]_��/_ޓ+�͓H��� ���p�q(E��B�`�a V^K��7}�Rp-�ـ�/G@���/h�C���<�h�z,_~'�/'��2`��0Wb8Zd>Qh>�o��k[ʶ^�r\� �@w��_O�\�nx-�R]ϲ�O����ϼO��m��Z�e�hE�_�p�h�2m�L�F�_�S��(W��+$�e"�J�ׯ�s	��,a��8 �_��b��k8�u<��r�Hܥ2�Q6@��"�o�����G4��v�L}D��#��`	��'T�{L�3:�1���J{N�ޣ3�y�`n�}:3�f�U`�S X]�F<~�#:��&i��c>����ϥ��d����:�{Z�3%�P�ԯ�-eߐ����7���6��EvJ˛U���)gR�S�F�auXNT�5�>�]MkQӚԔ:5�ZK��R��F�`�W�QD��?PjT�%�ZA T*�rB�\E�T�+��r5�HA��E�L=�,ٚ�5g���9tdv����˫�������ݺ���~׳G�o���ƍ�sw--�<�?���/>��ѧ�=�����7���T]�\u�f���Wn�\���r%w�j��k���^�[�����si9�ԩ�3g�Μ�8u2��������������ܮom�-/ۘ��9�25�B3�B�*�<��0�xf0�P�	x���+UL�/�`5>fB�$�SS>,/��J��5�]֢������ܶÇ�>\��o��?�������~�lJC�>��j̈��a�>�#_�T�M���
Pb��(�V��(��w�b��E��ڹ3t��w���f��wQ�HWp!B�'�k8`�i�d��`��k$�Ifb��Th�:�.F��Qꤗ�h��Eu��j���LMG��3_�^��(ԵiYSb8Pjꨰ�+��ʷ�fXʒ�yq��ܭ��b�C'I����t2�)"��' ��O~�s��^�f4:�A�X4�$�f�p��e�L r�>��Ǘ��X[��L"P)��iS$�I�cpQ�dT$����(F	ǩz��D�,7�X�j.˲V�X+2ͥ麒4mI��(ŕh՚�|��#�)�LD*4����DŠ�c01��\&K$�)�B�P*�`���`~���a(����###��V �t:0�/---///,,,)))**JOO����E"�X(��`"Ƥ34�Z�����Ш���Ȩ�00�����ckT�vBt��ᑝ2�O�HQQSU�t)]E�CJE� k5!U�K��AX'h�'֩1!�退�˚bkM�8Xe�5���8�2�����l����K��bj<��$Iu��!]U����IkSU���Y�C���L"��C�S1dL**<::r����F�;CC�S'�I�V��f�ۭ0�	��\.����Ba2�`�F���=�L��������{�����޽������spp&F�u{{{NNxMXi�V�:��� x��+�M�����թ	�~"����H%�TP��|�[P�o�PW�315�T��">��$^}��)C�;K�V�m-���W��@���_��P���)��Y�l+�7f����L�$�$��	-
�J@��|�G#�h� `R�,*	���9t
@�e	�0 ���L�d&M�a�Xt.���2|�P��x1_*��\�	 ��Qpr�.`PT��J��hF	ϭ�%Z5�$7*'^[��/J֗������٦�<s}�����U�(6��]�����9��BM�q��#f����BաRc_��`��3Oӑ���5ChI�4��v'	�|�F/��˪�0����'��íK�x�%Na������ -���h9EAQ"��X
C9R�@�˘b	](�	�d.��k$(�"��|�@H	HB��!p�b}�#9���;�J�F����B:�G���L.�*$0$T��)P�EJ�P����l&��ƓYx2O�c�%�D�"�s����2x�X)UXu��:��(������X�;�m���E��1��h��X���ٹ�������#GK�-;y�������_�|���ܿ3����W/�֭�֮�4\�����=7o�`���ͷ��ZÕ˵+�U�.V\8_{�ܮ#'���;��{bz�����������C�%yY�y)��d{�KS`��8d�VA�[T��W;x5.���m����$J���mIҎiW��`��'Sї����_�P�0����A�3��bj���w�<�d��3yډ�H�l8Q4/�v�;�Vބ�=�cN��J���2& s0C��a:z��!�#'��G�1���1�����C�+��o�-�p)��!��M�+��f�ό���?�q~��L.��T��"�x�@�'���MΤ>cP���Oh��T���9�k<%��y��k0��9�GD�?�	�{x�m�p���`a��`M����p�HF4��G_���<�r����I%��e(��=�k�DJ�Q	���M�V�5��S�쐝�KN8Ňㅣ^�W8�(<�$�U�S��)|��T~[
oЖȁ�f����`ek�~
��c��j�Nx9������8�~:��N��U�t�7���]��*Tw�4��bmo����௷�	]�ʮ"yw�p�D�S���W�Uh}��25 �_�Yw�%��Xl#��F�	#��F�~�J�)õ�H� �=A`����XQʚ�����q3�	�{=����>$�	I}:��oO��H��L��JE�L��Ț������ٮ�鮜Ɏ�������޺��֓ӽg�G�,��Y�<{d������m�g��7���b4�N(bj>zv15��+�{OL�^]�wea���݀չFhjY󕩩AL�B5३)��P���,Ondu��U���HF��hj���8�	�0�	�	\r|�w����D?��S'�2Oe��=3\pf���@љ��Ӈ��w9ۓN����;�W�:Rsm�iu��ܡ�}Ug���,9�Qp�@�����S��&۲'Z����9`=�7uhw``�gp�w�%y�5u�-e�=}�3g�1y�1u�)m�	�`3	0T�0X��v�W��X�mC��C��|yo��/_ڟ/(�����E�����K��0�oʵ�FK���QP�|SX�E�3���� �����d�0SbX(2�(4��7_̵�d�.gخg�o�9o�د�l7��2��$?O�>��?�w?q;�m����
�U��
_���.Q�K�
�q�̼Bb�k�J� VH�e"	�D .`q��8<�� w����Wt4P��"� w��M�M��!S�Q���G4�C*��~����< �������4�s���~��
4�9� �M S��� �B��z@�=d���O��'�3��X�\�_+xO�~��>W��Srޓ���8O��'
�=���}Y�^R�/�y'�y}V�:�eN��
ڄ�U�G��5�[�lS�v�h*j��Z��5(I��k��W��z�N�����#��/k�J��TiSS���	Y"B���e�%ŹɎ��#��N,��?sh�����Ϋ���vܻ���v۽k�n]=p������ˈ��{��'S���2����|p����>~P}�F�ʕ�+�j�<�]������|%��J��K���&�<�w�R΅�g��;�{�d�8�9;�{�7s�{V�5�ct�U0���Dt��i�s�J�� �
�E-�s��2A���3m�Ɗ._ש��k��Ӧ��	�e�)�S2t�����G���>�ީ�����x���y��C��N^��X-8��}�Pt� ��Hb�,c�*���)'�RI�D�:�ӆ��XZ��	��n趷cB��"wP�aBj�QL��t3/�oj�L�<1�D(0�-�B+��N-r�J�r�:S�t��,�i��3_05�ڎb�bj��JlMy��LKI�)ǭM2)\Z�V*ry4��őp�158 �ůUSY����c0�%~��zS��!����`��MX%I8�ϊ�&�@��D�1LUB�I)r��VUZ�>;�T�n+Ͳ�fZ��Ei��4K^��c�i���I���(thH����lD$&
)R��E�,��O���Ol$���o����l\��<,,� f��B�ә��_ZZ
օ��`���b��`�y�.���0�,�AY�?¡И���Ȩ�������H�#@��m�!�pѡR��Kr�^%=YI��&CI ���w15���Sh��,�b+�0.�� �v6���)w� .v������&�_� � �f�>`��x�~S#�J�ԧk��ԕ���TMm��ģ�qȽZ�YHU�	�Ԡ�#b�cBB���t�'�	��m�8��ݱ��0�L��24�����"
,.�+++������n���mmm]]]���� �EEE			�e�f�D"�	�XCS���uj��h%lj�Ǫ�G4��@4�FS�Z�	���B-45]�־JWo�����^�j)�צ
��vi��oW�u��K�3)�t_� ?� �1�4 l��!���(�M�1��z�<����l���5��[���F�Qi|:U�b�I�BhՈ�L2�]��Re$h�=�\��(�X�a��0�ʳ��Z��{s�{r�����kk�(�*5WZF��#���b-�ru���Sd�.�!S���2��}�ҽ���;��#]�E5{<�eIs&bt7b#�	F0�$R�2�$��9�"�s�9�d9�=��lO�3�}�:�����ΫFQ0L�k��:��o�* �n]?~�W��|��\qG��#�l��gg�-~��lˑ�f+j=�R��+Cu[�J��gS2ИTnt*�B8�d�0�r(�'�q�6)f`+� �;(Q�W+�����r2��D&�1ߙ���X�n��,7j�*Z �`�!#M�����ѨP�AD\T�EI6_�������I�"1�D�b��Tm3�3]��lsE���Ѿp��oйb�uͰe������7o+پ�|���]{�v�ݷ������ё_|����7��d��K�]\������Ϟi;sf����g�λxq����/]
w:.\ �N�j>~���іCG�w�?��c뮹��Y��c�ꅃ�K�55�U�U�{��]>C�[]�Q�8����fL#kڽ�y!Sә� ��*��U��E��ڕ%�5e��18�*�+��U& ����S������m���:&�D�>(ߐ%�HG��a�h�Ln��[���E��"�os7��MD�&��cmF3��X�I�h�5��"��o�c��y�����9���d_YD�1Q�6	�0`_��/��/���2�b�GB�R�gҝ��
?���0�35�$R�|���ŝ�������0���b����\�+iL-a@�HM�^�t�6\u�K�[(޼��I�#�䩔~�V�+W>S*���Ǫ�ջ�i���n�d7���f�5��S}ե��R�w*�����P6�9[�!G�&W�2W2
�	k���|agՕKuM�i �(k��i²��eMo����uM�d���M�W�ہZƭ�h`�'�(k�5aY5�$��Y����I/}��	�^�� &�5�f� �����LM�3.�fdQ 225�HS��7o�/dY025��Jw�BSS��Ԕ�W�WoYV�u�yd�ܽ{o_slצ����d��ݳ=2"���bj�{t���}�V�>�w��m��\|~�B(kΎv�dͤ�����3/L؞�;����h=�s4߱mRSsl=�]35ca5RZ�q�&�Ԭ�ٳ&�au6`�ܽ�����Pvt]y(����9��p|]͑��6֞��x|}��U����޺�tͬ�Mٽu��U�%��JKW���־va��Eek���_�ߞ����l�t6��48��K����Y��[R�iII_��! �jUK.���y{���e�卾�Z��
��
co�5�(�����խ�Ӯ�S��U���WTI+����*��*��j��jͺ*úJ�r��
����4��
��L��rEX����q�&,k��$T��#u����}��HSs��y��s5辒�^�S���iA��̻�M���tY�=�P��H#M�Y��B��	�p�s|hj"eM��@M�ϲ���LMX�\�a�q��;�h�w��0=�.*x �	��Ǆ�%~*  �t�+'t�@S3���ܣ�{b�T�P&~(=�P��� �HM�E�g&���"M�������C��Q��A�i�m��*|�߬����AѥAj^�ҡ~S��ݫLM�m�a��T�9%rN�NP�P�[嵅�-�>qp��C[O[}�Ț���_������{������K��]��w�B��3����ˏ����/?���_l���}�u\�:��yWn;tc�ͻͷ�κ}���ݖ���]��|���Ŧ���ϝ.?~Pu�h���[�+r�,�i�婩t��y~�ߦ��5�Z���M#vj$5�SC�uJ�E/QH1�\�YPڹn��+�>m��t�A��wg�t��/��~�}������v�vݩ�cO���v���Cw~�������\Y�����w��<Z~���>^v��Z}�ӱ){�p��-�֕Ά^k�|���#�q%:.)c��䔴�����(0��Ċ��!ǩ&�b���r+���y�� }c����FH�Lfj�:5!S�h��@Mc�n���x�4��V9[�����R�.ע��z������pAl���i"�ߎk!Q󝩁b4hd&k`�'h?�Ԁ���1h�\����IK�R	�CS�^!�B�E��T���\su��	kM�Ԕ^�N'�h�OrX�����Ĩ願�xP���~k�)�)'LӴB� StP~Ǆ��e^n1113f� �t�ש�銋�JKK���JJJrrr��_�р�T*��T&�He"13+�~��?x��3���Nz�L����8N9��F�Լ�Ԅe�65��������5MX�0�����\9��P65�%��lU�[0�245����ĸ����ؘ蘸�3�[�a��j���.����/*�
;���G [�$���l6���M&7`��tfff���TYYYSS������������������w8����<!8P��t�9	�apܡ��cV슎�9�E�S�N��Ӣ�a�W��5CM25p�'hjB|��˳r��AIG=�D65`MM_����6���or1��k\+�-�
�2h�y��MEj%����f  �#�����IJ( ��@S#���AocX�H$���q�_�*� !D�Q�<��p2$W)D-*�C'��h&�͡�U%�ڪ}m��9�o+2�.2��W�U�u����T�Wi�5�n��k��RgZU�d֘��`��S�	�]��*QE��PXcjf��f�$�e˚t�KRb�h�H��tI:�Hf�cS9ѩ��$�����\�&DlA�Hg���� s)��'r�TD���Y�kiD)�+Dl��%2������'/Ǒ�3���A�VQ2�@$E)Q.e
�H�IոL�I�Pʁb
��q!!2��t����H�� �#R�De�nCA�����P�\�ķb�w��c�yÈi���m;��(ݵ�b���}����;t��𑢡��W.�?w��ڕ����^���֍��G�|�Lөӭgϵ]�8��e �_���Νo9s�[�Dݱ�͇�����6��u�p��M-+V�Z����=�kqCsMyqvE��6�Y��CSS�xmS��D3!a_���!k��f͆*=�~��5�jL#���*#t4��՛��u9�u>��h�&�j!�p&�I��(�n�q6K�[��B�6�5D���mx�v,u'/��8���|j���~�c�s��y����m��ߚ��2_��_��5���s��S���B�#�xO�AS�D����8�]@�s��zș��&�$�f������@��k8�ˬP!��?G#���u8��R	e�c���T�D!�45���z�m�����f�_�*����f8��0KA�*���7�2�W���CŃ���aLM����9$�ucj�i��MM���.�#-�d|�lJ�PӼlj`<պ���T�-�Y���0w��fY�Ve���A;X�{MS3iL�d�X15kg/��W���e�k�¦�ՌU��@S��;Y���D�P34P9��v�@�����5��nYvtt݉=[N�>�s��P�S�Ԁ�a��2�aj>xr���}�[N�<<��ܮ�v-z!k�d��T�?���3La�(kNU�̙m�f?��jƙ�ck��9���Ԇ������H�C��=�:g���}+s �W�X<���Ⱥ��kK���ڊck+�������ꮹ�F��<k�ʆ��f���f.o	.k��,��ίpv��;ʭ̶�9�ڳ��7���\h���5��A��@_����U���2��z��z��*W{�uN�>��6'h��kj�꽊Z7]�7T��s��s�m���\��Z����&�F��:U�ԀΪJ ��R��B��\��̰|�T1�k aM3X.@_��eJ �5����r��!6�'k�V0�5[j�[k�k���M���G*m'˝�J�狜�
�W��k�E�wK�V�?�*|V��(��]6�/j����3����XzN <��FӜG��|F֜�cʚ�����u�û�Ǯ��/h^��a@Ss��="Eϥ��d�gb��lߗ*�Q�wI
ʚǡP�W��H;�wA4!As�˃Lfj���ߣ��"&��T��S
�(ѻ �PE<V��j%�t������L):%A��{��="�N)o�ݢ�oS!�l�V �[4����RG�h��l���ex-S����iRs�4H�m�b�j�F��P�,�
������s�.��:�q������ڹ��эW.o�s{۽���y�h��gC�l�qs��n\�p�������'���ѯ??��/�|��ڕ�k�V=~���Ö����^��p�����K��/_i�t�������۽+�oW�5'�V9��s{�����6_}����̱f��.�ΨЪ)��	�qj$�r�Ұ��pD���+����=�{�ᢣ��x����;��ܓ�n?�Y���|o��Gsvݭ�|a��'+.�b��O����ػ�wܜ��n���sv�Yp�a��g`�o�v�lͩ�ug�6��Zy��kG޼u��y�5_f�����
222�i�;�५D�E!��A���!��15��0�L��SO�����-�����k��6:��x;����BKu��إ�6)�:����I�a���Xl�Djhj�i�L@Mj�d��NSSSA��e��H�2a����M|��g��2Ry)(']�q�b�Q!�i�.�4Ӯ(�j�rL����|KM����Y�i��:	% B�����ij2RR�%���cJ���d�r��3Ň'n����Ƃ>�S&�������P�����|f�Y�ѨT*�R�Q(�r����b	8`Ό��ғS��I��������3#
����S��v��d;�h@��/�oj~Ę�q���ILMK���BÜRsC��ԩ�V	?ljҒ�S����fDEO}g:舅"�Ǖ�y�Sc0�Q��$�TcM�V�s��v�U��1; N0�u:�V�j,�������:p���Z��؁g�OZ�S�S���#�(�;	��d$F��Ԕ:��Q����ӚI��ud��i^650�j��Zc/�,k�4��5��jK*�%��<]��ε�?��UIhĨ��c
B1����y���p��P܀~dLx�"eh�f�ԄE�yL��\�D(��IJf'%`�b������D.�ث�t�SY�V��e^Y�_^�>I�_Қ+�(�,*�/-3�T1�fe=S�aeh��0/S�J}o�6,h ��r�S�1ou��1S^���7�a��iXB/6��Ɗ����O
�$[D�� ,� w�;��4=I���IjU`j)O��54"s$ZJ�7��\9�� 45FZ��Ԉ�,BƦ�\��/Q�R%*��jd!�\��a�, ���8�grʄ.�R2Sc������%��f�Ү�5k3�lw�t�F�w�+=p����Cǫ�?r��؉�=�n9rt�������u����o=�h�Ɠ�ZΜ�}�B��K �i�pt²��z���=�G��n�޼nS����˖5-]Һ������(�,�]����]�z���){]S��X=!��5����YS��P��Y�Ly�q�ʸ�޶���h���\z}�t�_��Elu��[�0�f�٬�mW\R�V1{H�q�)֐ }MF�w ���׵�w]�O&����\��Ɛ��k��(�B��A���@>�
�S�G$� C���P�P� ��C8w�Lm��35?^L�������H��^g�q��e6��� x�}��Dʚ{u�ާD�d�G
)�R��@i����;F�u}�$�ja�j��4����݅L��͞\�`Ͷ��l��h @�f�Ly�|&�	j�%���Y�-��3�Lhj �k?AM�~��,kzB�i&#�Ԍ�������	U�b4���@g�ʚ�Mz�w���1�����LS3?VL`BY3����Q�Ʒ}a&��5!Y��@S3��Ț�/d�h_�d15�5[��4���ط������7��3|x#Y���j��7_6/a^��|��ڝ+��.k:����h��ݝv-z!k�dͤ����ֳ���	��SC�P�D
�H&����	�j"LMX� "M$��W�X�ϰ*xhM�5EWCZUtxu�5�Gז��(=����ֶ���Y߾uiuoCvG�+�(�7����<��ce>=�R�}Z<�He�	��N�E0����b��>�Z�k.v�*ܺ2���,��Kru�-qI�9Z��&-�˂&"π�Du^)�,��ׯmaV�_ݨY^K�W��D�+��
�`�tE�|E�rU�fe�fE�
 t4��d,/�òfU#k"M͆��d��
&�fs�nK�n{�ag�1ljΗ�.�.�L�����e���)>�>�y��MԪ3r��TzJ$>-�I���!Ss%/`�E�:���0N� �q4�&�p��\ǈ�(1NǼ�=������'R�C���:Çj�{
��J��*�s��9%|*`r����<	ɚH;�C �}�� (k���������w�.)�+"��I��4~K�ޒ!�i���>�I���-�'f�=}M+:#���8����Crΰ�?�BG���&$kt�a�h��\�'�iѥjd��7O����^�Լ:��@��W#u*~��W!A�(�(α)�����i����۰�k��e;w�>z|��s��]�p��֫W�߼��ƭ-�.�����}t���o��7�~��_���o1�ޣ�s��<����7�.8wim�o�߸�p�F۵뭗/ͺtq��s�\�s�b���enYo�5/^`ojpUVZ��L��i�UJ�P)�
¢"�4�A#q�D�ĦU�FO ��vv�M��fm�4�໋��j���g��U����v<�}T7z�i�ݦ�k������ػ�>��)��9�i�M0غ�Nˮ۳���8�x���G��n�R��r�櫕����u�Ȟ�Z��lȭ�x
h���*�$�����B�

��,����(��Kmd)�>��15M��jfg�P�Lfjz��ucj�
P!Mc�m��69�f��4����AKe�X��d�N�����,����(h^�4�L���-lj�m�60}}Ec�u�cj�������|ဗ���He�jx�O%�ur¨$�`B�P���%#�k���AGa��k��i�R�K1L#Y��iq1ɱ���Ԥ�q�'�B	�S�j����_�15������P�@S���&�`�������G��	��Z�RkJ�����`��������~Hl\��谦��1=ꝷ��L͏S�=;am&35��2@[S����e��\M����S)�$#)=9!%%).!~�����NKHJ��e~�'7���.��j��t:��S��CM,���p���v��^/Le�Dо�s� ���8X��յ��MMM���---���eee�`��ê"��NKp�灵����13gF��vZ�t�o����D�ST�6e�[��	���9Th�r1L}Df?�/Q,��BS�]k�	�ʁ�v_�m���W�ꬶ-(��.2�e��;�m���B�J���4�RO�0���M2�5����D��x�@ol��[0)k�\���F�(�#0�Kaq�Rq[�!
R�F�*�Y���2-
�R���%nY�[R��f*Z�4s
t�t�u�Ku]Lp�@5J $p����S��.�--�t���E����\iG�dn��-���H�Ts@Zلyz�)�L*岰�Tn|'�Ŏc�ǰ�f�'�#��+79��%}�MOD�)�Jj�v�V	O.dKU�NMi��"Un�;`���^��aU��R���e�P̧$l��#�y9_�@dr��恛B��r"*H� 	� A
�dqd.2������ϵ]o����
U%��z����Ǻ��۝�{ݻe�9���pё��NV��9~�����CǪ���R����<Zq�~ϕ�K._i9s��̹��g�Ξ�u�r�嫳/]�9W��_���^��~���#':��5��e˖�u�[�5Ο]�X^\�+�q���B�F��Q58^�Ԭ(RM��R-`��	��a"�ׇ�3`��p�qW�m�¸%�\�-]3��C����N�U��L�!-�U��Fs���!1{T��G��!$y��4�Oً��4��{����o�&�����|���ol��Y�M���/5��U�O�Oi�#
�� >>���q�=}�3�� �����15���{�ﻘʏS�5�SS��w��q�q�j����mhj�8�8wp�@ ��~@�*�T2hj��7�4�	˚�e��x��`�vw�j4K�9 ]�)Z�I�Hf��ܱ�40��3� �nL�+4$R�t�Ʃ�0���\V0�cj����9P˸08��*��5���f]<��F� �����ҿ���CЇ�8�*�� w�"�_�����yY�0�f�wx��ׄd�XQ��p#k�_Ț�}���l^�S��qhE���=�Vݹ�Ȯ-wl>��Y�;�`�̓;�B�2�aj~��Ɲ+�Ww�߹��Ξ�.�^�B��ɚ���bjν05�F�Oל�Vw�qzk�d15�?��@YMM�� ��"��qte���p��C+�*8��h��"�P�l]�����kJ��(?����袳#���5�-���+jʔ��L�sJʌ��G���o)�?I��I���L�� Ң��)/A��IyI4�P,�^Z�3�;u9�A�*.K��$N�&ǈRb��	4+I�O5���AR$�Q
n�W%��*�*{*�+�k��+�'M��Z2P#�d"k�˄�JE���ي&@f���b�K%�e%≐./U ��YU�Ț5ej��ʾ�5[�6Uh�Vj�W�wV�WX�U�N�;/��.���8��ox�g?*�<)�}�x�v]5��+aMs�^J�15�Q�".��	/��T0���h�]`���o=N��ț�w���15��|ODJ��8�DJ���|j4f�>1[>2�3<I��	�(k&�9!�.�@�8Y�CL�!V� !n��M�)�ߔ�we�C%�T˘��f�S��IqM#9KNH�C���C���#2ވQa;�Ĩ�11�A�Փ˵X�Y��-T����}EL�����I�R�*��$.r(�ܺ�lWc]���:��m�ҿmd���+�\���ʃGW>����5�/߻oŁ�N�{���/>���_���S?��/������{*׮�ݸe޾Ý��w߸����E7�-�vkޥks�]�u�̬�'^�����+W�:Q�cĿr��s�yn����^T���T:�2�R��d�\�7(p��tj���:�b�RhS�,j:7;/;�,�������wGˆsM#��w>����b�{�;�W�~^������v=��]7z�u߃�CO�>��Y��V�;�{'��<���.9���箺�[v:oՅ��3�K��(���n�q�α�Uk�Y
�U��)�j�R��3K�x��l�"h�Z��A����&��i	��ۚ)P�	CG+'\c���k��u�к0�e���&g�����^j��3��tA�*S/w�ej���&8�Mز�ҡ���4L@MJj#d&h��LY��L��$v�U���jj�F�e�ad�N8�4KJ�i���&�1��Nm�W_�7�f��slA��c��i�7��`gp�3⠩��O�i<�)R#�A�cj���0�Rf�f�0������������@ �r�L&�a��(U����*Uj�B.���#�(�35��g@fN3����1�&�ife�"3�^aj���aS3��8��Ҕ�+q�3��E�d?I�t$#)#%����ӦGM}g:8�T
�����{|.���ˀ�&����6h�Z-8^������n�Ng��
�P7��*##D��
����*(((++����
5�X�ŢP(�� I<����G�����P���hp���x+5n�I4Ӽ\���%�vQ�k?�Ρ �rŀVF�0�������(��Wh:_T���l{뭃-��zwg�c^��5h�	(�,�حZ�"���R(�#��(&x�b PЄ����$�À1I1�k��w�6�T*�H@��}}�Qv*��B\��x���b+R\ '*!��
���"�UR���A���A��2��*�n�ѷ�텦�|ݜ�vn�fA�vI���0y��F�5]�Z(h�vq�raP>?O֑#��%j�2�V/����|�F���#+�����SNX�$��є^Mð4���s3Ĝ1�%�sd���$౥(O�b���6�V�q����Ȕ�N#2JQ��Һ�����;�Z�Ei�K5*J.���H̑�84���i���Id\1,|#���TM��ť��SB��'')�D��%r��V�T�1�e-jK��
��&բ��e}���,�F�;����=x��ة��K��.?v�����gK���dûm�����}����������|�B���-�/�]�
�̽v#�̿|uљ����gO����-[f�^�Խ�aެ����oI��&�Z��U;M?��YU��L�D�h�Z��4Wv�X����p��\�"�:�m�v�x�U4b����lX��q�K8#"�.g���Fx�;��C$��yϣ�<��U���<�7��|����ߘ��[�7�����Q_���ȧ4��C�!�>�0��8C8�IhY��������Y0^�@&��y���}o2Sn�e؂>���X�t1!S/���w��.I2���L���@�x`P�6�o�׌/d�Uyݡ��֜�����V��Rlϔm�W���
�@u�|O�,	��M�	M�'��0��fI�(�8Y�����/^*lj��ܯSק���7�|%08!�$�	d͏�i&��gg"�;@�/��L�i^��G�-d4� \jx)#k��Y3�B֌�LS���bcOզ����m��wض�ȎGwl94�z�H��#�����o?y��ݫVt���wrW��=K/�^�B�,x���15^�>5T}bk% t�9�0��ԀЇ����| �5���ВO Ƽ������Ȋ�C����r��f�-�=8<����@>�[Wvzs��-U�7W��Pvdmٕ=���Zrl��M]��y:�1cJ��)�oOI�����?M��YR����o%Ž��vj���3�H��Ӕ�odD�͍��K�@��i	Dz���fU�s�F�Z!�ӦM���$mڴ��S�g�#H��ғȴx~�v��xJ�^�d��5��(O�U��7�ժz*�=U�eՒ�JjY9����-&�QP�,/��/b�P� ��EzԘ�YY�ȚHS����5˵ hj6���Th�+t�++,��mgʜK]�J��
]7�ݷ�����Ks��Q0���k�]����L��Y�d��\��K�"N^@1@X�@/}M��@M�����@M�:5W�|�l��/Lp���
E�i���l_z<�����������sJ�@���Ț	'h�<#H �<<C8j2SsW��M�m��5��"��LpK�ݐ  F�(�GZ�S�D/{fR�kV>2�7բKr�vV�Q���N)gT��4���i��ECfj��X�A�T�N%g���H�^�:���15� 5M����eA�ER��TfY˲\�e����uu��kfϫn[X?ik�����V�]�j]������������o:p��O�_����Ϟ�{eɮᢥ���������A��^Ggľ�׾h�e�bK�Bmk�yN�{qgβe%�V��Y��ƢBcv����Tf�L�W�P���N-��PeS6eQʼ�?PZP9�n�ڶ���6]��|�d��ʑ��;�V�~^���#�~�y���]�w�o����г9G��=�؂��;���Ӽ�!Yr�Ӯ�����>�^κkξ3������u-�]��r�awˀ�j�����/�;�F��l��z�^e�J�FY��Y�%h&MX�)��&��i�P37O4�UT\M����`����3�'8��upw�!�ap������>$8�u.�M�޻����~����ݡ��s�:<Lβ-�n��%�É�x?R�]y�
�׉G���x�����涄�;�B~����r��p�T�f��r��8	�C��~Ӭ[(���a��#ޕ3�v2���&�7; �g븯 �����Q5����c�i�N��No���I�H�]l|��a�G�s�VJj��� 4�[ൗ��������~��Y݂M���a���iFu�_�?��W��*�l@4|x�Yự$~[��i�t��)��I��l|��&Ca����H,�@ҝY�Ϸ�/�S��h�9F\�p�:.�~�j*��8�Ü!�)q*���+i��h�ŞYR�y�r�-��b�0�>�s�?l��O��_��T�1P��������ǫ�������A���L�ϰ���^�O8&&f3�,�8;'�\�_��>����O����D���nuENS������JeU��U�_���Tw���7�Gb�l�%F�a����}mՑ$h�����]�d&e����IPR��U���'��.��6!��#<�����uX�/$�rLSc�գ���(���LɌ�K�H&~.����C92�1/3P!���(�8X�Xc�}M��w�w\#�>M������jV�*5Pð�84�f<�2���㒐��X"o.f�f�������^�7�\m�������N�&	�b��u���[�;�@�8x�$�8��CB_*�Si���H���H�Gd�$��d\�h�� q��Y�o�+�=GCL��:�t~T�Cc�&I��8��$J��M�6O�+�T����k�A�����\�f9�#FKF���BaK����)Z�gȪ"������?�1[yVO~,#�X�P�e��,��4�~�����eT3�_��+���3F��
�	�5��p�?�ѽ\͕���x���	'��8�͆���k�귈���x��)��G��w�	�}����^~z�;&L��*�a4L�p��&�
�i+@l�t�m)s7���[�h��1� ���܊����L!�;���O�~�����B�q�{�������@m2���(��O����?0�~Q��d�48/�w��C�T�-l9�)�U���T�r�q����v��?�V7+�=�����k�Gw�M�����=�c�m��їw]䆄[�(�g8�M��搏�_D�B�M��s\� Y���/fdw�ֹ$DFؐ�T�E�\۸�p=�2��W�
��H#K#�}����"kX$�}X��c��D�^�`����i��^��ǅѭvz�Lc5tHЮ�§���+�6�/0�]1��l�Jx���>�>�;�WÙ}�|_!�w���H�%Gu�@�Ʀq��
����D\�p�	�Q�1�X˪��:���^m�R
Y_��2;Ή�V�H6!�<��ؼ��r�����C&��<>Fu�K��`������)&�-���1,H��O��S�Grmg���g�F�����0w��|)H��^����������C�]��9����Փn$���_`��*����ٓ��g�Wd��n+$ivO���}�c[Q����}arF���o������lG�_[x����o�^Z�--YP������hDx�\�O��E} �!�N�fg/ī���<��{�"�h��8Z�ݧ���_�#�̤�'�o�;y�y4��=c
�?���n�Y�I�㱯y>S�	�Q|���b@WR��:�r�����k��O���)��P_b�+���{Qu����R9M��\��X��~쓏�1͕Q)M�Fi���j�c1�������Y�S�o(��;f��~�����P(6���ʬ����ف͏0��h$rV���_�<�-jk��<9�|�r
wZ�����Q]���Y�9��>�����^E�}KV��f8�p"���h����c��!	i�7(������n@o���=�K�,+��	�j�E�����ѝ~C8|�K�_��aOs��k;;�<tv�>����!����w�7�D���8�7Q�y7u0��o�.�o�Xn&`�Q����NQ=�J�(�$:1D�:}�=◳�h�ݺB�a��h��[��׻̳���hv��X�i7����~����Y�_w�8��x�TÇä���A)9�ؙ�66E�������xr�!Z
�tRb���ʘ
���g48��+8�j[�VNO����7�,^���}w�5`�hF)V�JGR�+H��D��s��{��&��3�զr��44����k@�����)V�3�-NUѪ���s�[���w�¥lЗᴈn4V���F1���v�ff]���և�u��dVč������_�w�������.��K�f��纾ti?�ג�,;^���[5���[C�Mq[K��&�g�t��S�f���Z�����wv+m�D~�i�aWO��<Pᠤ8��4ۨ/=���R�P4|<R�͙�J�t������07�V;J;��p���X�����fK&�S4��Z�>Ռ
�ev^]�֙�&�9,���[����٦K�LM�є�F�/3�@���!��J�(b��ۦ� %%���QTs;�Fb�i��@_	p��aL�_=_�;�a�zfD^�%���,!h帑$�c̄�|���H���ć�
�����*����/rjF6y۞�;�����2>Լ���ڎ+LA��,�LVhhh�0���Մd!��;�h�B�� 4�����F�Uɂ�W����3���Y8�hw ��'����S��'��v�|+��Z�;(`ʙ�:�|XOw7(����k�+�4���Ú?b$��󒧳g�Ib��BD2ؘ�����*�\P���Ӈ�c�@���|���^�?!..���(`�$���v+vs�9'^fN�3�9�l5��>H���ՈZ�L�&�$wL��#a�=
2?�(�}ӝM��N��j��)姙�ͤ���0N~���d����Å�ޅ�/��o�TaA�Z&j���gt��eV��)�d��Igڠ�ʫ�P��I�nb����IB��X��C0�e�S~�w���i��\�\d~K���� T����	6#�B�ҁ�*�fVyM�"L��$gW�J6�H��~���J:Kh>�	&�<#s4���ZĳF����/ K���( �l
b��ஞ�΍��YΝ����6��&X;�5
�����)��k	��C��{ܵcDW^r�b�^1�?T������B�߷Lga�EK)Zu��(B}Ǐ���O>Ni��!����9NtcR&S����mR��2�b3�K�2��FIG�i������#��Yk.��9G�^�
��`~��4ɏ�Jgv���/RY8��f�s?Y}v<�Zk��9�k�s~z��~ �o�$3>ݱ�,[����Api���!��Hj���5,zn7?y�	V����a��i��hN���6�W1�w!����Mx#���������ă���]ΓY��W2�N�����';z�Bb��W���ߚV��a���t�k|V����
�'�=��{��K�y�}&��y5�6�˓d���%�g����+��ق}L4���bAOE�c�;�*��
�&�-T���b�K�(d�wI
��$f�3B_�F��C�ީ�����8r�l���39LȔ�6�68�U�$Ԏfn63P�R���Db�@<��p[��x����pV4�4�5��&�Js簮�c��g�D�I�2������"3�k�zc�X�_ڞ;x�4�d�^�pς����}�4E�����L\��d�3�yr���I����]���x,�ۂD4�_ �T ���O�d_ܹ��L�����x�g��A�i�7[
@j6Da���Ͽ��B1P�G��]�0_}1�U:%��Y��( �?��v��nD}o�'Z��b��.>�i��L�{e6&t.Q[{���nKH����æ���~Ʋ�5����PRf`����M��YR}�j���B���b�=�N��"��%���BhG7vބ�����q�9Չ6�7٦{�M�y��T����ʄk|�Ƈ���Z������������<T�tS��80�TݪI-�p���ܯ߷C��B�����F��N:@���J�,z��<}b�h��>} Ǩ��Pi�ȩ		���&v�J�F�B�&�=~k����G�N˅��r�׈�	e�6|n
��A��,⮊��)@ݾD�ښ�eg�UU� ��.�)�+�T�Oҟt	�D^D"��de%�<[�8��E��I���,n��e�%�ǹ��n����,��x�����������8[5��O��!(�aa���������x�%�6�;n�T�3ź
�#�7����{T�O]���hv�:u	=�?�mm�dt���*m3&~�M�|��[u\OW��5��ܼ�X�C�7P;��^�6�?,_!`�`��|\b�;r�Y��.���
��"��R�	�	�D8~5�>aC&�mȒ�x��Iٝ�`��h��*����?>ԃ0Ȏrϴ��k2�3Jȗ��j&�7����U�S����iM�q*�Q����}i'Xc��l&6R\�H[U�1���͊b�=�F�I���������^!�����0Rc<{�R#��A; ��)�f'U�E�2��;N6D/��2&5�'��' ;f3�φ,���F^n����� Hq���lR"���G@����>��$L��%g�$����Fv���$H��i���`r� �gݥY�7�Z/�l&��Qy�W��5w/�\?�G"�A)�w���$y!e�Y��ʙ�4�T<����/���ѡ��ۣ2�zx����"W�n���e��ZU-�����r��TT�/�9_����Zߛ���5��}��ڡ�G<i2o��5��'��)�ӽ ������>�x�e������K�g
:�]��0�Μ��@���k�	����
m��ׇ_��9�PJ�������
mI��B@%�'Ɩ\x�]��K�!�w1wo8ۃ$�q��um�*?�	v�`m3k�������:Ů���m�YC�L6�Ʉ=�'�%����szgcD2�׎ɟkFk)� G�����j�jߺ|�̮���`�/����M��Dh΄e�/�Ss>�p���'�NI���T�S�81�����X�u����c|�HjU/��� +��F롁��B$շ�����J�@-�#��H��wU�{w�����܀d��?0�x�<uk��XU��/S캨�($o�;є��A��, Ñ���k�HA�j���>2/�`d3��(4��L�Ȍ++��@;��#9��mO��<�
��!
`P�Q�!84�)�ر6���Yc��@����S���L@2������j��/S�E=ێZ��z�U�q%;rs+bC��dU���~I9��a� )g���-��8�W��1�w9�;8t ������Q`6bA?�[��\��gv�|#�}.(8P��~m�R���/6R�F�V��X9����?�<ݎb��_�1�o��'BL ���T��l ^�
®	xUU��Hi׫�ȸȬ�s�nș�1L�0g](1-�=.;4���Ch� ���`��Dc5g��"���~�g��c��+��!��#�)��q\��8�d9�����L��H���Pӡs��?&ꛈ?���ݘ�#�ʲ{� ��ջ�o���1�#�v��2:+��MV׫�)y��^��eN�3����&Ԙ~����E[V��Tz�ϸ2���v�S˅5m4wz_5m�p�AP�v���s{�sQ>��T�c a-;�i��
t���æ<~x��Q�F�%��`-��T��,��O��$|o|_���GZ��+���q�8�����;�"�,��TU���R�c�����H�w�HANu��!K�W�J[@���v���sT��&��R��-W��(`%���ξo5YZ.*�Tȷ���`����CZ���E�l�Q���5���5����e����'��3�>W��6|�h.Aԃ����e�[��~D�1��Շf��g�n�Ȕ�q� 1�[6=-×��]a������]W\ܷ���x�	rm��%���i.U���<��t�%��Ŗ������9��`�B�'q�r�ʯ�Z��lj������[��@��^'�E}+�cf�c�;���4Ĥ�\���v�&)�yaH�p�i�v�&k�k���<�˴W��(2�W��)��l�:\�<YtW�y�t���M��@�����}�e���J忷i�Ly����8�^�b.G�6�C21)�/����J(�-|V�!hI}���4��7����v:�+ܳO��fs�J��_2(�>���x�i�a��h�0�z�J�uB�0L ��\/q��^x;��F�G(��g_?�\Q�mF�y)��[�	��O	�ꮮX�Q1��<����<{�ĻZ}N��מ�Vv��D��62BZ���d@9�5s%�Ni$�{<����V>jBa`�k���L>���5��T���+G������ǿ��s���S��2��3��DN�24��h�Ա��-0��M���]��@�c�V�BEX�%	����$�3�,��Fxs�����l=[�CA�Hp]urd��*�Ҩ#�C���IO����t��� ���s��!@�4� �o
*FZ��m�}b�Y���WN�rJ�^%�z�S��@_�9�nI�i6М��� �>^�s���W٧�s�Gi/�ƥ8�ex�l{��/���v���޽g�3F���G����e�IdZ �t���	��e��g.FF�<�+�L�H��
nJ0�M�[�7G��Gz)]�**�]V&*ʹ���/1!���s��xI�p\��O�&��/��37?���3&Fΐz���PV~P���%E)
|��I���U�Q���FM��
7k�����o�j'�e��l�?s/&�Q��1�ڥ���>���c�d�~�ty�s��o�.����,�&�r�,j`MR5���(Xqn~( RY'�b��6��;����V ���
jWU|m�m�PQ+^��^��Բ��0ҵlRݯ'sYv^�a�ы��e�+=+]�>�6��ω'������M���u�hc��Ϛñ�����_����v|��7�J��G��<%�i��!w�L�zB�陞���Lr��8v�˒�f)�����˂6��E���OL/��9���lK��2�t	Ijv�����KQx�o���4]�V4c#�7%��� r]n�����Wo!�sz��t_�����#�#?L��6�s�I&qt��F�[п�;7�]R\ƥJ꠰k�x����8�2ɨ�������)��8��)	�DM����� �&R�66^Rƪ^>c9'���}}���h�3!ק���o��)�����=1C1/�l<{dvLA�ʥr��3�e<��N�DS�w�U�~Oo�`���c0I�W:�^����
Q�I|�	HDK�D��7#����ٴ<*d`��y>	\S�k�껖>�j�2|��Y��q����%8mk��=�R�-��qޱ,\g�K�z٭���ˢ�7u������tt��z�d���*L2�,�IG��;��ṓy�$��Kؾ������n)��8
���
�i�=�N�E�Y(���d,S���,�̢)`�K�.�@#b5&��6]�J,<��<��1;����n!?�C���K�h4_%�l�����-�
WV��E��XÍ$I�Q�ɉ���Ps��)��O�{a��
��?p#�c��X
�;�M ��ʨM��=0e���%��b�70&+'#'���3C^�0�{�ZWse����:0P/���º>�\�k_��:�32��a�\뤩`�:A,!�J���L�J���R>����n��2Z���՜������J8�2;��2���!���
���@v�K̡Vbt�Cʠ�l�^�Y�Ջ����WTdMdK���?��9�	��M����j�	���U���YYY��ܜ����K��]�Nv�c���| �G���`�����Qv*�x��-+v����n��>0���.�!ǿ��Zņ�q�9Bh����L���[��2�h�eK�J�u��a�K���4:�8�7Ɵ(L�?��h[���1����^l^) �M�ߵ�;�`����rY��ş�� ��p���P�6�vBtٌ�K�%Y���;S��.X��{I|��`9�M�ZU�js�vZ�0��� T��~O�(�T5�)�uOz�9@s����Ţ�s"��Y���Z�+�Q;n/,ڶُ��Ԣ�B�P)�դ�/yl��=�ջ��O_:�k��\K7,�d���z�3�1-��$�P�W��'c�.m�h릑'uR�s1܋�:n�N�N�*�Q��]]b��2�-�����J/����G����OU�M��\�S�Z�Z�Ho6��g`k�$�EBN��	t�\f"ݷC8L���=[���]tC7$�ku>��5u�O�E7/m/c'�/e����7W]�agv��6w'��7��'з�����D�*/N[V_�O�e������Ar��Y��7��j���yK
~�7`��x������Jm�����t}ܵ�v���fLk)� ���5W�*�e)�5(4�H��2�F�����Bª�m�&��Z'lx>�b���>���E��ф8�G����4̧ˠ�bS>>R]5I�'��E���%�}�A�$�E@j��ƿ���|�Q��%V�w��5�u�K��;��'���?c/~#�H���8��N���B�H��N-������mq�Y�C���:p���1̤rxC�N�%��-�����m�[S���e�Q��3�d��B,��;�4r�v���&CC~9�Z�[�a�*��؋Fm�X����� W� /��T�.#���ix����h*�F`�?���n �W\�:�"�(idi�;��FF�XB�GVUg*���V�����Q��
���O�t�0">\ŅQ:�;q#��[�he{H��Y���muop��7�@(ϰ�g��HY^�)�0R���x�V s5S[/aKͶ'A+(�CA�	x'��p#�b�b2msHmYj��V���~����3��_�OL?޼ܮ4}`%Ym9l�9��1z|⽒�Z"z�cW#L��͜�W����B޳��5f��oD�,�,�E�Y��&m�4һ�Z8Mv��f�D*��ϳ������18N�@�'�d�}SR c��2�2S}��nr���p�D퐧�E�@����"�R�� ��Q�+Jh���ѣc�����3���y7$�w/�J5�R9��	��g$2�ss���cF갼?3���aZ+\w6�,E�\K�ʰ��Q]/"�I[)�>_kL���}AF������Yi��'8�A��7�h�$�PO��N��Ui5^ɒ�
GںCZ��ث�{!yHӻ��Y�
*�Kv�v_��gw���."I�'8 #䝃��4G=le#�,8�ZG������-4X,�89���[�P����
&z/"����o:�V�%���$�K᷺_F L����2���h��ۧ��>���r�� ������SA�FT�dGnל��@���-E�(���Ezd�b�`FJ<�6P��@��g��X�4�{/#o��iѳ����ѷ���?�����oV� �ыF�I���F���O��D ƴ�������_\T��ׅ��,��Ti�B��(�1�v:i��{z�Z�	[�����HKK#�JC���GM�G���g �<8n�!3h��ڽ�V���г����q�&�?H����®?�v^��]�����3ԭ �F�y��Na�y���_��?[p�zY���X�L��[�B�Q�h{��1����t
A�K�Iї��5�e�;u�\��7���;v�fXV���<w:�;��|����l��`eZ٬ڟGSX�cQ�v$I+C���u5YcBb(�c���X��f����S�yOkcM_3F��]U��ߑ5�r��b�j���O�o4#��r-t���EX�5����:yS�I�q$(���BN!��	f��ȡ�(p�0���X��E���}��{j�ϫy�Ecg����2!5��ȵwəa�Q�(P���{�DtR _~�������u���x���o��sIcr]�64�p\���FL�`	X\6��&I��fE�����Ycn�����D��ӥ�L��߮'li�G�'L�PڷC�G�Yp(,��l">����@G���h5���u|�)�w�h�/Q�C�+�b�r�n#sh+�[���&A����h�ǜ~b��x��
���mz��}ѹT�
nl�����J��������3��S����p B�����n?��x �N��x�o�0����>�F~�S�J7d�20u?}��FEE-TYhjh����)����f����D-//onnB������N	w�:��/���Ō��@�))�"��st�pZ":Ï�K�roU�(����l p�H�k��pώ����/�����H2[i�n���V)qw��c�dup>�PH,�.��`p	ϓ8��P�q�S��������֜j}jl�a��N/D�2PY.�,E#���[v�8�'�rGI;C�N�N�Y�[�A������#��CH��Z�G��p�V]�W�2�{�¿>�>n����H1Rm��@�dp� ��Տ#����^����8������J�o�?�L1m��Ku2ϧ�F���H�-�Y��u���J�yI}�_�b�bIVi�%�|/�u��Y,p��\��s"�Voo9u�DM�\�V��\~���=(q8⪂rV|�!a-��Õ�H�-s�5)@�5qI	���o�Պ�m������Z��̿�>/�iC
�Flon��ٯ��x�v���<�e&x3Cη豮��|-�yʺV�������ϗ=r������|�g��؛9�6��6��xW��NgK��v6��o]4�[�Q��Z�z��W�ܞ}�*���}�*��r�х��~m�T�1s1�9d�p"	MN�.�].)p�|���cf�Ae.}�9KZ٫�gV�j�:��h�җ�_D��6�������S����\��P�5,���p����M�	*G�[P/s��j���E\���Z&�nL��Zݶ(=�-�1���>C��=�/E�����ޡ��:����{������LvF�J��;F��A.�qywFiR��`�0�л�۲�DԏRп��c�)����CE�г��t��h_.� �O�����~lwMe�r��+�����C��҂��E�nG���2��xr�0�K���2Z�d��ǫ�!�7������;,���U�@�t�i�|E2�tBQ��(��)�#q��(AXP誓k.�39݉e�z�J�/�qM+}3�+M]ġ#��4&b=�q��&	A���:\��io�:9�Bޛ:si$ߚ�Ns�
��RE��" A�p#SP��{���ϕ�X�)�읣>����In8(��A2����`��f7k�bp���n �_,򵺧��蜬ZK����;M����G�7���pv�_ْB��������tBw���XBhc�/ܰ��F���7�ֽhP��dhS�+��N������Fj�j�{��6\�¼�X��[2mf:#\�\}�#�~�@��E����/V:N�����z�}��=ݎ11��J��)�Xzg��X6�ιi��ڵ9�A�U�T'��9��/9>4��P�D�5:��A,砷t`e\7
�'��`�Ѯ�̥ɱb0��HM4ϬaQ9�&v��������P�\�x��SZi*�$�S	\�'����E��}�Mo��n�`	��������AU�LC�LC�2�j��BA�bQK!u�F-�6�v����ձk��Ka4s�ё�ă֣ZQ��3k�Dz4fٮ��?��A��`5B*�������9�^�4(M�\�|�f<��J�W��5�O�A��s��y���j#��eu�|����q�����Pp����-��
k��鐣�H. /E����=���kk����(����t��3b\�6vz멧ۧ���<YW� �J���X�QDJ[\�Es��؇�i��2��>JsȬ���e?F�,�/�����nx]���`b� �ggj�'/\�4��ii���Z�W�vƔֻù��9(Sˑ���"¬%���cT��k~g�J���-���F2�b�,<��`$ƃ��(�|�L���H�ѥ	+{�ہ�
�
".cU���
��D�>����J)��(��Q����Q�ыsv�r�Ҥ
��-�m�i� u�����ꫫ[�+k2+Y��W������,�s���H`
]"|�-Y&͌���*��֯pA��Y6���s�5���f��sJ-�5�h\ԩ��":�k;�~�bL�g40d9+ǭIr*�J�p�<ή1P����:�F�ʅ3��74�L���!A4���L�ך���	��<w��8L!�d�HP�H�?ّB��i���?��`.�o�fC�封�Ԫ��C����r�GL��]t�@f. O�j�D�U���h$��fLV�7P m�wY�l��OJ�,�xY+�� ~�$hP"�>^j�w�� r�s�;�֯����4���`33��������J����$�49��}�)v��6�I ZD��C��D�M�]�g���Q���6N��J�Y�g��L�b��|�H�R���}��w8�fMy��!�"i�C��tw��|��mw����¯��aŢ�̩��DG��G�R�<ջ��W����
Y��������rH���[7b|t�*((������jm�坳���}{R�AΝO&
�@t��D�*����#��4n����8XdⱼՕ���/��`.A%�p�a���x_�ي:T)em[�F3>G*gíi
	RX�z(����匩��Q�{��@���NdtB��e@��S'�	�F��U����aH��E����Dj�G�q�C�hb�rxqZ�Ɵh^i�A,#ZV{"D��H,�<cv��7���v��gw, ��4S�<��#uBa4����W��YO ��J�%�+��gJ��<���y��mh����B0�����B��t�����2���m��Nu��2�8c�f���C����?E�k�kgEg`�{�wl^��y"%#��i�D�,��K�|����1^�1�{&�V�x��nd�@Zw����]֚�`����f�إ�<F)�p�P5)y�uL�~3�<�RIb\H�J�k��� ��aY��@G�P�%�q���KLo�ޞn�
������q�7��-�b�=]��?����!ߐ{z2Qʰo�4�$[��{���t���P߰�{��7�F*��?�(����U*��4wN�Jׯyh��&^l����YF]͖��� ����bf�����b�� �����f��9f65Ec��|u�<pi�ei�T�"�"�Ɂ�Y��?Bk�P�ҳ��i��X���dyZY�^a��܂7����t�-ņΟ��J����P>��]����{�m��)�e��)E�t���m?�_5�5:�@>����L�;��?�O�sƻ����ڥ���6s��]������,���n6�'�c��ID%��HhiA֬���/@�
� %fC|��C6-o��]�[�S�~�B���&�)Jq0ye�K�n�X=U�&��8�����`w�)�17�1f�&Ap�l��G�ۣ�+�A���?��i3�w�B?ᨨ��qE�Ą@Qu�	5�q2�g�QtBP�5���Vq���FKH1[%f��2�h���hx�Wh�?�0�gZ�A�f$�n�Ph9��:�2p�b6�����ʙ_�.$"a��i�Won�L��tθ�%MAeC�Lx���3X� We��}O��U��l�r����>߶u�:�C��	�`yi��>�/ѹ��-���O��e~&8�N%����.�b��M�i������𳇥�AV���7F렾����~�n���5���_,=����&$�� ����[x����|��cU���R��$R��<�N�n�Ñ)YZw�t��z�����A܌r*8����T'".� 2����5@AR�G1�sa�f�-Oض#����jLz�<h3�:|�-t���p����g"(���Ȫ�����)��݉��O�\�dg��ǐ0��d�(f�D�+fR+fS�aQ�ć'O�;W���;��=я�p�^���y> �!�m���M
?�.�g�v�%�$B�mb�"���m�_�.ht��[��zO������hm�	�_l�<������KYxA>�♽Ƴ���I�wQ�K���},�#]=�a�tY1��l��;򩉖�ls��r�.�a���2�ۈҖ�Qd��Q��u��ɱ���%ח�����4����
&��Ը���������:6m����7)=oK&���ߔ�kDp
Xi�	k�"U3i�OW3h��)`�w��S3�����`9R�q��\�揑�-�&�m-��|�6aV~�����-Cת�1����=���߭��%7k'K����U9���h=J�?p�A]�*��2� �č	a��W���m8|,i�!�9ƫ(83V\��R�44�˘�E9��}��.���N{�!��~ND��s�0:��A҂����<����Y��T�28t�*;�őD�C�ϋ�bO��&��b��Ǖ�T�6�!�J�1n�b���N��S���0�(��ɍ���۾��I(Y���H��+W$k�%7ŝ��r�ߘ�o���J���>]m�L�-\y�)��3v����	\�uW[� _J���TC�Ucܦ¿����k^����T��655�fJ*L�V��%�;M�t���]\� ,K��@�2q	�����A��R���@�P�,C1�(�sO"9������v�C_m.u~%g=}Zh�BLRv�!}7o|:`������O�̌��xxxXY�I�����~�r:ʃ��|��.D4��ŗ��=L��c_V#>fD��cj��Y�ļ����y%�����YT�TI>��g���O&�! &�! ���p�qJ~�-��O��Pd}vL�0�T	á8�,����]F]�Ytkm���g|}}M7:CIIImmm�,�P�K�pxCCCaaannni�{����@d��`d-����Jxx�GX�ow��� ��C��yX-<��n�*�Bl{�9t��O�3�ߖN�@ľg�E 	�M����}�w��ߝ�mo�;g���F]��XT3$�Tщ�dq%����F�ү���p��Ď֢5Q���Q�V+b�
9y�K�4F���sI��=��Br@6��\��d�WJ9J����
22zR���Mr��S(�6C������J���c��I(�=F�.��^��^" ����c����w�4%-N�5�Q���^gP���H3݌m�%խn���TЋ��S_볨�����T;ׂg��~��!�
�C���E���@�Hc���~- H���L�~�
mU3[��6��uf��;Ǯ�e�|�=6�j�6��+��R>��bO����	K@�dB�䯺nˎ�|"���5b�{��Ϡ	�$�$Y��e��0� �T�1|��2��&nѳ��i�CWJN=�󀅅���E5�����Y��	��GJ�O�ϛD�~�/�nj���6]X���j�^9�EE�
7������k{?��\b���sW���M�&��~�W�[������$�P���������MZ���J�O_#jM[}�l�}�4��
���oْ�3l�Sb�fe���-��8�K�����1�f(���S���2J��;%��zsꘂ�;�GӯM���(왻�q��Mr9s�˺أ8xԟ3���ia�.K4�Jt�K�����q�:F��?w��;�L�V��	�%�[�0�r���j��H0���?����l 1�^0�V7(�N�v+|���b(�KB���[q�m�X>]z< e���'�B���+s�=p����؟�"�Z�
��Cp��f�V�2Ȏ��/�C�Is�Y�V����C�?f;21ΜM�Ɋ�~w�Ci��?$������:䦡UQ+5�pR���Ն^Q)�sf���E�X
^^��T�؋Q#��f $��4��hY�T �'33�����i?�8��F�IJ��U�jm��/�͸���<^[S ��������`?jN�k��$XE���[2IJɧ�0R�e��Y��L�:��{8�]͊}+�V�󿻞��S$[v����⓯M<5r �ܹ;$:���}G<�q6�8�}��IA#��5�ҳ'ZՎF�m=�L���}��?2\�?���V��=2�W��p_:V~ڴ��>�b�驝J#�C�u������zf~�=��u�9�PV
��-âe�M-v������S�ʓ�@�pc����`\)���zI��Ȍ� x@���<6���i8'e%c�>.�b.��sL���Zݞ���K�˕�����Ϥ����~|I�`I.�2����|QoPeͲ`H�����A)`E�tep�׬-��+�o+R�(��+�.1/4�)0_)t�.t�/�>��<��?��<�<��<p���we�+1\��
)0�3���	���,`|�3����w����8S�Z��&JDڙH¦�*�]D��ج�<�9�ؤ�8�������W�{k���?��]WH�
���ˉ͹��=��wI
�����25�p����aR���	�� ��aSC^��Ă[4yO%~����?1ʿ0*�`������\ֿ���U1}L�q@��O�>�A��}�Qt�,9l�4�w)�Mrd���4�t�fj����� �X��T
�L	n�8Tz
;!L&��8)����ؤ��Ԍd?$f��LKk���o>~���O��œ�?���FO�2�LG|�-�6LIFb�LL<�O��B~�ʙ��:%.yJt<CT�O������� ����?���{c��SS��	.KE��p)H�w���p�G%�iȀQ�eSl��c|�A���̌��N��N���Dǲ��3��Hgz��i���Iۘ$|f�`F<�N��쟼�:��)���.�I&��[Q�i�H\���L��L§��	�˓�q����/T��)g�1.�YrL�
ڤS�u��7Ef�ԂVXx?VLͲJ{�k���k`L�d�7e-���-u6�Z*|�b�)פs+�����`!ap@��� ��cj`3U(Y�9[�A{�rI���4�������2�IL���h(A�D̺3�L%Th$
0<�Byi<n:45I�`�����������A����b�LN��*���I)���*%%%))	��A��5����K����^������Ԅ��WTT���M&�QoP�r�TD�`�&��#�&���9�%�)��@���*��1 iΖ5�(Zr�s���ˬm���,u�G�o��J�^ST(:jfLxWb�1��-�����f2��*񋀗HS#2�<�=���.//_�`�����7mڴj�*_����������s^���Ʋ�2p���GM�V��������?��Oy��̌�=#~&8^�HN�E�ϵK�T���1� �`�ZsD�r�P�@@?\���%���*]w����2�l���i�w6dvT��
�e>U����%�\� i.0y�Lcc^ej�5b�b�iDb -�.:�x���԰x� t�� �p8x~!��pB�R�Y�HB����'�v�"&Ć�ED���8G-B,rҫ�sl�"��̧����~Q�Y3�P�Q��ljj�T���4Ni���u+�<�
���o+��=6����}:�_i��LY2k��^&p6 �٨��|s	�9�,���؂��&Uqo���������":��*�c���ٍ_��K����۫�u,?RѶ1�f�[�	p�,��wh�jO��[k̬�f�ز*��|�ѣ���:�FoQk*�V��K��R�fꎫ5z@%����%�Ȍz��!sxDN�Г)�娂���2yn�4;(�f#Vw��+�)��p��O�����?�q���~��ؽ#���|nCA^mג�{vvm)[��(U��V��#v;0�@9��ߣd��y�ܲ���`QeaQYIQqYa~infu��6�655ni�dj`��	k�W�Ԭ/Ro.V�h��j�fӛ<�Mvb�٨�nR�7+�Cr�v9gX���Q��T��-B���#��='�]�nJ�O��/̲o�ڿ��4�կ�֫�֭��S��]�����F�'9�G)�;����k������ا�)����|�~b�B��=�!��eMdTd�HƉ�1؜�|,\��Q(�fB��q<��*�׮�
6�5�yȿS�5��:�\EyW.,0��?Q�O��Ż:�{�<�)�T���>��LéL��L�f��ń�@S�jz2�N?��O��5��5�h�EY��2�/9HX�@SN�ZZ������A4� (n@��g��LSì��B�D�X��e��j�5��J7L|M� M��M�y��"��˄�PӼ�Ԭ��.�n�-���ͺ>����Lhj�Ed<��Wh�m<c�fQ`4�iF�0�fdi�hO`{/L}b��&���޲�vS_���]��:�kӉ�C'�����~��/�~����G��9�vϖ�G�/~ݘ�s/L�������Ibj��#p���L͑5��5�TlZ�i0�*r*�Ta�[��j�e�
4"BI�?szZFr*'��px
��3���l��i��w[eIwKmWSyGevK�^�c �Jչ��*ߢ�������:�u�wϪi*��1���&Je�Ii�S��	7�j�R���NpRHn*�K���d����p-b�G��R����2#���m��Z�h���%���������ɧ²&ljY�/���5�5Azm��V��Y��_2������x������d��y��������*!�"_�d7��Rr�)�;.2[���JRW2lj`�S�Ԝbs aS����('|���D��8ig��]�#��
���q����H;�c?1>������U�U��Yu����,��G(v�ž���X �B)3!�ej��c��F�D���*
���Ţ��1uU�_����PI}`�nU�ʬ��I�7��9��ڍ��i���(�"���}D�>@s�+�t��ad��:l�6Ih�#:�K��+g͖���L�{�"�Ǌ�i�b�ZA�/��~1f�P%P��v��l��lN��k�fZ��ǫw�M�Y������o>y����?���}���������Es:p��r�Q�7�6��m�@���嘭I*M�D2���(��f���N���FFʔ��)q3�L���Է�cx�� 3�B�Z�US^��I��ͣD L��7J�����dU�IvJR�ԙo�1s�Ը��Ę$f5=a��$@܌�����XvZfT��V\/1MI����X�o�����$$�E�}��$jʔ�S~:cʛ3����N�3�ߞ�0-.1:T���z���o|G,�4J�M+u��aSSl�Z�r+�Ǌ�髰�U8z+�˪��j]}��__S`A�kV!SN�ĩZu��.�hHR��R�R���[hm"�L�W���65a��'4ƾ�&����@A����	���6��A �46��`\\�'H>)DE���"#q���x�\�S���K��ML�ONJf���1S�d�05��æ&TPx�j5�B/�R�L&S~~~]]L�������5��`����i�x|4
�c�9�f?M��N���0�G�hj���?S���9vS�����E����ܧʷ�n�@'�BS�����p��q�15v��l�)�N��
2������(�Db�X233��򚚚�/_�e˖U�V���uuu��e˺��a��s�̙;w.�b�~?\�<t(��~
��?����45�u��F�Ϝ��ɉ��yyVQ���j'^�B=45�Y45�Ѵ0�15m�⹅��"�VM�`�c�l_w�oI�n����T�Sf�d>��mV��T$ 	�Q*�P\FZNjj(\0.�F&��Sjୃ�
�&35|���, eq�i\^:�g	p>�,��#1�_�K0\���
��3�Bf�s��15�|��)ID+��
�k���u�.M�K\�&j��5-9��<S�(_	eMs�\��}�<T�[���պd5.e�[[��z����ju:�VW���M�Rc�15�r�ل��PO;�#�w����|*k�$o�0{!�í���ܰ�P�ZZ�+)Z�dΉQ����g���l���K�o�Z��n��`󚬚kp����R�H�?G�=K�٤ɬ���*Cf�%�Tm�K�6�Ƥ��j�\��h�
�Zo0�?&��h`�g��������4.7��&"x���
�s�� o��r���0��ĩ(��6R���������?�q�㟟~x��+v��4yˋs�J�Z2�ʌ9��`�Hl&�� 4�!�Q�j-�a�L�*&�R�ך�V{��U�s���C�[U�U��5nq�G�䕼���p(��+M�n}�bS�j�D;\�������z3�^�۠�l�������Q9wD��.d��Q�G�V'�)?-E΋�爌�4��Y��W���oӷ�������w����n�~k��U-�3M�YJ�QD�ND|C��%_��/p�c�A~�G?�a_ij �e�15�'|ٌ�)	�@8|��c�,���zL��:�;e#�_7���\��!� l��k.u���K���J���V��^�����Z���M��W{گ9P�E��Ub�gbj�LX��L�b0E���y���ʉ����4���Ź�Ey�		���������T��H��5]�갩	�Όզ�����r��º��诲`g�ƹ�� f�NF�':�pE�}U�sM�sy�	'k"�L�yG���j�k4 Ї�aM������L͆v�8;�+L�G^ij\#��aS3�$0�4��/]�0��֩�:P���fS_ö�m;�3���΍��l;�k��]�	���˯�?�x�ض���۲���?0����v6_i<7\f[��5g�U��97�L�x�U�:�&lj@�_35'7V��\�gE��l{[]���L��)�Ӧ����q��84=����� g��.��a.�8,6���ئQ�g��g�o잷a����e�ަks�mQkފEU{���[xv��S���\��*�Ԯ��0#��1�K���Т�B>2J���5"�G�90���Q��.cj0�B �BI��N�2`�va�G��C'�j��L�Y��#X�I,���/3Nм���A��@S3�'̗,��N֬Η��L9ᐩ9Rl8Yh:4_-p�)t��q��q>�r?��<���xn�m���;j�m��)��oJW)�����\
���,`
ּ05�E�8��9��,.�,���_A��|�:Wp��_�WQ�u\|K ��%���. t4W�0܆��A��lޑ��C))�YiOm��
�����ck�g����዆��3������<�aOq
�|��Ag2�	��w	�9)�GI ���>`�'��P@>��{(~�n��[<�. ���+�6I�P�E°hj��7e�9�H!��Q�k��f�7�_���b5��a���𞊼���ŒO�X'���r�~%ʘ-�WG�7�$G��cF���WΙO�f�S s�M���۴ �,525�%j�q�&���N�V���E�Y��R���TT�6�T�j/i��]Ue/(j��ߺ�ei�Mg�=x��_~��W����?�=x�VˊՖ�Za (�+�V!���$���D?�(��&�z�ˉ���&c�Q��U')�qR*�Bf`����Ĵ$�*���u�WO{Ք[�9d<��(���ee�3��M���15j�Qo���;QoOg'�3Y��I3�f�&MOM����8NB79IM� ���ȏ�e�&�Y�8��!�I@z:��ʏJ�x{f���Ę��TN|JFlbʌ�PvF\��'�'d��0\!ڵR�V��RYz225eV����25h��65���
kw�����S��s�6�{}sKmMy�r�.hSe�TL9a�HfY,f����D�27ئ%%GڙH^mj%#� g�`
7a�3[��Π�G����4�|�	�d�&-%���E9� e�|&� ���<n:���f�ם�����e���''�)�����0'O^RJJ
��O��|�`+���z}NN�����������L�ժR��엙�RB0C�x`�ρ���L��1=n���U����|MM���35EڌbP�g�8Ї�~��(7� �S󯚚 �gjČ�s�lEG�aA����P�W��6�GEBS>�	1QQ�g̜MM8��n6Xz��*45���hj�^��竨����^�~��e�/^�`���K�vuu-Z�h��:mmm0����*++�n�k4�$���r_,p��r�'�j��!�	V�}S�5���3����a2��ɖlrBS��R�Ucbj	��V���������^U�U�1�n�R#I�8!����p
A_���
S~ePCi�ڤ�� 8C�Ԥ>�x� |E $~&�0���k���I�1A�'BHJ��\L*����T���6��o���4�a�CP�$��T�WT�4dM��Вa�\%�0^��zD�I���qɫ��2��ة.t�s�f���v��.���W��2�_aͥ�儧	��|���FF������M"s�i��-1ԮQ����~"w������:[d�Kt���:���Ԯ*[8Z4g����^ڭ�uwi��5������E�٬��kܕjG�+����:�Tm��FZ��Uj�F���V���Y�f�A��c('&zZ\�̨�oO��o�L��;3���$�lƔ�	SމcR�g$����N
���7R��1���������_����އ�o�]9<�t�ZSf����ֶv.*n�W��JΗKS,�ϙ���Vb`zrbTjr�rHb�$�c�����ԟ�,5&V�g�h�EU`��,�2���Ƅ25{$�}�f'�� Z��l���C��
;|��>����*B��15������˓����A�@�b0�iV�¦fm�v]� ~�P��R�)֎ia!�M6�f�Y�ۢ�l�Y�4{T����${��T&8�^P�+���B�94�>�|nW�%��9ֿg��#��_��o��;������dUØ��b���oI��C?Aџ#ȧ���eS�~Hքs�������?�����V�8��B��� �J�.�^E������H|����XLp�k�G��1571&�&|�{S ��aW1��w�d҇
��J�T�z�W��S=�)�j�z��Uy٥>���T�pK�zDk�ԠG�25K}X��X"Y���3��5#b^h �6�X�#'h�t�*�05���Aiw!�[��)Qv�K��]%���\t:K��Ku_�͚_�[Xj\TfꪰC�+=UN@o� o�ո��z �C#/�u����[e��Z��Ϫf��V�@��������Wg��uW��*U]���*eo%@�� z�bj&`y���z@���f,[j���ׁ
���u�������nl�cl�� l�p-�n�����	�-�L�����E��ř0�fG'�i ��w-+ ��g�+��"�f���޵�����Gwn<�{��(A3.�&R�����������3�7��9xrg��#���v��ʡ��{;��^pzG���m'�fASsnt6�Ss~���H3����#��7�����\����% �i&45��c�j�	�0���̑5E�V�l�ڸ8��b[֖Y�M9�p��k
���%�2R��<f�p� �$��J�����-ZY���3�i���wo8�o������s��4��[���Ԟ����9��֞�O����ɳk�j,��kl*JK�3X8g�r�\x�� ���x$�P(
���s� �Ya
������P%�	R�`"6�LKT#Z~���D�J�*uɭv���0]����h@�\��)�iS3&k��r��OaV�IW�I�Kԣ��]A���t��r��z��v��YQ�������+�b��d{o��]�k���Tz],�,��DW��k���H��K��ސ���	�F�A��v���C�sq!y�6q.?����׹�:}��Ϣ����8�".q�WY�m��>&�����\���6*��J��*?��:�ʺ"�<�Y�����겿/���z�5��?����:?,κ%��W��a������	02!�pr��y_(�| ��N���=b <' � ����P|��bA���֋�.�-�AbL�5
�)�nK�{R�#9�L!�H-�LGmP�ɬ�������_}��;����)�N��g��!	g;��Oä>�H���9d��k�E��Yxt�0q.��&K�M�whymj6��hW2�	m[��fC���y���*V�^�╙�EVE�US�婪,m�3����yi��k�^��?и��u�y[��o�ݽw���sϞ=�����/_�����ߞx������+=}���k6d�^��|E����s����(+�
�т"$/����򂠥�\�����l�P���Z-�dbT&�%��f�vЈK��r�GA���l�2Ϫ�q��.J�Gǽ�ִi�̌����;#>96=-��N�YIxZ<��O�F��Q&�&MJ����I��dn\";::��SSy|�a�`�!+0>93*>)���$����8�����������ӣ�x��)S��ߦ�t�(���N�0�&st�-4�ev��Yxv^��Sm�j�H�̍�Z'����}hc&����s"`���E�jXmL�z�l}�.��1w��zZ<]��Eu��#�˕��y�נ0���?woǑ��;`3C�03�F�̶$[�-�df���ْ,YdKf�vh�-��Y���,����S�D���f�����{>?��������3]����R |��0R(���F��S����l����2��z�G8��@\�V@�΁������ ,&`yILHNM�3l.�ާ� �R�#��K8�P���K� $�	��R��l6�N~QQ�헔����\.�N'��`�tq�r�rM@��r�珍��������計��H���!9.����@���A�U�S�g��XA^4���5fN������r�m\ �4H~��w�@���t�2A43�i��In��2��LPS�hf�tF�hf��%_4#G1=SY�|j
����N�H�M��W%,"<2*&!1�&�H�Q+M:�Ѡip����$`|>b��T*�v���X,�!33���☦���@8�������Ԕ���[�v�Ay�\n���<�}�Ɓ;n���وx�bc�##B�"����	V�A�H7`�Na�G}j���i�4k��SW�1iL�7e 3���l�%�������9e��������O������rgC��*�X��e��N�ܠ�*eB1�F`8�' �Rs?'0ȳ��K�� 0LL,�x�A��Q�h���A%�
�K|�A��L@��(DU�S��:�'@�"BD�"����צN"������&A�+r�%.a�[T�T�+�5U~9H�f��2�e�_Z��y�>Y�OQ�U�xE.Y���O*ǡ�۴�.���v�<F�Gc�h��*w��W+����g4K2[dYmҜv 2}� c� �]�9G�5W�;_�� HW�T�%�l�-f���m�KNثVJ|͚����%�������E����ּ9��o��Ө�4|�M�z��6����*Q�=�Y�0���\�P�,&�Qo�[j�����=|���:%|�s�_���s�{q��'L}~RdX,=<�9%:����bx��q^��|hQu�?��/��kw_�q�D��/�<��B8(Y��<c�<on�7?_�p�`CH�r��b"&�N�F�E�E�O�<),$<2$"62*>22><4!|
?)J�O�k�<���"��K�ۅ��ɂ5Y�F��Λ��7��V��%�	祑��$�3%K��˲d+r+s���T�
ԋ�WLu���
+
Faͪ|ź�i���
�@���ۊu;
�{���
{2���#g���[��)c�1�HػŬ]"�}+��K:��t��WĹ��o��*�K��_7
?��~���]��7>�\�߸t���;��76���R8�ӧJ�"�'��8�>�����G�E��P�x�
�	�a@��I�����@�B.��}忊!@ V�|�����/>$�WB�~Z�x�k��.�-���X:��KH��R�V���5����R1h�^G�ہ6�0�w����Q�c�r�p$�8< � ��h��Wq,�!bTWIhHH\��R�M��V��^sK+��W\7*��}&Y�U��Qwg�O�U���~��4�j/5Ԓ4j��i�B?9VйfA���,�_��Lr^�hn�ƒ������\Т<��|�bВ��,.Qw�j����rT�k|#��962�&�w�]�b���!+w)���4m}�az��!�<#�63�Քk��i���}��|ˌkK����5�ڷ�.}ٴ��ӳ��פ-��-����1{ucƒ��R˜rSG�m�t��&����z��:��zyG�hQ�xy�|e�zu�nU�~E�nY�&0TJY���
�8�)�i��Y3�\��z�los1M��ح;������=Ϸk�{�|Ю^���{:ҁ.����WTxpY���e�YV�oy��%�W��ZY�sU�K��7.�ڹ���֥Ч�ܑ]O���C	�xeN�=�����ׯw�r����{���\7pre��%W�/�9J���mc}j ����b4L�te��=ӁzvO�����:��[�)����1�:R�_b�oHjή/����s����s�69;=�N���\Ĕ	1S�b�L�ŦpQ���<�z���2��q5r	#9�kӹM�y3k��\s����C�.��;���ȺK���|i���3N�7xb����Ww�}��zv��W���V�#-|��KI�qP��(��ҩC�9`̕ � �p�@0���$"�Q9A�	�
y8�ࠩt��`%k�1^d�0�\��h����fp!�� ��|q� �%ٔ�fQ���*R�+P���<S_��j��F��A~�ky���3���f���\�ٯ��
ِD2 5A(�/���ӰbHjz1����A��|�2��㉆���M��`��d�u���\�yB�#�w!���*Gz�'���obbʃ�ǽ�"׸��\�M�$�R�Rٽ����iM��������K�k��/6/���ٟ��]�����E�n�0�z%���(��B��^%%�	�P�e@0�a�{� ��B��]��{+��o�a� !ț$y���	��\%x�H���]�ܕ���7T�w���T?��?��~�0�ơ��S���7����&��i�I�	��
?a���NY�g��KNU�Cq�.�f��SZ��V2�M��"y��P�F��X6*��2_�z5�F�*W�*�h�]V�T�MŹͭM����z���ή�W��q����@Gn���۷��{C��#�n���O>~�׿�����/�p��޽������]��:��X0r}�s�g�L?z�h���5k=�V�-s.Xdj�e���՚5��^U*��V��eИ��T� T2T/ǬJܮ�\
�"52�-'�JQ�F�i�d���v�����	�)�!�q����QIqѴ�vj"���Ғ��"9�H�%�c�C��F���@Q��:��@SyLIcR�V$R)Uz�T��4:'.�D�QNe��9�4vb=&61&:!"<fʔ�^�8y┘�X�+#0��T��FI��,4a%6�"56n��Sn��� �������U��u�%���u��jc�Ը5��km�%�)� �1�Dr!��(c�gr��n��� �`M�`�:h T��p���&66�pP�腂�#욂�-���� �`�*����`_�F��xrssA�???���Z�V��W*�����#e�����������H��A��*��P�~-����X�@L$5%z��*5��ʌ�r���5`����ǒ��\����lyK�rV��5O=3[ѐ�����r��pى�1a������%5l��(2�Z�W�D���iR#�J�57��N��b��f2���������JOO���,Xvv6����m6�V���堙!
!��O<x��탤ܵ��&.6::<Hjb�WI�S3�ã�����G���32��,l,�i+Q�-�ί2-�6u�XNs.i�Ϋv�.u4�+3�ߦ�z�L!��$��8�>��">B�A{��!5`_`�j�+ �|���guԀ���ǅ���4cHM ��8A�6F�p�Z$5�U�,�$̶Q��R�[\�U��ir��NW�d(��2MVx$%>y�OY�Uz�Ni�C�����Nm�ǜ���y�V�Ggukm^�3G�꥾YZ�,�I�1S��,�lU�ɲ���´fA�,I�y�u�"��U�;�֒�z�V��%���"W�*c����Q��V�ؘ?_�ݮ͚eɚm��4xM�f�L�o���`s׻��B�£T8T*�R���{2i�z��b��J������	n
3i&Lzn��&�8���!��FM���K��g��Ѐ���#@�	��3�+���g���_�^�a�����II6o�9{�5ye���L��&�j�X�����C&�N�:9$d
t)6:9>!16.1::%>:5.��K��0b��x������m�F�`�	�iB���&+��Ι��6����h���FR�&C�8S�4�"5�r�s�k�T��TK�I�ʗ)�*V*W|j��+��7i7i_�Wo�Sm.�l+�R��"�|žt�NJak���W��+aw������$m+��M�!wD�^��G�-qC�����7K>��m�m���n�o\�߹���6 ��o���t�OT����~*&�Y�0,@jP��,�(8�SPЛ�!�KA�2��@F�Ὂ!��(H��<��Sa�Ll
�?$�'�=.�:*z����8��ڙ�r!%�5��e��U����pK�	o��\ ��#l>h�B(�ג�Q�$	�1$\����䷴�;z�-��Qyä%5Y�K��מ�)��w�I^�
�x��Ԥ��Ƞ�&5A��҉^s2����99���g��d�;�$��@�rd@�
�ˊ+J���tK��%�yE��"sK��&K���zҡX4�Y��td�N��f�9f)x���v%\:T�.H��<���o�L7We�k���9�i���y��|Gs�����Rd�[���-�N�_�i+�7��g�۫,��K�,˚�K���˗�J��HV��W�*WըWU�VV�V��WVQAm�V�V��Vי��g*�q�Mj��Ԍ2���	��յm�h�lH�̱[��v�yw���v�I�=Ϸc�{�|
֌�����Ғ��*>��l,�	����+*v�%5�V7�2Jj.�}���,�_ӓ��?~���/��v��ړ;�_u����c{�v\>���М�����gu�k}&�	o��1$5�su?h�:���i��XԹ��{o�U�+�=m5�4#7%fBؤ	��!f
��\��|�
�p!h����J)G�\B&�E�9�i��꼃;V��;����ׯ�{���w�^z�a�;�v>�~��[G?|p��;�~~��_޼�����s:�t%Z̆҈�hv|<���ƥH" �2AR�g�(O�R�F�b">FrP��FRh"&ML�����!~"�T�h��z������/��	Hj���Z�C<���85�s���l�l���|��\��\ͅCo��Z��f��a������f�Y��j^����:`1�˥CI�Px�${p�2��U��@XC����ԀL���+M�����!LvS�}����u>����ARq����+J��a��\C7Q�ˤ�)�C���*����jD�L��� E��+J������?,�����޾��E�X�~�� �M�_Cj��S�2� 5o��@ca�5H1��.����!���.2�n{��zk�[�&�S1k(���\���r�\�R��Z�c��S��s��7N��f�o}�,һBf/�'�0�|R�V�Ǎ�Sv�i��[��7��:���v����H�$��Yv��`�(���oHj�i9�z^�UX�V�yueY��5�֯ܰ{��ӧ�����?pu���/�����[���|uh�@��/���'��ͯ���o����^����￹����K�tw��o�zu��`���%�G_k��q�b��s���4;Y�mg����[�T�Z����.1�i�V��d��t:�^M�ՄCC85�[M���(p�R���f蕙F��b�I�������0!d��Ȱ���D^R/!����%&	ѱXX4?�.�g�c���T<2�C�bR�	l.�Hf(�p�r3s˴FJHQB�G�M�f�Ja�i���0jV��а����)SB�B��b�9���3�YZ��&/�I��x�-��˝�r;�1�	��`5�;��� �%5p^��u� ����\G�mq�k�tg[����R�o*�0�4��$+0��ĥ�/%5�]@�Z��Kصǂ@b` ���
���W	�� �僤X�s`�Ԍ�&$�pt�˵Z���酅�pܓ�`���J�Tj�� �g��`�g������ZR<�NU������sķDj��4�
���! ��3IMK��9W֜�h�S�.��䪚�ԕ>u�Uj�r��Hj�#bc�)P����`1q���J�H&B�A�����0\p`���n��n(n1��ؤ�h�F�-`&�	��F"����@P'�>W��~���w�5Hj(�'
�D��SS� O�t/?Hj�k����@ff��YXKٚKj/Uϫ�AFCa�Z�鮥���U��R{}��ܯ�si}�U'Ӫ�1)8�����&�|p��:�	^pA����Le��=40Pj
��Xk��FD�"��5�=K�"�N"��~#�c#����--�� �����'����++���P��46Q�M�m����\�%'ݛ����gڼ�V_��W�M�V�MS��)ӧ+�)e6)3f���9���&��@x���ܹ�����]���-b�4�- �[*3��ic^����\0W��,�L�8�4�iW-��]o�5X}��4���d+Wk�dr�Ji�h,J�V*�K��B��kM�B&��,i����9�^�0a�C&�2��)S��:)4:$"��и�ѩ!q�)14 �x>,���٥=�/��k����˦�r���x"�/li��n�֒�Z��!����tڔ��ᡑ�Q��S_x~BD�T�ںz*#%�roO�I~b� %�1�L�BR��4!3-��Y�-��fe�jI��
�Z�XV�\^�\Q�Z]�^3��X�R��Bͦ<��\��<����"��B���n�p�٦a�TP��IY���}"�m7I�AҀ�a)=b�-9~G#����I��R�u��Y��C�������^�/�ڀC���.����p�mQQ�F!�XN除�={���.��y_�U����(���Ӏd4Л�5}��� �y����|�0x"�h�D{��@��!��+|�&�*�s2"����� ｌ���ҿ�v���ޖ�n��w"К��A���AW�e��OH͐T4����(!��iV�0�����e���.������G��{|��>�Z/�܇-����б�� 5�d[֨@: !��J�2%@��eI�S�4��t+*� �JL��3r�Ӳ�E.�W�[�\�5�0��+E�Z�aЁ�B�I�2�Y@�f��J4_=< j̾� ��izQ�^��%)�V���p�2�_���ayF(׈��b��6S1�ܸ�ѱ�ٱ�ɴd�fE�ve�zE�jE�bE�ry�fE�vE��\ݐԌ�5A4�U��S�h ��,ft��WMPp+d1O����|�>5p$��z����?}p��ʙ��G�yiN���/�������|`6�w�S�LL�MI͹%'�]�YbS��y٭�&��ŧOa&�2ScPS�Qc�yL.�AD�@B�%"�\.W�
�����X��mk��xt�;�޹�����۽��l�|l�͞]��֎�_�r�gV�}i��#���C-yK�L�f�_�&p�P8L�C�Hd��90�	�ZBG��
y|!p1��Gi,$�FҒIђ����4<�\������e�`x����汰E�dP��(-ɤ�LR�>K�#W�'Oq$O}2Ws>[9�0�a��a{5��Va�;�y���0�^�o�i�3jd�5�э�]r��i�'xM��	d��|,HjzQP*��#�������yOa�.�^��e�3b�%�y��P����!T5������U���"�(2�^g��s�׸�+,�
��!W��t}V[�떦�7�����7-�{��W��ys�6�h�������iݣ���Ra$5@����	��|��4��a���*�%��I��� Q���_p���;2�e��B�}��G:ŧf�/��ߺ,���~�f��K�0��� I'��a9rL'8e����/:UARsأX�d��ѳ��6I�,qr����|+>5�v���_unu��P��_�`����w=|�����.]��ٹ{dx�����6_����s����n����w���O���@o���{~������/��8��kzwW]Wg�����+�Wg4_��ze��g`v �@^�W��#�[O�n=|���Me�;rg�pV�2��4�ͮ7�F�Ȭ�դC���(�4�S�}j�_�L�kӌF!&f0����ɓ�'L��|dHXrT;<��	��E�cqDH�BgB$��X�s1�	�	���"@B�"R�T�Tk�,�i)����
��@=1<iJTjx#&�O��%3�c���EO�:ir�)!��$D�3Si�a XYA�K[�T[�"Rf�W8�o�SӚ/�n5�Ŋ��*j��Ұ��
I������Zai*����Ӎ�N��8Jj��V��4��}H
Ռ1�jg��4����A� ��=L��5��			�<(B� �a�=O����z�~���2��:�N�T
�BP!(?�����lz&��2t�"@O	c���4���Sc�&���SSe�f"{�|�>5-yrJ���<U[��+��,���"�-L����B@EG�F���'$1,��H\Lb"��C�����t@"�(
p����sss������>2a0Ee2jvv�$AP|f�c �.������ ��kARC�����|j�s?�85��5!�2����LJ-�x�Ԁ;��i���
{K�uZ��,M���x�J�V�UH�B\A���J!9\����H���%z��2�������L�C`�5G8)���%�
3��v;̀g[yvq�ST�H��<M^�&��� �)�K��"���-�0�S�k�X��Q�E�iUd:�^�?͛��r�s��<{z��S��V�|5*_-��W�Io��M�kIG��]'Ik�����rGQ;O�����3������msf���������ٺ�F��Z`)�e�R��Te-�;�͞z����1Z+��2�.S!w�6��(��d�R*���`��$f���u 8'��=5,6,<6rRdĄIS&�8��)Q�"�&��_��?�:!2qBD��	�)�l��i�,\�}��m�r�ff�4���]Y�
�E(P46�^�nKIe�D�'d���|&�G�ŅDD�o!�I���sS��L<Q|��e!l:'5��$E���*,_�W��z+�`�LH��?����,L-�/ɠ`͗�&W��P�8�i�����y�X�%@j6�*��f��@�j_�t���a�mW3��;%t�Ԉ{��D�.,uA�+d0d�]��e�䦒0�Iư�sO������O��W�3������T�u���6��e�#X:����>�H?�>��@���PAj�M>��!��qj�P5ȗz�?Dx�c�ว������ 	
֠�C��S^�&�������`4P����l���6�K��<��P�_�[;���*J�������Z��\qW(��;����f����I͠�����j�-��AMM�dQ���i�Q�e�^t��z�|�>ɶ4�:	I�B/�4�$�����y���m���Q�t@�9�@"��� ���ϒ�͒w�閗�WT�����3�5^e��K�j4I����Q
�R�!d%�7��$`��� �
���j��!�Z���u�e���O��R�$J�D��c��$�*b9�\��)�4%j�Zũ�n�_>�ڶ�%mu�{y�ym�mM�qe�vE�jY�hE�&Hj��5�i<��'\i �
��'I�3a�wIj�s��'���$���g?�9pv�������k�x`qס]��AAR�s�m<R�5��2����Ԇ<�' MPO�{
���C+�/���3s��Җ
�Gǒ�r!�È%P�G�y�� !$�X*��F�Z��P�D��FLIw��J2f7�]:���o��~y��H�����]2���ȥ����xk`盝�ܻ���O?z�o�t�<��J�gH�JF��h.������@0I��QQ\��&�,*�0�K�y���Xh*�HM�"�	S�̐,QL����f���!����
�@p�e��$5+sDTP��/�&K�6K�%G�;W~$O}"G}>C��;  ��IDAT�����7�m�秿]��^I>Л�9w��!��O��Qc��h�����^d�/�X Ճ�`��\i������<�2���	ٰHu]��!Ձ�Xs]��o:�7|�^�Hf��k��~��W��#��:!��f �o���l�51�����*��3��������������犎���xtl����n:==�Ms>S���@F3��2���eB�� Ǣ0�zuQ�� ���b�ah�$P�<PB誀tK�ߓd�����䟘u�;̿s����1���S�^|_E^&����'D�#�q5q�(>e���ɻ<�n��G}*S�N�oCcfa1��QR�����P��|S��Z%�Zͮ1�Y�GW_��b��#��8��`����5g�,?{f�`�����{�w]j?~����m��>��{�Ӈ����G��ѣ�?�d���{�Z�/N�X�y���R��SU=��zj._����ꪽp��������9:}���M��,�ikv�V�}��j���b��4*1��)�v9ϥ@<Jԫ$|*�O-I��|�G���r�+����ь���/N�	g�$a�#X�"��x����	�D��x��qĄHބrb�d*C��&
�)b[��B	M����ڶ��&[f�Ԕ��_���E��O�F'�8�q�����'��8q�IS&O�2ejld-)��R�FKV��_!5.�7�������&�V 5u�%�vН�w,��Sgo.35���M%�l��mT��R9�l��V����p_
Ռ�5���V��?�v�4j����X͓��9(+	�������f�9�ݮ��@wT.(����	T�LR3y���pzr$5ӫB���S3ޠ��|j�Ij��4��I�-� ��#:6&ܫ��T:��e��E) �I�x�Ql�@����������l���h<@^	p��u�)@*�<��
��	9x��஁[nQ82|<��7^1��r�i�C���Fj���\��<!d�_Cj������R���hV�5�BL�(FP5��.�8�����"��� �j\`��=��2� ���3�`M ��XR#�S���AxR~��L�*�>=�i�:�Eny�_Y��,�)ʽ�2���-.s��rԛ�)�s�l�� ��4��-�I�0R���:�Bk����E��4 B�'��>�g�̐��Qc>b���r��l�:��瑺l��#��9 �V2��mCI����fCZ��Y�ʬE`)�*,E*[��Ye��ټ�g��^�p����r�M"ҋ�r��j�jJ�J�Sjm&�L*��T6���MIb�E%FF&DN�	.4d���&O}."nr=���q�>	!l4�GDc�XB��*�[��r��Ҷ�-w�&-���PB^]7c��M�3Z.*��<^T*�JN����>���$����sa\&3!�5E�m"��*�@�BR3�2Jj�Lܯ!5@���K3�+��@Rj�&5p�Ӧ��Ŧ�|ͮB���l�n�x��	����0�,y��M�OҎH�g$Tl��hD7e�K�ASnȸ��%f�?��>��>v�fU�ܦ��K����G�q�Ԙ���%����"��S�O�;ȗ�>J�-��5����^Ġ��5O{ӌ%5`�}�c߀��;L�.q����0��8�J�h��G�;�}����j�<�����D���$�m��!$5��5�dD)�����ˡ[�u�r�(�5H�M�K6�Y���Gv�'��mL���}h���M}jƂ���t|v���*%2 !P[��-]Ҟ!��)j�R����/4-*�-,s�Z�5�vY�Qh�S��M2�<���J	�a#��-���M��$E�W+!�F��V"�L��@(=�-�͊�e'ıb��	Q��h~B$+:��ʊ��
�Ċx�5�5�L�$���q~5oZ�fA�kE�oe�k]�km�m�4ӊjͲ
��rX.��,��=k��5_�S�H���;&5߹O��&�'I�/>}����K��Ooٱ��입]IM��v8�� ���<Ӝ\����ZWtr]Q���gX[�Zi�x:]-�"�d!����NMHa�0&H�R�/�\J |������wk���*.��ڍ���?�z��[߼y���C����\���=?����?���ˑ���sju�n���+LI#:f� 1N�`���S���Ho� �a�дx�P���Pq,8,Jl���,>��at6Fc�Idb�<9̆D�hh3���t�������	*k�%daԢLJ�3(�����R�3�k3��3��rd�OM���_��S��n�m�禽�������r3_IO��^1h.+d����P7��ù�b�g2�x<�
��	 J�y��<���C���!R>"V��5Ce&�D��:�M�����wg�9�����o7��RX9bI���� _r"d?�"�uD<�1�~��@y��U�wܾOKJ~�0���M��z�iգ���l�qN� ����|*<���e*H�IT���b@` P!�	+Hj(`�2
k���*ƿF�#B|X���%��J��R���}��c��N˿{l�q������C����=��'�Gż*�^IM�Ww9M{ާ��o�l�砱mh�ar` T�,9c�|��RF/W�*͒J���${��#��l:�o��S�Ο]v���ӧV�tm�[�׻�ʕg�,8ur�ȵ����߾�飿���~���?~wi��󧦝;Uu�tٹ3e�.V�ԏL���)�x�������ܶ�`���mۋ׭���j�7��2�n�ɬ�j�Z%aP�f9j��mNӤ�%>�ԧ�{TԈ�d��ɱ��HzhH��)�S�ّ��)q��dI8S�Մsu@�)�е�ls1j+Gl%|k1b)d�sh�4�!�Y:�`�
Oy�.�N�Q-us��0�04�M��T"��'��D��:5,l����Hzb"ΠY�,��̦���'�����j���0k,��s.��s��Ӝs��3JE��Si�!ۮ���|�,��V��#���c %9Y&�hF����O81Pl�8M���KX��`+�t>!��Z�΀i�Z�A]z�(Iѝ��4�����<��L�:52",%!a&��4���U�9z��򩩶��4���z��g�~�H�Ib$�$=4sS�"��#�#bb� ���\6Ex�M���� ��n�J�r8�^x�޴���Z��D`�H��nx0�K���x�@��	P,Ax�;»n$5��E����SS�!�=�t/��\��Y��l���������O@�~�>5�Y��O�Y#���R�(�t��u�X�� 2�0x��=k �<�`���O��P���p��h�Nİ*xn�i�ei�R���+/s�J\"(p�)��h��!�!s,�� ��i*1J \p'S��	��8z��2�	LI[��Q$q�I|U*�O%�t��&���x���F�)�.,��g)p�$�ʢ��e�e�����u�b�!K�ː���<�� $@�̘�6�meF{��Zb4��y*�WH�	T����Z�ܠ��j��(�Z��d�0��I�1a�!S����bTĤ��p3�G��d��n0�4Yv�$3qz�6'X�g�T,Y���\0wAVk�8#�W����:�9��rMqc���1��"��F���'G ��w�Bi0�Tj�H�!�Tz\8+6T�N�ʑ?_�T�:QoƦ�x�M�3���lR��BR�$C���[͊��*B��"��B��B��"��B����B�&��Un�V����V��Wjޟ�ݛ.�� ��[��*�)Ejv���������E��H����Q���):@Ё�i��=�˱�n�ȭ�Ȫ��"��]�{���>�.㟝�/����?W�?�?b@㑚�0"�wpJo��DQ�7z�RpX�5c1�3I�k�#���'.v���M���CLΞ'�U*m��h���~T\���РE�%5I�oc�Ӑ���f@L��VH���#j�����
U3d���%=FI�Uv�!;��Jw�ě�>|�Y�F���$5�i�7S�3I�if��m钶L9P{��R�fN�yn�mN�}v��!�Pf�g�����HY�$#	�'b�����L�E����j�`J3)��MO���G�L��)��Iѡ���#�#"�"�R��A�͈�a�Ɛt��II@O�����h$.
��f�Of�MFb�*9q��.C=�ܾ�޵j�we�}E�iy�~Y�(�Y������)F3����'G?=Q,k�cR��Ԝ3�i��$5��^���]��l}iq��]�wt��uh^���T8�m]�Z;�R��;����4�|�9�.�i�\�a[�m5�O߻�bN���'���r!]��eb���l5�l2���
�\.�~����UHp�Seq��������͛oݽ�ƍ�oݾ�p���K;�^��ʕ�������o^Z��o�X�`�����j=�O'�VMAK��r>_��B� ��ℿ�@^I�ņS��D` ����$8,��Ƙ�����"R��1*f�O�\gC�d�:r��y�IM���Hoa�ϓ�5����RHjN�����A����J���t�ki�n�m�e@�/��E.���`j��N6�"�u��̽M	�C4]iF�M�| ӌ��T8��	�)$WY7&>�	o���
��>����?۴�[�|�a����_qۖ>$���AD��ï�~z�C^c�Cl���1�2�
n�T�s8>*,|�lѣ�/=Z�����}���	}��IMp���|�=S�����h`B��� �B����E!��o�� �B�ǰ��P���aI@R���)�nI�{R�U����C��s��?��߻u_����>��~�4ܔ���Y!礈wF-8o���+����\��{_���Ľ�$����F���n5O��%�hZ�%RT!��(@�NP�3�(�Y�|��7ܷ���ݗ��m�6�exh���Kׯ��:�����v����Go���?|��?}�?o=�˹����Z���W��{z{���^뫻9Tw�ji������]�;y6���]{r��(ڲ�tӦ�ys5eE�l�!7��2�
�F�U�jQ ��n�󨙹UX�Z�����J�RH�r��Mr���Xv|4'2��MD�Q<C����f���4]N�>�i+B�5��ҼY��vQv3�Ʋ�ǩ�CI�2��^ݑ1suv�o�s�,iZj)`�=)K_Õ' J�@��LB�Y �"�������G�G$DE�R���C�fj�B��+���o�S�VI�c���j$5k����i��Ֆ�"��BSu������������V��g�@4��4�G�]kh�f��$''�s�k�@�[aa�v$5��@y���j�N�����n�ժP(@O�e�{1<����ƒ`���	��
�a��*4C���|j��M�̷Bj�Ƨf����~m�I�#R	Z4;1�k����C�>5)�T������x<j�����S�!G?�l6p;|>������@hg4``G�T���A� ����VP-L��	b���� �e�Ԁ�ϧ��CL��&��4#�h��85��cR3+OI;|���s*��ֺ���~�(%b�WG?!(���#5�DQx�6p���4���x���f�`�� ACK�Q#� (
� <�&�hJ]/f��\��ȴI=�R��ԫ,uI��b���!,uR>5��8�A����&�"J3��rTȣӒ��j!��O��0)⅐�I!	�C�D��D����	܈$^T2���%aS�I����/D�^gL�?9��BL���/�YP�l���b��XP�	�_d�
���#M��N��B�K(�I�W�X"�E les�(��H�R�F&��t�V�M&��L���&EGђ��é҈�N�Ë;��<qa�����4��8�P7,����/Y6m˶�����^[�lE�y���ܺ�_�Xױx멳�_�{����*�-�3�SSi+-4�d��<*�Me1�g������(���N��i�:���@2�B�ʈ�Y�z2�ěf�L3�m��H�"���V�"G�,O�$�ɉ�����)��6�)7�(6f+��w���e�w�%[��-o���S��%g�3v��;y��YQ�Q����.2��l��U��d�):"�ސ�߰�>�q|���Y��#��#��gVů�?���Y���
��X�@��Ɛ�wj�'8���8Ի�wHJ��5���`�WPj$TЛ&ƒ��G�cT a�*�0y����np�.���I�њ��V-�����b3�7�^�j�$70�.y<��5ԯ��RD� ��$�B�\�K�U�!�pX#�iP�0)G�A��� ��/�dg��#��䥴Ǥ����>5O���U�k���2���	%��!��)��)���hˢ��l��<۬<Ws�cz��ԡJWf����E�$;U���L:?5����c0P���� �h���$FJ"=9����r�*H$�E�GS??�%5�ELBRtPrl"-6�G�M�D�n�%$0�"�CC�NI�:���Jy�5UɌ�+�ui������e���u��5�պ���e�E�����_���@O ��ק�E[����|�>5��IR����>����Ãg�m�>�c^0N$5�����g� ���b��!5���=Ck
.m�>������m�6y��iv�L���*�H)�\����J��Ke�y!�W��	ѡiCE��i}����k�=��kC|���n�������7Ϯxpq��s+o�ӿ��LG��׶*o����K�^��e�*�4)�-A11)�
E2�$ �y&�-!�ˆ>58�}jp�d�IZ�85Nώ˔3fx�K
%s�yR��g����@��}j:2�fPZ�Ni<��M~rw��h��D��Oyɩ����{�\֗��;&�U��W"�@�g��s,�%��C񚱤�3����ǣ�m��^.�
�c�@Ä�.¤W0q&�!�=��Hv;7�a]�+��v���=�ũ�<z��/m{wZ�Ì��j�����D/�����3�!~���I��Jb_Jf^f�n��o��?/+�ˬ��5�]UJ��E��0أ��Θ�4��i�Ij`>�4�Ѽ��@7�(d4PARC)@j�_^������ԌH�tCJ����U��m��C��.�����4���[��o��i�)F/�i]b�9�uZ��n�@��fiڽꌛU�e��fQ�Ώ�/xLjd�o��4h8URz��Ua��̳*W/��d��/-߳k��S��v\����k�K/]X�׷������y���?|�߾��<zt�O�=��kK����v��m��U}�\مŗ/�tS���Bι�g/��Pt�LށCy�w�n�Y�m[��y��L��%5&��1*	���s?A��4�ȯ���R�R�Km2�MiV�zW��5��V���Rd�(2��raf�(g&�>��>M\8K[�XY��Ҹ�׾3s��������j��Z^4W�7�>me��c�7�J��^�5wW��2�>'U�IX�+��(��Fw�Փ�3:H���B��c��T	��*"W+�Ѡ��Y�K��,��ȧ.� �免.�s-��/�st�9�*���i��,S�G�i�8�
�qQ�����S�w�_Cj@>8P�~�'�Jj`a`�� u����'@j@�S�������,��c0@�tP��AП�8�R���#5��
v��x%ƴ��
�+�ߖOx���f,��VH����P�tgKfdA��XR�e�q�WHMh�����'��}j�l�쏍�x�0���^��Z�>�/;;xV(�@b� @I���}A�`GXU�J�2�4�T���;p�-w��D�������|�XR33�l�%5�rɱ���=��8��yMG�c�tϜJGk�mzΗ�a�����f4�0��}�&�XF^����4ip�Q�1���z@�po��
�	J��5(_Fr$G!`���c_�Fa�C^��{TE.Y�]Td>k���B;Y`#�-d�Y�ӑz1c&��G�DEGFŅF%�D$Nx!�B'N��2%&$<!<*9"���aL�L������	/�Mx!v�ĸ	�'L�x~R��c�&L����[YP2�d�P��B�%�DFc	b�!Q�x:��F��#��1�Db�09E��,�%Rf2�O�&�19�7	��T�&�JL ��bT�9�,v*�p0_*�:lւBwU���ZYPj�٢ihPM��ml�55Yf��_�f�C�۷�8xp��nݚw���K��>�~�ؚ��ݸ~���o�4����,>yd�C�W5���~����&[i�9/�Y��Q^4cN�?�G�\Fj�+��,v���%���Uz��L��z#����gH��t�XR�4W�$��5���+���k���ks�sr��/e)��i����U8���v;�[�Kj�V5w���W��+an��n�D�E�G��^0���-��U��JpS�ޖ�w��j�=���%��猒�O��Ϭ��:u_xL�Z��0��a��M�{��r��B�� ��H�lR�B�{$�w��#5�Yf,���4 t��e��+z��?9K�]v�O%ү���Q|ۄ	�l֣E-����9�ܷǒ�����t�R�/ 5��ʄ���z9k��a���1˻,�sN�1�l�O�%M��G,� �]� ��.HМ�'H͓�fV�hv��-Gߚk�U���癞���rLJ�W�BF2?1g�6��)��T:[q�Zt�h����S�8,6�rR��?1	$@~J���HM�S���ƥ�cSi�I�D:h��8����hNB'.�Ǎ�a���L��<i7r����g6d�V��8���!�YV�Y\&_X"_Z���V3>�ק&(k�!��[a��[�wOj�s�� �O�Ej>�ɛ��/�t�>����Ч��м�����}ao+P׾��F?��i��� M��:��5@��+/m��8����[�.m/����7 5Ox�yH�Z�wrM��9�We]�}nK���e���n����-��̖ᒺ�R�Nl5i�$F���D�|��$��4�@�C��#��H��;*��+6�;��W�����O�z���������{������v�Y\xvU���U�W�_T�����VJ�~��%�n�⨖@��B"U��R%���A
0	}��f�O�f`,:�f�O,�`�iln���LҒ�7C�׸��K����Xp��z�ьjA� ��ġO�S�,����Y�`����ҝ��}�#�3>e�G=���t��4׵�k
��L�/�^�/�E��r/���s4��TH ���L
�t�9]n�\Fʭ����𮰐Av�+����4�&��6J�=�lXg�����U_��������_�;�_=]�}����|��aPc����^6v1�~)�ٓ��KA�(P�N�\�O=�4���*T�[���>=CK�f3����S�!��)z �<P㛞�3���@wy8P��u�G	�������2{y��}��x�"dH̿&An��;r�
U�V�������n�\�?:uM�����#��LpM�]��g�JA�E9�7�*I{P�{�*}���[�<��n�s�p�fq)��9RF�$�YN�)gĂ��`5�9�t5h��U�dB���@u
X��F-�B�Z"e��e3s��y�5oܺa����N��z���+�;������0�֫C{{w\�z������;���?������gz�����9��{�f_��?0k�j]_OUWYϥ���rO��9q���鲓gg\�\�w_��-5۶�/]�)-���Y>��`0��jR��
Ԧ�jԥB�>5~�ا�x�b�\l��b�ӈ1�\�ҙ
����%��W���͚��h�ђ�'�6���ziڮ��]�����k�O�2��y���>rs�ξʍ���)Yu�igO���;zJVs�l2U/!��|k1�T(t�볧��[�Lo_�[V��Wn���d�i(�)B�R�Lr�N�+4
��R���)�2�l�Jk@?�Ήջ�:7��=��TxQ�s���H1�4�\���:����꜋�Q�[���UYڲt]�K�5ȍ2�Äl�#��SCa������
��8�c8�3��F�{����a��`�
�ؐ� K
�gƠXl�@W`�Cj��^:0��G�j����^���v[,�L�l�%�y8`�#��@1��XTdxr|��(G�p�f��2A4��	��WY)F�LA@�DB�Q���33]Ԝ!��)l�$ƈ"5��"��9Җ\es�bv�v^�iN��9WW���0
�x���I�ũ_ �b�b��c��i:�7:���a�� ��b���%0�A;\p��'��	�K�H$`+ExNF9��� d�>T�+�j�Qƹ_!�aSb�'�ƅa����ף�v��Eָ���0N�(�IЧ�	R�4�� 4��>�m��|cy�2�!˴*�F�I-VʄR�@,P����@מC�,�O�0�H�#50�@�~�
$@&�\FP�^:xݨO���	5��&�B1!J�/.A	)F�pBF�%8[�Ѐ�8C+��T�G'̱�������))uJJ�+Yh%�$P�� *���V<�B�Z�^-ns$��JINJ����܄I/<7���L~14djddD\LLJ|<=:��:5<��)�^���\8%*D��	/���s/�թ���H��֖BG��i��nL<#<*yrH싓�&L��09��ɱ��OI	KcD�ѣ�ia���^�L�H�2�\��4"�Q)SJ*��	tr�RB�ĘLF�"Ta�X2�i���:ma���:k��Y'N��??�����{����w7޺�|`���[r���w���ƾ7^�~�ƪ��{�.�=7�쑎sGZ�yie��v�ں�bnkM�Қ����ip��^�$]Md)���DԘ�:3��̫�p��8@㑚ř8�S0N��l��,��l���\��\��<��\��\К,��t��t�KY��y���ݹڽ^��p�٤`�$en�0��Rw�)뒧leD�aD�G�FGt��]��<�׌�������j�}��u��}��,�^�Gn݇6�&���������z������W����?�_�D���)��G)L���G��Ű�p|<���E����w�·��o	�7I� �	
�h�`��C�p�{z�����osy@AG�`>�t��H��ٷ����c	q�WW��������J_uX����*�-RH���}dsX��9@�Pa1�A�ׅ��pX(���<&5T�!�/U��R
��D#j�u��V6��i%Wt�^���C~�#��ot+��R/������ǒ����LJ���h�j��2'����TP¶lYK��5��4��Z��Y����cc��:�U�0��2�Sc\)�%b1QZ
BKE���g��,x�����f�Yt&#�NK���U�	r��f&��7H*=��G��NI�KMM�'ǥ�ƥ2�h�D�N�,�`,6�T&McEE�""�ё����R_���G�D�Y�م�y��y��%�ŕ�e5���j�S� 7��D� �	"�P�D�	��n��d��������6��+��v��v�y!�K��{�������s�^�0�´�3�-�ϧ����KJ�-��wY��Ż���\Q�iQ�e[���^�zh�ғ�ן޿����gS�g��� �쑽0 M0���@��'ʏ-	4�g|����=Gz�o<�m����-�:4�ҁ9��]��zq5E��ĩ����؛���@Xsj�觱t�
:Ԝ\�{ru��%�^�8��t���e�ӊL�^E����&-�p��� �3`P�@�D@���c�����T�C��;���6���Ԟw>����ׯ��HM��C�kv���ޞ~tii�Ɔ��3�V��ZѴ�"m�K�/��0����I\%)$R�L��+�R�T(���AR�a0!���
������8��2�ARC�&qN��vJ:
�K�����Y��&�' �c�b��!5С���Y��9��Y���c~�9��۩�bU]5���~15�S/�]ƈ.���gs;��N6g,����<��5й�x���2�������A5^i�'��t�r�p�u�P�#R�uzߪ��p��_���Ӈ�:��כ��=���C�����CG�2�#��vKn��J{��>&�7�ןJa��'�ۙ@?��Kg_��{2�-���ǽDK�Ӯ��7�Ϙ�i<R3��G�4ߔ���x=\�Ӥ��a�e������v��ۯ��?:r���n�����^��LxKJ�H��T��͊^��Z��F��Z��r��'�~ګ۪A;��ٜ�6<�M��,N�%g�(�
V@l��J�?$5pbP�FF+&���uY��ܐ����y���k�nY�gϺ�G7�9��¥�.�8wv���s�\q��ޫ��^}��+Ͻ���/?��ѣ������_[~�����9�.�uu�<��̹�˝��+.�):u"��Ѽ��)9x����ҝ�J6n�X�6�c���T��a����I�ш��S�{�ƣ��2�Li���
�Ü��3��zQY󆪎}��O/>qU��7�h������M7>x��O�r޹7f�~���k�_�s浶g�9}��YGn��3��9��i�y�vKW�K��V�+��8���-�k\Zּ��meìE�g�),*�k�KpXR��&x6�'Cr��"���B[�+���+���ʧ��z՝����Ӑ��)�l���4_CjT�;*�k���]�k�-%��<Ej��y�W'7K%
��P�>��O���/ܗ�� ��ɳn���� ��a�f���<4�c'|{��(v��j�YYY�Ԙ�f��X�	��}������?t���&).�GO��i	קƾ=R���<�' MPA��'<h��f,���I��y,��|j��se-�J��B]��Ԥ�2�B-�
���Y��bb�s?Q�t��1�I��Bx# 7�b��P����0l,�IOO���	RD��?&5�a!��AR�1�Jj���ƒ���x>5cIͼJ#�\ 5s*3�Ui����J��R!!�$N�|ׇͥ~:b��)�	`Ӏ���`1`A^�3��z�KG}��e���3�;~��b��Ą���$ʐ�l��oV�N�0�*ͱJ�m�";�i��+I}��GIM��(������~=i��dc��&&DDDM�*,z�S�<?i��C&��O���ZB|\JlLRTTRXXܤ�1/L�|��	�G�������C��BIR.��t>��KI�$&2ccS#"BBb�L�z~r8���&N��4%nꔄЩ��S�"�$L}."�����x~
C��H\/R�D��:�$�"�Ԩ�2��b����T�769�5�gϯݶ�����3�Z/��u��ܞ��C@ ��j�@Ԣ�~JC=[^������Xy�����v.�|��Ȏ�om}yh���U=g7�_��{~�٣��[�ʫ��s��^S�MS`���FA���5~Ij�m���'I�\$5p�Y2kƒ�e9��9�U9�59r�������5~�z�ds�b[�z{�fw�f�K��,�M2�f	s���C��M�neG���`Ee�t��z�[v����7�����W��j��������OҌ��|jQ�֭�[��Q��Q������_�U���!~��?O���S�Լ�0A��S�H�N �@Ra�ӌꙤ�}�Q�i���e�Ij��*�7B��2��xl����
�����Ƕ�ˋ^�8X���u�!}#@(ئ����,aDa�>�����D�*�u���F��I�V�o�w;g���f�ʃQ�&�X��Ri�@}È�O1�'IͨOM�tf��9Sٚ�m�14g�2u��4Cy���iM7iJ�N�*���"XL�NC�>3���C�|���x��p���"�Fg��@t���)�t��&��KMb&'��,z3%6%9&��59���388�E����4eJҤ�Sّ��S�O|a3�J����l�����"UG�rI�fi��	@�8���5���f} �Ϳ@j��URCa���& kJw-/߲�d�⊭����m=�e�=��rf�����%/O�R���}�v�+�zNl:��#�S�yp�s.��5��z����1�����P����'5�E~���LputH���#�sOo�<��z粒e���Ƃme�7?�e��9�T�����UI2���AC�"5B�2H����*���Z��uz�_y8|�� �@L���7o]8��ʉ��fell�}fMݕmm���.��qjQ���.}��,η㘍��B!$5J�H&
̨��
���?k�*�Rǧ�HM2���r����%R3�O��,PС�ҽ=G�'[v0K~<]�/X$]Z�e�������<>5���t��K<���8��v2Xi��)4��t �s����Y
�p�AO��'��ar���&r�E�p׸�n�����R�#W����Q��nX��3~q���2�������ȣ�_}���>w������Ի���0Y/���B��� ��D��T~o�+�q1.�'�	_}f���bq���<�i��� �	��;\��n/�u����8W^���'�H�Э��)F���)�Zu��,�p�����١�O���i���7��2ѐ�	�h��Fy�]ݗa�Z�(�_�4vf�ϥ��D+ȔvNt+/��Hl$}SR�i�:��2U��J�F�N�ɪ���L�ܦ�M׮X�nՖmk��x����W9�h��y���t�ҊG�<��rO�����;�~��7�]���/��>r��ȑ�]ݫ���]��?������ړ'�.ڷ�x�����+v�+ݾ�|���uk�/̚5�[Wi-�1���NʧF�S�5s?yU�R�T��Z{����bV뜍�+��;3{kO��-n��|mι7g�y������ZOݛq�vӱ��_�~�^Ñ{3�ޟy�Aӑ�M�n�=���ӯ��zy֑[3�7����j���%Gr��ə��x��ʅ��l����a��ֵً�[^]3�as�q\�c+�UF��X�/0��"8�S��[jg��SS���x�u>��t���=G=�GjV�V9U��y:��s��M�ƺ]e��ħ˶��:�A*����� �q�~=�ojpG_��$��3���V���O�huϲ ��ҭva&�
�-xh�ǆl�3�	,��b�+l<Rs@I�;8�N�����z�p�n�\:����Q�;4�
6��A���:����pi	R^�Y��\�˧f�0��s�XG� ���!��=V��$P-y��<��i~���j�t��hA�f%P�c#è����Lg2x<��1��e��S�a��������L��g��
�X>�_��'��M��0�D�����S36N�:��z׼jWs��*CS�RdX�.�L���h	H���@[�r�e���&�bF-Hd@��d2p��kQ��Ps��峍�{&B���"QL�P���-�H1N�I��c\�p�R��M)H3J2L��8�&*�	�lBHj�lD�*��V���囱<3�a$�[C��n*-)|�&��O��6i
P���ȩ��aQq��q1�1Q�Q���a1S�FO�9iR�ĉ�/�8u��	^|���`	��b��x:'%����KE���85��hr���1!�c�&ń<9i��&%�D#)4)��!P�X`��4RR-��2R'%TB��Ji��>�=7�SU��ܚ�>�d톶��J��:q���9�i��4^<?��bӥ�z/;������e�@������W������߻�q���+n�λq��V�ܫw.��9��D�ɽ͇v�?�o�����,l_���6}Z]Qe~Zy��ڭ�w����CM��3��̜:+��Ϊ���٨P3ܙN�,7:ۃAR�(C���~��hi�hy�te�tu�h]�<Hj^ʔo�V��Q��T�w�[��f)g���]��)�H�><� ?�0'�,?���Y��U��Q��Q��A�r�yE+��IIͧ~Ӈ�f���?g9��������bP�Q#��J���c��1��LH|, ??&���p�����@�CR��J�	)AR�n �|_8�VD3Oh<��8� ��
yT0�������}�TX�K�)zʛi�_5�������"�~h���oI$C
��v�(�	�g
}m�&�cRC��oBj���9I��Q���$��R �҈M���[q�+���vc�|�b?�ȇ?���KÁ �iO���7A=�h��9�@<k�2�Ydk��%]��5�e32�3s�3���ҵ5u�K�nV�*�Zj�
$"�s	t�����vC.��C���/c���g�, �f(:Cc@d�`�8�I� qV*3%.!!*&9*|�$���R�1II�%'��cQ�IS_L�<!9�v�Tf�ĔIءD	!iRN�[:�ĺ��<�H5�X��B��Iͷ�S3������8������8j�\���iߖO͖�e[�Tn[>mϺY��-;�w�C���9�OM0���g��>8_��_|���w�n��=�����3�;.^#
S:��y��kH��85c`t����^9��t�(��Y����iX��
���St��Xt~c��9'6��X�ge�������B[}evuy��nJI�O�T �1�B$JI� �� �p��b��loUaF[C���[?}���~��w�uw]�o]����-s�-+��Rs����kf�m��4�`iI�t�![��1���8a!	�HI��XB�t��AX��A���������6�<����L�[����&�iV��f�7dK��H�f�g)N��g��sF�y9~Q����
������ J�~\ rz8�.&��y!�>��a��5聤�����1�a&1�"��2L�2��Ľb�����ϖ,�������=���~�ޣ�z��O���^���E�n��k�#}?GЕ��Nb1��L�� ����h*�J2�+>�r|job�$Z*}�����px��~!��i��O������A��Aj�F�����i��+|n�Kj��<�!1D�\�n�����-�O���m�?9����f����A�R��BzSL�c�ʯ��W��,�H��j��'�֙n�L7s(�KYs91ͬ�f$n&�8[��BՌ�SԬ�|=�y�P%��iZ�t�����v�Jݖ�����U�׮����;��>�f�ᕻ.۱oɶ�m�6�,�0w�֗��>}�z�o������΁�e'��ܵ�e����O-8y����C�6����[���~����gf?4�����֯/[�4���U]�,����n�֢��d*�@��
ܢ��r�.��G�{��J�SK�4
�F���3�Ey�3f.�X�o��S-��7n�i�s�f�H���u�U�Q�g�b����E[z��ި�}�l�H鎫廆�v_��{�n�͚=כݞu�Aۉ�-G�L�;T���⥮��r;���_��p������5.�3k�κYK+�[��:��$�8
^�.�$M-�щ�L���KRc��SS��V�9�^�4Н�$@�F���V9�x��z��yպ�+�3
Mu9��tm�G�cU�5r�X,C��GR��djJ���<���� y	v����3�ˏ=��i�埶���7ص��)N���
k {���^������|.��d2�>-���e�y8h`lu�EGGC�Hjc��)qn�I��VI�7���k �	&���	x���d0�pk�bV����OMU�Ư%��d<5�6Jj��cb�b��R�Lj�i��|¡�����o1xB��(�1��n�;===++���;�N�)��VH.�0
i���S�(<:�S�����r�s��j�5Ny�E��ItrR*�DJP���
���Ԁe�@&$5��&p�T*�&`j�Z�T��;0P	�����AR��5\A��k ����"�ʱ�hwΓ�7��V��e�yfQ�ETl���b^ 5�6|����f4τg��N%�p�<:#%12<b򔰩S�#��GM��HMhdlDL\dltd\TDlDxlXhtH�k�L��414djĄ	/N|q*X>��$.�!��g�9�I��ؤ�ȸ��������а�АȐ����>1*����&�Lx19$MJ���j���z�P#%��h�	�BE�UBD-�-�1�d����Z[3,,ٸ�����ݻ*Nk�0����3'+O�=w�θ�9���������־�Y����������-￶���s�w���{ڇ;[�϶\>��u���Gw���8���5��ݴ�cM��E�-3��K��3�^C�G[p��7P������&;g����Bf{�9�Hj�s?a��ǘfY�dE����ՙ�uY���ui�~ɖ��,��L��4�N�h���*�os�I8���!������#��N4���|Ϧ��E�}��m�׵�Wu�7͊�u�-��h��@+��C��<���Gٞ�r��j��I���R�r�/���(�c�LH��H��P�P�S��'Bя�	�����d4?������E_�q�+(<��W�/g}���&�ks����9���WR��+(r��x�i�eC�f����������Owd2*�	��i���ؘ5Э&��kHT?I��KH�2rX!����VI�@bD-2Ȯ���ʣ^��p��>5�xP|��4ׇ�R��
��'4ۋ<K�v?N:�=��AM�ԚN�L#��D�n��+��WNKWץ��]�B�$�$1)H�B���BNbB�GP��X(��fB��K|�Q��Q��k8���b�8))4�@��4 '����O�l.�Obb"##R�"�q1��X~b����&�<%K���Me�N�'��	a��I��瑨t��"39�Ա��1�L?�X��R�����	�����`���ϐ���85���w��}[>5;�Ul[V�}��}�g۶�̾M�o�xd��q|j`���'5��~���~��f���cN��8���򑅗�,��݇�\>0h<��QX��a��"
w���Qui;D3�CM�β�]�1��&5cyM� A
�Ij�n*>�2��ڢCkJ��9��q킊�������E>�-!&���$yL��E2�X��K�|�����<MYVs}��=�~����n\��w�sߞ����״dl�_pdU��ͧ��ܷ�vm}ނߜ\_�͘)�I�N�B d�UB�\,	�������g�5`�}jt(�+�Y�99�y�9��S#
1͚\ɺ	$5{�e����姜�3z�=Op���8��C��P�0!H���>��EzX�N�b
�B2
���1����`_fr@�'HM�+�f�/����^��匬�/���Cy8��7o<���G��ɣ_��ѿ�ۣ��K�/^z--g@m�*��2�K	���U&	IU!�������A�?�՟��K��'ӯ�2G��L��;ޠ�o�S�4���A��!���!�^�Ӌs!��򮈹}".5J̿&�\'8��M*���uq�Ӯ��4�_������+d�S��HE#2�5��M7�n�S�0-�δ�k�i���L�i��%%o>/��قƷ�ImcHM��b4@3��� �e�f�:�J�V�Fi�Fb����/���
�T-��*�Dg�]J�'=�Je򊵶���u{����}��ҽ�L�Ŧ�2W���y���oi�~p����Nu�,Y�;�wf�eZ����R?�\��ۋ�wd��4���U��b
B�H�D�SHx:��d�q�J4T8M#M�)2�ɔ��SPT?�yY��=-��կ:]��r���MG_k:�V㩷ꏽ:��æ���\s�fٞ����.�~�`�P����ת����1��9��Xx��y�^�y�vͮ���=��/f/:�1�@ނ%�T.�?}���5{J��I�)��-2�\-�"�BdW
2t�<���,�
�ߧ����H�S��ַ|Z����u޶
{S�yZ��ܯ�V952-�h�q���R8��o��@��S�d|ŀ�]�.p�g,���V���=ػ�l���	�1����.��h4���j�3G��8�WH<7�	�|�Ԁ� +9V�N2
Y�w}j��&5O8�}j�`����YJHjfh��
u3�5Ui�4�Bǒp1�cc �a����1�@@����qj�f3��^dee�����LF�$5 ��B�ç��D#
w�X�ۗNw.��>53�,���|�,�,�k�).�$����-� �	Lw�/ĩ	��i��\L�J���	�Z2aPO��P�3�	��i(xJ���)�V	����pv�ܛ�(���@B�V�X��K��G%�@�I�K)6�E�QFSl�Yx�fn��_`B�Lh��t���#F�lZrtdԔ��S��F��EO���ԄF��ǄG�F�D�S��`MxX\Xh,�kB"'M��f�䰉/NK!y\����i�D$5���"����>��152rJT�Ĉ�	S"��B��RR�L���Vc\�� 7T/�AQ'A�$G)�S�����k�˱WU���ӗ,�Y���ࡼ}{�O�h��j��x���ɺK��{�*Ќ+�g���U���+��������w����������~��������m�O�>d��c�Ol;�k�ѽkO��i����;f4�(�-N�ʰԸt�e���7`�F
��ZX�6f��Q�`�[��Q��'5 
����"8K7вǰ�
[��,�/Ϥ�"C�*Cj��D����-�-~�6�l�N�CAl� [�ܭb�s���O�Ήޙz�q���j�С��E�^��I��I�}��M��{z��f%$5y��h��*���Z�����g��E�g��OJ�d���~%$��?���Ă��E�JDK$���%?�H~$�P$��P�E� ���D��`��"a��y� ��D��ϧ�!�CR󄂼�	��$~U,�I��0Y}z��y=��ﳚ>o��QI�k>�C����F}S,�IƂ� ��1���XRVaD����
�+l@J\�	n(�w�R��*�U���"��T��#\���x��>d��F��)��Q=�h��mi�v?7@j��X�o�b��D���r���
���*��>%hg�$G.�bH."�7� �c(�)!<�D}=��
9�+*0/!|�@Ë�
� �^#  _֔o�����MM��F�b#8��V�DC�$�� �$+Q�gi�NH�"qfɈ�#��0~̋���)!�Zln�sY�oa���T�VN3/~��@}�>5`���L�_3�	h�7'Li����ٱ�j��+���ud;Ej.�q�؞�|j p	
 �Ԝ;��쑽0�"5����:�yx����/�|xq�ю�c)��sd^����HM�ަ��3���mk� ���Q~i{����&�~���
�����ά+:�"���#����u����.�W��PR_]���	�gM�� ��K)�[���s��4�_U�1wF����_>v����Kgl[1sACv]�va�c}k֎��][��7�(^V�Ӟ�6��.32�2�X�K���D��I���N�M����1�@F����S��$��W�)1�mY���R��0/y���y�q}j���rF1$5�s�s�Ч�P��x��Cz�(�� �EX/�`� B�aLt����⫘p��yh/��Eg]Je�%5Ӏ|�i@��PR����3�W�������;�b���״����������x��o�έQR�?��Ǐ�~�O=��_��Zz��1"�pD=��?Hj(X 5ט�5:r���QCp�Ӏط���M��E�)L3���� ���b *�>�?2Fc�~zڧ��]���8����HM��3�Ԍ���}��c�S�n�ߝ�Gi������Q�/�~O.�+_	G���>��⌷K�i�~���fMVo��J��W�E�_�Oh�ƴ�I�E��JV��5K�iUqZ�\���א� ����Q�m�q�i9�Jf���'��E<#���BBh	T̳��ԘZl<;9e��\�,1�1�Z��ܤBϓ)	�N�r�uz�l{���Cq��t���-�e���Z��/��	�wzIW:�N�]>UN�>�@���uJ��J����I��L>�@Q��`��<��)P���S�>�S	�L�e��XL�vg�??���r�¦�;g�>1}å�;�5~�r������X��n��;u���U��Z��ە�eٞ�;��*v�T�9��ݦc���ߟy��ƃ7jwUn���_�e�`ե���r�_��h��ʎm����ͱ�Hz�DnV+��M)�J�,�8W/.2I�͢"3�KP����ϧ����F?Q>5K��V6d-�O�S�j-��(���4E.M�Y�TIu����4>/��m��P���4X�5�p��O,���V���甁t Ό������@$ j���On�{,�Ղ��<0��9�*P! ���T�Fb���h0���Ԍ7��	FӜ!jɔ|�OMk�
���^���LU�_��h�����b�cbc�����SY,��8J \�G�m���F�[.c�)`�$�T*�f�����|�v���R�T(��y�GI�㘸� ���j T�aa�uY�ky�{q�����^ao�3Vx�6I�Qbӈ(RC B��&��@����a�������F&���Xo�ֈDj�<��y��^�W�T�ن%A%��PX���,����_��XRC�(XC���5�"�()�/�qb|)�S<������9z��@�"Zl�==�4������#�V!z1W�1���D���EN��<%r�T��)!Q!RG����Ȉ8HjBn5�'GN|1�~
��!�8&�q1:����LJ���%�D'���ԄGǄEESѦ"�#�B#�C�c�D�N��|~j�SYQ�]�f�x,��JpʡFNP?�%�R�|�B�r�<����BW]]ւ٫Vg��T�sWށ}�'�M����Kŀ�HE�kj��e�
Ej��8���~����[vkh����W��{���=�~�Ĭ�ێ�[p���#�:��Z�{˼�Kۖ�n�]SS�_U�J7W945&I�����ʜna�%5����pa����t���cR�,C�<]�(M1ͺǤ�%�d�C�C#�%l#[E�m"�vk+������#i�qf�����E���ŏ���ͪw͚w,��To��XT?r�>J3��_M�#Gn��W����/��|O�(��I�(�^*��H�o�3��D��X�3 ����#����������(�zSH}O@�3��}�R�rA@�
)���O�>W4w{i�>�'Uv����迗.����*�^��XM��,�������)�x��XX�>E��x�����J����/������BrO)� u�(��O�e;�µnl�����tx���{)�蛒�Y��ě�㶥q@_�=���f��7����a�V�ЄeiQ��k0th���(�
p�D��Ą\B��IP�}(������"�7x��A=%���x\6��G���Z��I.��0v2�L��q�bHv���V�x�iF�W/���tB�A�1 V5C/NV�	J~���'L�E<'���Wrg�@kpQ���Ҵ�Ƹ���Iͷ�SL�5 �=0x<AR�%����s����ٵ�"5�WL�qj ��<�o<�����4�,���sG�7M�����_������U'vttZ�stQﱅW�/�tlA�����ڿƧ��>����k��& k(RsyWM��걤�{W���T��H�XXs�q��s��� �������kr,�<��������W�>rp�¶m��ͭ�,���IO���4�

��I�\$�s?�����"\!��<Y��u��+�o^�n���
����e����"��Z������2��r���̶��Z��Ƞ�P(�r�G��
�\�%�rB(P��'$� ��"�D����S��%f�Y�y9��Ԍ�S�2G�4k���ȕ�ɖ�ϐ�IO;�-��:ɀR<$�o��]��T}W��%����!��c�l^7�=��1ȇ��
���D�eq��5&z�E�����Śa\�G���N�z���p���;�~������?����?��ɣ�}�_o=���η/H��WۮI��|I�hx���85�a��t��]Mf_��n���L��s�ƾ���f��<���o�S�4���F��!��~�i���5"Р�&A�	8��e�cR�������.ӣ4�_]�OU�wE��I�w䐐�aԼ��}���'s����jk������@��K�Y�[�%�����d�v
ӰZ�iR�4����VŬ�?�b�'+i�HldRHH\�����ѡSbæ$D���F�㣙,�c��l���%3#�S���?�G#yh$J&��,�7����΢��&%�R��hSR�aL~	a��pA,�Dr�)�!���aQI�щ�I�1)�h#'#d��|�
q�P��H�~�0]+�4(s-��%����*�.�/���a񮖗�5�l:pg��7k�^y�{�_/�������#���S�k�t�����+��.�w�Kv�T�^{�v����o��Q��Z�ނM���.䭽X��JΊ���N�,<�;n���ֵ��Vy��t�\�R�m:�C���$N� C#����B� �
��R���ϧ���"
:*K��W7e����x�^�{V����]�����f85I�����$��-��S�&�D(&�L��)N�ݐ�5�I�
��	��}�o�Ԁ^:�	P���0�pvv6��t}A��	8
(���'N�z@�ARNO�0�$ëB���-��'\i��f����P�&KڒM�.?�iɓ��*gf�%�V���5�t�@�%��(KE���OLN�1�,�8�\�!|�I������3 T*��d����F������f�J�`S�Ԁ� ��˧�r�)�/��.ot���]���s��������l�ȫY�B������P.��� �$�UR#�������z��h�X�5K��T*�L�Ԁ���~�il.�B5XC�R`8g�s9@j��QX$5.DQto(��#C�:!�"�;�|���a��Ph@�LԈ�"o��9@�Fn���c.%� ��qИ�%��R.�a��DL�:q2��6��D��E�DDBXX�ԩѓ&EM���Đ�S�(��������p��Nr
()�����F����S(�M	��=%<frx��S�&�pbb�L���0�^�׈�3*H�R�!�l��N)�����l{a���*}����k27l�ޱ+{�����ϝ����p����X�߸�v��쑡YÃ��Z��7�Q���_;������[^������WW�\5ҿj��k}��{V_<����m�7�=����[V�^6�����"���W�m�qi���>̀<Mj�,��ʭ���ivP��=Pp�n HjF��@R��/\�.O�N�N���֧�)R�&��m�	wjE{��t���U��J�6#��91[{����:���X�?1J?0+~hV�oսgѾcR�mV�kU��E��O}��u����/��e8��1�ޢ��A�g����$5���g�W2ɿ���JD�H���e��AR3��I�?�H���wĢ �yK$ ��5����{<���Qjf���k�����f,�����9H�u�O''ua�?̞�h�G+6��U��e��{ۛV�}��:)p� ����[!5=�G��1Hj�>&5�U�A��G/�d�wIw����B'w����A�����̗z��@�fy9�}� �Af��3��4'ReC�mԷG�����H��%HE�By�x.��<��q�� �|���l>�A0.��0�����|)�}\`|!��TLbb*%8">�`'�D�'�$dH�]�X��\��^_�����<��o*vS�y�yD�>a�[�`n�(�K��H�D,�E��Քm�t-��-�0.��/�6�����d�Ý ���!5p�����%R�|j�-��kM��-KN��x�Ȏ�����Ssb���� �yf�'I��?~���������[qr{G���=G]9���آ����w<��t������$5��j�uRs�n5_Cj�$5cg�޷4��抾�s޸�㧯��?p�Ȏ�뗵���J�2Rb&M��HIE8\	)��e$N(dr�H`�j4
�Z&�Iwg���Y��\Ϫ��%�k���[jr���fUg���g�;�+��yֺtsC�cf�fnF�ݚ���U�F�Q��"����!�D3��׌�AA�\.Ƣ��Ɛf��$R������E�5]:7[������=h�Kg�h\��g��M����=ي���#>�)���M�cVU�j�-��F������
�/�t��ʫ9��W8��vg*�b2���즳@&t�����r���p�+,d�I}���d�op��%�!Lօ���t畚a���u�u��_߹������?|�ŧ���G��ѻo������u��2.+LmGx%���	b @W$h���0��8�p*��E��He�f�U�n ӌu���H�4O��L�kT�]cS��>5W0��!x�$?k�d(EjH�U���� 5.�����1?����L._ xS �C�CB�����_��q�{߰b[�Zf�i�ffZf�j���d˒���YZ��-Y�%̜8v��I<�I���Z��+8���=��^�}���j������.��zM�Cz2y��S_�p�)t�.�V����/QIgyS���J�D������<)�l���E�f��)�yNq������S������IYI9\��ܴ�9@�]���y������ҚL.��PY�bV�!��X�T^H�dJ'c��K��\�3��]ҞN�J�*�����.	�]����駺<�.ݻ<սK���2{�e&ef��#�5%��1������*6P%Fy�IYn�W�,u>Wm(TS�PU��{ �"X9~��1+O_un��K�6^��F󚫽W�ֲ���o��~�����=R��dӊӽ��n\�ִ�d��gZW�����u/�~����皗����r排)[��6EƬ����j����W�U=`��W�4��F��;��N�5��,�"=]fd���jUm�j�H�����i�����01��V*Y�]�S��ӱ5�q��	����I�&���r�h��R>h�́�ZBc�G�-���\><�V��(F���bq���Ej8.�p�H��O��X�%`y�Р��
����X6�8�cI��
4S�(�����`�b���,hĂ� 6HKK{��@�7�Xւ��}~Oj�S ��� 5�X���=5�ݝb& h���є*�F��F�+��3߫��J	4�T1�\5�\3�T5�L;�� ��aUK���"7��Q����ρ�F$�piM���1��a �q�\>�&xv8
���i�r�"QR�G��F9��I�D$��%Pb�H�����������VfzF��~����^J�,�����4QRc�d���5kp`��ȴA����A��>��j�2b��ͬC�%��<����Ba(�cOJj��T�����v�A5�L&M473X����@��ۍ���Ԁ��$5�@g�D�$E�)'�(��r� rTƢb=�Z�K��ۡ�DT��j+Qk�k@\zNVY�EZeE�,h�	�e6F�#���-?;+-%(�=���M�&$uOL홖�����5�)9@���=zp����vK��yj��)(w��S(���������@�y|�T�KR�����=�gמ	@ݓ8����-1�kb�3��]�fw�ffk$+�;i­ -jU�Ndb&���p�ʊ�e%��*��ae3fT�_P��ҥ/��\V�e��{�>0��ޡG�?{j���'_<7�����O�=�6��Q���9qlƙS�>���/>_v��3m�]8���˫^u��=�Μ\y���ݻ�o{iٞ=/l�1k������6��CS]q����*�����m���F�␴���.O̓�ft�VI��0k�߷� ��4����"���ӳB�ܰ|^�y6(_d���˂��^f��^e�Wk�J�V�D.ZB.�f/槮��$�lcD7�������
0}�ix�i���q�ƥ��g�<l�e��E����y��m�����U�9��VN}E�_��o��_ȩ����B��L��D���e?���eh�1$5@���U|k�f�[���\��������"�tǮ����/�ī(q�.��e��B0WI9(@Ro��F������9#� ��ϜҾnE����p-����o�]���38q'�bݝbh,��:!�i�$��v}:Mt��s�G��� �9&'��9��V��V�Nݦb�����n�J3ߍOv�ƹ%���{j�ä́�Q8�T8�N�&�~��s�����-���ht��f<�Y�|� ��M�et��d��*�H��q.�7���'*F��j���/��߽�š �D��p %M�RC:WabV�S��l��Wbe�U���'�]1wԆ�',�<��۷�:��ѧ\�Rk��`�[e��,�	/��Ѵ��4�9����dO�������-O�3@?�Ԁ)L$����W����]9f=���z��f錾/�h]9w���n_�l�S�fGjV���%��Dj ���f禵@�6���� m߰z��UP{^ܰ{���]������^<{h�������wͤ����<�Ȧ��6M<�qБ��8L�~��Ïlqd���Z?�к�W����U��W�ڷ�h��^Q5rZQ�oy}�<D� ���%�����v<[�/ͫ�4@��҂���opa��KG\:��¾����Z�`��^e�a-�f� b���x�Ҩ�Z�
&�թ�F��j48-���~���n�*/�{Jޚ�HcE�WY�W��>���J]����m��:J��0�<:�[�q�UVVn�i%E�I��	� 4���0m(�{j�hWpT"&1�i����q������l� � �x��
���C<�+��+�v4�6 _"�P�@M)#��QPSK9AR������<5��ٕ%�u%�ME���~����p��^R�nU�;e����׽�7�K�YZq��K�Å����Ky�ㅢ�Q�u��C"�A	7�77�����9�}S_µ�	�e�tW�UY1ڃz�>�m�����8����j��f�������?}���/�o]���Z������$�)Ty����"�@�Ɠ�,��=#����s"���2��s����m ��� �q��:��D�3�(��P Hm8ps?U��ցi�$���8Ñ�QXs���Q=&G�h���.<CI/)��z��.��aϷ~�����p{u������s���9��o�E����yc^X}o���g��د��ڷϯ���l�Ո&���y�5�1z�(�p�A<�(�I
5�(lz���bF�ZP��:�P+1��ԩ�~��,�������������������������	$)��yR�,�{CE�����1&�6��HeZfA>�͕v���Si=zduO���3��]{�w���9�y�\.�����l�EW�711�g?뒑�,(̑f3������~Zb�KMt�UQ�P�8u�.c��T沇]���ރ�L7y�ؙkG��8x�����Xzv�C��2|�k#V]����k�����g��:=t�!�NX|�u�������m�W���ܤu'��0fY۠�g���n�����zMX�k�Һ�sK{�WT}j�K��X��� �FM�IYa�COM���Jk��G�i�\� 6 ���\��R.'+�5@�ju�M��7Ln2�lqOk��^0�t����K�����������cRZ�r5E���

5�ӣ�Qd�(@��k}E���g�� `�h?w�� ���`� ��?!:�@��x`��(��DL���F1������$5�� ��4V�F#l(�l6�J~��{�;������<.8�4�=���������*��Q�"��'x�,7J+M�*���$�Q�(��!uV��"i��T'@�ׅ6��f7��A�yQ bb��:�B@�)���C��a%��R�,(�,���`�@̂�C��!%$��R�<�H��"fX�jx�zh�jL�q|�ep��Υ	YH��Ź)�����LP+\秜��B�@$�HD�L�˸LRiG6"x����Ig�`08�N����z}>�:�^�P(��h�<g��k�?���@ɢ�^6�n�����p�K ���9R��#5�GVj� 7���XX���{薠|@D>0Lp�&������47fy1GjF�ӣ+����|D�jx�z,��{['��s��A�9C����k��*7Ֆ��C��W�shlzV-'i��n���p!�(9�|R0�H���њ`|��.W0�A�� kAui4�Vk�X`e��v�$3�ēp ��Mj���|? ��>�L\·���@����4&c��@,,���#Yj&ˍP�IZnA8&n���8��ƊW[�r3�.j $�L"+��gfg$�w�ڣ[�ݻ't�أ;�c�gBJτTn�������Ԭ��i=R�vK|晤. �@]�?����N?��T�$pk���N���KNJ�_�$==\�	=�y�k�=z��8%�grb��=����gO���tzׄ�]��u�ge$2�Tb�H8�e'��I�BH�$b��\6S����ˋK�4���m����\<zd��顩S"�g�̛W4gNx֬���W��es���8rߞ	ǎL>y|҉cc}`߼�gw���^q���ݻ�8�������޳{�֭}n箥���\�zĜ�C�N�<s�С��4���/o�)�q6�5}]�f;�bǢCts�t�8�$�R8J�P�,��	hB���'���ab�Q���D5��C���s��avQX�BD�*�^P�����J3�FO,���cϳ�Er�BYּ��3�م�Cy���|��\��l��\�{N��~�;~��.�M��m��}��c��#��3��C#�s��76�,�9�t���g����I��NN��B�!�_����7J�/Y��V��?g�O��
�#��M܍�m�C�k@���(��,uGN�M�h�-��N˯2�7�2�_�c�S�URv�Do��-��`�d�8yY�|�`��2�G�2�k��U�}�P�%׽I��`�U�y���Q`J^���r�d�c*x�=��I�yF����c�W.na�W���,��)/z���-��e����H�8�����K6���P�4������}Fðg��iF�j�h��$t�$��O�dC�d�6sZÞ�)/�կ�5g��6���N��,_o���Yl����'ǩ��d��"G	�Q\o#|(Le�9+��62��SCt?Qo�ʵH���%�P%�&��e9��̞��=
s2��h�a\{(�Kp�����&G羵��9	Z�8���L�bH�+	TM�9mR�Fe�3Z���M(���9�R��*��X7k���s��[��̗����ܨϏ?�v��M3��{���e�WNׯԯC�4���`���,��rӤ>�ѵ���̤��z͔-��Fд&=$5�<��iv�en?�414���l@ځOj`nPxn�L!�Y:��CA�f�����G7\��Q�F���r-�]1ַzBp��$5�����Z�fJ��i���U��^�vFͦY��f�Z?�	h��z�Y>�qռ�����3h����Lۺr��u�wlX�}��a9�Kk�Ea�Jb�oX��CML]����3G��>�f�ⱻ�L۽jM���fБc�b�����^�U��uP{���zj�O 5�T�4��Ź�Ԁ�+^|�fϺ�ӻ&�~l�ͳ��<����Y�g\h)8�,*�����`�\����gC�Tj�Fk���z���.+*�*+/
��nO�(/.�.--r;#Nk�j��tn��cԂ2XvX@̺�j�NeS�f��II2�&:f�����v����h^a(\"�dNR%"17�~!7�Y���x�Hj�$�)�f:�R��0͏$5KK5�J��K��t���m>�>���r���V]ջ�jj�.+��\v�_6Z�ȕ��`v��\����BN�xbHj��D�$��8���*Jj�1�k����4�DT'�R�Wm�e��s�>�5����������y��~���ߴ���wn�vמ�}��T��I�Ә�?+&���IOt�P
`��P�Y���D���1P<�z��(�Ej^r��Xvah�i��N�:0�I�	����g�cr贚<� '(�Jz�Ů�������}߆�����%����?٬3�w�yS�\4)_bDw���b�ث�{�`���G�n�z?���{�[<�(�Ɍ�����<������k��#�p;ۨ�e�&^�"/���x晴�	)=�R�C�f�d�g�f�����]PSU;i��%��oܴu򔙑H%�����LAfZaFjAjr^JzAbj^�䜤��������l/W��U����������нg�n	=����gr2�ż|/_�=:�Ȭk�=Uf�+,�j��ڡ�q�*�r��2��h��g萁��5d��ç�={��NNXrj��3c��������:3eͅ�kN�_qb��ã�?4~�ik�������'���h�����G����o��cV��i��&�0qe�����O/��/�7uF��`��n��o�����Yˑ3[cU���<r�'������azh�|x���&���TjGWh�U�'7X�&��tV�{v����e���X<�O`p��_���ƬbT$�KEb>�W���'�Y(�\��#�����ek���(��0���(s��?Oj�����y���`�O����Kj@��`0D"����@ `�Z�I�-�O�SÀ���!�I��i�����(���4��T��*���$�1K!��`�E�`�B+M'=��`-�H͠0I��RzDIԃ�&q������fX1;�L3�\;�D=��<��6��P�RD���ЂLi~�0/���]���8;'���$�.���2)"� +�t� Uf!�q�\���~Pp:��H� 8�C0#5`9�l�Bp�*!�Z���s22�����~Hj(q�Y.��8RC��fh	3�� 5j�#5Q˥�Ҍi0��e���1��=c`p��Ȥ~ޡ��rse��$hyt.�ڬS(<��|QRa�T��e(GC8TP�����Ԁx�ԀY�Z�\̐�8P�`!��3��T�����*6Z�?� ���cIܸݨA��� A^� *5��KC�d��,1�eY�	)3�\g(�Yl�x���6�5Vy���I�����g��L��yd�NL�Ii�)i�9��i��)�1�L΂JH�鞘ե{z�gR~�5��`mf??_������������KMM�b)I�ɉ)=Rz�&�L���tO�Zx�%?�-�g�t���3*;�"E��R���$�"dvLj�3� `������5�Ez7z5�6��_9vTd����Z^X:b���[�M޹k�����մC'��7v���[_�q}�5+_�|���~���W_]|����?zl�K/�۾s���C�/��ّ���<��q�O3a���M�UM��}J�MA[_�a@���A�؉~���@6�\�$5@�Bt���)h�f��D��&$>�XR�	��{���5r�_��^`D�҅��������K���圔�6(~��ֿgS�s�n9�w�z�[N�u+��]%5��=�/\��L�-�����t�t�ڝ���ӲVѿg��P��7$�C|Ò_�)k�`���4�',�K�әx��f��U��)�,��M�o��MR~�R\e�˩WY�59v��]%e7p�-���o��W��(N^Tk�X��7��+Ǜ�+���L~QF�ᣗd��u����U����
x9F_�����`Cr�y���SƵ/�_f�|p�[��E�W����_Q���H�)�e4�H�4E��)�e�)��'5'�s���I�nS�Oigt�s:��:�YV~Z�ײ���&+󂓚�Ƨz��\k:��#H(<DdT���ɊWi�"%bQ7��Q�ZT����4QfbaZ/'G�ヶl�)�Z�PE�5$Ep�ցf#�r$ -CihRC⠍ib)��S#�85V��qa
��ĕ��ـ/Vs`��s��?��Į��v�;���Wv�pe��W�.�qjݝ����]�dڠ��6�B����y)v�_i'WZ&�uO�7��)M�'$5�y�����1���·�II�J��&ӌ�/�]:µl�k�h��1!5��r�f����3���N��4����Y7�q���53�Vͨ_1�q�ܖ�sZW��v�-/�ؾ�ٝ��ް|ǆ�o�k��~�2��kwlX�s�zP~���xu��W�:��mߪu�Fm_9y��7N:�a<�����sh��kG X;��������:�f�CIͮ��Q�sZVӞ�\�����hۂ���+9@������\�||��+'���Ҧ{6�<g��*���V6��,ɑ�7 ���J���H�ր)�6jVa��F��l�=špY8�6�:�U%��Eɀ�Ϭ��1R�8�J��QNj)��"��
A�I�e
`6�PMU#��|Jƣdh���@�y����h��n��\'��	HF����<��fE�~u�a]�aC�nKH�3h8��*r��]�n���{�z���^U��Ҳ˞�9��B}�dNH�Å��ù������B�i���G���B�PsP&:��GP�J�F��1�˸�5\�*���돊�G	�)�������<��H�_._h��n�7������?~�����o^��K���uGȍ�E�LyR����OJj��L�b���x[T��@��e8�51RsN$��A�4��4:~�9)C����L����g�r�8�s=uU�);%����gH�+r���Mi������ �o�����iSM�bUncE��5|�p��i��\:��9�O�ڪ�{��m�F�b�V4����S��0�p���f���0U�@Ra�p3>������@_�Af��RR�����윬������N�,JD1�*����Q�v�����W.]]�fc���(�葘�-!#1%7!1��gҞ��TBf���I��n�����523�2�Srt|S�@��3	(!!1�{��/�q�W//����HO��r��Ң�����m�R���l(��W�:���~�[Lo�p���C'm4qˀ�[Z�m�3jc��{[�4tUi������MX;d���3^4iC�5ͣW��	h��̓'oKz�XV;��~��>�0xA��ufU7O.��5ڜ�&K�d�v���9vG�n[M?�S���Il�Ɠ�I�fHjf4��-Z������˧����X�j.w���A��eTU4� �"�৐�@İB�p�hz� �08�d��4`c���(�v���	�|�p�@X�������yJӀ� 3�� �
���p8�D`F��3R�yj�R�s3�d�&v*� x���8׀��pt�����*���,jx��@�{<5QCM.�,�CX����1R�r�����3��Aat�nL�~T�nR�mZ/׈
s�[1S�ϊsP^��0[X���p�&T�/��BHj0T���x5�4I�4�����t�8R���h4��,��q����h�����œ���Ό%5��R�ebx!#�#<5\er��R5�J��U�����}����g���Tk�-5�#~�ߩvX�F�\A�f�@�=��OjĠn�g�X� ���>�k��@���I��Uz��b�8�NP�6����l�	j(Vo`�Ј���axI|�wO84�VFj�F�B�
10�CE��DD����D++1��F�ҌU[��j3^i"j��
�"�W8U���	��0#;-1�g�D���������������HS3y@�YN٢���e�R�&��L/쑚��Q�͓
�mټ�D(B22s��XvV~n�6)5+9%3)1-�gjr�$��3=zv�إK��]��+F8p܁bnw�2!�cR!52-��^��KR�1j)����I�����`@_]˖W��"��W�p���v{����T+��}���S6cZ���}�_�����}��ڵ���:uf�ɶ�+V��1c�s�Ϟ=l��1揜=�y�ئa�ZF�4xhs��u�e�E�*��ڥ���AR���Z~�iGj��	!
�~���C?$5@�S3?�,
�˂�UA�Z�r��Ye�W�Е*d	-|�,x��=K,D2�V���%�<%+xפ�&���gzǦ|��^�ҷ��[N���M3s��BR�[��K���S�g��oNc�����Ӥ�/��/j���q�/	�/)���4�,�������>b���;y�az_)O�����':��Kw(���"�oQ�kQO�k�&Jj���R���-d�i��h4\�?�l�WT�NQ�_�e������O8_�+��}#��p .��]A�|nD�#<�����F�'�nn�������Fe�Ne����|�W5�ǐ.���N������2�fβ
���)���5'�8N E�a	����
����5g���:�i�9�������	R�p�e#����`����~4��"F�#�^R�$%\��	�<<?C���KO��f�x|���P��?����� ��\eY �B��sV =�a�S#��qV�C�<��/(�eQn��uZ˵�K�:����-�ֶ���M��6�{z��?~s�o�x��]�gO�_]�R;R�$˭�T��Af��4Y�֪��2<��r�N���?Jj�G������.Q#=ODj�̬Y?�a�� �<5+f�/�ٸrn��9�+�^�ܘ��f�X���KwmZ�4!5�;�|�z9�ܸ~צP� ML����7�|����㻗�]8b��ۖ�>�~B�ь;�n�������)Jj�vx�ph�9�n�����y(�ٳ�����IIͶU��@[Ԗy���W����ȖW�?��+�o�Z}x���S[G6Ef�nӿ�c���<�~~�	\�* ����	0��I XQ�Y�N�q8�^_���[��֮Q��,�4a���m�8�A�)��BC�,�݄ht��N�'w�7ԀU�L�d�S� �22���(��	��<�$�C�i��Nɰ 2�X����,,W��1��2�/7n,ֿ1쉘O�z.To�mx�O�;�wkk�V�ܩ�|�:o0_P�����R�_t0�$�,O t�':Ηt��͍�$�A�c(݆2��\�ԯb�W$5�1�61��R����_̝���������n��A���ۿ��_W^��歧�z��P��<�M&?�GO�'%5��_��p��@FS��@@��!�� �$5�ēhm�:�)����I �<!�J�~�"ڔ�iz���D�I��m���w���������]��Z~��أ������)������Ss�ʻۣy��ntʟՈ&Q������'��@FOj����6f���U�<�|]a���KJ�ޥ�3]�<�����RR�s�
�"��D2�@ �X���S��X}����|��[����~�F�K��3�
{��u�ڥkJ���]2��H��5)�䧺'?�=�grx\NNᔒ���zLJ��H虓�.�φ�ƣc�F6���x��(5��&y�EYnV��5E&]��Q�/i��3�����G4Տ��R\2,\<"X4��	w��:<���vW��;��`u�3�����v�`ɨ���������q��	����ʱ��1��Q��!��A��!EUC���K[��:���b�N��j7Z�{��9���I=5ր���@hَ*W��mZ3������Z08�pX	Gj��M���n���.����a��e`�

4i0�P�����}Rc
Q���0����]�k��h�AR__�`�=� e�%�]�<�F����wAL'R>i�p�4`-�0�@����`���	ڴ�hx�^�Q4zA�����su��=5���9�P��,78}���\�+Oj���F�,>1ML�.O͐"��o���5��I�@E7`�b10[eWmSi�����3����Q��\����p�K�B� �q��%"1"���D9�9G&�l5�"�(
������� 8�#5������V����]�X$��􇊟_P�����IMvzFFJjj"��&+5������4Gj����=5��g�Ԍ�э�Տm4��e��>��cJ?���1��������Ұ!�V{l
�Q�W�,�=�<�S?P�$I:�NO�B�U����I� ��`�F��i2��f��h��U��`o`,j������ ۀ�_�%o�~�����	N.� ొB@����j0���b�A�XԣB�j4���%��(1�&�VSm�Te�*�x�MQna#F�W�4+�,�Ix�����Ԭ���̼�|A.O��G󄄘�	5S�#�\�2K����y�L�R���|)��/�����]��"%58�%�z���	Q0* y���AVf~fgM뙒�����)~�$�@� i7E�	�M.uЈ�B�$��V&"�����Ҳ2���s�����$� A 쒝�@�!W�\eI���JQ\JB��/�xg�՚e0�h5=��D��h���om<sn���V���ju٠!��`S/Gy�1Ը\J�]�ry��j������.�(/
�z�%6]����{9�'���HM�(�\�L=5�4$5�S��F�4b+���
�bJ�,���*x��{V��D�������yV��Ȫ�}��K��]��m��M3u��ް)�Y@���3����wn�?����X�=�v��ݢ��^�W��

���0�/	�����RN��!?c�Oh�c����ߧ�N��b��&� �&�ۄ���N˯0���:�]�d���L��DrU�\�8Pr�a^�y�����C�}���~P���;x��nv]Q�\*����%z�F�� 5R�b��;�_�6)�A���C�8u��c��R���vUɻ%�|�״�����"�!P��DVq�(NLGV ���,�8�PAXBAX��~�b�c~C��1�8.�N(�65{Z�8�V����,}T���3-���Ԁk���I�{�}m�-/��{�|�,߉���FȌ�X))$
2%����~n��/ �=h������'5��
Z�&�Ƭ՚�J��5��E�ɬ��M��l�.���������I�E�~~y�gW��}a���K�>�����N���柿��WwO���s�~��E�F����Z\'��eU�_�nB/��&��Z�O����o��
����<��<JOJj ��'%5k��m�Ѵa:�i:2
O�]9�n��U����Ӻjސ��n]>{׺��lZ�w��Gyj`b����4�6mؽy#О-�:��:��_y�ā��v-[�p�����к�QL3&�iFX3|��a�����������A������l�_S���eK��/�>�q�kg�qd�m�v-�f֠��{-�>r�����ӄ�u�fc�Hj��1#�A�?D4�5ju��mw�����[�f#(��%^7(�Y����k�Z�E��3�:�;����L�-
wf�8L�A���,.RR%�*p<�eR����u�<'�W��5;%��������l����U��5捕�ͥ��%��e����k����+o�U�]S}���ve���W��ͶW���r�	��r*)���$'���@���O�0��N��9���)^��1�ˤ9��vH�=�j��p���r���;�Kg�߿����_}�%����˯�jӖS5��Z}q���Iu4��MsF(}"R�,�x�4@14�k�:���*�*k���;�}R��#����}��:H�q�<�$���H�q��eT}��&���g�k��g��+��S��}��9����Ϧ�������)��yy`ͩJ�N�j��Y�d�ē��'���kP���4�}�X�\��xfI�B����&N�L A
��|�8�/��y(�'K��}���8�ʍ�?��Ƈ�z���ISy�� L�L�%#�'_�#_�=O�5��5��̼g�s��g�H��ҽ�Ϻ�|�G"�ر�{�G��=z�HJLHKM��I��Մȩ��Z«��4h4Yud��.1�K��^֩C]��Q�)�TV{�"�2�>bR��lH#����
hɀ���?-vꨰ�Xr�	:z�5ZE��
�EzM��\c�֙�5FS��Rc��YlUVG��]�ԇ�M�P}�W�vF��^e�+�f��i0������Aj��S����jb�fb�	���}��G-^0�t���	������2k�b��8�rKИ�W�O 5Q��=��Xl��������e�`���G�?P���3���D~�@�aM���� :a�A�y ��`
?�
�N������xRӱ�'��$%���f����岀�s�9�zQoC��3�F=5�0����d!���ә���n�l� �1P<�[e���5��7����Ӕ�Y�J��x�$�f*���A5�����y"�@&���e00�vP��t���\��:�Nh����~RFs<Ǹ@,�l�J�;ᮛ(�yP���p�Hj�8�DBfJ�¬$���'�Y���b㩁�#P?�j�c���z['�qD;@y���j���몊t�A��ź,r���))�-�Q��h�֠(
���Zi��$517�Z��h4�Ɠ�=�q�р���`���bg�&�}��u��KF�:���2Bp��LZV��nV�WJJq�)6r�A���*MD�/3��+|z�S�5*�,��RB*F�ܿ��O)E)�1�WXBrs�2�qcч�ڠH��<ƚOp�U�sm�Gj��,��g��lA�#�1{UF7�s`r�4�E	)"�<ANZVFBRj�n�=eY�:����n9�9R�UP%�V�v9��$��@������������=��3�I��3zde����.E���dp)��ӟ�-H�R1Bd0I,V��$�������B�cqٺ�����j�n�[=p�����p>N�
��j3�]:���ji��Uk�j�Yo���.��oT��j�`���S3.@����̴8L� ����p���>��,�#˔���`��P��B���(s� �eL�s����ᯂ�w��[V�M3y�B_����#����c+�������ψ�>[��Α���ߴ�wJ��4�+B=5_�ؗr�r�3�����!��G����(�yP��.�Mb�I�.��+n��ku�¯��U���7�U��u��5�j��ݍ��_Ϙ��s5cƗ&�ׯ�jq��`�m��q�/>�_J_�"oȐ7Q�B\�q����'+ge���_k�威��h}���V]��{eEoy\�4���\�%5�H
�,EŒ�g�@�ԜS(/��@� I�BR5�0�(�E�#r�Ď0�E�(�~O��cꈊ��f����!���f�G�y%�܂�Q�K�d�*r�x�C�m��Ze|!uP��@�>V�%�N�ev���̘�����v�Q.�;$5�)j���F�M��hT&����E�E-O�!�
��.R�\*I<�r�7on����O�ly��ʷO��ul�;'V�ڮ?~p��������~�����8�O�3h���l�JRlA}�5���qu����f~�S3�,7���;��v��~Z3�f݌��9L�45˧�-�Ѱ|v��Z8R����V�ٽ~�M�vo^�(O�i��u@1L�R�I]�������ݹt͂�;VN޹b��܇5ߓ�}���_34���_3p���[��h�5[�m�S�x�oݼ�}��mwl㘝Ko^0�Ņ�7-�z޸����&^n&??/�T���S�?-��Q�Yp� ����j49,V��Q��D\���
��_U8X
���%^w�i�YLn�ޡ�X�J����i���D D%Rp���� �TԿ6V�(��&44�&)A*PD�H5�� �w�%���tdW�>9�ybO͊j���*ˋ���C���5�W�K^�,z����ʊeeo�rz3X������z^�:�p�|�㉏����xN�I��Xt�n8��q� j��g�"��(�#ʗI�q	s�����h�A��������q���q���������O��E�'�_z����O��ѻ��{r%'���<8ⓒX��&��@�k:�A�3�l�xR�Qʍb�>u���Mӑ��8F���q�<����T�I���Ԇ�ΐ�7���˗�7.�}������k5�������C���8Oͬ�X4��#��|�һݡ�`!�٨��򼉊�1��'����N�<(�h`���E'�U*$R3�¢R��:���7�t6���2�=&����!Z�����ƶ7^���;@o}���7�1wb�
�fmq9�h�&ArT�d�H��=%hw��;O�-��ם[�%9�Kbr��ğuK�Y�O=��駟NINLOI��H��Ʈ����SHCj$��"�XG��-P˃J6�Ԅ�WZ�(UeZf2�6� 2N aw�6'��/7�a�$qiEv�2!�����R���n�0�"
�+'�r�I�0��I�Xu
�Fnb�w��U�*%�*0ZC0f��e0�,��OO⩉�2h�Pր�-t"@R3�Z�3�8���;�hf���^��ն�%�"k�G��:F��"AD�y	�?�����c�h���le����xR��Ƀׂ ��!~Bp�E��1���4�!5`'`{0�T�V�0+
$5�'TX��IMJτ�I�
Zi�_Ñ詁����	�i�#��<=���fp�K�A�5�r���� ���bT�� pU��Ѝ�2@O$5��
�ʫ�􄀑`�1��_������+���@$BRCa\c4�A��s���B�Z�p8|>8���`��~
a1�^Ƣ��A��y�Cp�D1TfjZzr$5��(/CG���8R�pOM~�(W���p���K'<��}b_'$5#,�e�ʈ�(��9m�Q:%���£<5�� eH^ ���X��'5�m��1XCF@��% ��@u�=����G�=��p�d\'5�*�ڹ/�R�H�􇤆�N�$
L�#�Jꠥ��Ǌ��x�	+7�V�n�BU��r37P`HG�r�^�1��Yc֨�:�I�3���ަ18�&���[�jw��[��5(���>�P�2�OnALE�1�rW��D�.�=b������?fNI�PwI����������+�f��6��z�[����F
g�<IAzNAj�4+W.Q���=���P��ū�}jګa�
J��0^^7BU��Ğ={$<ӵ�Sݺ?���=)�{jP��IO%�uM�욖�Ljf���.=�t��%5�����s���{*+�KzF���.�rdذ�S�L�mp������reZv^bZfbjZ������?���3O'$$d�e�/����Dv9ZbV48U?�S3���j�$5��4�\�E�xO�yj���C��ͺ�v�_I�R�h�R{?-��H3
�V
2��s���� �_���UY�� Gj޶�o���,`�������<��������ԧF�;�����/����x���[�Ԁ}�����/��M|Ba�8�&���n��S��t��x����	�-��ˍq�Gob�b�%�
-oS��x\�Ѿ}�vl�����,Z���o�վY^�f t^�?̗��s����}C�]EPN2�M�z��=����Z��pΪ�zԠ_�������N��5�o�9�T�0n짗��2�op�P�(Rs�U�&�E��,\a$5�A��2�aTvGGa�1�:�`N�����'��Jj�����i>��[H�P��A�˲�K0�-luIM�by��H�]�oG�
u���Db��)�J�g�
��@3����h�:*Hj�<�h�85h�����Z�VmV��Ԙ��!��
9��e�J�L�R!�qv��/^^��[>����־s~՝�>�������������~p�7�^8�n�ܱC��]Z�(�Ŋ�:q�Z���h�X��ܨ�i����ƙ}�Z=(<�����?!5p	�j��I=5����L�_5�hŴ�e��MoZ6�y�����}�\Hj�l\�(O$5�S�cHͶuk���W?�s|��c���}n���S���xh�ć�~�����!�ud�ٿf���yhF�hR�ι����Լ4�"Fj� ��8�dՌ�u�*�-�wŀ�[��n�0����G�0{�ܑ���*��%�����?v��h��h�@���T��M�W�`4��5�v���E^w��S]�]S�\_۫�����4��x\~��m6:�zprM4�0�bR�,����
�kb�F�%���ePFmP0:9��h�)Q��|;�S�*hqIG��ː�<5K+t����j��j컫���=��¯֗�\�Z]v���FE����W���F.�����*5Gj��#B�	��x��p.�_
I�I1r\���1��a���)yNB��2ge�yLuTD���{��R���3X?�8��G������wo��N�g��a�;��Ϟ�Ţe����"j_�謐l��΋�'%5p�����X�M<�y#�c8�%���{��K�����t\&;�"���<��(ōPx���ʉ�
褚8&G�1�6Fz���g�74�]��#��K��w�v��:�W&�gV�5s٩=��}<���sG8s�WK�~<k��1-m�mvv��Xm#��S��yO��߇51L�� ������j-ZmV4���µ��P(P\�/+��Wz+*]����sq��P;n�s�>�g��:|���_~q��o~�ն��fo��in�����2,ɵ�d� �b�l�K�ΐ��f(�<�$3q"]*M��{f��HNԭ{b��	��i�=s2�Pa���8�8h�yU��
	��(�!9��J�S�~�	r��0�d�|�� 3��6��$-��l~�$-!�&�E��V�q�~�+�z|��!������[*�\uak�MP`R�#DjY>!+@�P��Q�@&����	��1���H5$eSq큐���q�����&�gdB���i}3[���fMi�jt���)65F,eMЮ������3&�
��k �f��m-ظS����2h����k!���y0�Z�;�O�h�!ѱ�� G���b@!k~$���R��x�`��g�&�G����I�B�7�"�ZVj䆶��auVn��:;
��@� 41�[<5���C3
�g��̂�p3Hm �]����"��2P֍��Oit���Sc�2T��>f�DrY!*������σ���W(p��ITʍ��eG�ң�V#�Up"
��f�z��Ԁ��n��K3N
���`M��.�[ǅ�C@8#�$5�YMU�=���h�\�N�?zj ��I��z#7�~_���fД~��-��澥��"]Q@�s�c�Fɀ��(O���|jh��SHj@E���Hj��X�p�&Jg ��1����7p�E��R��K@�:���'|�("�����J�a)�$Fʸ�T�T�����A�݌��D��r+]i��l�*�T��.3��F֯c�z��dtYlN��fvY�N��e��-N���xJL�JC�Vl҄z��-���ҡ���ʑ��`��נ�7JE��|̼uk��9k��)�jL�4	7�W��7{�z;���`��W��y�e�9�jr+(���3b��-$�)��q�)'�9�KI�ԴCI�I�_���֣k���t{�gO�쩟q�nOw��#1-1%3+������-H�������͓HsŒ,�(��O���LF�3�鉙9r��hs�
5B�@�4+;71)%==����HKMIJ��$6ݞ�ؽGJB�ܔF��uv�O�Ԍ�a1R3�LIʹ�0��,ɗDT��u�����v��Ujt�\��*|ϛ/J_�KZ�O�%�9-��d��\�]U����Uyǡ��Tܰ�o:T@7l���{��n�;V���PO��g�W����V.O���/�&�NIs�?�د���O�V1ѮO����0�{��*��Jn��[�Ct�@�=�x����w�m�x���nb(���*E^E�
��Q����%�ۯ^l��?���n��Ϟ�}w��ۭ�W�����a1��ϋ��$�2���5�2���=#sMZ���O3��v��_�������7ޮ)��^�Y^Q*Ϣ�cHͣz?�e���F
����P����J�$1�A=�=���\�'��|HA��R�Կ��qI�2[��^I�G�d��yn4˅�9	�����G�XH\.�I�3��|0���;Z|1����j����	�B�|Z�8���2��I�i1[X�%���$�VT��I�2�*��s��'������^^����޿��ݶ��xy�?�;��;<5��l�zj��������U�+�k�ef��2��>��}��z��S�` (�g�5��0��IM'F�bL��1<.���k�L���fŴ�e�j�N�_<���}V��~�ؗV�ٵ�����ܸ�Q��X�'�����	���HR���Q{�N߷v��M'<
f~(�y���?=Jw�Ԁr�)ۼ�fü�Mj_z�צ����7��k��S���=\�e~+&*���F�i�c�iTr��A���S��h5�L:��b�%�`Y�_U�S[=����`گ�,,���br�6�ƨd���;���P1R��8�U%#���-�I�4�V��5��0D���H��� 5EĄr|B�����sO͒2ͪJæ��z�Z��Z����������*�4�߬��ZT�z(�z ����р/�C"�Q��Hv4�Ԝʀ�DH�=!�^`��=+&��Ih��R�� ?�*�����r?�:�4|2r�_vl�Ӊ��W_m4�UT\]ӭ_ 4���	��Xp���=�;tpo\�wָ 8w~�q����c�V�3k�������K��vݾ�{�	3�����9%T���"�C���X�?��o����&�r�7"a���	����2a9i�Ct3�.)�+/�M���r$����?B�
�qt8N�@�y�㇎n�t^�2�cN��x�ü�}U�U��c��S뜯2[vm�e�)���t#��ߓ(��_�.>�]?P&���}��Ú��]|������of��-�4Z5�8)L��D���%��5�`��|C$\�u���F*j
����AT�|�b�Bg ���抦��:����*����s����.G�����˟��~w���������%%{���aFM豫�Q(%E�F߼:"�ՠ.ؼ!r�����cÿ�'�2s���.bX��?���R�% ��Ʌ�ki��Z�DdH_����X�nQ��T��德�	��W�Dr2ǚ�V�*�����+״dK�1���F��&��h�(��V�/�.Uxf%�#_��Q��H1�r�J���Aƒ��_K���*īp��4D0�� C����%���V7�����	��s���� Mۗ���x
���Tg�^`�~B۰��Y�alu��lmF���\^��'$o߯�Ĉ�"�EIGwȣ	��6�;���f�M�^�ƙ{�P"qmOr2��-��ػ*��xX�S�`G��Z���q�M^���q;�I�$j���ޅ��D��2���˝IĿ�\ra�ގ����Z�dZ��WMr�WDږ�q��<]���ˣS���gg7Л%���6�c�;Rak��B@R)I�׫�ڇߣ	�3iX�lP)E�ȓ��#C.~'ܙ�w�����+�-,��Tq��_�3$��6k��z��<	l@�GW#����Е~��}{��-���&-�GlB�:����^�xp�X-<����`��;o�JA5��3t�<4#xB
�M����r��%����Ms� 2z��8BtN��ԸZf�̶JņFv_��m/PX��52S�:zg�b��~x��ר8L{G���~7���P�Q�+
�����`4�|,lD1l��fx{�uZM���O���n�b<��=�����n<�
��Z������[F�/:^5my���3���ki����X��V]�tsV���]�.�����{X�lYh��n���GXL� �9!$3'3#a����ޤ�[?���Hy�L�M��)��<o�Z�<2���NQ�"7Re��_i"ğ�?�aO�h䢲��q5��] S<��3f�Z	�##c�!�tt��~%C<��*���XN�{�����v�v��"�E9�Lr�����K�QЊ�r�N�r>J$z+G��י�����26Kg�� .��ZpM�۝ (aW�3L���၍�a�y����"� >L��|ǘ[a�`+}`k��ӸΑ��Q����gzVS|Z7���V��6Vqi��RM�A��H���^���^��QE��wC�(��R�$�]�r��+������v�gv���f�`���$�$�&����L7�29Z6�˶H*��<�z,;<-'|l�����{�5Y�Բ4�(��Y����P鶩��b1{Rf��B��n���ʈ��2]�%��<&��I(z�'��0�bp�nܜad���?+ꀺ�@B�#��QR�ε���0���h�)R�1�fB�#�������q�_��t��FD-�c��x��m�r�'�-Ó�)�C,8v�����4<���	B��;Rn���c�X��!}�ꆪW��w��[���¦��>�B�����f�c���ɷ��Q7>�"m��#��YG�^��6D:�ggY�|l^��1��<T��`�>����j"�@vm<�c��\��L��v��eî� ��,���ω�o{7�z	�������[YJ�k2��]�k�#nѥ7z�|6ä͛��)���>)��O�tO\�j�yWx^�s�<v�׻�N;EL{?����N��"�BW
#Qz>M���#�����:~G%t��'ƍ�rk��m�Z�M�+t�Q⹳�-�c�PB��l'$�%�V
:rM�����At���O�Bݾ���f�;�<�y����_kw���L�>fc��d`�Q�a��qN�`�8�g߭��Elꤚ���L<���R�P����ddfF��D��f�M/��������O��@��,��3��p����C�DM�2x�2�fe���=ZG`\�_���ӳ�i��;nW)�|<"c�)K�D%)aAVxx�<�� dopIڬ��X&�E�n֞f���ؒ>J�}�h(��W���q6�#ەCR�Z8�c��kEp:X�f>m��]�v(#}?���4E[0���
/�/4[z�3FMz򟛰��`r��R�Ek" Uw#� �5��W��
�S
�(]~J��}���?�Vr�) &�?�u�Rk��8�r�`�g��a�V4 ��u�6L��&�C��֟�+]8wnc�z1G����9eq����b��j�b��V՜��s�P�R�s-�8�Jk�Z �������Izc���K�\�8{"���t��|+|$Z���l ���;�_�G�+p[�x��&M�iA쵷�U1�,�8_�q՘��Ck�����s�9�;Ҙ�<t�h�<�>�~��4��I0�P|�4��JU�A�}�V�+h(�=yQ���-��
�H�ui����\|��z���R�	�����f�hR��:��1��݈�s��˧���稗���iih!��{���鑃}����N�*�6���t�f{=Q�*>4�f��r-�IvdU�	���ʪ�����wѿa��TjV�Z�l�\����ޖ_��P���tu#��[�% B� �NU�g�B�K�4������\�v�*���9�����q,�k��4��QfM�HAf.U�S&	R��6�6)��~�J�4�����ݛ�<*�T!�����_��eѵ�ߴ��/�f*�s�F�JK�xx搷g�$ʭ��t���lxB��0�5w>�];E�x3�2��f��U��cw��b�f�ˀ*���֍*_��Ƹ:�|�<��
�O�Po>�,RY�wXΗ��F:�=e��	D�wju��A�@�۬���D��Q��1w{��E���m��x�)�����1=S((6��Dr=D�c�-di��c�^Yus`��Z �[$���k����=��C����C�'mLD�?c�礥�����K����DOO�J�:��44��*~�K��t�V&	6�~b>�E��;L�P��<�.,i �w�&A�@��>	���c��Z�k@Ɍ�	�̓s Ns�y[�%�n/z]��U�J�X�F�*����[�[fZ��b�э�~� 
 �w��D~+x�C��46Ʃ�&XA��y�{���B����w���R���m��Q�VP�TR��WVUURU9S�����4,?�\������Wd�m��^�R��2�а�XV�1��ҷ�d��c9��c����5t]�Y�a��ð��������21~L�y~���.f�gZE)�Ww`� �D��:�ߊp�� ��r�/
�<
b�

l�Ʉ)��� j�0�Հ	"�`6K15�ۨS�h����|����2?p���W�b��w���ɸ`��Q6�a��/�!��MZ&�֠Zǧ}��>��� f��01{h�"�-�9�7��x�.�.���5�_��ɮ�Y��*?ӳ}r��9���u�9��v*R^���Ϣv���~r�fT�u��B	�S'",��Z֝���x`�)�lL��p��w_�*D�\�j�ඉ�+�(8;��̪z�r*ۋ�YM��T?KPe(�f����X�%�rU�^t%�@*�z��w���E�z�
��������i�_Z�b���[z���5��|�/]oKs_�$���U=~c@ 0*&*Q6��yÑI����Tm�
3�Nq����J��]���I~b��2�Lhj+#P��}	ce��fᩎ���Y����n�تQ�/�"`\�wڃ�?�]�����Y��u��1d�>=��&�^�glt���]�g��_z��v��p��H�'�sC�7.$��k��]�ׯ��WS�g-�WהӍ���+@H�j�!K�+>�Kj�F�\�)j���T�����aM拘#�,���0�3<Y�y�\�gH�?ݾ��J	�	RK6����8y���m�ء�w}G�p����+˷4`,ɆY7x����O�b0&p�'V1�����Smd1�Lg�"iy�:!I{������6�9lV�K���!��A$������J�=~v�I5V�%H%-�*�Ţ%V�(�����~�1riobm[���jg<���?N�!��g�-y��B���� ��q����-x7����ݣ(`��-]���l�_�=l���|	��f>G`�ƾ�A~#��'���{IY��/H���&<X��$���i.6�!�r1���pcsh����lÚ&kͬ���+�j:u�8�]ڤ����nJ�K�3���دn���-�ܯ�q�ߨ�->��W>���w�֟|_	��gy�����=?��~���q��S�7��C$ǯY�$6(ə߆,M~�@iE��Y��Skx��ב*����]3�ሇ�ͬJ�)�^j��@����|sa��;���b��"T-`3��Y/��j��P����
)�5�t�u�iR�Z�Ϧ��Ϡ�>t�����K���n��e����C�-.-���7G|�`�����-s��i��Ƥ*�:�>j�D�B���A���32�}�\ ��>����A�h�%�.�1x9p9�D����Y�������~)Z����%�ׁ���7�F���s���~;��vB����;�o�Dˊ�[��%%��崄������J�U�5; ͐�0���AR ���[�[*��BB��JtZh�`�_�����������c�/��mYjq�,�b/o�4a�����2gB3�xŸ��l�[�ʽQi�s��� <Z=`�X�@2d����h���w�x �]4����O6���y������;ԁRD��-ë́ia9����o�m1*��xr�d����]{���J덆[�Ǜ�f�?���[f���O�{����9�6��C�pQd���CbK7�7/�)�W?��5SLX&aZL\�R��1����o�{�E�cW"Џ�r�I���ʚ>|�a]��tU���Ï_�E�׺x�N�Ra\�c�sc�h�k=�]�c�:د��̝]y<4���_z�}ٲ�wN{-ʁ�� �����6ܦ�4�#~��7Y�������.�����\��KxJ�~:ڏ�7بfv:����}|��,���yQ���b���ew���7���ڪ��`ܡ��U���AN��hB->�u!q䐖����p۵��هΊ��O�y��bFug%�Љ@|VjE��,�\�t �.�h�(繘Ţ1��t����2��b���*���6��n�6�y2cv�z�wÌ*���$�{,��v��m��Ө��	qV��=ޟ�n�`�bl��w �֙�d5�q3���Y6����y+Jちt�)fQ�y���)_�~{�ʹ�Q�i%%BSD���j�k��٢�����6'RUU
G�I��X���ҽOP8t�dT��#�G��%o�HS��N�q~��߀���8I�l��4�ȡ�}������~E!�:~( ��6�3�_��*�o��Y
 �Ӥ��,H�C�Ả:�VR\L��p{��LR�)��ppP���lk�d{���V+u��G��(Åm��I���� �$@�#��2༪0I�iZ���F2d�	���^�-�.�_��D�N1�3��gf���KJ��sdf݉~'��&/�7���ҍ��^؃�[sC�I���Po�{Yc�x`�.=AC����C�� ��tb7�8���g��n3�'т����r��tH��tl��~�>`��kk�d;�����$����Z"�*�UpK��:����F�e�=�(Е�bͫM��/��_A��s���R!�.F��WP[��;G<P��o�HM!�(,�AK�̪���R�h� wA0��#2��F�lm33���bt�ꤵl�d*�#;S���տ���*�߀��:x*=҉���LB�We�O+�nͣu��Iؚ#����Z�ihx��ΩT�k��[��Ư�{�l���΂/��C��>�HHG�H���~[F=rgj�5be���%��6YO8Z��1Jl��@ÇhYP,�gi��,��vop��[V���8�y���WU��%zH�{U7�㜔���4���I���,�����5�V�X��������y�#��qt�N塪n������L���#���H��$��d����L�F��e	�"z���Pk��:G�~U���"��o�=�Ap��d���=-0�/�*�����Dzk~����~a ���ј�M�� 1	�pfN��n�ZJkBz� �=����j��Оs�pa)��|&��?<:���Ɏ\Ǡ�����&Q_�^Z��m���O0$c`O��p~�E�j��UYwaT�����x�G4\1}�_��V|j�/����բ�D�≔o�8�0�H'�`�|伞���|�r���r~��y��_5�c���������"��E��I�B,h��??2S�t,�4�N�ݑ��A�&��O��^;��-����Ӎ�>�6��+�n���Q�0Wj i��;h�Ԟxv4""�ׂ��I�/x ���@Ƙ�9�;�$�=�o�7�����=J�E{�L�W	����1O���N��υ�|��Q#�X�o|��9Gʝ�'D�q<���L�
!���"� �-�z�$���[1�E�����É��Q�T������V"�2֚�Gq������R���ɿ_�،�8_oV~����0�?o?�c����6��,����/�f�U긴�=�#�*A�%�
��K|�5-2�W����啑*��ŴOe���2Bu�:�O�Tނ](puQuR��x�K�z�;�N���K�D%�ǟ�]��(s��x�n)��@�+�O��l΢J:XHL�J�Ǝ6U���u_�Sf�܉5ب�I^[�4�����8~U�	�z��B�s�o|W�g	T��M��=w�P�� ǆ.ā�$�v�9bJ;�%�c|�$03����PY�hƼ�B
Az�7�\�Ϳ���s�\���L�ωE��m�dٛ�V���B�` F�|�We�`���8H��1&1b�W8���R}�E �!�T�Ϡ��0 �����-[3N��!?�R1�:�R�66^u�͋Z��Z17�%Ђ����a��0�H��:n��x��ͧ����m�z4����&<�)DǷs�}ū�&�`=,��ˢ|>Z�wk0.b���5��¸���k=����2U�ac�;Aj1��	}�f��#�(0��K	�6�:=tV8��6��tf	N��d���s�0j�R~���p#�l4�>���τq�[�0f�q5��J"������*E ��ƈ�a��@X?!����Х�<��z?���'�R>��d��'� �����瓤���Ӏ�+��Soe{aG��L}��#�����������7�w�Bd�����5��ɺ)��R�w���0�(�3�8��%���!�i\�<��պm���'+��k-�!�:���j�1�4f{�,� ����@zW.�}��k�����|���z-��x���l���s��G��~���R*�-(xsI�gRI���g�q���b�H#\�l�2���@s<$�ev��[�@��P^ɇ�I8T+�i�Cc�b/ȓF`�����U����fyf=*"$�h�������+�G�� �#�*(�g.Q��e�a�����U���1����M�	͂����Ԛ:��g5w�	ы�S������V) ���Z�$x�N/	ڊ�&Fdy���,K�X]�vĳ�gʫ�h��/g"���'6�4�m�B3�3E(>���'�K�N�=$0Y��VR�}Ӥ;n`d��J��/�W !4'�H����
��u uo_���s�'/�T=ػ%�֏:����qNLIK2JH�>GM�
�y����IK"�����y�1�a���qۉ�3,�=�9�����Y*�+�1f�h�-x���QW�V�]�Ĥ�e����KD�YN}���6-j�8y8TԸ"�R���\)u��V�l���H�7��5ޔ�+Ϳ��qe�q��5��I��q�<��Dp9	��HM
��KX�c�@��g�Ag��Ï��c���Mo�,o����Z�l����M=�r�AH�C^`��0ڞd�nտa�ʼ��p6�yU� �Metx_���?����(-.�x�-V_"��#���#�ƹH�i�pH�E1	��h���i�H�4yN�}��4cѰ-�V�lM��_�^}��kΌ�-�@��"k}S^%��!wļp_~�mW��<��6���d&Qi�UF����G��FȺ�q���~&��04�nh������'3El���y��A,�5��V20�_��Ȅv�JG�#d�Dl�+Y�ʸ˗��U�D��Ap(�(���rQ?;3����&��;3��lH��U�ddT"�)�`���>6"?<y���@����"Vl���b��ė�j%�g��z�������u�o]L}@�/��
Fˡ4fU��A$p����J�L�G�Ep�A��8�ɹ��IΦ�*�6	7uT����K�b�E�y��X�o;�����6.�"Drf��犎�bC'a?�����Vq�5(�N�K�BY��i��x�%�p�r|���7r�\1�E?� ����p/�Ү�kXpl3�x�2.��?�*݋g���XD�W����	 ��k��_�L��@�<w��;�9�*�����L�#dR�w�g��S��$ԅOQ�=���~�/4�9T=�~��ɞ�Tx�0n|ݽ���������8��{����-.���U6tqD ���0@R�Hz_Q��w�^x�)��Ff���E����wB���t,D�``��>[qh�v��|�{C-ޡ0������+�U�aUM�<~�Jfq����C�$����'Rz�(� �K\S��������~�~��&���*�a�~{��6󰛃ٛt{-��>9�8�|��3�O����2s��o���H҄6��Ҕ
��<\V%��R ������$��z3�p�z󴭮�y�	6����|jiܞHv�w ��^h�aw��\��0\��\l6^��}�N��e:��vMU��e]�e�ŴU��`��#�G�x�q}�Z����#�N�y�Xl+�������z���_e�Z
�SN�k?!� �<�:}���ɽ�^���aBU��D$k^��_k�c�0��nE�� 3�{{�� ���;j�b�nmV�w[��
����ӏ��҂4#��RBH~�Cu���������N�~.5�&z� ��'{�ϧnm|�|G�Z�43���N�Vx
��es�}�}u�ǖѳ�7BJ���9OLF	�{<���3x���+?��*��FA@�C���+��l&�t�β|T�iH��m`�w)�2�|��\�"X������N|��`�S�9i�mvzNF��ƅ����!��:-Ո��'� P�iP���G�|��O"ʙƅ �_��c^�e�q��+�W,K� ��ɟ{��e 	Ţ�hQ�N�wIs������1��a��`�,�u���^�Q4�Y !c6mH����,*?S�lG\����[ί���!�-��)엛`b�(�W���!v�������9�����֧"�\�3�^�19c��~���CH\��˾�k�mK��Q�4]g6��Z���X�Q~�]�d�Z���O c ��
(��� ���勐!��QN�"K�C�q�	(���#̘P��7=+�i�7�/��n����=E�]�<Y2l�p���ڽ���cr����dE�v�P�k\��}����J��͂����D�VM����4�M�'�~(M�
�����bO>���FG�kg�d�1���Y޳��٢f���u�G���ت��FiY�:ED`�B,��h�`�p�.>u�μ�8�,8�)
'��`�nWi�3�K��v��U��GÈ��q��ʅM���Ұ�.�֙��`Ӣ��$g����߾T��"mdg]W�9�P�<E����ۛ�"o,ʷ%�-�ES�,� V��H�n��r�JJ�ST���J��Г.V6�Ә[Nqs��H.�؊�/�f{��[^_N���o�T�u����w/!�/��y�d�<$OM3�����`|����$�@�9�����m:Q(;{�*@�!�1跼rʌ� o��[��TU63s6SUSM�����$�]�������诮����6��o�I�_YJ]�����Zd��%�nAނ4^?��Qj�1����5�ے�(]0�)-�m^]k�*����&�]����ٙ�����A\�[�+�x��}��@�~�C��km<f�UOq��9b-K-E-�)�.�p�5�˥I$<	r���b�e�����E#p�� B�^�˪�%И�f��f@��(�e�d_+��]jK��A6ʼ]l����S�Ls�m�VyK�}ɘ�l��{���L�Qlȥ��L�f~yoLD��t������~�'��5b0�@0�L�'K���ʊk0���Ȭ�qjչ�1�JͣaQ@-S?,E�}���ߔ��3_{��a�`�V�s�yRM�>f��e���C��e5���ᇏ��o�eI=����S/��s��)�hŇ���K��l����Ӯr[�����j�����?|���oh.�e�"8=B�u��y�״ÊꈴdP~���Ǧʰ��K)^�SU@C+)�����abcm��sV0��
�����㐦��Z�R��+���$�[;=�p{&d>�M�B�r"
�$�K������I���_kv�m�j��s�)�5}�=�Q�?ʁ䤐w��;��8�44�x|n䔎�iX�PJ`b�ov:)(�fB*����B֎�����-w�6��>^�_�x<��1/M���k���\�X���B��{0ZX��L��FuE�[k�+��ޣĦ#��d]��G*SQZ�����~<]���{���7��q�x�P�/�G�r�!��o@�_�\�S�2��>Q���a��I��`W�ҫ�Ks�"� �'_��C�ދ�5����y�L��%� 焐�{<���"zLK�i�#��)����Ψ��"J�o����B��ѶٗR��ח/�g��+��>�w*ǯg��]>�K5᱾k����(��+̶�bڢ�j΋jv���Q�K�����(J�E�@�"�"��i���?Wn�%���6�F|�=S��kI�
��Ig>��Bw�!!�E�~,N�	y�;��Mu/~*?uv}�ncG�����p0L	[��n��k��4�Q
� �T�ݭ�����dv�k��l�h��S"�?.%�K��]�M�ɢee_B_�����=��wr`��wt��q�Ђ,d,Z sb���`�*����TZ��C�뤏lZ�{.�RG�Ɓ!��Y��J��J���������h�d5���v��챭E��bm����x(>��di;gy��X�rZن\������u{��-��]�.wqg���z�^7v��x!���.<
w���:=�@��B�w_MR}��4���M��a��e�2����ٟ�U�`v���X�2�8(�,�1ps;�׀1���'�z`U��W]�����ʟ?�J�R㠄�Ə���`���H]�c�@����#��D�,�&<�d*欂K���:T�7N�{��5���~�gh~V����r���+��e�@�,��Rʠ��Q�@�'��>gJ�oDA1#�Ę�d��q.*�S֨0�,���9l�)�I
C����%A.�%�zZףQ6��:c��l^<x���~W�@�m�y������-?{᭿���B)��<)�"�R�~'*g���I�Ӊm
l��U�.b����s�V������Kԃ^��~.*���Oz�_�)���q{�X��x�q��(C�@�5q�0�a���[��OG����D(]�&GX��p�\4C(�)I�=(�ԡC�[?�V�nhR�g֬�l<�u��tq��-Gҙjq������!]t������XA�pC8��ᅴ�С��1�͑5�Z�FY��7NV�$ʘ�ޒ��K�������ɖL��kl���{�~&{��l��n��O<���b��,��O��|���-��.���wۿY�^ײ�^���P46S�x��^�:^z����z [^s~;����~��\q�n�����Mr7�����z�g��\RX�$P�9�l��X��Xڰ��:I��!}a�|Y�w�bAڢN�1��Vh[�M4m_9*�d�M�	4< n�*�%��^,���~h��]Ӱ��
C@_"n/��!�B��!�Y�9�����d��c̈́�^�f]F:[jo�|/�U/nX�&�U�w�5Îh��+����M���4�=[`��g���U���i�TT��q`0�b��x_?�N�<Y��֏T固m68u�JhBK�݊��9��_8���S��o��]��O1[$��F��KJ!Ƅ���`>N������sYP���n��_=A ���i̊Qr��׎}�1��'W�? q��p�C,=��+ǌ�B�HK>Jw��A�����۪�!�r�4h"O��imz�����a�6�K�cK�B����M6���SS'����;cR�P���l"1'"��g�&іڬp���΂փcX��[�vh�L � Xj`���Bb[�I4'Q&}Su�0��x�l�qd�� R�jf�K���� ��mn��SI 7Q������p(���uU.%K
I��n9���9���I`�(�&ն|,����;�L5j�hU0��(E�"%�MP0^a���:��G��j�=aJzA��@��z�r�y�v��1�w#s�
%��T�7�FD��g��Q��M�k=Q��d�)}��
 �ۅ�����+^�S�H��-+.�b��hOá�8ۑh��"b��D�0ݪ��ִ�	���ڭ ����h\Z:xuoW@�W��dr���\Z��S���t�ǌˍ�9K�+`�S'�0����LM����7:�ط %��W/�d\���?<Z:d.����>�Ǘ�D��z���;��M�[?�Xҵ&rL��&E�a)kB�vk�sQ�$���,�|>� kd�w$�4�3�5c�w������D����=`^U�:�u�t��T����s��X�b�P��f�K�g4>��S���܆�~9t$�^W�	�ن^Z 	��rӧ]�x0jB�aU�|��g�e�qj�*z�dR/	�s���M��-�σ��~�@�ه���Ӊ��Mydge�g�E;ƜƮ��M��?��_�)	�d}u͠����Z�ս��e��x��rE󶜖�]1�����<���ɒ~�. ������`e�#��C�F�zr����N�}�^����F��L���'��vt�UЯ�yj���v�d��m��v.b���>��9 �ؘ=�'���_V�2_	-������Џ3��1���u��3�.&��Q��g qE��zL��Sd %�;`H �*��7b@���傘��^*��k0��y�~��I��Bq�48, �;�?T/�edR�K�*���ܸ�T!q�O�����;"��t���/
�xk��i;f�%*H��"��Zu������=Xe����bp��2�� '9p7�j��:��*�{rm�f��\��$� ����5N;G�����2���X��͝�]�!���{s�FT�����ǧn�v�7��'"�&}Y}�I�x��@$����Q���:�T�^6~X�1���	��x��޿V�Z�mȁ�9[��Ƴm�
]t�s/`�r��G��g�>�"��S�>�s�H�1������H��K�.$Ɛ��'H�e�DG�'��t��{k1*�9:������[����5��
w���duѲ:�Xp1S�T��F��HY�L��0P�o5GLW�6�{���:R6��&>pX�$�Q�r�_p ��u�s��gR�o���u�v��qo���|�ח�_9�Q����K-2O���e9�&4`N,~S�~�K��L�	O��{�fWMLX�P��VM>/��[��Y�Xl,�/.�/�틬n��j�����qv!���)��l5ҽ��2��?x��|�_��[G�^0�.	W��_߭�i��Q�q֖	:?q�]��\$,Kn�j����D`���E1R�;Y��ˢ�͇2�{E=���*��K�(e��&��/l���I>~�������sd,���6����M�	˼AP�H�=C��D�q���d�yQ�c�[n����Ud�eP�s*v��|�1������xWN�Z� �T�����п\c#I�@~�ӷf��˟�~A��i��X��v�Mk��)\�<Z�\��ʃ�d�z6����MS��ji�"� �a�L�H� P����q/��X��F��ަ������g����0~	�;nu���5<`��z>\q�\���>��ί�������犺XªC<ά��;�מU)�ˮ�_�d1��gm6~D�E�U��5x��]�=V/��Y���j|��ʫ��E���9S�H�/Or��|PfP���)������A����m�մE������������l���Z
����S�J��`'C���Ɣ͂�赵c�2Vk�N�z���Ӆi�d�eu�
��S��W�X�_�]3G�93a=K�2�o%)3�~bz��?BN։a����Q�m��\����RK������ͤ�� *���d�*���l=	�(y.�-��{�c�)��*��<�	u¼���H�!����ˠZ2��i���&�Z._�!S�8a�s���@���p��[�I�r�b�����I��p��L���3Z5�E���rQm��!H&辢o����d="�$յ>�\Rg���\K��ޑmN( �<���I��>���NZ10��mկ[���Z[�L!us����~���k��g�Y5ɝ�'�?�ױ�G��]���S�NI�C &��众W6"_�y�D,��R��?`�h�`��*?:��3og��l�]%Um�j:��ӘANڃ�m:�V��Ϙ��ޚ7^�ϖC�����SՌ�}a4����"F�'Ψ�>TP��i���ƌ,/�V��_�9�"%�l`z$蚴�piq/���,P6���D!Ǌ���:H�:� ��>��:le��D���@�e7���Rj�bb,)�)�|q<�s*�al1�=��q8�fȮ��n������`�\�ͦE�-�D_ܥ�ec�묊����xb'Ɔ�v!�7�VM�� �n���/�B<{ԍ�(�{S*�Nc�� �р;	6��1�]�Tb7�&������ʄ!��Դ���R����E����rD�Ztz��7
�c
�¿:c�_&p��'2�?�x�e�Ρ�iO��L��2��<��?�ޟ/]���}�ݟ�lP!#�w����ο�����fⓗ�E�ys������Hr`|��i�fU�^ʱ}�.C"]�'Nc��z���o9e߷ڄ#�,s�.	U�?�z�r�l�-+,%і���<V��1��OhVY��X�CK���2�	d���O,b"�F�������Ԫ�H�F	:ӳF�e�C�d��;/P"rȣ�+�:��v�ft�}���<��#kx���5�ﾋO�&m8�������c�4I��h����\TM�5�_��Z��k��u��f��7����4%�.��_^��sh�j���~� ��ۺ�z&?�I{%D��W�QPKj��H3������!j��Lp�P��q��2���C�5��B���x�=�㬎o�Lζ)��;�1���OÈlV,[yU���D���jۍ�Ê?]"�gp׹hv/o���x��DLĚ���d\���A���рy�NQ�ˌ��`����Q�C\\2d�sMfY�sz�/�+P*~��]���>��qjɽ�P����ˇ߬79U���;:��N�$��6v�+�����"98���zA�LwMcJ�ww�����M�I�h��
�����a����33<�K�3�n5|�G~��7�;t4!h�jT�Ƭ�`;0�p����zP!T�Jbu�Ϝ)�z|7���dZ�0�����u����L��(�!|�l����:l��_�W������k?�d�YosQ7�y�`�S���e/,�nֻ�����	[�(��夠�{����C�S��Oק����܇��0o!�T箨��qpWqQ|m�	EAB�[��]RB�f��S@j���V��ka��RJb�]����������|ιy����3���˿�&5�z"�n��<ތ�U<�}��H�y|f�Z��m�B��l��)�	��n\-ە��_��.�M�D����H%ģʠ��n<�v:W���Ls/�,�<�+�Ȍ�u�o�l�r����g?@��cO)� ��8a�R��T��!\Q�9����f��DO*t�g�5&������?���/e �z���$�F��N�B��j��ۑ�X@�`����h󖰛��kc���w�ǏQ�~D�䟴>�� [خ�5Q�5±#~��ѬN�2�b�������v�( �x,z��Ą$k�iM�L�t��榦E�[�Q�9pa5��$�z�-��Ś����0X��AͩǐB��F[&�	����/�%]��ƱW���ʧ^�%��@��V�ks�X�"��Z�k ��S��w�-H��1������<j��gOz�|��j:1mf3����:c��,�"�o��pm���{S6Y���t�&-t�3�}��X�J�r²�м��-��2M�΅5�|LS�x��"˵��/���!�d�b����*�I��R*�]?��ib{|�D��=�����:E��q����S~%�KL���v�fU |�9�/�q���E34/����OT�m�|�
S��x��ۆ���q��oΘZ�l�6lEj�ЯP��))Q��j�[̩?�/����0��H����/a?I������p#����U_D7�
��u9�G�?d��n��á��m7����^�_������h	'��3��L�f'�?`Δ�@��z����YMg+ٓ NFb��&�P2c���`IF3�{>c���t$JEIi�8)j�%!Xn3�_)�"|���.�ߐ[�J��63�1�
t����~����O�o�=�/�<'b���O�M���2��q��2߅�*��ֺ�(S�]�X���a��FDF���oL��}HfcQ��rYs+��⌐���@����wB�5;G���)������:(�Ar�o9�o9��o��~K�q�h��m�mm���8��Jty�HJ�N�,/��^�v�w���)�Oꆙfs�ˋ^P(�K�c�
��H��"����ϡ�Qo�����\a������'�V2Zx|L��XEXC���ܬ �A>�����#�f���V8:�w�PR�E_<��4��5�DOG߅��&Oy=��xOa@0���v:Ec�-#�9(��e�P�Xњ�S�DC�������?�XIk�'V'l���n��>�;�l�sh�%�[h��و�K�b޸h&3�2
��}S�H�Aë�,���j/�#L�!0?[Cag:�Ù�#�x�����e+  TE���z�S��U,&Д���_o��&dQ����a�k����?K�5��8W��:D���U����`�o#պ�S[9�\ �����%S�5�g50�§�b�'��W3��߾���J����N�>�~|�9��\Ј!��ȑ�S���ـ1���zRU��:�G3���פ�|C)*?�k��[B�7/sV�'s�T�t��O�s��
��op0Xk2�Z�"�Y�4�1ؤ^eyl�-FŤj��`h�FG(+�Ɵm$IEgg8��@�mu��$67]:�$|J���LW�Kr��ϫ��£��j����ԇR��2@߮c��:	ԕ� dR��G�t�lƔȤPX�!���;�^����a����:Q��h�[6�6UieT_�u�>�1*2��B���y{�'s��t�뻌�9�^��k��8��?���W|0�{���s�e�=�����son����bk�߿����ѻ:S���2sW?�����Sa���sͫ�p�~
�5z<G9xG#$�zۂ[�a���݌�U���c����#��j�糗�� ���@�7K(���:��:�V��sz�"���䪩����[��䍭l���3��y���UR�!څ,�� �[�e�]�S+	���G��s��� l�ye������E�B����������������� ����.)ՉK�=��9	��#8�ˊ	!��0��d�Ce�.��d���]���ˣ�g��Ʊ�3������>�켞�3�?���$��w�-�o�?����w�%@����dβ��oO�̂���?���#���O�f����m��N�<��,���]f�[=؝w�L���TBZ�G�����0#�e�Ь ��me�o���iP}o)���#3x@����A�`�=W���u�ؖ.uR]���7��4�\]�+�~�ө]�TP�bkS���J�Iv�ئT��ǐ����r̄�Iӽ���f9��ף.T��㏏���Y��&Z�r�b�D�p��q�A(���~�d��sW��Z��
���K�]��*=�5�Alo��SP���<�������M:�V}��j-eE�9��Ef�:ɨ��ڋ�c���t��.Jֈ�M�r�/�Y-����m6���)�R�ǃBS�AܰM�~T�d��{+�{�^T�mi̢;�IT�
�o�Wn
񿾩E��6�s�d�oy����v�Vf����e�@�ܙ������O�����m$����j�P�֭bK��0��dn����Nq��+"ܑ��VB�RQ��r��n�[�~+ݑ�����I"Q	1��ƺ�AR��<�W%�=�{��<f��Y��&I���헃a�J�.�U-���ң���~~WO����~9�%����wH�[����$X���Q�[O#�l�3��������:1%D��ޮ�|��ݭ�V��t����򯖕���4�~Ԥ����nNV2�87�we��CM��s��'��z�-�QT�F�u��F�D����O|�u������5�M$�o*��K0�9�G_%M��]c73|�����}6�\"V:�)�g<_�X���%W����4�I��-�H,�I�񵑔��(�z��"nL�L uK:tڑ ���>��c��3�>rӵ�/a�Z+bܑ__��� �ӡ�5�M�'����O�}�[��]���l��2��èP.Q�tOʛ��M?�UE߼"	�#-�p�T�UǾ\� �~y�A5��2`P��h��x�=i��tEC���|�diqD^���R])ښ��>�N�YA�?��d�*2�����ښ7�f%.[J��N��b�W�b5�A��"��iI���b�+�'7Eq�BwS�	�[�}����'q�����|���d?���2����nq*_V�hQ�1^����}~�
�����rҳ�٪puT������cBj>����Z���b/�B��(I��W��>��!;� o�)}��PL����G�>�W�='�yM�%U-�P��_I�����^zK�̆k��A��R.ec'��ȡ@k�J4��6���)Mm=mC�eo�_�6Q�hC^�����-��/s5k��a'�~��4�ɯ�*�mwVx�;tS��7���u�t���^�S	��UK��H׷��tǹ�����k�vJSǵ�g��l)mK��W��0�@%:.^@L*T�m$�"�!��}��h��W��7�P����(���L�4u��H��|�Ɠ�y��"��7�J����9S���ix �t��A�}FVpQ�ą��cUQ�\��0>���\{���-��cZ����9��HT	'��_3�/ڕ`�FӾ��T�M/<�;�ұ�lʅ�	(�C6��03���O��H �ە�,����60���"�r�.�`�P9Ժv���x�gZ��`�� �k��%�1/��̐��JHo��J���F��;�1�n�c�q��� ��DQ���|������3NCl���g����MMֺ2�H�=������qof�"r�^��ɩG����|��P���^qo9������>�;�)F8B�s|{Q,�me}(�$�:�&Z!�Tb�L�G��kz����0&�F�p=�s�X]w<�k|[�T�S��k���cm&S�
�^�%����kv/"�;�����i�QU���(����7*�QN7�iU�������W��������Y^�'���)!�R'���9��Skx���Wkʒ<9�@^M�0��%ϋR��␏�s�1h�pK�Z�=�����﬒��)kP�&�H����uX��]m͌��㒉�{�HS��xw��j��͒�����!rC��w��uz��(�eop=��b��oc���t����ies�Q��S(�b�:�UUZ��h��3����H�8҂�V��Oq�Tx=��6��4��v}�������Ea�<,Va������}��Xk�2ޞ`��"*�$�"d��A�1f�F��I��غ����c����<����;���ٙQ��s)y�pv��B�[C���$���߸����[��.qN�-Z7��uR�p7V�r�.}���?.߆W�I���m��0y-K'[{�*��U��8��Ժ�q�G���@+ �+��旧�_�櫘{�
��+�G�-C+��I'g�a~�_�����Y�9������]r��{HX� ���d#��q���q��b|�+��qep���os��T����}'j�t���w{��\0�\��O6vlJ�zK�Gם������5��o�iA��Rob|Q���~D5|���{F��A���`�X�&�L��6�ʠ�����
B؅�$-�B�wϧu�(d�2�ѸmX��	���x�\Bѷ��Y��r)�*	j^�ϸ�����S|gQ���{F����F����x�1�uS�ɩI�e I�>���ۚ/Uc[.��h��Z�V�U��*z��B~`��PR�A��O �#�V|U��8�sH���}�C��\Xx��������f�*c��M� _jN�K�Lb��Hj!�,>+��L�oͽi�\�ff�Cb{�p��hYC�`����fZ{:��֫w%�� JcXxNĉ���F����|Ze`�X�����&q������oð P^`����"#��$v����q��f�(���?X8�#AS�<|�'1G�����ʇF������UR] [�`Ѣ��ԥ5s��xu����S}??��chh�7�L�5��&w�����H��ũ����Z6�ި<%�@#��	ɜ��Ʀs`�����Sw.���b�*Kk�&��(�l]��U);��X��a%ĩ�ajЉ�d⟊�K(�G�|��)Hk�XF�ȉ�5������uuu��,��ܢ����j����\��pW>����k�膔�$����\�_�a�9�i�#�ƺ/�<�)�i�F�YE���X�(!��e}����~��E��):o����!��4��]���������F��ȴf������<>N����A7�0�Iq}r���.r{ilevbe~iey�ha�LD�TD�R\?����NFz�f���k4�l�s$����b�B���T��r?g�OZ�ȟ�ۅ#Y?�px͛P�U)ۂL�x�Y���1�J	n:B����f����#���/C-�i��|�4�5w��u{H}?C�I�N�H�H�}�� ��������?��:"_r�����F�h��W��~�H݋&�~�R�>kl����5�[��%����̖O��	ff�+`����+�o�zǪp��V�H�	!^�2���-@�pXi��]z�o2q|�|*w�(ڭ��Y��-*����S��5�Z��T��N�c�&���o̢Vye�5�o�5��c����+P�e���d7$�o�P;e�bC��Q���H���9��:�ZL[��8��x��i��������KA�PR:����V�2>mM�rg�Ů;,S?�a����̔��'���!{�6����/�*ŽmG/(S:.V/F;\N�i�o�ii��ڗ�/�����3��~�NQj�9,�z���Dm��J��{��f�k��k�.�X��mj2�k	� �>��#1c@A�埽;�z:�4�di?���#s��5dqKޕ�B�sbO n�#�@o���r���@��>�������N�ם�7{q�����V��e��M����n�e����TA����|��~e̢31a�rj��T⢇��~��T���M��'"Xj��2yd�'����X�R�@@o�>4�b�dĨ ((���K�c�`إ��A�S�#�����R׊Y�e8Lc�F�nRY>S_�觀�y��W�1���g��V.&����x��2����O�jÞ�q��)�5��@�n�}���l7�&�q��g�̸��2E�i�U�r@�rh__&�I�?�X�l}�Ok���:�8�_^ͬa�.~�&w���K�����he�zH���:c�7(�V>���4���_6�O	/�	I%L�z]��o�hSTY��b�bPqL�����\�DǹgZ)L�G��9�8q"?p���U���?(Ho�_�{��G���mӦS/۝N��6�Z�2�va�"�n}
'uo�vd�I"�g�FM�#Z���m������Y��t���]��bV���3��3����R���,=%Ce)�	��P��N�9�;;���}��3#5ձ`}�����d�)h�� 
o�7T����
=Ƶ\{wa(s�H�iTN�|�q���c|�2����N�O��A�
�����(VrE@,�k����-^,��;�/�߂,.e{#�e�zJ15�~��������������������ގoP�A%�-��U��l*�҃���O@�Ӹ�K	T��ݥ�Hɂ���9�X�	n��������������αJXa+<�9�B�Kq�:���r0}w�~� F�K�����Z)�̹I=���W��p���.�׎h+�C���h�J�4�򧭂-�(T�6gw|�Wr��*Y�jl�R�ꪞɞ&�~���F��/�N���Ux���ٟ���lu�����8+�| ��ג"|,�@�L�w�L:O<䗷�%�-y*�A:��?�L�q������^� �5s'�7��>}}����K���6�B��iJ�V�"s�yL�￺��|��W_�@	��~Ņ7�Dw�Uu�0|���O�'G�Z"NGm���m�6�@�T�n���	���G456W=���Ԣׇ���ݹ����b�c'�K�[I[��w�%�G6��k���p�;��~M�R�2�F���T�����DD��ٌ�Ť�iU�����!ּ�EW��㔋U3ڙ xU���3vW�/xZ!���p�3�L�y��)�Q�P'$8����F62)&���S
1\�+|�,�c����;��ZT�̤Wߤn�$�{R��ô(A�^>�i�!�̙	ѫRd�@G���M��gkӸ����ɣM�]�G$��>3ͽ>�_��K;ʫ����V��pq���C}��V��K�01��
	h���w�-7G�Ĭ������u��֮��}6�:s�m�aǦ��)��\�2B�2M�"���qN�j���M'Q�g}H�w�ᧄ̞X��#`�'�]t��t��p&̤P����6*টT��ߓǯzG��E>wG�4>N�פ��~�>˻ސ���Y�^͟�Y�q�I��t��i�ΰc9�ߺ���]��p��l�����M[$HQ�n���e��@x��.!5�!��'���&p��C(έ�PPR�e�+�����۴Ρ�� s�5ږ�=nL�E�+7�!���t*�s�-lq;����O�����=t����C�fMl�-,N����^4$e���qR�Ӵ��l#]ƻ��C<��	O�c�q����E�����Ș*�7t�z;f�^#}��g-.��L	C�=;i��ۄG��8�ѳ�JF�ȅ%V�p(�{��2IJ#̒)n�Ϭ�|����!��z����_eb�>�����4�������BY��A>
�oֲ��p�Q�]p�/�g�M/�d!9Z��ѯCs�������^�$M_�K�*"��N��&�-=)���,��F+��Z�b�����=���}w�Ox��BR��X�w⸕g��V,iN�Ա	�=���#���RT����2��m�V�B�ϱ���d�T�y�֢����-I�4�������"��� v+����`��%�l���Ѕ�N��jzN��S�LS���nϸ�OJ��~���|���|v��Y�!��)/ܭ�ҧ��5��P�g�v6QiY���r��@F���o�(;�A���k��Z�<�ŋ�ט�x�qy����,��v�w��+�KN��ֺ�u������i�����ާH���u���0&�0:4�>y�u��.g�v]]2}= ��Q�vi�*�A�����~x7���;Q�\�vW�A$�r�E�< '�)�&l�3��� �-����k$�n���J����Zҷ�6�Xy'�u�o�-v,�`}"��i�"`��j��ؿ�g��Z���|.*�F�����-ʆ�X��,+i,�����9F�n�4��	�ъk����y��+�;�_��
o��&�}t���u�n!����Ǡqx�F� ����}�����&��a�ҏwӟKJ�ס��R�h^Lc��V|��kK3HP��wv���%#S6P�ϝ�r���	��T��I�E��bB8Gg�K�z�zć��wEfy��Ĉ�D��Ѕ�`́�'tWzh�Ck!��Q��.�1I�K�_�M� 0p���6�V��F������Ƃxv��&���s�g,�*��Q��?�%�Wl�H��	�r��ab�[���He��򇘖iv��a���i�Y���I�lӿ[��OٻJ!�E��J�sPЫ�k���Q�/
�����6�T�vXηd�Oͷ�\�Ro)�7;�_M�rgϹ�L:�	�����-��ܞ C<���]��E]�-�3���Gˢ�'¤�í��#��ݗ��Wǘ>�BV����4d| ������/�T9�~s�k�b�$��g�t7:Z+��:4"��-�G5���jF+Z�qi�GD,vA����z�Z��$���ֹ;�&��Mr�����v�|̞�te�n��������M��;����C��+�~3F;ܶ	#�[��a��e�r��ac~oڠ��	f�3�7T�l��Of=��=�O�ſM�������J��v���#/^�����d�x�Ѓ�A<uV}u���G�t��YT�@U��c� F���q4��Ptm�?���� �9�����~rYZw-� �&�-ǹ�g�����k(X?ѧ( ���(���1ȳ�H���+�A�]}�i�Ԁ��e}�JwL ��w�� ���'�'*ښ�
�P
�@��JsH�	�o������T�ƺQǹ�^ώ�#u��v9�&���� ��9����܍r>;W���~����V.n��n�M.�N��s3��
_10W�}�W��)/�`A����
����O��Ŕ��Y���rڒx����g�� �3�T�WQ���/���q�� Dq*�5�H�
��l�Բ���]�I}@B�(�#%`��~K<!�;�Y cz-�B�y�宛-�>w�E���4�H����+�k��I
3^�G��|bS��l�镏�Pd���>�)�}���H����>���_�㙠C�?&����ʧ��m�:�N�ɢ�������ǥ��d�\��_�J����w���p{���H�c1�4���<z0��K����OK/�|��i8�!�Ņʀ��2��nFbjQv��lh�ND���ݓ��֖��r�^��w�U -<����1�;�{�Q՘����}|6J�6��v3z�6� 3�K���㦵������ԪY��A����")w��~����MBx��}�����+�����)��r�#q�����ݢ��K���]�R�D��nQ�k���Ԇu{��`��ׁ�4Be*=����6g�����F��1����)�~�ǪֆU�i��@'�Z��9��=n5e�{U'ɒ�2M7	��YN7��L��������T�$���EoiS^q�}Vyy��t��p�}�ȴ�Pˁ����������.=L����X��<����]''��5�{�}@���U�Y��Z�{��vNb����E�a��-)��h�&s����d��dqG�8xPB.��>�s�����~�B/lR���x̘��ް�ۥ󙶟ΕeS𸛋�~Lv��Gu>�������҂]<�+��C�w[�L[�9GYx3+xQj̇�[�ЛE{9�m�F�"����%�ax��&�R[s�F3�DP�?/�-*�@-�LV!|1�;�cӎ"��LL6��)�#탅zW��ץc;`@�G|Wj�ٌ?J��9T�=���绊�%��
=Ag U���Z��$��M��a�g�
(T1��sHTE5�\�#N3�U��֍n�sV<o�6���A��5�k�$%� �%@�1��Χ�hqx����1/�I�
���x
�����T�(��f���_�}��a�;R�2���&.���8P3{���}־UQqw���X����n�Q�CфD�ഞu��9z���� �e7�n���d
cb�72���V�vZC�@��Y���_���.F�t4��e����0&
cp���dj�>��uI�Q)Z'J"�LH��[W& ��~)D;���Վ��Μ��]w�K�1U�[F�ژ`�5��VJC��_�y�������<�!!�� �,�&ݥ htNgZ�]dSpYO��288��j\����	�#�z��҂��rڃ���me�{h�Y�n�喺��պ��|���!aQ;	y�ք�CY���al�@ ��/]4/�	��#pn�ss�������ox3%*��	�����5�wh��僚����T�R�."z��{���-N3��'M<�� I�:��E���Ӏ�au�R[OD��(�P���vv�G�8�6���/�ˆD�3��ٜ[?�V�t�.E��t�����Zgo����f������-߾���F�s�K&��ծ9�$`�=�&�jv����������%����,�5R�ki�����"Mu�Ab5pH�8��Kq#�p���"�u����~�1�.���R�gϦ&�I
0�խ>��������(�{�v��Ɂ���>�� yukU�+�b_���ɯ2h��x���'�Z��_`��?d�{ȓQ�A9񢂰�2��B��Bƥ	� U�}޳���o�x�Q;o�b��R��%�RE��o��jݾU��Y2��t�2���=-ι3d'e��^���PT�N���n�;�܁z�}�İU�h�o���h������a������>UF����b+�pYt�+(��*f����f v8A�h[�F��0ݦ��|�*���J�_t�N��X��NE+vr�T'�E�(V�����v�kK�fn�ɔ?dU�߆���SU�[�w�V&���w�Cs��Ul�^cr
�O�h�:u@f�#c��Ʃ�թ�~���q+嚪1n<�z��дI70�g�E��^�7���U�h"�E�����΋��L%��溰�6{��;R��/��e���c��W6��*(����U�FDH��q����K�ч`cL�x��Q=�!a[�^D��"�;�yX��z�~z��nV_��V7W�n%;�4�6l�r|�+�Wz�d�����|�d2]bѫϏ����ڜ�ǋ-�����Ə�	�Kݐ}0�ĂJ(�p�?c3d�~rR
)	&��`���r�9Lu�������9��k��*C�$S�$��`O	��z����D7(U�VI����D:Pz�|DMd�����џ^J���x��&�I#W��!���|�ĵEo�e�b�������R���l��iJ�p�q���v�<H���q���WJ�ĳ-���#�����{b3�S���!w�kÚ6��Z����m����t�ģ�Mjv��B?���i��Ǉ>�����;X���c/���L�@��1���tV�Q���:��ז0�����ѿ����Vq�{�e���J�� ��><�T!O���_����s� ��!�[�Q�5�C~y?��Á�r'��ň�Gy�!��w����JӛuU�j��|�'!�Oڊ�L�
Dg}�c�ܣ��\^	zxыG���%P=u�T!=�ʩ84^_�9D-��[� ӯ��,*�3���oq>����8ZX��q��y�?}8�_�qtܸT2�\k�uy�y7�nK�r�J"X���-�?��mye��*p�;�����d�PtT�{4���A"�R�w`q�����=�`���9�K�ҽqF9��[�0�����a��l��\z}@|��JD)����R!M�D��w�w:t'[/JM��,⹉��7�t�`�ER�����K��T`�ݺ�V561�d���!�0�C���ǭ�W!�j�w��&O�2|��ؘ�r��W	���砻3j��"������u��4�gq@[�@*��B �ؙ�j��{���Gq��-1wx���7����Sc٫s*��w��~
&��ۖD����+G��b�^�XbFF��{����I��I%���W�:[�6{K�m�U�@w3�W���˫�)�g��Ũ�7����?߶3��)��e8����}��j�|�;˃�����Q����;�3�"�R�j�O�G �2���3�PPn��� ��wG������tdV�!#?��c?�rY���]&'��֬�*�ϟ'�����q�Ge~�پ|	d�n4_-_L%^]�P(��/� Dj D��	E��R�b�@؈�D�:�����.�s��WR���bR��=c��I:��	!~h8�d��kOJ��0)�
q,�����ְ�t�u����o���p6k����y����!��A�#��zE-g�N<�8dNg��˽@�t^cu��3N�r���$|g��2��|P��76������FG�,�P0�x ��&��,��l1�;�25'���ޑy�	Kg���<	�D��p��V�<hS�ZJ]	A�֭D��l�V3�}���57(�ۥ̵V���v߽��~���z/-�&\��������O��XF����
Z��"E�-���
�ʾ�,ir��KL����hd�;�wZW}�,T'�[#�^�{�ګ��*���d�*���"�&�����j��1ؾֺ�uL�2�ֹ���I�S���%���d�f�d��:�xf`R%����T����v�j`����Ք��}%��<��L�5������2.��v[��.rEoy��mtM!+��@�<��{F�P�^�_)��G�˄��[ҳ���z�F�Orr�y���k�l\�׷��c'�R� d�R�~#�:�C�@ >S����8�c��RZ�1�]��B��"�f�9�����u�2�F�Q�|c�p���L����L��r�9�O�QE>�_ȅv5\|Q�]
c���2�Pa�;��TF��8��!t�M��Z�@��)N]�4�Y�����v�{��8��:�z�&��֗p��)��sڙ�#o[K���k�!$1��kf�dF�xF7�M��:׸�+�W^�v�Ρ�@mv(����9�`1�D" �V���{�3a)Q�'�/VǍ��:��ַ�M�]ѫQ��hV��DP�%�p{S�ŭ��;��x`G}��1n��W"����oaY�5;Lڻ:Z�=�.yxAr4�8�W4W�4���lh����Mmwx�mֿE-�����g��t��V��Sw�F�`%�mz���'G��򂱬���șE����f�]��4�f��J�o��xNL_7?0�#��g1��t��կ"���VcM���kݨ��R2��JL6�Z6�JR2+��t��5n��I��Z�Ƶ?]L����zu����M1.��m){(��,{�O ;�-��4=��y�p�*8�E�-F���mc�O�7Xq
h�m
T&E�>W��M�t�)T����l�?����d1,��u�EsD���5_w�wAP�͞���٢Pj��nD7��\�����R�,��H���
��{Q]��S�����KͫRr*N^]���۷��x�'Nm��Q��j|A!���P-�Ԯ�B�@��/WA��qI�S=�H�1��~��E�Q�����4�6 ��2GC��(������ T�	�o�28��]�k��S�e^�rRS1��u�&��Q��ͬ���#�,� (�	��nr��5ȱBxT��aX�&�n����:��K�Y/���L��� S�sa^[q�P���9�L�T�M�E�.uD�^ޏ����m�U�x�6аfsJ!Z~��vL��w�ƽdl��y��T{S0�<:��NAp�z�7��ۇ�e�����c��>����㷦 ���=x��<�
�{��TEr����.i��0f�������P�!�=�.��K)d�&�*�!�S"˘�tP����;? �>B|\	�jw�t�C���qϛ2�,�5"�\2�0M#�z��E?՛��[��U�
��$l�f�cl� �s�N.�aFJ�IZ!U�/�ߑE����΢Õ��v�2Yb���;>���W�m̍���";s;�*�6���EƸ#./G��n�!�%#�������lo��,�3�Cc�������qk���Xi~mW%�����̬]����UL��_���*� cv͸ ���z�����\�m\�U]��?K��)(;F��<~���\0!�d����?���j�������s�W�Lu[�A� Q�%���*k�d�������6�(�Ғ"���;�Zgٸa�ݴ�9	��T��]���7EꞾ��{�f(���d{TE����i�2fǣ,��lZ�(���|U�>�蹛̤�֐6V����.�J�lg�w\�Y^8�����M�ݕ����3ߊZ�/�m���U��7xi����� �\8�W�ke]�ͫEFw�q�'3�͖+]�ETW���4�R�|���"�oFb�%aX~x�/2&hW���b�ۚ���5{ka��6�l���ݪХS��Ԥ����l鎾'A(�o�l9�K����?P�{ [���
�ŏ�)�����B3{���f��<	�;�Xr\2��ʗyYO�����J3m5>�j�{Oo�_?����Tʭ9h�{#�:۩΢�q|J7	���do)�-����
���i��s�d7� !$�^N����X[�o[/,�f-�g�K˟�6%�,�衁<�ʸVS6�>�����S��Of�h3>dkϹ�	� �?������H�gz8���L�.���s"ƥ�\�O�Gx���,�暇=�ܜ��h�5a�}��/r��)���g��0�s-��k��Fu6&�҅hV|NJg׋T�r����B#���ܿDN�x:U�{��7D�?�lx�~?��Yi�0|��-ݐK�e�#�3����J�}�	�<KNVC�%���F�:j�MKن���� t�F���m5�*b|RO*)� ^҆e�L����: ���=����`��p�H��D�s����}������ogCV��o�q����K��'a��M����)⋆$�K͘X<D������F��uӅ�[dCF��R}
�,�F�#3dͅU���F���)��>��Y�����w^���W��-m~�i��c3';�s��SS��mrb��|n�?`�m}���m���2���	��UM�^^6ӽ��v��  y��ie��Cγ�1p/9�8�,Y2?��X�K��@��Jk���z=Xb���:\�4�X(�`�S�%zsw�'�o&D��h/��7�pƼZ�$0�W��j#��|\{�pHݺ�6����"��,M�I�D�/�!);8�͆e��E�h��IM:��zH[���s������gPh1L�t���g�$fQ�e������d۵TK�\K9�������5Y�,���z�Y_�ĄƼ����d<z({:%�bO/��\�_<�ڭ׈���+��T�5f2+�m��]Xq�`��^0��g�µ���4����&�=�&��T;E���s�-�E=ν��S�Ax)'��Ѯ�\ηc&�׀;���3&���-U�`�@���N{����)�/ eBj����/ؕe�%�EhICʚ�����ꩍs-�$'�4�F�GD�P�S�;/>%����]Օ��1�%��J��{�h�y~ְ�H�3���c�:S�d4U%R���}e��()��(�#�o��'_u�]�I<�t�p��5���lj���������ͤ�?Wi��Iݺ��㣞�F�~4�a5���Rx�L���o��C��I��]���g�3�-���G��2v5g�(�ЙN�V-)�2eoj`蒲HC�qķڱ ^?o�t:��*z ʽSa���)�Rv���1s,&��v�.�t�Z~��8���Bb�U*����JPĀ���K>s>l �B���������fgg��"wj]�*լ����CoGk��EL�>�i��:;�f� ������g�S8a�V��(=���L�uP������'��XpYlqwY��5X�����	�aq��n�ɛ��ݷ�f��fjz����ӧ��k9�5�J���
�{%�}��Z��*��`�r�
�<��2�6������Ѥr֫��òvlƧ3%�]��4�3Nj��Q�OR���4����P�o���x�����Mղ��v��N#_D� 3�D�e*�f�5ط�qtZ���9��?M��7��ZF[Zb�C���ԓU������33�I�6k����㲵�����d7����z�RK�Qm�V��(c��s��.l�Px�66	h:-h6ڹ]M�6����>�㧞���9<8�x>�T͝����.��к�pv]�[v46�;{��k���3ۧ3����x?��h:Q��N~�t:�Q���Ժ����M|���2�^�L��>+å:�o��L񆼌�+[�Vɘ���}�+ц��G��KH�Ӡ����Y�ϕx&eZ��t��}Mi�Ţ���	�����Ut����:]fK��M{J}�����u�뗨�������M�}S�������q����G�P7G?7G����Y�Һ^K ��/�2P�0(�ܹK��W.��G
�'���?�X �F0�����>�3�PH�u%.��)����+��|&�x���\ބu�z���K�4o���<�=�|���x�6]˿��Z &���8)�𨎉��J{�3�,s��d��6�
��f^�T��,<�B0@��❷���<�1�ohy��7� �Q0jU����X(�U��Q�/�Lb�����N���(G����s�\:3V6��|�V�ub�{���>��oV��]Y33u�3ן�/6�����T�(>��H����T���s*�x�R�ܼ��� ���61�l���.�m+�I����Z�/>��2��+��>��g���`a��H�J�}�C�3�8�oG[If��y]��#�����ۇЌOx�n�L1�]�;�k�������/�e!��������9�/?�N�~���F������[�M_O�䵩�<��Wx�E?��F|N7�a���$�_��P_l�8�GP/�G��J���'��\��N�9��o���th�� ����+��Nme���Y���|�bs��bB��(;J�k�7)^~�i����K߬�6�X��(� e*�B�e�1.��$x]ǰR�7�Gf���/��S�������'��8yB޹$Jbʄ�bJ0}	�a�z���6���=i�tc9������j2F�ʧ,y� �� U,�y����a��ԡZ��ő����22��p�0��[��T8kGY���@�%��;n@9Z�O�ژt�x����1��:��9�@ �����wfA�c�_d�3##�pm�8Qo�OS/���1��*����e^U��W���d�ּ���;��^iV�\&�0N�۴���U������iA�+��ާ�?֎5sn7p����%��_f��X�!_5*�z�G�(�EV@��'����w��P�N|U\�i�x5Ii��by�q�P�ʀF}���,�1_�N �P"���@�S�{���ܰ]�P��S��뱒�����Tϯӷ��oÌ�U	����k���8;j���/���C�We��Ax�+���%��=�����˼���ɧ5I�Y����i%^
p���&Z�W��G(�:K��� nw�����4�U�<�6{����^U�k����K�er��/ ��w���vL�%ML0W|������s��Pz.1� ���+W��W�[[�u�u�+�eÇOe"٫�����l��+y&�56X�c�렳G���w7��T��'���P�����������B�8vg�P��`��F�ttVD�//��/�+�;�g��q�U�9���W���U�9$�?��g�ꃢwL�2�P�4�Ƒ� ��i�%.MqV#g��Ak�|��[|��-�<2�� ����E-^t���W��Y��69�9V��
����P�|ɘ�>6�rmhpa.$듻q�����?�[��� p5	[��ӵJŗ�*g<�/@r_�+����2Ő�BM�Ae��O�䌰�D�0���`T?��W]�������g�2�TT�&
�B$����xB�:yEn���*���6q��},tD��L�}N]�ih���-�ڏpuy��꫱>S�ַ]�:�񢞾6+��[kܚ7(��~�wBn������~3�~��NKOǕ���Ĵ$b�~�kaST�����xM�)�پ~|'<�2�u`�vٻg�������"�8*hw����U���Uyfl�\�o@�׸w��Bj��p� 䟸���]�?�����O���J�z������77u�o�� �y��)�����:_P1:�r�����~��i�B�`�>�� �ywm�K�>@����1���ܹ8�ef+C��C4խ�y8s�.��D��ŌQI��QQ=��b句B�����	�}��*J��h�/����#�&Q�?e�Z+m��v�����u��zx�h;|��o5S2˩���٭,�8��u�[c�qDpF���,��B� ��r:9�w��t�-?"��v�H�j�� �C��t�!?�ڶ�fo�O+}�}fcp&���|]o� G�9F_�>t�P�sl�^W��fX�}ڄQ���Vk\܎��b\���}��rr�=�ژ1nqD�K;a�2c����rMU:r�9�ӡ��c��6�a�JH�[�(��i����i��K�o/�31A��~�c7/"7��s����w��m��K,�	�>�V�]��S��Xn�)�� N�M��S�c,�x�~�i�� ���>�ߏ]�D�����!�"̂T�b=/���^H��2zWXp�[�C���Zq������"���~_�����x|Ǉy��������m�Jdϐ�db�1����iU�?�p�����:��V�d��rڲ��74q���or�=�Vh�|�V�J�I�s�N-�d���l�� ~`��k����}_�X<��S��Z���(!�5>)�\G#�eR�������3!q��R}b樧���~���.)qa��BY8γv��=�?��I�g$�(�t��3�h���П뢃&���Y������*~�=U�[6��N/�M�KP���]C����gi$z�
�cɧ������VJ�m�iOm���<pnT)�����{5hV�?_x���Q]q����G���#�3��+������D�����d$�3d��HQ�o���.�0@�k���F�~o��Fk�f^��?.{����),b�����ip.9e��� v�TG���`�/r0f�-6t�U���t��\#�*���|СYm�\Cž���9WS�^�(�ݥ�`��=��w����>7����̶����ӿ����:,��^������j�}����X���x���i��hg��f`�*�%D���j�K��#5�`�N�#Q��0�HH�M��ƽ��f`%j�C&=g�\d����]*��E-z�۩�VO W�?����@�d�'
?fq�!��[��	{M��o3��'G>�(���OIuvꡑY߫s�!PuH��0���`��f�4�Pj��S�S� �����������z��B�p����	���g"��Tb��;�������y{�+�,?��ݣ������TxjA�X� %��,�h�x�a�m���b��މ|O�{�;��;�ԇw�^߉*V��TDj����T��Q�(�B!��3���2�W�`���ئU\���HnU2Ns���%��<�x�n��)g�n,R+���'Ć�.�Ѧ�/rq����\VS��hK��JW�C��)��g��rsv>��
����\~C��F?�秼��'��z�d�T��\�?�_֡C(��p.2&��ZS')q�C�Hh�~[�Vm����mx}��M3��f���!&/�N�EQ�"+�n]8����:ѿ����V�.'�F@�,8.]v��!!���e�M��v�~�ks��ʧ*
��/Z\|Z��¶�[[��y	�t[�����l�c��1�]�QR�9�qcf _DX�1�ᳰ�P&}J�@Q��`e0�H�1���`ϳ��#��+;�>�Rn��&G�kH�2��*!3K48�	nW�[ ��J��nEƾww�(�p�^`�?f��b�7�9V��Tf�VU�$��[���9�:�by��á�^a�w?L�Ǯ�U�P�w�Zge�������C��Xq�\�}U����H����D��m����Q�;#�ۖ~G�8�={�#�>�:é:�OV���g%Tl�p�v�����^䚬z*�~~O�C�޵��ҽ��>�'q�Br��E��+�H��Rl��g�S��WY^��ۀX�<�v�i,��'c�Aq<@��D6EО����Q�'�ZC����	ފ�������K����1ݨ��1�W��?WQP�[X�=4�����^�4��L�G�A)H#(Rڸ�c:��EbZm0$K�1G����s��z�h���l��ª�@ȭ��I	%����e�5+5��#]���H!2o� +n�Lw#�g�f`�E����
�U����ż[/h�5�R�(���-޸�[�/^�����:n�)��g��,K�#����(��F~����_w`j��{C\+,�C#`����΄���	�\k� 4+���T�%g]�������]/N����y�QϏ}?�wM%sű���sYw�B�{ }�� �}x�cV���'e�Ϡ���(��@���w
�
��6��󳖖��f�r	T�8�sb&8�N�L���h�#�U1�0B��e���K>��%�$�Kޙ�������-þ1�jWS�4�����?�Zn�B\�r����x�,Cp�{w~��$��t���|wE�������q�ש�rcRLU����4�����϶��{�=�
Q7��E�L�E�ÅC���Zә6��4e�:����&����dk�r�����;�?O��Dk��*xTb4n�Ơ���� _��;��Ujt���7U�|�Z�S��W�S͟GSj�jW/t�]�]�3��'�W�SeN�����pN#x�*��AȈ�/HKx��R�<���"^���/J��U������4���C���]4P�����iX�Ev�>�K���'���d��������-���>*�c��=�Vg唨Y�l���y���+_��5<�Śk��΅��u}��\��g��>@.��^T{9f�4®`�N��+)��C$����e$&�n���b���3>��M5������;yDg �_��-�Y�4'γO�\�!iv��럐����a�m���l.���J9}@A���W=��2�o��?�����j��e�u��:!f��{KgR��������3(X%clP��z~�֒� zS��Ւ�.p$bn`ꌇt-EXt��D�(��U��ӏ�����8�d����_'��i��|�;��u,eI߮E�`��%���L�P@�Я���!Bu~#'m1S�y�D����*�A��R�fA���v{J~��������Y�4؁#dC���Ŏ��D�"����"\�Ӿ�U����E�	��1%�c��5;���6^�c�c,�:J��	�Q��y��jo�v}�4���)#kM����h�M`e:eK����H٩K�r���,����t/��x}Q�N��l�s��ɻ�I4	Ŭ}g�]1=l(�����EJ|�e����xK���K�"^�����œ�蝲0FGX�������	�H��lHJW��/6r����~�2.Ah�۴���4ӝ9v),�G��!JK�M+��H����R�gl�ڷ!�� �g��o1K3Lƚ��ɴ��� �sz����s�W��)D�²����������25������o	���i��}>�'���G;	���qt���@Y���\sS��{����5�=���GIQ�_�Z3I|�d�5
���cLH\њ{�1��"v�����V�u��穹�b)�[��>zakd�|V���}�%����o?4~��O��]Vm95C��yct;���Wf�2��!����彔�+ȍ��{et7��I��2�k���+ց����m��.���a�l��b3��wĨ�9����l�������E�\p��pvN.�����҂�57c����,Y�%�-c�h�Nqƀl�,j�b���1;�!Խ>���N\�R�
�:J�ʮ���sJJ�g~s�Yf�B _l*�e���ύ��}|��s]	QD-�����?%3*����}�HP y��w�p�
�&F���J;�RH+%�������%ʸ�6�(��x&�7l(^@����Ҫ^�Zm�����qف���)��W�mw�Sk$�.ۉ��r��H��WW��b_b19vZ�~���ߢ���V#�)�-��OJ1�ܢF5�ʎ�C��S�GfGCs���<�/�I�6��z� ���I8�߫�-jr���l�z� ���"g~_p�sMȑ.����Dh.j�z,��@0�	�� �
�%!k�{f��\�HDJKf�?P�J�y��M��=�:�/��=�шn��_n:ٝ��/�]u�����}ʇ�В�������A�fCO���<���=�x��C��!���X�d����z�iЊq 3���l(���(��1,ژe#������- �~uҀGL��he���&&L�+N/.^;�(����\HI�L���O⭡�N�����헺�f����N����avL#�`_����`֊�V�)���V��)�z�����]�з������V��+J�f�j����e=b1Ãy���N��ѲV_�2L�������T���N?8��w�>��{�u��>�� ��
*���x���,X��I�E�����LB�G�81�8b�MR��i�Ƭ�D�߀�ʂ@+y?]��o�rE�M�s�M5����]B�('U91�y��9���B��G�)�4��^��?��sY����9��*8ʀ67���5�Ӎ���E�mU���dR
TP�;�-��. /&�x}���<����p�:��k�uTL��<N7���u�Zkv���:�U��fc)nG�����6�S���eߦ9�����D����|����Ᏸ�2w�IM}�����y��y�#H֠��9dWn���񴨿'�~I��9o$�p}����͂y������a@�F����ˤ�ߌ�{���Gn�?&��8?�f�O������b ܌��a��A�i��\��(߸�:�Cr����4�������_0<S��j�	2���>�����$��G������Z3h<���N��K�~��^�]�g���E���Ā��Z߽_A���뭻�����l�ف�큿_�����v1�H>�ru�ilߒ�����W_��V<-��p<~�w�\@��)���I�T3��n�ރ�l9C��R��J�0}�X�Fi&u�z�+b� 0��$�`k��>j��H�&☇��4x:>�i��i؛�r-���g'���UD��'�:[��յ3�I��F����}��-�����%���)Z�UI)&e;CtuS�Z�I�'�-�7S6���nɼGE��q"�9 74~ RdNm-c�º���,P��u]f}�vZ��U2�0��M�B_�"�ŅX��5d�.YCe8<V�N���[~�Z�Z��AMo�Aѡ��y���Ҩ�����KN�K=D��}����Im�;���S�4*�k��t
���%��gbm~����e2�E���*Y�9���Q'`��b�-�3N��&YK|��`b���4|_����L�9AY�p���2��Ǆ*�闳"����R���yu�
{�jy(����K?���
�i�b�'�/�V�ކL?ǔp:,���8Zy�[㏼U?�x�d�ľ	�V�c�|J�������	�� �`Oa����T�T��ه���M�쏻�:�ռ)�m�$yR�U�I��2��b�Jx�`�}�㭗��Q���)Ǹ�LlE����.��R�d��@^q"�P��}2�4�T^�EN# �st1�x1� �������V�t�U�����1�^�~+��z�ϧ�S�<u�JJ^�+���*���~o}�:�>����p-%3U�(n��v{K"�����(����O�7��c��c�A�M���#���?V7�w�Yٌ�D������<B�3�A�/�؟q SoT�j�P���蟊z�o��_�� �2sS��噏&G�%�9l}�ڇ��aO+��(�L��-tj�#j9�\Q����j/�>"��4���ʽ�s�_��W3���v*�O$m=Qv1f�`H�ITQ���̞q�պ��/�*�-����B��&g�h���|T�D�SO-8$ ���>2<:�9j��Я�����ёf��q�C��\����5��.:�t����8���!o��q�|%�r]�a�/R��
��s@Z�M*')˻Κ'W���·�]�t�ͳ@���9�aB�
\��"cy�F �39P2A��P\x�C����Ob$��)���Hm��m�R���-v�5���l
b=*g��c�l�۲<��(C��9TY��Z���إ�-٥���0ar�%8�S���<��3D��"At.����C0?��$�G໺��G�e����Z�Y޼�,��d�S=}�j8[`�3A�)�ղa)���'Ig��Ӑ�Ч�t��	��Jr-Q�[���C�ǅ�PY̽��o.�y�6��֭�'7�W{4Xcةk��3��,����M=����z5v.y��-�VF[G�����K��k�vh�f�O�2�,G�-����6WO����W	^2P��Q# -�c��Pw|�J�$������_"�ط���8T
���Y���	��5 hpi����b�{��!"�ܤ���Qd�2��ge�j����0`���CyA;��L��3��NO3a�6y��'�5�I�Y��c�������c�5����%�@�B0~�	�>�D����E�D�m���e̍���6��Ç�[�J�l����~��RQϨ��h��RM?x�?m�&~t	E�UQ���h��C5-)�����]-��xA��oA)T��Tϟ8����6� 2�w�Hm����o��T-ŏH���Y����#�=�f�	���{Ppn��>�3��
�w2�ϦU���b���4)Ņ��s�6Fq##�%���4 ֣\,�n��֏rî�������Ĕ-����qq}��Σ={[�N��k	�)M��dr�6�8����W+[:		�؟TU@�(6��_ݡ�gI<�c�E����CC؆Sr+�,d,��K�.x��C�������_���ζeĥ¿�ai���j�}���:�ѯb�_�է��,�.H��3�N9����d@�A�Qq���6��^�j]�t�i1����ܹ�_S�2�4��4��{�A�?�X��N��G���`7}W�᳃V�� �|�MH�X%�������O5_}�!���+����u��.������iI�z��?�U/���dh0�/�$�V4HD�q(� �����!�E������y���!�;�\�-0�v��C�#�17y�-o�Ld�{i�̊~�I�>���Zb�s^u�̜����܆����8��a��*��ƥ?-�l�E�\�~;dp:D���Y�����J�|f�zs��`_Ҽ��qrZ�T���}ݼ�x��g��G��ekܞ����\����z��Ւ�9��){iM����?Ms����N�o��DK�'����Z��1l��Ƹ��M�ؐ``�Ƞ�*��Lμ��i�����5�Sߚ����P)�g�˼2w����?8����B���S�I���i*a�MSZ�?�iS��8	��K-W���k�H��̺�2��]��43h���������y��n����"���ɾ��ݱ?��ߒ����$�[_����3��f��Cr�n�;�Q�ʽ^���-?��`������}��<�+]���u}��0�ݛ�e�cT\_Zydڍ��79��j��[���v.S1'��+?/��ȗ��z(<v67??��妥��d�%��g]i��Ӳ�<��Ρ��C�j�Ǔ���'�~t��]�1��=�]c�zK�apw�������C?�l��X����3��8�[mE�*f���}N��=��8�j:
�Ɲm����<����wOT�p]�>~��P�=���=W�@���U�R�-�u%[ʄ#��ai�y1���q�n5֨H��a2�n!q��
�� Ir
#�إ"�ŴRs��J���\��ж[����#eM4kr[�,�g[琭�����!�zh�~��g9N[�eP^��u�������6�6��u�5�P�Tɘ��G>�����_�z�0�l�&Oe����ˮ@�t3D��~%��n�:Fw���o\��ޠJ�Q0j/�m`�CYy�:�\����G(�+Ĩ��B�.�k�`[�m��oxm�b�K��|Sjuf_}���Z��x����ޕ~wn����Q��qW��C���t�'c7'��!�{�D1U��䡘<� ��Y��O�l�^n�_�S�ˋ�o�y���@���,ߴ�+Ep���ANx_�rJ�����ɥ.^���U��cc�Z��?�����W��ʠ2JT��K햃��7J%�co���y5���ZX���f��Z��y�I&攒�1���ґ�t�3����	�A2���AY��{_]~2�L�����m��D6P���B��2AN̡`ˆ��j������_��Q�m(����a����S>ua��M���pe�"n�ȗ�bF�\�&WWc��<��R�Ζ��}E�O����T�E����0룖,����ef������P*��;�o�]�/����W��.�	)���>j9�5����C*0���/�rve��B^"���g≦9��1�a�M�O�q5�A�z?yZ�ޖI��Mec�e��I�.Q;��y4s8%A-�7CX�	�8ٞ���}����F9�,��e�A2?mIN���%���?%b���H��Fk����L�5��?�՗6����Qn��]v����͟:e,И^�5��J,[��I��;.�b�c�<����`��g}�}_�;A<����+	y�1V�F��,�^�^e�J4�R���`��|�uE�v�|�9)5��м��3��&�?Y�7fX�\c1���\T�a�e8��1p����z��W�S����]&��[ħ��dKv���H�H�\��#����'�#�q#1�����C{Or�N�у�B-_��t��U�"��ɜ� ��KY�Ą�9y� LR�Y�3x^�)*~g.1G�5.�H,ʥ������a.�G� +Y<uG���b�Pqș���X�gb�G �s�Vu6_R�Y��I�OaR�Ns7�4���yOjϝRݪ���74\/;�:����׹��tk{'>b��zt�!��O�:��/�W�i�Zu�CgQS�[\*��n5���Go�i|TG��_8c��5���1Ԙ.P6��?K�-'����2��Xۖ#�m�љg���|3qV��W�j������`c!�ɼ�x9���;�Yk�g�z�ͽ�����7��/�J�Ӧ�{�������S�1�������R�/m�U>g͋kp{p5��Fov�|P��F�q�e�ll�D̤��P�"�uY9�G�;q[��C�1E��gF*A0�M�IRp���嗣�ی�(���jy���"� ���@�o̰�������m��+(@�'pS��_m		O�GE��F]�piz1�p=NK���i���]���.�m�2ʀ��_c�M"Jw�&�"YH8�	��I���+W	"{���eee����{A�|���GH�-Bf����W��O	\ያ�-���p�9q�Y�Q�`��;�<kM*S�;ř�|��Z>�7���f4r�/��jy�!��1��T�e�0�ف���#@�V�)�{��L̻�-@�R��&���[@���c�6����^P1�2Z��2Z�Iz��(=Y��	>0�Ҁ�P�רӱ�,�v�P���-Q�4�2,#�A�DQl�w���u︤��9���EE�[8�x4c�v�o]�����8�S��v��9�1���';viqq�Nm�h�liW.I}2
U`�HG�%:�Ϥ�U�9|A;}�Z]1h��gw�J~��L�-ԇ���J�[�	T�-���d_5;@;z�z}u��Z_~�Dz�.ֹ�ݸ�:{����状����T�1juګHQb��Xuge��5}i�Л��� ��Qݽ� %�����SPjey�g���TFt���T�N���f�Pn�i��nc|�?����kU���iiyRa��Jl҄��$׊q�d)��/y^�}��^d�K��u��"c�z��ܑ��������Բx�1�~1@�������,�W,�G��G�m�~�R�}v�#`��Z����x���5��$�q�a�n@lT��Ua�����|�w��aJ���}9#��Pכ)�)�+3Pg:�y}���r���8���`& �3*�9(&w�,�!s���j9�Wv3)�ɢ%񽐀�zc�A�A��=���'��˟����v<]���j��!����^�%��f�(��B7�X�<���y�Z�v[-���rPʠ��5e�Ȳ�'�F�C6�(��k�ou:�b�C�O�������ǔr�3���D�&y���uD�T���h�׸��w�3]�7�Jo�P���h��~۴��{ao��/���ʕ�Y��V�e������-f��<�Eŕ�sf�����}��R4�3.d߂7"(��XH������j�j
m<�����>��{�#�z�ÿ/���W&���)/�G\��Y�3 �R>e�¢2�����#ӈ.Q O��c�n���"W��?��B�C�~��S*��{�OL� �P�˸��q��֭��{��1�v��(�J�Q�V}O����G$~`I�p,�B��e!�κ�{i���/D��-�C>R�$ˤ�Aőc���U_�>�����(����5J�(�*Hc,�~6mf�Y�=��K��{�=4�G�h�|MZr^'�����ɘa�5�E� Q���F˿�̇uW��Y�t��Pr�L�z��m�=L1��!�uf��֭$T �mLU��|���s�h��k��8�A�G��U�� Ŋ�2j7v�+�8�w�{>�I�/^�?�*�Z��<왞��Ͱ��#��>�]'����f�G���on+����Iup]��sf��0��-�����_��)�wU��\ܵa0���gk5��[�q&��;��4��4X�t\��?�LK��J<W�4"�mn�0d��*PяdJ��d��i�	�@iy�m0O��/X���̤>\�����+�y�q��v����U|?�7u����j� �Š,����q�봾;����ż'�nD�F79���=��Z��t��E�������&JQ�eIAUQ���sad��C(�~���ʝ�J+�3����	�Ì��
��a|�5V���p���9��^"�:���KFWu�o�Ď����3
��aN�nE�Ks�?�C�-C�aC��/r������'̒Y��.0f���Mc���n��`�-z��#�=ށm5g^�fz��� ��nn�́����S��{���P�d��ӹ�~���)܊_���� ������@�k���t��s���c��uY����*ISr$(�t��7��v�Pn	[� D3I[��Q=E��ZZ�.B-��a��?���rpfT���*������Jsi���o����j8�ǃ��(aa2u,cu�M�!)yL+H!�}�a�q�(LϣrSF���A%�RH���rx��l.��F��U�U�Vq$�,M�%�)N��H׀����������f��&�y���,��P� TȊE�>�Q�#rj��UZ� 5c�1�~"m��̰�0eIH.tϾ˵E�\p�6;��W5G���T��N ]�I�h�J=�}ee�iT������F#eI���ق�ϓޕƒ�c�r���jS����&:F�)���P�ø�����9ͣ�9�����N��o�@Lq�k�� p2���+�>���� ���	�u<w#.!�?�~����~<��0�Z�c�D�s{;��}w:��%L
���C�\�A�8�5�� ­�����;��x�7s9w�E��y4�WAO7b������� �[��{�y~ p�|��EP(�Y�:*�IO�	����8�t�G�P?}b�PWW������<��V����Z�����%H��[�J���~��"&�ff)p��P�i�/)��Dהjo�p/�	J b���2ￋtTDɽ�O��GmyT�x��y�IG�[��(\��8�<r�������rf^����9InT����Կl`��yA"O��w��8��7* f�nX.�>�l�@/,�����H\�v�zK��:K� V��A�owY�hw��R���3S�N��.ƾ��~w5v>:�Ynu^!�$���Y��dfk��0w�$�O2�|.�a(E6�/
�C_�����Ii$�񲉉sy�w�����~/*6�NH���Y����y�X-Z�a3L^�Vhd��R���`o��PHb����Q,.$,�溌g�	`a��&�b����$M���#)�xg%;����n$��fc���8��ۘ}S��\�c_�NL��R��r��1v&d8b.E@k���Q�Z�{��A}	(K৕����������芩���N{:���3d#��"�`_��p���N�Hf�;R�H�w��1<�v^�Cl�٘�a˯���n)=V�S�Q�6rz�k^���ٗ��'�uZW�@̿Ut��_��gP��R=GWPo&?���O�-y��9=�{�K4�K8�4���?�߇<���˿�����A���vN^���
a�[P������r�� ����?_���գ���x��۝}_�����)9�\���.�\�/�Kѹ�O�n3�)b�g��[�B�â�DE�b�U�M"Ŀ�G�0��VF�rVH�emO����C�ҩ���p(���?��������O��]�a0ft�g�+DGb��	�	�;?���|Z� ���@xa��d+*�4��p��QkGq����Z+�W�#��� `��Y�6DƆm*���o�. ������{m9�ۑ���E��*��`3rЩYl�8�D�
�@��lF�u����J��>�:}\��)3 �1Y��/}�X��}[��>�|�
����v�9 �yY*�vdHkj�P4ڤv���v���vzF?�����8��p�ζ��k̈́�H��Co�Ѓ4���Fz̴�
6�R��Qq��o6O�mͯ��x�⽢�)����J�3H�˾5��.�j3H��js� Խ�CN���h���L�إZ�Ü���&�57ݫG�y���z��5�h����+���N��EU�\T^2p�?h,i��څ���/�Pő�b��"�����Z]"as4O�-/��[�����R�Tl�B��.`��^�~X�h����14��U�}���px���Zj7ҳ��F��M�N{����8Q@-�"�p�E,?��;���̌�{E��y/���
�DCi&\5�HKx5�D��҄��DE��fL=5�DRo4eY����Q��^h���$��Cjs��J�J��m�u���N�M��C�E&�lev"P�(�H�>�ԛ�JQ׭���xvK0������������� �x�~|� }��)�;*��s�򂉜Yk�q��.T����Z���V3�+��0�[{.8�O�|���jѯ	�Ua�IG��eݺ݁Ǹ���r�=�D��XZJ���(5����ϴ̇#�������z��ZϞ�ؖ]��9�َ76|:���~Z�c�4�y܎� �����/ng���K���=d�W�u��u+�4w�&y�0��p2P��.�}���/R� Pm�P'_��P	;`�����g�\T�����S7l>�:C����""�����i��\��8��OSqn�e���u>m��";��i��+e��et�?%�+��>%���I�n�n����M�Z�<y��P+2�v�i�� ���B�G̙�}��)
��w+P;G�Ȭ�b�;�� `��I�û?���f�[Bӈ�}v���0��y�6P�LA���u̚��z}��g��c̐�Cz�+$�ݠ"���9�i��oy���=�d
��$,�1�F��D�w��*t�����$�H.1az �����y O��ZM#�BƏ�b:AX�OGu�b�k�x�ޕ�Z�����W�^���L	�X�r������VCQ	J���B@��!z����b��G5���ց��R	���炤�?:�K�zK����b��4�Ϻ�(=i]r琡�p�<i��]U���@\���U55�vZv������yi�F|���3۴&���Z#.�FG�~*��UvU�S��Q}ݘ��fr�ez�cf��75��Qe��|geȖ�0xu�t���Jƛe <eb���aO�����)��	�Q���-���� p	�OT^x��M(�q��Wze��>�`u�'�o�G�~�+MM��W���{35�����?�z��t:����3�L|OX��P���� �J��I ��A@��09��Qi�QS�aj�t����⼬��j��D�k
�/k��L`t�J)[�[&3�Wj���L��M��v�<`�!fj�WZs<s��K�_7�F!�/6P����pp����
��p$q�\:�jP@�^����U��x����Lw2S�b��[X���A����SS�C�ljD9*�V6�OLC�)f���P�����5�Y������2��"m]��4����!x�6=m�5�F�QJ�BS
�I��<Z���h`��25�
� pR�yy���{G*�P�P�pB�A���,�k%�d6�^=��4F
!��D��L�)�d�T�)4z9f��z�B�!eҤl�B'D��&!�"̞�X���Y�8e�WN���_�ԔW�9�*�\cC(��� �]�6����tD"��JF��eR4#U��������HD"�2�GOz���U�i���y(��R���蕙�(Y�'L��fR����̤���aj�B(@�#Q(�D5���ҠRp�0�UJU�Yku�-NJ�1m�8r��e����h�^�T_P_U�\��Iq���U���.���w����^�zS�M[lc�L��l~UL����ik��YrV������0�4­/�tx��٦�.r)X��/�ŭH�F�y��^J�W���2�n��Tv�|������}V֋¼%y_f�2���C�}��S��[��6�S���>u�Ϝ��o���8��9u?��~�������щ���4~g3�֬��	k����@�05�*��A?C5�15 P��杨�� �?B�o+�o)������Zu�@��U�~�t|;�$���y��w�h�s�~�$�ȰG�H}O��/A Īb�C�W|����Lu_��S!����(��Dj^oj�k��Ow9�C���rWo}H��¯�^�m2�0�����ړf���>��vy�M��$5ryM3'�n�%OMo�fB�JY3�+��Gx$Ü�!vi�IY�W��lBԈ=�Љ�l�̦Q9���	"+B>�F��|�����-��pBn� (�Q4�יlV��iw:l6��br�� ���[�63Vc5pF-���Ƥ��6 8�0�^�9Ra�-�Sp ���.d$���*��y&5��5xf�;��kMs�l]���k�F'45�Q�Ff������M�)�aX�����C�Ā�����_zh�u�"��{ 3� ���j 1S�5�f�����j6��e��+��^7���ڿc]w/�2yLt4�7��45�n�:�}ف�sw��zj{�ٝ�^�(|r�x��Oo�pf�8�Q�%Y�������JSspi�j ;��CS�s~X�à ��gq�iV�XX�}Aٮ`c��E�WXTq`I��%�5�XԼ���cj����a�!��$�)�"��	������s֤$R�i���q�H* 
�T,m�W�&���ݹ�P�5p�bL�ĔM�;�DC0�P��".[i��X�DȤ%��t����˵�i���u��u�U�yUܼ*�e�k��u�%��e͖�l+����|�c�0�ˬl��]=ҷvt`��Іq�M"����4.gݨ���aVsxt��q�W'UߙZRݝQ���֗<�.zX������(�75�9O�"�"᧡��������(��^'�+�O[�� �i�Qp#o��-��}�j�#�僡־��٫�=�����^<��_x�ϛ.�z�[?��욽���r]e<���( .������g�g�U�2��3UW��)zI���&V��"��b`F����aj��{��aL�y� MM,����9�w��9�4g)�����r��@Ss�B`@�nT�S-ީ��)��Ԋs��Mݠ��u��.��iJs �oQV�R��Җ(�*��*�����s5�E�j�[i�W94K���zq�6s�1Y�9�,�l�M�)&9��Ȥ�����gz�^j�����d?Ϥ@� ���"�M+�O)r�/t��s�e�+��e��Ң�@��{=��//�/��J�å9��\Sة;t!�6��	� ��W�0^'�Xr"������HM���5��٪"5Ű��f7���VzӠ���)ɉ�i)�)	I��A'M-�J��T�uD��5`��H�������-�7�mn���4�e�S֌��i���cgoݺcČ�MS6�O\W:b9��ecVU�]W9n}���U7���X;}]��5USV�L[�غi��m#�ji�	*Cڶ@�gn(���p�"W�8g�w�(ɘp��@A��S�Fs@�uh��6)��`�4�3�#&�N:)hj*���(�nLͨB}�e�Zc�V��_�^��s�-����M$����:oj�"�Id�qf� �S�����w��^S7SV�����Ԁձ/J����������v���3A�j��=�W3��
؞�����Z�����L&M�����K�h�}J��ۛ��~�fj�YF���4��� ����Ȧ9$��i`zX���5bD6�LwG�L�Չ%,`Ri�AO=�LO�k����Ֆ)��֙��U����9����S#����Up0�����.����������	T�����aH4W�*�����_]����Q8VMMr|\�/��SSb�d��s�ѡO��25cK����պ�����&~�Ә2}s!W�˖��/p#iђz
�Q�F�Oc�(��15�Ϋ�n�pb�&�ibI���75�>��c��ٯkj�,�������V�`���r�X#Gxtrր16B�MAΚ�9r[6i��!������X�-���YO)�(���R&,c#265����1޼aO%c-�:���R����.���H]%]a�(A�@�1#]����O��ZBm�n#�5�n-j��vRꦤ���q�2p��2pāV�83!##!-=>]�*T�*q�R�!��*�$PL�FAC1D�(	J���8=�32x�h�BI2N)�̜t��ɑ3&���ꪊj˵��Fv��a2;�f��l� v������0S��@\$�"Ycg��X�����UL_�"f��Yl�kQY���"�f{�m����I�Y�i��rG�g���� K��u�̽�y��!��7����cv��������]���;~�'^�N�s����{�d���У���}ץ�'��W^˿����x;c�^8/<�n������~�����~L�?��?$5?�0�����0O����fz55� M�;���845��ɏ��y���R�
�Ic�4?�6?�6��`�)5���Q���x���FM�C1�ej��Er�C��X�#U�����{R%�51Ys��S�ل-g��%|O�{d4=�Z�z����i_���A˨��X�,�S6�w�����6��UY�lf~.='�nͣ��P�r�e��\�טHwY�5�2�/镶���\�Z��Ҍ�T9�4����(jj$VTf@�Z��T�42	m>)��F�K)ӭC5*��iΠ�8�v���rZ����pZ���f�#�-�.���(�`6� &�b� �^��iY�cX�f���8-�r$/n���1�B-d$�q��+|����3���Cl�u�hn�i\��it�q ���:&�i����445��v�;=M��j�aj�ס�����A�t�1S�yV!45��5�fݬ���k7��u�hj�l�طm�k�Z15�7��ڰʚo<�~�~ڳb��-���wz׬ӻftʚ.Ssb�3;&�l���	��9���KY�i(�S350I`W{�y�0����\P�}a����;V�ZP�gA45���G��Zڰ��q߲�{��l�װxjՌ1�u����q!Q���)� (QJ4�&�75�T'�b�@*�@�o�T`6@�6>D�(��hP����k������u��A�zL���YNm(��M�!#ɐ2Б9��M��/��-��.�4ͯ�ίf_���h2-j]9ܾ���5��ݯd�HߚQ�����7�o��iBd�����s�L��2)������֍
o��ut���uɑ&�{�{���*��J�,ffF13�Xj1K����L���nt��c�������xt"+�eYR{������x�':T���̊x��͡cM��-Y�u��Uz{q��֢ۋ�T�?*�}X�u� r77� '�0;�05o��oy=o��o��w���J����x�aF� �(��+��5�l����KO)-��Y��×~���O�]���oM��ۉ���ˋ���8p��o:K/	M׸�c_�|�E����=�"nd`�e�9k^�o!�W!��|<.ka5t��i�&�kf557��N�5� N�ID�\g���s�$4��\��\��\�}�y)8#�NQB&���=�A�#�»�!�Q�M��5��U��E)uMB�#�Cg;/u7i� u��
c�#iC��a(m	�[-C7�Eu�Ft�Z��MM�2�G�٭�v�]f�ۂtY�n�g'��!�d�)�\���'oh�C����>d���b���hiY����E�m��]M#}-c-K������zF��G��;k;��;�{�K�ZK:[*�J{��vVt�]5�wW��5�E�L�,�ϧt:5.�=�e���r��L�F�Xz+=����MMOIMY��3eB�I�zԢ���i�l	�)EFm�ٖ����'�]S�U_V�^\�QR�(*�,(�嶆b��pC �����B9���š��p~O��+�j(��?Z�.ꊕ���҆��-+���v����qpN�`1��b�Μ�@QG��3V�̮����ƀ��թ-Z�+U�X.Ĵa�K�:I�(�6I��OEF����ޘ���&�������V�\�m-��]��Q	~���M�g�;�C��|�?SÌ���3��A=	�a~̈����d��)�9gf�<<�$��ٟ��⣼Y
�1h�=�|�q�83m����Q@����aj@͜ 
8<%0ĵƋ�f�N�K��{�<>(S�;`�����$�f�����k���گ���*��	P��%��Jj���L�4~2�`MS�bhϚ]��t4̚M3�i�4�A���D9	hӀ���RC_�v��4\f*5/�v&L�犩�t8�`^C�b�7Z*��\����������������P(�w��G�O,�T�?���v��##��/8+��i	Y�L�J�� y�<�+��Jf�387�,�g٨r��6 mK��b&��-[ܞ#i��2@ʘ�����j�5����Ko��5_U����9^q�Ax,"�J�,"F�	S^�����b6�����*O55�S
^�������] �yG��>��'����񪱠�����1�4ۦ��%��oӻ�F��^�Po�k,A�5K���{
�b��$N��2�k�Y� S���ׇ�)[	i)�M
gE����}MQ�2_~�+�ř��d7xs=Y�����j��l!�ѭRAW�p!F�\9�iĸI.rj$.�ء"�R�15
 �Q�H��HN� m/}nFʳ���fd.��\\���<M"�_��dP��*���݅�(_����b�cs��/���m�����q_N�PHE*��f�iel�� �#l� ��I�)s�|9m��Iv�����e�ALE�e�L՛����Ԍ�I�Ԭ��WY�1�F3��H��r[S���B�Ŋ���F���ڔ�v��{	'��(��4Y����=������}����ۏ���{l�r߱��4�ߴ�޲ʿ�Vӡ��M�E�S���m�����4~l�MX54��4N��6i�������������e���	E�X$�>N&�
FL���S��m�|GD��oc��������o�I�6��1�=�x�'x�Ž��}��-�|,  o�G<�a\� hYÆ阚'��!yċg���wy�=>�Ț;p���S:̀���LNN}�jjGøИ�l�qG���V��UѦƨ�bR��)�;��݊�>���lU��G������̌�aL��5�N~�����L�-�%G��Epm8ׄ�@��j��DH�!ɐ�'`�>#{)�f@��d
j�?aj�����uZ��h���fT&��lPZ�*�Ik5[,&��h1�M��^"C�Ө�j��R��r@!Sʥ
�R��e�Xr�L"�(�
X��_�i��<[[����2Z�_d��3�&�il�����5�%ajh)��� A3�i�&�4A��i���j��l��X�Yx��cj�j��0!6�mj�������:M�L���9�c���[�1ij.�tf����������ᩦ���΋���v]=�ym��}����N35W�42���5O75�DL3���4��=1���a����4Kc��f�[^�oe��EWYY0SC���S�J��)=���ĆE���^߸}Y���꾖��"_ԣ��	��O
�av27m'=����I�`��8�lN:��1����10m��`zϠ�ţ�A'��͙�l��$�7�V6|��"tRҬ��R��2b��\}f�.�Ys�W�����bM�k]�ci��75����0��Ih&�扩	no������Z���������:�>�9��ڞw�������%o4=�)xT���t2��15of��}���߻�{~�[n�C����p_����ܒ�_!�/�"F��I�&���ץ�����K��e}�g�]��z�/~��?�x�7o��n��'����߮?w�S}Fh��U��9����k8�W!�=R�Xf�G��`�Waы\4V�9k������aL#kf55�NF弈���!�*�<����4�,�a�=1��T4��\xcjN�>	�9����0礐�@_�P��e�I�7���;�C{[�I��qS�e�"8K��C��!8m)�_#�6j�Mzj�^�ЦF��S����n����5�M�m�{�P㢆��!���%�{B����C3��V���.�w���wKi��������o�-����x����G7�9��䁕Gv/=�}݉�N�|����Ƕ^8����玭;}l�S�.��z����W�����7��y�ޝ��MẺpuM��&��.��6��&��2��g������ 0�`�yn�8�,üZ2�#��x���9jQ�I�k0f���X�;?l�����B����_a̝t����^K�MX��I�1�!`���yVk��Q���|��H}NNsAA{nnK0X�t���Evg�+Z�o�*��)��*lD�ݾ�;�lp�,����L��r��MN����DLF�|TBg�ޘ����9K֚�`LMg���H�Ul\\dmʳU�L%C�S�7(���� 6���e�8l.���fr�M��ycj�13�bFP�`)>x�:�K���	�4p>�A��:��R�sf���3�ԣ��(�`ofa�0S�{�O1�C��g�P2�	�&%%=�Ԁ~� 
x@�L���f���f����z0 /����2����:��|bj�Ι3����~�o�T�>y����j����. ����NS�#h��9$n	KZ"�h/��2�i����)��?�i�j�O���rS�n��2Vi)�.�q�W�����2���*x%��ޅ@ PUUUQQQZZZYYYRR
�\.�TS>����O/�ob�򴘚�B݉	PqY3/y��'�f�Y�˲Q~y]P��6G�<�t�SӞ.��f�B;Zm���W��
ԵY�OL��2�H��T��b�NR�P�=��<^����F��45��2UӀ�4S���ff�jjZ�15Q�$�I��Nq[���Iǻ�>�3[�*й��"�����Dk�Y���:S����h�iXr[hr�t�&C�������eu۫z6gU�֍eU��zå]��޼�������ܚh���9]~��E����Z��H��0))�V�֋]�U���|:�Fĵ�t^a�H�E�/Θ�I{�M����@I����(�a�Z�ԩD2�PP\HS�b%!׊P�OH0�J�̳�t'Ο�h���2�V��h�$��KG0� �DQ.A��Ӹ���s�i�D�LQF�$#� �H�-Y�GKu�SC7f�~Zs��E+u�^�f�
jM�ןn�`������!�R���y�/x� I�_�(~����j������o"'������_\?z~�w~�efL�c����k�7]��ؕY?6�aQ��A��	W|�n�~�i�p�S��Z��iY�s)-k~*!����&�L"��X�C�bd��S�阚'����P�c��{0�M��zG(����Ǒ���(vW ���>����O�.L��'���o�����=��8��4or��<! ���u����À��k�i15��ķH�H�:%y]*{C����<����\�L������15���aR]���;�ǜ��^���IR3��) h,K@�`,B�٦f����nhe���$�vY���Ѡ!�J���[H���DK�*��~��&�EN�#k@��	)b|�@0�ll2�7P�\��j��ɨ3h�z�7@��i �^n4*mf�ݢ�Y��-X�Ng�ht*�F�T'P(T �\	PȔJ�J!V�$�����pҞ�j�eY����2��&׊�H�~�ʼ��ʘZ�T[�Ʋ��� ���P�Ś��2
Ϫi SU�T6u� SM͞'��Mä���5#yO���:T�}�z����}Q15�o=�m 4hSs����O��w��9zy�����W^9�+���15v�];�E���&njYsuoӕ=����e���bj��No)a4�?aj�Ƨ8��ɵ���5�(F�г�ƣ����[^x`E��t@�ѕ��W��gB�^�why��u�g�6�ܼ���E놪V���6�F-~�خ��"�H�.H_��H⧧p���鴬dҝ�L��`3NFZ: =5�z��iq迏�-HJ_�����JIc��r���cBl6�k�|>�$� @C�"¦��Z�Za��f�`+�3rR鴩�Q����JךJ�h��i��f55O�4����15[[����a h�h�n�k�k��iͺܑ�Rwɭ���{���,�W���:�^y�ݒ�������� mj��IS
����=�笹o4���nɕ/S��
�
)~U$�����X��D�WD�q�E\�VE�Ö�o<2���{?������O'����������3���M_�i�rMh<�Px-�z�%��P/B��"�c����2�-��T����An���8��y�����V3��yU�30�楸�y^�N����4���)���4W%��pYNsq
�L�%�4� �ԜBI�y����5��%��TtV���������셫!�Ԭ&�Kь!(yNYJr�(Q:��@��A�u�%ް�ӯa�iٴ��s{�B@�����!�x�-�sKz�PO�5 &���5���� �^Ek@������[+֍u�ڶ����g�_\wp��G6�?�����Wέ<w|����;o�пg����+��p���k�7]� Xs�ܦ���¶W^���K������{vT�XQ�ly��X��`QWwnK[΢�����ֶ`~��j�T�\��(z�=,�a���Y�GG/�Ӌr�D�F�����\�>�6�}QCЧ�MQ��d�tRcĔZ�\K5��덄ހ��Q�3�!�1�P����EE��u�ˡ�l� �>˪�8tY{�ɜm��C�@�Ֆm���z���5�mF�^/�^J�H�%�R��P��6P�^���5��15�^����i�fj��T��Ņ��"Cg����ژc���}��.`T�R���y��s38�0�b�Et�*�(��gfLŌ��A�1�7P�O�^����������`�(���Z���� �	6�σƙ3M�. �̷ �ՐB�t̛?�ys��y�Y h�M�s���p |�p�A:lv��:av�ͨ7�$R!������d�g ��t�f&��b�)�9,x���IM�HI^�p�����ʜ�y�����t��5~Y���t��jY�4$	MØ���&�hM���F?����ef�4��)����"�`�
0T�f3���l�f��8Xj���W�ƪ���K��ٟ��(iHڼ��_I~S�$�ebj�>C��O� �{�����[ F�8�EBẚڲ����"Ш����n�[��&mj��5ajJ���b>!��9VZ:#k��N�?/e����N������Cr�����m٢�\��<:Icj�K⦦T5X��ԍ՘���U��B}mL]T�x�A��c��"����()��IR#D����L(`}�>�5���ijd2��YS^|P�g˔��!�4��	�F�����E�r�!C\��B��T5T�$�Y�N�[+qh�1�+/�{V���i]Jw��U
P{*��ZcV�)�Mm�ĚU�U�UkSe-��tis�M=��a�ҡh�ʪ�]}۲-/�X�׸<R=�̩-lZZҺ��eI0V��Z��5��6����jJ��PLL�G'�jI�Bh�R�]�5�l3�5�\-�qS��yp�83���0m�I�IOKB��B�����M�TP3�/�"�E2�(�R�(ŗ�	�\� ��Hp�ġ��6�˦1�,n���'$bAB6"���KF	rR�d�qz����&��*�T�V葧��4�Z���V;��D�fj���� 53��x�'���^b��Z���n�ȶ�4�Jޡ�u����͝x������k�U�L�m(|D?G�����d�_錿����M��&Jr'J�v�*��i��=��=��M��-��=��kn�7]�o�5X��7+~jQ�֩���2�1ӂ�m��a��Q�;���5�V�)%%�Z.��B��T�3���"�H�#�# �ÉY'@�������x'�T�]��T�F~��GQ_Ä������L֛B�1J�	a�
E�!���}��->�6��5��#�����c�x�d��'�4�7�( 4����<Z���A���q���ܦ$ Z�L15��Z�Լ�$1ͫR9��P�zr&��FE/�dP]7�/��gܚC��rk@�.H����x(nj�"�ؙ#ѧ��� >����s�h��ܲ
��@�FP@�(�!q�H�"\K�*�����pc��ubL�$�0�khM#�I(�X$�:��Jɤr5�@�ΠgL�F��h�\��e�ɨ�Z�v��j�M��d�덌�a���M�B)QѾFFoJ(�C0��K�k�`%!}M���ĸ�ٷ��_��8��&>��4�k��jLqY�J�$�0�kY�9&�f��I0��$�z4!k ���=!f�L6.�e��L�΁(�	 ��l�c4Ͷ!��ds2�������k?�Yw���SwLS3���cjMØ��;��˝�Ν?����e�u]�3~��kGF�\;2t�P|����;[/�i\�����������/�YtqWåݵ��ԝ�V�ihe8����F��
O�/ �S���'�0����#+���1�&�n�� �4�L �k�e^�wlM��Յq5C��9�<7;�`��5�'֖�\Wzb}͹]���7���vV����e�G�+�������g���gR��^���HOfe�r9|K�gә�@G/���{�q�F`7��,L���ϝ�2���B��Z�s��\8岔�W���
Ҥ;�*�N�թ}�[)��1.0YV$Cǚc�<c�|�ϩ�
W�9��z�
�cE��b�P)���ɖV*�W��zU�nm�qC�ec���ٺ�չ��=���.P�l��^������h�mm�2lo����������=�8�<�>��ԙs�'����W���h+�ߐ�FM�vY�va��\��lߛفA�������~�?����ox�����N���5���B}S�xU��Iю�X}�TеH}��]��/k����;��?�\�����t����ߛ�������{�O�O\x��e/�r�
����sxW2��b&~Kj�����s~���CO�D}�+<�\bC�؂l�u��s/��!�M{%��f�u�����	�7���0���C������»,�_��k$rU$�D!%�KR���� �*�+j���LpAE Ϊ�*�:�$�K�#|���G�'��|�DΑ$z^���8zB�"�]o?s7m-/m� }%��B��D�:�$��)cd�29{�ZoD�j�cڸ�QqzU�5�[���q�,p/���;�>��&<�/��z}�>�d�K3�1x䴯qɺ<�N���#ktR56�ޣ��:+bC�����;vo8�����l�pb��+.�Yz�k��=c��/���ºW�[���5/\^v�����N�=�w����s�o\Z���5��X�ҵ��_]r������v�hع�d���=�[vn�*����]�^��3����Q�m
�A&U�A/E�Rآ!�Fi�D�x�P15S��q35�q-�TeP�B��l\�%5|J/�a�U���nB��4.�ʉ(]��-Ty1�ך!��Xq����٫�F���16f�1�&l��U�Y�(���ŐL�(��F'6e�Ԩ��L�p����clH
ZRn��B:y�I�g��D9$� (�A�a��Sj�ٸ�v^��v��.�������:?R�C��آ ^$�YҦlYk���@�Q������K��������g�9�=��T)I�H�Gx>��V<>�ǋՀ�߬#����i��D���g�=P3�c-�|����_W"t��le���2y�)e��gFz3
��>�q .[  �IzjFZJzJRr�¤�)����V`�Q�l�.\�4o. ���yv�W�<��9;=���9�+s@-`�I!ᶹj��d�,F�A-SII	������w!����t�Lz���~z*75����J��h��5u�W��|)陯,xf^�W�<�,{�<���'�>5�c���b:0�̸�z�ȅ7��7��M~�9�Z�8�5D��I@{D�� �cb��l�+Gܝ+��\�%�͗�J_M�|�H,V�JT#e�p����(8�.�ga�������ں�޹��1V��]Z%e.�S�gΟ�px��^lx��ۖ����B�W7��/w�- �
���sUV�TU���T �J�
�sss�
�c8	j����-�$ p�A��˧�մ�Hی'���>����vRR�h�>@I.�� .�@c�9��W~�\��u+�=�JU"�xk��u�:�����|qk���@�Q$�eM�f�J?\c��TY�����lc�_si�V�U'�(%R	E�(�fh;C��O9�i��3O���d��⅊��0���0W1(���F�y|�e��o�y�LA�0�"$
�P�B$��|	
+�&']
ܣ"�j2�G��,�*ˢ�YuA��k6yl���v��6��T�ˤ���NZ�
7�����Ū�nyv�,�O�3 ���R���%��mɈ�r̳h��i��yU�eM�}]n�Ƃ�M%�[J�7v��6.��j���Fc�]��o���)�;rmְ��6i-JR��DF1i�`6��&�lb�M�u* 3Ŷ�9n5�T�*�E����g������N^��`n���<[.���&�N���ej�T%V��|�
��`�DIa��R�/9�\+��]6RQ[i���H���,�I)RS,8��d
_��R��t�V�̕��%�Zn���媰b-R���S:�6�ц ��p�i�#m!�ۋz}X���!r(,���|�_�#>bԋ�{��^b}T�-G7�l��d�V[ecj|���^�x|�RSɑl�	�y�{ͨ�����`��J��t"��.��4�����~r��k����]��=���U�]����5��N�w�o���I~l��!h��g�p����+vۍӄ��w��c��/����?j�L�{��?��_�a5T<�0��|~��`�G��C��CR����KI�I�ߧ�wD�cR���K�we�{r�;"��"�}R��{��~G�F�w���#�6,�Ci��;|�]��>��~���� ,xC@�~��e�T���y��������ۈ�5���!�-!�:J�<���#��!��W�hG�Z}[��S�(�[
9.�ݒ�^��ܖ}����N��V��Nz� �`��q)���ªŦ�luX�,B-�R�1j,K:�-��X�|("f�n�&�l�C�LU6	&M"��7z�Z7
�[�$O�D�G�8DB�Td�H-��L%B�@ON"R��D�PH�(�cbbrƓ��(�(%�H&"�`7����D(�X"�J�2��I��P(&��HŠ�R)�Z�^�U���F��h�^�Z�R)�J�#��d��#ӹ�AwBB�e"�l�(
8�I��_����טc�-��n�Y�_���J��ӊ:h3KqO]扞�2�����>I-6��u͎�M�5�6�f�������������n��f�o��k�0�i2�6�`lhsL�0�݁��S3�ܝ�9;�s;G�v�����1V�}�d��ʭKj�/mڻ���֥'�l8�o۩�;���~b��Sw�>� ��aڀ��;��<����ơۘ$5Gw�'�˭�O�=���G7�^ڳ�������YtyO��djh�o�`Bi�43Mh_�{luca���4S�Y=�,8�$zxy����PG��k>mjr�9���Z_qfK둵�;�*Wu����r�9�G���sE��RKPT��80��c���������Z8�K)���`N�¹�I�i.�HJ�LNe��s�ټ?�+`qP6G�ʄ3�i� (=�HCX���$a�Z�4�z�M+�׬��a�>j҅*����<=��e�1��8�y.dN�Jj��+*'M�H�b�D2\,��J���˪T˫ՠ^Q�Y]�_�h��b��jln�oo����f���3M�tw뤩9��?�8�:��Й}�;�jO�=��:��4��n�ݩ	�Q�_x�x�󉩹�w?��w��;~�]������|ˠM�}U�~M�yMB;�˸�R��H}��^�8^�V�d��n;��}7&^��ĭ����{����t���ӯ�th��oo��,Oq*�Ρn�DX��j���W�ê�o�5|T��8Vx]m:�9�Et�]��S���zI����
�ivf*�P�ua����TSs��	������Ҧ�
�\��%��E)zI�]R�U�e�芖��.�I�958��Ϩȓ*�?"A�p�A�w8�1\p�hSC��E4�=""���`������75ˑ�q$eY8�%/�Җ+�k��:36��F��A�15}jN��ӣ���~+�o2�f�C�{	��M���{"k=�a�0����݌��Z��:.TR�7����5K;W��_�s�γן޿��%�N_:=p�\����ׯ>��Ћ/?m��+�7.]�8p�|��s}���^:`84�⵱��<w�3|�b��#mGWo��u�xǑ��kWWm\W8>�kj���Fk9���6�^oת�*�R&F5
Ԣ��F�� �kE�((#BR�'��̆��BC&�O'�鸆Mh9��G��lB�S(u\��~��+��,�#BeS�a�Szp��81�Gd*�Y�@�!3F�G0��JD/��\9��S�����y":`�����<���t�Sy[(G�:�^�*�囤�&Q�Q�k��lP�-��m��T9��� �ܵn��+����>�f��i�cL��Z�o-4v;[�QK����:�VJI	G�`��@���щ2��.�E�f���;������lڀm�2yxF�<��2��3#���[��
9B>�aFր�w\��#�Ԕ$FӰ�Ry������` |q�̛���g���_�[ì5����LJ�m�A�s�lV�٨֫�J���1a���<����H& gdB�i AZ
?5��2��<��pN������R�_Myv^�32���/�GqSL/���T�[T�ƫ�X\Ӡ�.�م5��&/mj��(cjM`4�,�&KԙMu�Jz� ��MM�0P$,��J��2`�T	��~p�@�b��I0T���/�2�W���y�"��z�h��6�eL��I�Ϛ?7�YڈѩX�'�$Ѧ��I'��0>���ŏ��=��@���~��^YZTUV�PZ�WX����%�+!X�"��pyAi'L��6����d�9q2��B�	SC��ybj&���Y�M75t0Ԃg��O�kS����Oֆ��075DgѕOv����BI{� �@9���D�]�bL�P�i��:X���v�x�b�|�1�2x�*��NZ ��ࢋ{��K\z����|S�_��aډ�����iO�(nj R( a��a�ѦFNz��_M�tҨQ�e�dYt��o4��&���v�Ψ�R��2{	�{j��E�`�<�&�v�b�Ҭ>*{��压�
�S��ą�4�㖪%�E��+}��C��:6�tn�����X�ױ.�eUpј�f�_3�˭����G��J���j��^�Ʀ�t��$٤�C�ڥ�]·KxN�,�X$\�ZhS��$��I�&<L_݂x�{;�'�Q&�)��E}�Ek�2���J��c~o���;�9eEᜨ��2��z�Ec׋rTI�lJ#�	�i����sҒ�
nA2�����ҽ"~�/գ�:x֘@��6ؑF��فf��� 1$GB":��_4�븩�G����K��F���no�{O�w��:q���oߟ���5}7:�.E���M��Ē��/4�_�4?�>'*��R��׊��������c���n�w\温ѽiӿ�.����o��?t��+��������7��c���N���FZ�X�7��jP�Y���Z����J�e�������!�W��!�~&d�G���5�x���ЦF,{��ޥ�w(�J��~O
}M��%�/�ޗ ���(�u�6)�I}�����k<=��ȷx�;|�k��]75�#�Cwa���Ŀ�L35wy�534�݆�����S��5��Q~bj^��o�hM�#W$�+��^1J���S��ɟ3Ȯ�e�����roD�5�X���L���͒��PD�Ț��h�����ajY�� 75�E^A�*�@�Z(�xD|;%"Ihq�CT�!JR '!� O����_�4$��HB H)���(���q�L*27Rp�e�0��X�T*��j�R��F��d2�(��I�z(�XJJ�,aj .+e��6m[i���9Pb_��__�ZQa����j=�]@��Ɛ05	����\���y��Ih����y������ɬ�Y39;sv�bj��Wl]R�mY��5}G�,?�{��}�N��qb��25t(ͬ0��Y��65�\;~f���W��6ty�����	Sseo=cj.�fL`��Ipf�伧��aH���O&@[�H�����8F�X��'�p$>+��h����_M'*>������k��li?�������݅=���lCYH�RCfߡ��F�M+�h��TF�?���?|灯v�����GB|�e{=��E���ŪGA�&Q-��ĘU%��1�kݦ�]��u�&۪ϵr�ڰ^����BUƿ���AqJ�"�����Wպ��9G�5�%��R)�x��	�YQ�YY�]]�gjhG�f���v���s���V�'�^�M����f��'a5���ޕ�����m�w�s�6f߯�zPyTy�z�>���iSs?���>��a5��;f���F[���пD�^&�/b�H���D�W�_���zա�n>���'n}o���������#7w��?�����CB���9��b&��z�\���oy���tQ�Gխ�j�fQ�+�Y!75�k\�u.�Z&gZX�+0z���>��P�Լ��/�M�s���������D�\��3M��輆<��k5~Z�W`Get@�!Rp�@�������1�s���"�=��3�f7}?m��J��G�I�D�2I�*5o�Yo��u���Ih�=�ߊ�촩�w�b�G2��g������-�q˻<��>U�O��V9ċ¦���>�Оumٰ{����W�ܻ�����GΟ�x�����˗_��}�J祳ݗ� z.��^9��y�������k�p���ɎS����{�t��#��67��Q�|����[W��t��[�A��c2;�Z�\&Ҩp��r�^�ī�d���)܍"Vda	,�����Y"#��p	�	;D:ʍJ��4�*"�&��C�2�(*"Tg��(��a
/��	5�'1FT�,�7��6�#��G�1&%��r�����%�B&�
�H��)Lf�4.���Y��]�
���@�XHد@r�d�I�o���p�*uA�6�S3S�ϙ��"Gc��2l*��"6�C+�HD�?!��O[	v&M�g���_��a�|�p�G���"f�
�[g+��g���O)3�?3қQ&cj�0��ё5|� @����i) �`e��Yib�/#��696399u����$�S��ԔUU��<���gљ�F+�f���^�U��bL�C(¥�	�LL g�hXPf:��&�H�%sR糒�f,|6}�W��5m�ܴg�gΝ�,�
��RA�B��%���Ma-�`n�Ѵ��f/�4E���5�Y������ILXMB�|��0��15��aL�p��!!k �X�L�Jԣ庱
=`i5��W�Y�+��Am�SC�V�� s�܅�>��`!mj�&'���grX\�O�)A`H����7�ǥcf�!���鰕��� 
�
�� ����H�x�m�!J/�
j2�&>A���J��2��!5��fJ`M򔐚y�]0g�/	��Ѧ�)-������,�����,�/�k��ru�v�R7Te���8�k�e�*��\�>��3�F��'(��.�1&�T�1��E��35����\����	\h�rK\ڟmj�F�N���
a��<~\��C�G	S#B���'���lrҩ =*��v:%�&lR�Z���1;�)H���Ԙ�Ke+;�d�j:�&ب��+b��X�4�W��/���I��ɊV(������Kܵ�ܵK�+s:6�l����_i\�ռ<Ұ$P=���WDk�K���K�C�-.��Q`1GM:�IeՈz��,��v�1�v�)�!����kS�f9,�X/f'��tVZ2��%''��'NIe*�Rg�:,��Ǒ�ym�Fnӛ�.O^��ڢ>�Ϯr��#�WUb�E�qX�~�3����C�ЉL
�(��-:����ٽf��q4
�d
Ӓ���x�<'�C���x������S�M�㴬�ѦfE��Qlwb������gj
����w_�����v�����rU�j�}JF�$����P���T�J�g�{�8��%���g�W��K���N�G.ӷ��wm�7-�GV�[.�;.�7|����s�>�����&`����7��c�����n�ߝ��m�'��*ٟ��?)���R�!&�C)��B�s)�S��e�|�!�C�H@���#k���k�MQ�ߠ�o��oIi�!F�A	���a�w��D�rz���P�!�[0Eg�b�Aķ	�bjn#�[vk��af?�&�۔���L���7T��15����P ���m���V��NqӠx�$�l��w(Nz��C�=Qն��651ɲ�iĀ�,�HL:����*k�BdO�f����la5�)��_f�ru����q-8�F	�8�Fa�R����D���b�JPD�6B!�D1 &�q���Fa8%DI! =#���k���c���܄�NpkM��+�Hd�"�g
;�MP�&aj�U����D,�!"���~)��vUgw���J�+j�`���ֲ�R��Jǘ��4M��0RԠ����\�dgL 4&MM\��jj�i�'�ƶ�s2U�4�	���&eͶ�д��ge�`�TS�c,�x�%%[�Tl�޾�y���[W0���>ڿ|S�����CBӀ6mj^�|������=�s�ځW��}^Ssu_㕽��v�^�Y���&O�4.l����f������@���5��aL��e��KB�ƃ	��G-�b��4S��5Lf⸬)=����k{z/��9��~�����2wWU�Ы��p���r�c���ݩ�F���C�5�Aۡ���m�ӱ0V�Ϭ��4��mи:�Q�ߢF�W��Ӛ*�I���6]��Zr�g�ʳ=�G�ߘ��r]�<�6סɵ+��TH��t�pnL�.2p�mHK�)6�m W�}�T5^�/�/�P,�T2q4+k���tk�5�64[6�ٷ�;�v8A��͵��?+��aL���ݷ���`sw�oO�oo�o_��@�9�9�;�8����;s_]�w{q�����M���r�g=.�>�<�z�=��A��P p?�{�u?�:����&�=����r_c~E�xU�~Y�zI�~I��B�/��紎��?���kO�~Ǖ�k�M\}��O�1q������g4��Vd�>�b��E��J��	���+�sF��)�eK�ϛz��k��eu7�γ0q*�.�s�ͽ��N55LX�ː��5��*�ބ�W:��H�Ŀ�¼|����K(�"&�L�WE«b��M��˪��'-uU'��� SM�ivJ����%�!Rp ��r ��C(�J�՜	ϋ��gH�$!܏";Qd���g��e�䥯�.�Җ����q,e	�N�h�M��<S3���k�}Zn���g$j�X���A��~Q_@�����~頏f�+z�Y�[��Ut�Ռ��vJ�æ�u�����-���sb��{V�޷���᳇���:r����϶_8h=w�v�L����-�t�y��d ��W/�^�Bs�b�Í�T���v�p��][66�ٙ32d��pTW���\���H���.��$��*9�S�@�֣����_��)$ B�B���9'u�I�@p�17�pL�Q��0i��Hu�����P���&�e� ��j��E��S�r��<�?���|^�Ì��|��-��($Q(����(y��-$R���L��T޼� ha
��!���C�N/�!�M��oA�lP���bjZl�ٶ�����Y�6�TE�?Ʊ|����3����a�#Lmf,Nc�g�g�ŭ]��:[�<<�L~J�����ތ��c����@홬1��`Ӊ|����d8�(�?+B�Q60�C/(���MO;1<�?���]�SP^X����^�Ic�+�L@��t�l� bsQ��!�3	�e�2R�<k�I�y�Is�|%}�3is�Mv.{�$e���j���d�GR��Y��X�o�����C�x�f>UӴ������S�&���ԝ+饃e�4��́b6g���)M�4ӈUM4	�Jԉ6cj��Zˬ5~]�Sg� bv�0}!k��p~҂�)��$gd�s�lx1A!>��S5�=x�Pi)�N����5��������B��zŠ�L"Ы�px�E�xT
��|f����ɤ?���)�2�&3�%LM"��15�4F��MY07e��y`������ U"�"X[�8���'�D]���B��L�]����UҚf�J?Xi��׸@Ǧ��]1�uA��mR5trЕ�1�X���.��5FO35���C8�Lf0����喸���<5�� }�2�)(��<���@	yb�/'5%���d[�QБ3|&���tۼ[�fl1�)[b)��K��r��FlЄ[4�6u�C�ե��U��F��K��K�%K�ec��q��j<�iME��ݥݛc��V�7��Y4������b�����DsZ��J���b���Qe�J���";"��p)P�v�!p�[$<��k�Az)��b��0�%)L�Ӛ�.[ h�n����k�/�h���j�Z��s�R��i�)�j���]4�ײd ��ܷ�y��}�pǊ������=͕}���m�°3�猺}1w$����]��� �b�s��d'��Ua&��F�nj>L�P��K�:S3��F=B�r�hO�m�W��%ٕ�x����ޖ_�90��ŉ�_����om}iq�f�_$�&&o
�䪟HU?�*�vO���,��y���Z~�40�����Y�Т}�4��4}�g�0��~�����#���~�ｖ�y-�D��w��c��cV�W˓�O*�\���o���d�VI)���D�c
�����t��O�P_$�!)��'>aP�����#�����d4|�a&�F:r����c�`ѻ���z��'L�mmj@�=Hp�,SsB�`�7�'���x]H0�f2UA耚O���J�
�Ԙ����g �$��Ԫ^�+^2*�3+�ؕ�\�~ա�zoL�5K�>K�2&Y/���d�ǳe�Q�g0S��E	Y�ħ���|2ʇ4��T�*�H���y.�eA�f���9rK�g����(IXAbt�a����(N�#BT �!!P!	@������Z�-p+74�j�I���4�	D|>��+�ϓb����I���Y,��
�T)�ґ5b���B����s�W̡���-��[�+l+���j�K��U��L�3	��&jf��a�h���4�$�yJL�LMw:�i�&��'�uO#���԰��������c�[�k�/oݷ��ض���l>�w멽ۿ�����w&4mj^�r���u��;�k�ʁ�����&Ps~G��5�M��I�v���	e�X�i�6GWe3s�.������������P���&V�5�'V��Y_{qk�g7�XV��3glQpMwQO�Q��:�Z��� Ce��,f-
ѓ�E!SY�V��n*�6Gk������4�	{
��|�3�g���AGq�UsU�j�š�"U��4f+�
�������̲��LD��ȳ�V���9��~�#[��+k-��k�-K+�YNLͪ:��z��E��F��&3���;�ù��ض�ڻ��L�iL�3	v���/�v�COΞv��V��&��&��f����S�����]9���ʿ�Yp���^S�Ú�7+��,�>�	���'MY��>����]��7m�G�#������B���|Km��2���>�2\�k�׻�*w�|p��7�������~�������W����;��_P�d�N����$WRы�����D�o�;ޜǾ�_���v��;��UX��|��Og�N�<�ɺ�bѲ�û����	��CSׁ�:7�Ÿ�y�45�>cj.c���K$|�^�b��9vQA�\R�W���pIOsQG1��
;�B�+�G��
>H��c\��@��#8�	���$8�������lG�Mg������Y
��AI�H�R"m���J�[�����tT����<F����A�	�	S���t@M�|�Q�O75}^y�G��WҦ&�j��*]R�a�/,lڶe���[\8����Gw���?x�P�#]�O,>��ܙ���ϝ�9�t�C�ٓ�֋���g�/��q�繫��r�v���=ۋ���ݷ�t˺�-�����.�6T�j*����"{V���әmj�A,!�RL)��*�W/da�($�Bb܏	=��^� *��H �aB����$*�f���jjb�>J�B"��T����������]yFO��պ�R�SixR%�R�	�0 2="6%FT�C�*&�"dO�@�ҐI����Xr*�����VD%���q
�����<K}��,��s�&�E)}`����ae�+@1��XS��s0=p8�9?>@���� �`��+��>=e� 0���B�C <;����F�l(3]�a� ت�n\�r���4'wQyEYn^��q�:�LM�eN����r�q)��Bj�O�:i��Jp3R�iI�)�ғ��a5Ϥ?�l�ϲ�|N�#�'Y%�-v��~Q�����>�ه���v���O4��4O���ʖ�yOqC'	f�9�O4cj)35���L0Z�-��d����a�e5�5��uցRSe@]��Y%�I�3S2Ο��:Ne~�¤������!=,�LO�C\>�͝\�!��r�]%e�E%�����������%�P�3��(⺎���j�a��YL�i �e��))��� �A/Y@όJ�������_0g��g��s�-��6�65V�m#��U����(>ij
iMX\$�P��5M�i������p�{���^�,����M�2*��B.]yp��=�'Cfs�0���M?�s���Ǚ�s91�x���lS�|�i��>�:�,����M�$L�(DB��)'���i>�S�m�f[�YVc�fX�n��n�ۭ!�-�6�T�<��@�,�y*�Zc��n����c��.}N�1��P0`�����G���ᢖ�M#�Z���l)m]S�NSҸ,�r0T�	�*�.�).���i�*ܮ|�%d�9�
pP�R�\�PR.%�V
�
ة�l2�U�7�9:���Bz%�Q�29�5i�.�=�w�f+�*{�Gv��v�|��Ս��U/�hX��{�ƾ�[��nh^��`�g����� K������/\�u���'מ>����eGv,=�}١mk��ٲ���=�<�t��֠ϙ��%�A�I�F�>��Ɗ�h�	���|���� �P�����^l؃���jo�}MH��Fn��i����w�����͉���K'><����C�r=�U�szÿ!��X���Z��.�DA�De�Dm�s��	�~�62��ޱj�5��G.�c��k~�Q���L?�~�7��k�k�6�Ldy'Bο{�u����b��I���F�G���
�IiS�J�o��xX9V�	?Đ����5q_�)�1!�)N���~B�~,"~(¿O�Q�d�w!�K�5\���j��E�G��u��6y��a��1黐�]�u!55�&aj�
>���#D_⷟D� ���R�5�T~O�dLͤ��+3��00�6Ӹ�V���_2ȟ7+�۔�\�s>����`D�;K�-[�>K�*K�"&Y/͖,ɑ��S��L�ʚ���7B3M�$�&k�|H�j��^��%,1�Yj�W̶�l�&禉�)�{��2�W%�ԔP#�U$.ń�@��G@�*�<`Dߊ��	!�!|�Ԁ��%��[1h�]"�;-b�H憜(�3]$�X΄��M��$(��3��k�]�[�/���GJ�Kʌ+k�K�tK�L�5+ⓛ�i��V&vfM�l���!F�$LMB�д�5����4��bj�ڙ�0k?m��3�&V�T�S�i����ٷ~���U��9�g��/(����4'������O�;�������_޻��05W�60�����s�+���6Ӹ�����R���f3�'����$�׀��e��c��#> cj���.��g�9_
��5LXM�ԜXStfm�ե�V��[W{qs�������m��]�]�]�}�~]Oyk��"��ϵ5�����E��B;�[�<�U၆��梡���E]��m����@cA��� �(?R����zQ~��(�Tn+�Ɖ����J|���[e�X�{$1���hu@Ҕ�l�Q���3@�te�u�|7YW�W�j���7�����N��l[�������5�X�����=��4��y2j��t�bj����	P[�l5��B'��';hYs�;�zW�]�//�}�=�vK����G�yoU�Y{������||��n:����~�r��p�ew�iq=2;�魏��7��[z�m�������u�]�����#?���z�q�ڏ��ӱ�[���,��8���K/�ϳdW��R�#��"ͻ�Л��Cg����6��ڶ����u'8�ci�g22.�X��l:U�M�05O� `�i��*¿N W	�]$h.Q�	�E���梂�a�=]щ��%��������W`t"a�05P�A�8.�O��gd�y9yV��"��B����n�6
�����y+�i�y)K)K��%x�rq�j%o�V�� �6���ȨV��Z��x���5�n��KƗT�R}AIOH���dِ_6�S �|�~��׫��+���T�e9ECEl�g�ؒ�5ۗ�8�g��=��7��wb_����g���=�~�d�S�gN7�;�t�l�3gOן>Yw����q����._�~�:��ʥ�s���ڽ�d��=ۋ6��ڹ���AOO����V[i)-�Zb1��-7�:�XJIĸ\�U�נ�U1�,� �"H`^�	� ����0.�b� 
�> Q�BD� 1TA�!X�� �	�!L �^\�F%\�h�U�\�#����wL��KMT�H�<��G�a��h!@S�� ��8�C�g���DR
�0OZg���j�Xa%�k ���SӔk����|���oT���@��;�\6�i2��D�Τ'@}Q�&�� ��	s2(�1��yS#��?4!F/'F�AG茤`�G��q (�Ņ|��a�τ����ok����x��(+�y���ŝ��%�%�9�C�b 1"$���EXl h`\��q�A��0���J��:tz5>+����N[��2��;�3gw�W���ʸ�⌨*�c5��/Z�#��d�� ���� �2ۤ'����D���r��;�ؙOO!<]� �i��ru-3�i&��q�Id��Z˺f��z�@��§�sjmR�����Rӓ��{���s,\@�ʘ����	�p>���}D�hsb�i�j6��L6�H�=�¢���"@Aaqv����r(�� ��A\����LM�d��X� vzZzrR*���%-mVJ'-���⃇����L�J_��:aҜy��K����J�g2�	͜k���D1��C��mjڳ��<��tQ��bIO��15մ��5��Z���u��Z[��,d��U>��i��R�L��ࢣ53 (��%~����l��SM��Aa.(p��W?qi���� >�H�2�y���y|����
��j�(_�C*1���O15�\�>�n���~�ݩwXt.��k6��֒����Fg��Sj�U�|�_��_����`�.ج��C-�p�'��W�*�h]۷�p�C��7T5��i]]ۼ��n,��'���i��u��D��B�
�;�a	�4�Jऩabj�J̭@�r�&���V�Q�l���d���6;#�����κ����ၺU+��ִe���c�^z~�͗6?}����^���^��Vb粳���;����v߼���+�o\�t����g�\82zt�����/�q���c�Vl]�=�]�PUVZPZ�S��U�,	8��\�<�@�O[��ycjFB�����5~rć��72�W�${��ª%Vb�K��+�/�9�9�÷'~��=����۹�zC�N����I�-��P�����;�{"7{��t���o���E=����豾k�=0k�[4o�M��w=������Z0�"h�O��Q�D~p"?4���8�c��^��\����2���S�I���Rʘ�_˨�S���~.%&&"�D`�Ǆ?$�����$"k��O0�O1�g8�3R��#����ߣ�o��7��?f��)���C�?�?&����|��O��A�w �=�H�Լ)��	P�=�L��Gh�
��o��S4��i ���)�ɕ��5�l&��i��Y�i�4�u���V�5���Ws&�9��iv�h����(Ve˖eIhr�˲�3�=Me���}M��&k����0���/l��-!��l��N��G�|����R���$�$K�L)�I�z���4)�Q���8�;�p.�(_�O"k&MD˗�;דPDpL�����xwc:�M<�&aj@�ߞg�?'d�TDR��EWg�)_]����@�g��:Zf/5,�4-�2.���j���3	M��F�$Lh$�#h�O4M|�����0�f��������&h$����S"��15�i���������#���jv�h;�~��Ssb���Ssbߞ����ًG6_<�����{��9S�L}:75	Yè����J����&aj0�7L|M��0� �[�shy�75���a5���][rre��%�'��]Wq~}ݩ55GWV�.ڿ�����=��õ��so9?<�(4T��hcdiK�ʎ�՝%K[��s��b}��� ��"�[��������^\��ꪎu�d�Ԃ:�U�.�
��{������,M���6�s��r/ޒ��)3T�K��6�g}C�cc�mM�a�"��:���<u�J�h�]=>�������doW�����Y�Iښ�rݓ�v�����������;��?�8�:�>�\�ɾԝ}�3�jG셶�WZr�4<h,x��䭪��{Q�ݠ��s��z���v2��m����m������zhq���߳{^3�o9<�X��t�+:�+���M��s�j~!��N��c�ʆ��Y|Q��?Su"Mz�#�%y.���^�㗹�]������3�����ִ~����7|]�<���d]�p��x�x�|��9xB /�Bfs:���$4�e!��\&��t��.��b�^�I�ӦF�_T�5�4�+:�e�i�������i�S�	�9�@�Pcj�t�����?LNH�S2���<�����E���������(����3Wqӗ�Җ�G��KѴed�*g�Z�����:�2=X���iG����j-ȀM8`G5}OjB�i�&.k���ϯ��)���AM{P��W�e�1[CunOW�ҕ}�v�Z�o���uC6u���qp{��='��<�v�X�ɣ�'�-:s���i@��S��S'�'O0m������7��_�Z�L��C�vU��Z�mC��my���������l�����s�Ѱ�唙L
��^�P.V�DF��kP�M�V��1��a,p���	?J�*����0��!�aX�%>H�( ^H�A�T��vTjE�L�겵�<�+���5�s�����譸H &D���~R�Ej��D��@��$�%NˠR�E�)Dr�4]0�����j'�a%���s�B&OM���bj��5c�W�mSx�2���b
ѓA8,Z�0�����bM(��	���9�ɠ0]���օ.�o��L�Q&?��|��HoZ�M� �p<�,cFh-B�c<��H��@� �0.�	$(,΂Eİ����	x�E�8`MQ������Ɔ������p0䰡�L��5�A�
��S��t�#8�K�(��$B�v:�0�&� ���j�KC8)��$
%�G�E��!ҞQ	:��1Td�)� �� �$[d{P }�i�f�IO�����2���Yv2�f�	h�^f���c�'L&���x�a�\ǘ������U����
��15/a%g$ϟ��W��[�`ajRrzj+�E���1�`!�'������2����!Dq�ۛ������+�/(
Gb^��粫b�B>�˄�t8+=	��Hd�.HY8gἯ��=�����t�X��7 h�=��4VJJFRR���Is�К�_Nz�_3����K8����mAK]x}�j��Q�Y���H�,�af?1�f��4VoY�ȱ��=��;X�k+v����kV:�2:�����3(�����Y��K5.j>��0�S���.����s���
~
����Z��:�y���`>cj L #`�#+�s*�%�}<�EM��"ۢα겭ƈ���M
�Vj�),:��h�!�1l4E��,�9�`��[�t���Hm-T[���"��Xf)R��Ԗ�o�+���n\9�����ڦ�%�eU�U�E%ݱ��`��ԇ�u�Pu8X���[Ĭ��$�Dj��-2�]!r)E.��d��f)�$8ba�R�8݆HN(\s�G��űֆ���X_gᒑ�m�z��߾e�у��N��<�q� ��\�����G/�[v�2`�����|q�+/l����wn��¶ןc��ڍM/_\s����׎�n]�r�֍�v�۹yh|�~QuQ~Vk}esuI}QVe�]�՗�e�ʂ�X��&��獩KGB��h(@��!:䆇���tg�yCL��A�pȿ�}ţ��W�������?���n~���w��|m�i�]��^��"�
����Z���'�J&�J'�����m�����C��=��15�=�N�[.�7���E��?�~��&h�k�g�4:Q�5Q�8��[�N���N�-�?T�)������������B��R�~!!~Ja?&���@c2�f2����(�c�)��DD���PD~H��!D_'ŏ��o(-��UL����f�w����Y ��Z�#TL�!�B��������7P�6J0�t��4qS�H`L�}��15L@M��0Yi����ժ����W��)o�W̲+v�e��B@{*�=�������l�U3�fy��15Kse�ٳ'�*k9k"T_�&!kS�`��i�[Hkm��!�"��܆���Z`DS�P���$��0�A�ZՔC+7*�Z	!Ǆ$�r2aV�����_��D nK$L��@nz�6�������&�r���ܐ�[1sOfbm@I�gn�)��JB��� ]
��9s
=��
�H�wi�kY�}i�iy�qy<�*:�0����i����Y�<��0q4L�	��������I�4S���ih�S3M�$ظ؛�5S�jf���i15GK7�U�X�r`�б�O��rrϖc����15'�>���ȿ�}���c[��[udC���������gcjM�05�riG���e�mjA� 1j��9�"v��Cˣ�ƃ�G|��':g��45g��Z�wlIֱ%9'��[[qyS��-M/��9��n�PѦ���&�������z߲�����X�w��=T��rT� +[r�5���#5����Xmt��eM�K��ƛ�G���� �e�4��#u!@m��&�U��(�6f++�x��Sd�Ն��B�@�a��8V�[Z��-��M���U�4k�����3g9%�iv���v��@otV���]~F�|���i��@�oj�Y>�9�8r�/�\O����������ٯ��m-z���ͺ�{ű;1�����}����s9oz�oy=o{|�]�G�C������7x��}�L���m�KZ�E��s쑯����E[��@�u�뾆G�/�o.)��2'R��,���9��%6r|!�e����7�ߪZ>*��nn����Hq�+8��^�o ���鎆�;�in� z��k�'��^�D.���"��:O�$�K2:���Ss9P3��\4���D��9�@��ѣb�^�)�����9L '��i9qNEN��#$����M��cm�s��3��3W�&M�/i9��\�^������*=�\�Ws�u�O����u���O�����7,�䀁�|0((�U��t��mAu�O^�/��m�/��Y�q��='v-ٹ�g��e�v��Xۺ{S���m���=�v�`�MG՝8^{�Dݩ���ӧ �ΜT? ��/�_|�j��K`�d���};*wl*ݲ�j����u{��?��l�v6��4�Y�ܘ>R:R�Ye6�z�Z��KL*�W�	4~��+!|"̍�6�΅<�"\0�I	p @�+����G��"?,��r�@n��vH�u�֎���� �m��/5���\�����t��ᕚ��ڄ* \��5�LKu�T/��IY#N��eHRS�))��Ăyؼg�s�l�3$7�D�u�Jw|�2������MM�P�QgY��#3H	�Ԁ�����d������aj��`��8�9�x���E�&�B�3'����%�P��6�D9��|!�����&cj J���4;�ո�������� /?��yp.�L��Sy)I����d8#�$�\	"H������1�� 5*�aI�\
f��t��F�R��d�<2u��5G�wK�s����4��5@��5�M3��0�fj@cj5C%j h�M�s����5�?IO���ij@�p�r��I�����R�h�n�"��6���@��ܧ�w��xU�KF�I�����9s.LNNNMK�`��L"� ����0������\�SR�p�t:��hV(�����+B6���v�R0�� .����(�T��2��'�{f�3_$=�eNJ/%JOC23P6�A�/ו�MNb/\�1on��$�+I_�R�3�W���,����_u��9fa�m��iSO'ܕOuIz��]%��Ų�ReW�*aj�Y�68�7y���mE���.aj�*�TS�\��|�O+�4���ɟmj�����0�'(��	
��g-�Q�@��O�s����*1�u�?ejr���&ˤ�.�VO���JAj�R�Q�1j}�'uA�>�Ӈ���FVk#*MX�
K�!�2�*cFk��]5��-�74���v4/��0��8�=/�!��K�������)	xK���H�$�����V�E/Q�~[eb&��K�;�B��Ȅ&)*'�8�!��ހ=�<?��,Z_���T6>X�ne��U[7Vn�X�mS����k>zh����./{���W�Ξ�xn��EP�_:?r�
�A{���o\Xr���Ӄ���=4|����'V_?E�ל9����延�޾y��5�KF�{:j*Kj��
"�1w��X��T{䋼�+=׉�5���玩KGCr&�����F�]��f{�qsL��-]i�w��V�\�k�ݣ&~��ď����'�{v�7w��Z�u�c�@a7	�r����_�,�&�K&j�&��?. �@Y���W��W����f��c��C�Щ����ݐ탐�!��"�_����NTfOT�L�?�r�5��{��w��.ӟl�?��4�����N!����9��0����b�g$�#����&Y�05�F����9�#J�}�]��:)z���#�|�����O�#�^9���Z4�ך����w�؃�B��!��0ɘ�w�[|�M�P x(�?��<��<Dp�!�=�	B�.*J�Z�<15���O}�jj^�N��S�8�W�4��T����E��Os&�;���������n�S��S2���59��9
fM�$d��9PSd�԰�YMM\� �!tq�舀�J�ƅY�=d#ShY�$���J`W���Ϣ�(�:)I�>egB�itF9vYC�Fpx�� �;S�}�!陴))�=l���4p��7P�����{2�f����FoG�  ��IDAT�F�F�ܥE)Q2J$!P��:�T�����4��r�|��;^�[��_�ȵ�ڼ�frM�i�fՓ�M���a4cj��ώ�a4M��l^�&hL�3S���ij 3��f�W�5�f�p	Ssp�Љ'����-�7��ԁ}�2�Լy�څÛN�Xrj����]�3|�����W\=<x�Pߕ��W�u^޻������M��;�Pn�'�f*S�C�v���V6��9O8���t<ms��4�(&��Q6�������%! �h�����4����O��>�"��ʜ�+�Ϭ*8����꒳kJ/o�;����]9��"��kZ}�����U���>���ű��9:sW�F�u�m�����V6ǖ6D�5�6dԄ��5���5�E�+6���+^�^����7��[�c��Os�$ߔV`No�"F��K�-�U�e����u-�M��[��[��[;�[۶�ӎ�Q3�;݌��*h���'��'r�/v�? `s_wxZLMb��K8���oqpg����o���m�=���c��-�SM��͑�[s_m+��\x�&�vi�nQ�~n�n$p��y�G��x�sө�ݞG.�C������}���ux_wz^��_��^�9���_��n�
�pW��߉4��x5�~3�����EG�M�y�r:C|>}.�)�^�2��R98���=�����}Mg}I����/��%�2�w�Ϲ�c߀�02�kh6hMs��긦ar�\��	�� F.H��etz�J��4j�N|�(�aU>gS=�P�YW-�f�9uJK�PcǞ��!'��e�?,��P�	vL"<D
����p�.(c� }� s3����>IR�L��NG�VP��*w���Z'X��V�K�!=o� `�i�MРr`CN|�Cz��H����3��'"�O�Z�КF9��5}am�O���4���aM{�c��z��uٲ�5���ݹz���#����\ӱ}m���{�����~pw��=��v/ڷ���Ѻ�,:u�����3�A]{�X��C����}8�d�����
�-/ڸ�d���]kv��_1�i1Ֆj
b�ܨ>��l�An4�tz�FkШ-�S��hU>��/��"+��2�������!��g��)/wrh<�ď+�"]Dj�@��a��3�SlS�������5��B�[i�������.WF��]1��f&�R�l�N�Ȥ<J	�4�����*xB%g���l�"9�X0O8�+�/����X�̠��ay&4߂ZEv^���t
�\P����^��<	S�@�Dc�üƨ�)[F��l��,.6v��ڊ������ܯ�w*�f�[+aL�P���ī̊���O� ������H��(P@���@c�p������0Gg��Y�'Lkz�3��B 	J��H	�SR����8W�q�GFreO�AJQB5�@[�B2� ��G	8$����R�o�����°�����8��(��*���`nҼ�9_�%χҒ���gqK�@2��
��yp)	y2�� ��B@����$Y�<Y�o��H*Y�n��[��B�!i�-�5���Ț��aL�i�a5�i"&�P�:b�l��i�*t��y"b��;�D�LgI�a��0�� ���ʘ`i�iu�c]�{Y���PWP�Z%v_*H�3�qS�'�K]8/i����$��e�2 �.`����-����I���B!l2b�H~~na<�����i�v����<���"V�\v�<X)���t��yܴ��$ ؃d���:$��&x�e	x���&/̘7�^L�������_���~�_x��Eƛ�Up
mh��ysk��s��qo���L�[��)W�j�5��Z�h�yi�}E�ge[`E[���^Ֆt�}���i%z�DL�/ࢣ-F���QzaN�[�OL�̑ 3`|h�C�4�.+pq�+�� Aa��ɍe���\��]㉑�Y���L{�O358" �9Pp	CJ
�^F��b�Q6�# #�6I�|�6�W�dR#N�!g	��|�|��Ca<		�ňZ���A!2�(�7�I���]�L┊�.�E�s�R�5*e������{�;�d7F��NK�Y2��Vuخ{��!ga�U�E��Q_��5*-2T�s`��$b�RbW���j�WM8�("j(��D8O�����hi^��ʬ�������c�W�nZ[�i]������U�SypOա�5G��?�t�X빓�N:.�m���쉮+���:����熯��zj��Ɂ���.�;wh�́�����\rh��}ۖm�8�n������ё���ʲ�`q�Q�T�t.i���u�vl�m����1!�&��315�a�mu�mnb�t{�1$���h���A=m:�4���� 1�'���V�$[�u;���T+���m��o����_߾��oޞ�շ&~����xk��w7��(/*����B��R�s��������겉�¿��#��e�����kN�;.��!��c�坠����!�wB����_DL��q��8����ߊ�v�5��q�{"��8h����W��oV=����jٯ%�/%�_�P�JBG��\�����"~$�~��Ɨ��#� C��B�����E|�"�&"�QoK��(��ܿt���o����~T;����/�����-���2�(�H�?`�X�TS�/`L��y8�C���ǁ�wy�}��|��܃ф��+���[�z<�0cj�Ĳ��])�qn�>�u��df��8ot�;z�-��5��U���V��^qŦ��Q_hχ�'#�Ca���bSH�)[�>W�&W�*O�"OX�+[�+ˑMs4S�k�d���TL<�%�eY�93�f*}YTW��]��-m�H�<x�	ky�vm�r�R�KC�m�<�� ��&�Hq��(#|M0K4��R��z�H.�I~'���wE�Τ��3���d��s����"S�ݖ���an��n��M"�(�rR���b�|3��Ws*}��R�zߒ�X�qy�y]�sɓ<5�HdN���0�f&Sg<1�m��m�2"�g�b��/`˓���%��cj��OL4ͮAz����i��o�`�H�Α<��%���n_R�e�h�`�Ƒ��+[n>�uőmkO��v��!F�̄�439��^�{&�Mͣׯ�?�����Sۆ^8���ޑ��XSôtXͶʋ��/l�E�0"f��ad��LMbTB�0LS3�x���ѦfU�'�fM��u�gV�]Z�8oW_lgo��/��+��;��'��7��/��?��/osWֺ�������9�۳���*�5P���pM{��%�"�#k;����ؿ�v�Қ#%��� ۆ��l��Y�^���ԏT�V6��G*���;����[��z��z�[�mۺl[;��;'�i�fj���u��qS6w�����00�&am�wG�v������O��.�E�u佼������ͅ���<*˿�}#�����^s�n�m��lw��7���;�k@��{��y���p��p�l��j��a+��|iz3��q~��ۡ�ہ�ۮ�W����U��{��<ᗸ�yt���H(^So���)-/I�ωW��+r��ׅ��0�s���tE���4�����9K
�1rN*<'G�h��OL͍�l��l�v�i��
="��H�#<��9.��m��������A���U���IS�D�N�)w���J#X��4@���h� ���g��	ؐ��{z��3�)�i�=�IS��5����H{�����#�l�:b��b�P]l��b��}������ڶj���#;V�X߻kc��-���w��sp/�{�����������G5;�x�(��ı�}{���*ݵԠ]�/�+w�(ް�h�Ң��y�F֌��w7�Z댕E���>7����.��bT�M*�V��h�*�BiU*�J�K!s�en�Ԃ�:�t�X�ȴ|�Y ��$f��j��&�8H����5��66��P�-���w����vu,i��(�T�z���!k�Gti�s$��	Y��]\��/��_Au"�^d�:�T@��Gggr��4,)�HN"���=C�V�<O�K��������X�UX�SS��:x~��qat4�����u^a�Y��A�),bLMs�|VSS�V�4�OL�^�KP��O�&��05�p�c��C$4�L�Mp�9����I13��CL�<����&���	C|!�CB|	�ė�D��N!��B�U�a�H #�����x
�'�9R�/
���h">�� 7�d��M�6hr|���XEU��eE^�NK�j�.d/��'3S�OI`����`��� �"TG�M��kp^N5���2�p�^���Zх>Yz��Sh�Ϣ 
>!L��� �"ڞ��$4cj�f��S�P3�H����H�x�4f15���ؙYM��ze�mm�kY���PS��YI���,�2�����c�-�d�p3��LD�&��NM�G`�����JK�d���t*���(�ˮ,-*/.�ˊDް���Ѵl����-��5��t�5b\I
1n����� �@9� ��Lp�)^���)�d0G�pB@
��~4#I�<��������"H�
��%2�+:taD'(uP�"["t:��<QO!�O��*��4��Z#`��8\GO}bL����pg��&�/�ks=z�U������r��W�|����9�ґ>�(d�"fq�$�2����B�&ߪ��T.�Ĉr>Nf
I|�|.���$�S�Vʄj9���Z
V�קB���q��h(̒���F�ȝ^�jlWo�ʼ`M�U�4D����0������Z���g�z
��TSg�0j�DvS�n�Q�9fU�4b��y$	��2���/�זGZE�[���r���^��am�֍E���ڗ������GΜ`r��^<�s�����o\�q��ʙ��gz/��p����γ��N�9���Ȯ�C;��ݳud놁5+{�����67T��#����"���Ȫ]Ԭ����|����S����eM@4 �|ĸ��nlU@�9�]���_߸��[W�8���&~����<������;;W����l�qŤ��"�e�o�T?����!�(/�(˟(��.;���C��k.�;�c������S����A�����X�#�����DE���_
|��|���{��q��7��N0l���b"k�CN�Z���BhY#�hY#&����MD09k>B�����C?��ob�7Eȷ(���w��7��{���zB��4?)���0�z�m�^Ӓ��-����k*����(�&߆����wy4o�!�c��!�����?bj�ccjk?%bjS����^��!�i��Wu�Wtt@���C}Χ>Ԟ���t����ưtc��������옚Y�Nj����ĽQw�`�kf��D��ѝ%���o�z?Q�f�A5�)g9���Y�9nS�ϖ�z�j�� =��e$�RS#����<ʇ!�#B��7I���i�������}���,�;7]��AwH.��0����K��f>��ӃA���ˬ�O�%����������t���<-��4A� !h��a�B��NF��)�i���o�p�H>S�k�`���E[G�6o�ڱ��𦑓;לܽ������;���a�&h��g��I0��<x����m=�����k���|ppR��M��=��.����i�����$�����*�m���$�0ؼ��������&�iS��5O35�>�T"Ćq13y���=�28�*pjU.���ӫ�N�*<���_sh4��H��Ѽ��G�m����7�hi�奇��/�?Z|p�t�@���l����C�U�W�]�h�H���M��r7t�m�/�5V�oYՑ5uG��^]�y��U�G�U^S�oi���ㅇ��ZZx`<��x�內ה��������so�um�u��q�����0"&�� v���bj ����h�d�3��Ә���o1�����Б�A�ԴN���/κڙ�|w���}�����������UE�
b���/�l/�-�;���/YL�Z̷m�{v�}��o�=���[qY'p���*|3\�^A�7*�Y3����7{�-��Za�Ѫ����Uv!�}M�\ � �P�*}�?O*_����+u¯����B�<=�	�#�u��e>6x�!�%�`4�B�	�'hMs���J��2�9`4�%��Ar�,�nS&�bS\��ϛ$g����>(�����eAsXDg�9"���.����
�o�Ҷ��z���M�JA�2(c)�>�e��pV�x+U�U:��15K���`�ѓ�LP���L@͐O�D�Є�	�/"�ʺc�ި�/���T���7���c��������6���x��aŒ�M�Vlݱ~ݎ�+ {6�8�}`׆��[zvo���ѻwg߾==�7���x�@��#��w�9���	�h?y���޺�{@�phӑ� Ю߽�z��ڍkvl�߶�lݒ�5cEˇB=���2cy��0f̍�#^�۪���6�\�R�Uj�B'��2�Lf���r�\��xB%,6Qz��n��M2�U�w�CneХ��>��c��S/r�t���8�((�iZ9�c��S;��:q��ζŅN{�Y�m5f��1�*��{��ߞ0k|r�(��_�q�
�6�N�iU�F�*�%�`dKNG&��)x�Bt�\b�<I�7ٌ�d����R�J�\@��W�T;YCБ5>4ajCdSX��0��&W�V�M���CmD���DL`� �Kp�B����Bbj�-��M�N�@����9�7��/��Vf���x��&ʴ����A
�2R�P���*�#j1����AAr�"0&�0Cq0&�q0Dq�	v*�����b�kPŜ��ͭ��ݕ9�����ֺ���kP���JB�扸�gS)^�B�Q	���&B�)��a�`����47`s�-�El7����u�\���І�B[Bhkc�LGX�6�)�i;���\9�7O`��̄15	�E�F˵#���D���������~�ߟ�w�3����4333�Z�L���Ͳ,&3�2C��$��0�$�������#w��Nv���{��<�ԩs�%[:��>�ַ�!�\bg�)�G:EM8�ȒGM�;����6,ʷ���3+F��1#�_(q?"�^ �W��4��g�	b�J`��8"j>~ ��"	Ä��:�4g�}�Y)9�!��r[��r������|��Ów�Ֆ9rR�
!���*k@�����Xv��%��H	|% �ET�����a��$� �<G\�c �#&�yf������+�R\��Z�b�{en�:/�2H�Mbק��2�u�" bj�r��y
x�S��t�Zڋ���L� jjTB��K��15��W���w ��,p��n�������|� gAY����N'̡ɸ��b�RJ�SEw)�^3��%�D!��%��Yt)	⢉�<�ET�1/`�+����@�c�,�ab��IXMƼHD=�Ǯ �P�8/��pDh�Li}-�kK�}�T�ү♄/�'���(����$:�C���0L
�J�'�Ⱔ�x+��Tl��CְI:.Y�#)�D��gCt:�΀�"�ܤ�\��DGI����P^j�����x����6��nJ��L�O�M����RwLe��ٿ+��^����
��/:z�d�P������+�O�k���;W�g�b�T�������&����m�6����,om)o���[���Xݺ�*�&�4s�M�\5O�uZ"kHyr�w���X��6jSD�<�5S����5�6*,k,P�j7�;L�g�C�(��4�\m,�i�ٮڅ^]��O>�������m[{6�sޤ>D�ߤ3�X�5�~o6/�C���T���ύ�w4�7�ʇ&�-���Iqע|զ|͡~ӡz�)�){�!��K��������g�����{�㯉���>��ƪ��A�l�or�ż��ʁ~��M���N�9��D�Ds�|L&|�?$�>"�'ޤ�ߠޤ#@���i���+$�*�_�j��.�_�9�����s�?����>�_c_����G�!�rMx�"<@æ�U4�e�
u;����x� !��5H�$��
�&��O�D�,55���+GsQk����r�o�U��!���=�z[���.�z?o bjz��������ۼ�/��4�>6`iX���I��*'��:/���.k�9�$H��F!d���j�K+M��|F%���ITt.����k^ĬY	���x15�Db��T����$� ��@AV?�N��F�j�F����qiA���3��#~���)..f���������q�+mb��[���RemYʮlug�Е�ֶ�Q��f���05�(�����̰�ܸy��	�����$�25��������ġ���-�[R64�m�(���r`rӡ��S���4�'�"�lLͭ�G�O�mnڱ���L�����EM�����j���A�:J��4H���ǆ3�n{��AtLT�,婦f)��Yt7�4Q�jj �{}�����{L`oopWW`g���7���������&�D��#qGw�=���{a����6�V�Ǜ���ҦZҧ�2f:�&[�G���C�uAИlK��H�jO��J��N��J�ٛ�w}������L+�����3�����Ͷvv��%��̴y&��c���z`��<�`�jtL6�L����lc���R;e��>��x�}���O��A�De��!��IS�0��6��4�eP�p���
�N�Ҝ�jG�;ݕ�w�{����ܗ��n�=/yL���&�	��BrF&9/W\V�nh�7պk*�U���pMc��3]�Y�<wl���d�~T��IYߧ��v~\��iA�Ge���k�q�@L�Q�$�t��<Oa�&�N�I�s��6�#��H'�3�,��9ID���N��O򄣁9���"���Av�F�/�48$D��S�,��2�	焊��� ��"52�^e�8��N2�4��J� ����Oұc�6b,�i ��1�A
65��.\L>���A��e�����Gk�ԴI��
B�G�,	�i6њ,�F+���@4M���s�jݜj���ԹxN^�C h�H[�򖀪>���+�u�����7n�Էe��ލ=��:�{&�5o��4��~�����u۷5�noo�������1S�gg��= � ��f�*���LVLO @ /���8P�y���me#[�;�z[S������MF�65�I�*�V�I+�*�j%�'rB6W��L)����|����A]��"��kpI@���~�$Q�L�kҌ��^��V'�L�Oqe������Go:r�̅7v��ڵ��U���L�%�f/p����Ng�ј�R�b�H�`�u$����x�x#`a_�&p�Xy��b���V���܏��g�z65�+CJrX��H��d*U�J����3�5����qҋ�,@��55��)��$bj���Ԉ���'$�P15�Ç%s-d而!��8K�H���4�<�i�o/Z�~������(f�	GELH@s)�����Ԣ���riq|*JLË�!��AX$t���E��n �^�q�!���gw�U4W��5���&��0ً!ǽ��ǁ��GBI)X�dbBf6� �ab�L���3s�f`�b V��ź��|"l���m$�Y�;T�)s���Y�d�t4�Z'�� ��6�ԅ����YFc$m�i���H�`xY"b�6`Yp�c�Yr�ȴF�� �t"�9Ɣ=yj�٘$*ur2�d'7V=/�?'"���$��I�pH
U-�k%�$c`�T4��ǲ��lRh�q1|*Vɧl�D�!=`/�
�|un�wbK��o���[�?y��7n_�w���c�[j,r���? .1Ԡ-�`��K���D�x15ABC��(g�[� �\"�A� ��Vs� <�
~%���c5�E�0!MG*��J]40%��3j¬�nc��1KҐӘ+4�)Z����"mW����ܚg*MT�[a��g��|0�rh�զ� =�,�2���������SC��*N'̥�yT��j�QJ�[��A;Y/L3JC*�[�50h<��@���^@���1�"���D���Q�	j �a���X:i%D\A5y5�C'�s�<QA�c۴���m���~S�^d�3��D@r�<F<�C�_C%�!aW�Q/�P/�cW$�W�Ak�h		|^��(Yd5�r`d,��G�s�,6��e�B�Q��:��9/G���*,Ь]kkiu����i������v�ض��0h����3��o'R�ܓho�݀���+��^�g���s�f�ds;&K�&Jg�J&�KG��n�T�����������������,;7)�%z��.U�]�a��Z8��ђY���|xVLM��Rc�6�iMNF��	��P�[\����m6Z���n!���>�����n�+Ĺd��T���ڃk�߳��݅/���;����i[w!3��q"^"S_��ߤ�~����`Z��ޅ�����O��7��w,�G��Y�gUܷ+9�o9�o;��;基?h~�j�K�{!���L�?R�H�.-�?��X�7*����E%����g	��<�/�������M��M�	�!!��#�
�m*��[ *�M
���B�K�����kF�Bk����C/-L�eu������7��7x�T�C��:��O���<@�`Y�¾��܋O���,S�DL�]���VC��$�n<�%�Ϙ��\�p�p9����<��'���Tp^�?'�9���3	w�;]�Y�h�+�
6{��=�� �/��	~��<;��Y4y`M��� Y��� �k���A����7��K������>f�JҒ\2�E�7� ��i�r�2~Ȭ�T�T�c� 1v~�
B�*|�j*�&��T2�F���
�ohx�SLL̚5k��4�ƪU�@g�� ��D�ҧ%(�A����/!����^|���_����5&�aV��)��ES��ڕ���U���sA�2O�L�,�2O�5J���y�Z~����$�25�NO�?�m
lk����58�nM�Ҝ8Ԗ��1}s[���c�C�;�L��Y�4��(K5 �(|`j��-�S��ǧ��O��m:>� ������UG�*��=���'�y�C���[�@7���������@��,S��D���t�ej�eyz����5]�����L�'�k�:����v?`�#0��ٗ�g k���Sc�o)�������x@cK�w�1<՞2ٖ<֜8�D��5&ZC����}��}f�w�����'Z�;;�sm����T�o��=��n�δx�[=�ͮ��h�u��2�`�hrL����\�M��F'"k���O�15�FL�e�45�p�x���$��L�e�f�ܺ�±g��@��Pe�BK֫nm�xc�ݵ�5U<�Ƚ��t+3p-�}�g9mU���O*�gd�s2�u��Z{M��*���J�5���z����x=��Â��*zR���̀����v�����r�>�%]Ui��i��	�Ѩ�D�"�s��=Oa�!��A܋4�)<�$�
���I���81�>v�����(�2O�>�G&���G"5�h�c�Q����9�#P	��E��8��q9��rQ�U��(X��LX�H����4?�ƌ1Q���*fǷM�f�����C�[�1��7�V�5>f=>a ���æ��M���:��}L	���Hq�2\lj0-J|��ؠ$�DjM�d�7�l8aG��f���Z��ǫ�
꽂L�[h��ۂʶ��1���Sy�޵)�k��j{��z;Z�j��j{Z7��N�L�tM���'zf&{gf�w̶��ѺoW��=����ݸk�ff�rr��&F�F�J�ou��6��C%�חn^�v���I�u��Jom��(ې�j�K3g���~�߮q���D)��@�勘�%fp�<�N�q�Z�U)sj�!�:�#����,�
P�iM��U�Ji����l�)��hq%�Tn�0vb�����]����[�<�ta��wʛg]�mF_��_cպ�2��s�R��,��,��s��6�J (I9� ���0[���Yd1�ȃ∸�(��p/��?���ϑ^x��z���S㓐U�ES��鱩�,��)�EMM�����b��υ	����U���$Yi�65VQP�u�:]H�7)�&��� 15`��t*�G��#�)p2� �G�i?@Ú��B�\td�|�o�[�'��#�cX���ٻJ@W�2$e�$,���2P|Z|�X=J	� ��"�6>���ebc@��l�נ���r��NC~�k�؆��Lo=<7<�����,Ѯ�14�\R,��_-�$(x3�`g�\���xD'�`�`ll�[�x�X�W��Ip~)�/!�Ā�����1�E�=�P�*sB�.r���2, "h�:$����:��D�R#�D�,u4#e����<�h�d4\�5QMә�@ �#K�nN�T��zX�vpW[81>�&%۔��b�3m*�S�wi�N%I��b���W��j.��S@�F1í���D�*ũ+J��BeU^�c����?~���=z���g^;}`��Ѧ�I�8�'��T���P$�89#V��S��������0 ��d�h�~;az������|@��ԓ���Zu�Yb�%s3M��f8�F֘+o�S ZTm��Bbj:�Mٺ��8��	�^�Ȥ��yT>���cj�K�����#��ݖ���͸x�DAnϥwh���˲o�Y��c���K#
Y)����2�EIw�^˯e&��p\�,I�w��U�%��0�Uh�	��c��^$R�P�	,�`�9,��� 0���85�BYM$�"�VB�UTb<���WQl*__��ڒ�=M/�ș*!Y""	�D�d��,�G&��+���������_C\C����2:�`�_Z��j�$���!��0yR�P#�Z�*�G��eg�sr4�E�wG��w���g��J�O��
�n5h�͍g��Ύ���ۿ#����=3�������ٳ�r���;g��Kg'JfƋ�G�Ɔ
�o*�2�?Г�ٞ�ژ�T�[WUPY����!�!ŭFLM�������(�Zr�*TAE
R����X��驦��Jk�Ӛ#�汬��&_c����Jn��{��A7w�G0T��p�F�&��]���*�`����������5�I�I��%�_�(������7z�Ϸ��Y�
/����h���߷�Y4���[F�-���Ev�&`�?rH�r����>�H?�+�d�]���9���B,k��A�?܆ص͂I�w��/J�_��?��aC����$��M���%��s6��HΚO��O �k���h�wh�;»���M"�u��#�$Pn���֟�[�^ؾ�7խ������xW�}[�x��> �^'3���P�Gh�kX�C�I@}���5^���D�܄�7)��G��ih��tX�<���ds�>P\x�n�e���-S#��	�Ʌ�Ղ}��S8�NFv���7yy�>��SMͳcj�|�'i�sM��"�Cd�3�W;���M��P�|�*?�*ĨL���Vj@CrȈV	�"�[�l���T�]j�]!���|KA�)� ���I���T��g�l<6�<}���ʚիW�G%x`�Fbm@AdMdDxL���O�< �g/h�~py���ǽ�"�;!�Y�擂^�OV����3vf���jGlgz�՝���l�c�E���D��~O15��'\̿óbj��S����f�`�55��B[[C��C[;2�7�nj͛��rtn��]������w�gcjn\8thf㮡��u��;���N�5" ����Y���H.��f��ٷ%u�ִ��� >�%������Z�ej�45�Y@T�,��55��A.��vt�g۽3m���t�{�م����h3�Z�;w����:�1�`�`��)C�Wb��R�Xs�Xc`��?V���Dp�ջ�<cΩ�t�o�ճ�3��7��;4���ە4��qn����;��<�����@�4ӭn�� ��5��'��[�2O55H��Hd�"e�HD� ��3���9�Hբ��Q�5v��
��
��ƴW֯�h���mm�lh������ks�˹_�~';t5��4�7i�i�/)U�u�kꈦ���H�W��kr�U���ۓ�zZ��͟��ո��M� �l��q�g�-�d���]Rk�2h{���X�I��q��9Oa�#�/@�KT�y�s�@?����pp5O�;�]�Lx�C8�a�bj�xD�eC��pb$�氈vDL?"e �e��r6��I	k�y���yH��'���i��>q��CLSC���p^ad��$��F�	[I��	k6�V6�W�'��15=��I��w�Q<\� �'��I	�2|��.��T�f�QElА�P���b�7[aM��`5:YM.v�����4z�>n��_�����>a���#�9�^I�_�Ԅ�Mi��B�@U�@S冎�M�]��m�u�u�M�}���[�G�����M��OL ��'��'��?�g��^P��չg�u�d��X��p��P��P7L�4ώZ��:v�4���l�Z�םXW�*��+6䥛rS-Y)���9�%z���b���b�@�J9|!�ͥ�t��'�Ɍ�M�7�$n��ğ��M��f��K��Uϥ���n�_�z���Pi'�@I��u=�K��GOO�7y�����8��O�]��؍�m�}���`j�hr������F�+G�g�5�H���)ӰT��)���d�2I�
+�~���c8%�.g��P�*��2��b5������$�X%��#����$k	�Z|��x��iW?�[�EMc'9h%.F��(�SS�T�(�R��(y�K�a%FL��OP	,
�C��D��S4�2�::�#0� O����扂|P�N�e��	�q�O�+xT����r@�35"�J@Q��rA��I9����2&15� 6>� ���mmNJe^Z�C_��|�����_�|b�K�vٱ}n��"'� a��i?�e,��Ct�>��'$�_���q^:$&���D	!,�'�	)JB��������$	��,�	��3㊝$�RSS�bFd�b2���A��DMJ�h���p��Y
bj����0�#����$��.] �m��!:&jj���?�� Y�ʉ��1,�t�L�t5>ECJ32ӭ�t�<h&��IVi�]���6Q��6��:�W�t"�V��BI�]ԋ�@a�V��I������_���W,������go�}����WN��m,���)
ADA	�xP�8%���������iy�z� DE�k�Va)v�B)9 ''�)�FZ��]��Ԇ��avC*�%S���ۙ�US��9_	k�bmgQ�B}g��6M��%9`,��	�r��K�2��jSjp��� w�������� �ғ9
h/���]S� �$5rK%d��,���ֱ�:NP�N�q����+b�	ώASW�H�����{KZ	���� �X͡���kȴ
���D]I�^����PI	l2����k��5��YU��L�̮�Ő���q1Lz,�
�L�O�b	����8܋����V��V���Ј�Qq�j.E�&��&������D%��tj�]
��L����[e���=�3�����u�$�m�oKu�����ь����ٻ�S�F�a�޹��;�!h�=�����փ���ٳgݎe�S%�%Sc�c��7�m����loIonLoj�i�Ϋ,��K
';�AS�G�l��Y��6.bj
t�" �@~�5�X	�d@���155j����7���n "k@�is�Z��6��No��:�@���ogڸ#U��گ��$�o�T_5�w���X�{鏗��|gs�����]�KTګL�=�c�65~?lj��B���4}�2=�h��7��F����Y�U��!{�%�%��#��+�<��E�񏙎�e{��;�R����i�eX��,��׈�������{�7l�_9�o�d8s���<�/���Yԟ�H�QH���"~D�|H!�> ���a ��p��o�7�gVşF�_Q��Pްй���~�����=�15�!&��	K����&��%��#=�b����Qw��Ss�ޥ�Ss�D�Keݎ�(7��=S�5�yܗ��uO2���B��Љ��Ĉ��
����>�Fo���~���e�&J��4-A^k��&?Y�,j]�:��K��P�<P��R��nH���nf���W��2�M�0�XF�$�%\Pkyt	��%���aP�(`ЄL���qY|&�A!��Ћ���A�R��<0AtFO��d�䢵�D6�I�<uA���W=����=���ؕ:ީ�;$%~yUXޕ��]��PU�櫻�`Y����h�i��05��Y�����C��D���=W?�ƚ�#���/,k"{?575��g�oL�ؒ?������c;ƾ;�f����Yjg��Sstǖ=���k��k:��e�.�p@��75H�RS����۞�Q�41MԼ<�� z%*k�)䲨�YƳL͎��l?�\���7��Lwyv�� ;z��]��5ӭ��6�x�w�m����Dgh�3i�+y�;u�7��*���,EK��-O7֜���F<R��u������.�D���N�uy���s-��F�D�{��5Y�j�N6��띀�p1l��Z܀	����G��i ��,s4Q�Sݨ;�eS3��6^��*�d�Ԁ��o���P͖Yv�¦f��<Sj�*�L�ئ���ko��?������7��dc�ǽ�o6���\�V}ѣu9���I��;�۬�M��:����T}I��(T\)�Hԗ���Z�eG蕔���?��Y��ם� �����������x�ժ�Lh{�D8��BԳ�,�q� j�"�%�4�r�?�B��P'���x8��9��>�2q�p��=�O8����晤cl��|�G9§�l�}T�8*c���lD� 랐O�d��R�.>i'�8�#�r��3�BO0PSd�����A���񈩙��G�	ä8$�f=n%`�j�&jjzq=��n(�����@���BB��+#�ȣ�ݦ&6k X� 5j���bc���&��͉j�F0I��z���5�D-^	��%j �O^�U��U���lkgibOuiGmu[]uC�ڵ%�ey�E��s*��j*��Z��[[K�����skkK{:�z)�i/�n��j��l�nk�����۷�O�u�Mv̌�N��N��ݸ>��%X]a+ʁ%��R5)M�_p��NG�ϗ�8��H��I9|1�˥ЙD*bI�R�ܬQ�x�\��Z�Sݽ�v�X��SuCW�߻���]o��<��S��Jņ3e�'�6�Ꝼ�~��M�n͜y���v_|s���[��>yw݆�U��6]���?{w��Wj�w_h:S�0m7I��S��Vfv��|��Z��P�N���E)�R�MEC�x<9�����rQ	rb���v�i�����$�Ia5.�A�ha"�q�zb4�p�����b��IGLM��S���aIU��:M�6E���hL��GP	dL*6懊�Y6�Z:�58��,RD�e?XF��/�D�%͒I <��|�O�>���K#JِF�4�yf%?ע�Y�0�3�izU'� �r
8�	:>Cå���� h �����U����r�*sS�܆���o�����^�t���o�>x�����ʠY��`ί�S4<�^H���19,�����,#�%�D16I�O��R��T!]E��3��,-%CKMSQ���,�g�7�-�<��I �:YC���� �q4K��<SӔ"|*QS�,Yzlj���Ҏ,���H�S�ʁg�� PƔ�ѓ���� g��1��;[ّ&mI�WyYe.v�WP�����Ƃ�6?��	h���|�,�+�u��|�t�2�&u�[��R�<�4��$ٖ0�L�iNp��(�������~���o�v�콗����ͳ�9:UJ�
�	b*Z�&���IJ5�&�,F[$�g��
��$\*�GC�j)~=0��zN���m��;�%~ePX��Dސ��<]К#i�Ռ��Hh�W��ڋ4�%��b0&i/4T�*rݼ$#3��ztB��#�9t���A�)pxxgpg�����x�fj��B�V��Vۥg{�쀑2p�G$�&9bjtT��f�AQV$ �����1�X>/p�\v���˚�$ e���  =L,/�f��^9��ڒ��`~�;ͮt��*��`��x2u�O�%Qc��<�MX�}~��ϑV�BL����T65��shB�Pa�h�VC�kMK���x��}յ���pGOb�@b�����[�7�F7'M�NoO���1��s��o6mfP����.pXrxwә��N�͟�82�r�`ݞ=�vΖ�L�L����nߒ�q ��+��5��1��!��65�Ii�pȜ�Q���T'���5����PC~,k(J8��MMKD�<�5SÂ�ktX��`SӢ#�9X�F�_��*��Rw�����n5��IO�N=�6����g��?�{:�'5����d>���H�s���	���O�ޅ��_�B�I�}�<�h�dWu��:���Ax�,�o�햾畾���|P�:��oY.8�&�˚$�B���6.86]$�F�w9����?���~ǧ�+��6�[��|��ٴ��P$��	D�"~N�~
�?!?��?F�?A�?E�>B>����[	�K(�U��������)�Er�F��R�kɫT�+D�k$�},tMxCz�M �A�ሯ�1��ϊ��5^��2�v�s�L�E�ܡ�����������M�y�k|�>ﲀwQȃ	K�墋J��ZrA+=i��v����	�p�+��7��H��� �7��
r�LLM���$m^T�  a5��O���7��~Z��\�%V���dVs��*�W��fؘA=ݭb8d,��m�L�Q���`T��R%t�����0��(�S�t��I�pXB�àCDxցg���<5b["�6��f��A�7�3��@'�i��Y�/�\�&v5��3��)nuaHS��iJ� )�{r������mO�fي�(QM��D�k�ڙ� �15Q6�i�p1�ϊ����e<�Ԁ���6�uGM�pkpKKpcSpK{:S3��a����S۾;O��f��S3�kh�H�D��ۛ�6,55��5G&*���5��� �h$g�f��<�i�?ޓ{���=x�����ʚ������ bjf��3� bjvuwv`_��ir���&۽3]!�TGh�-0�N%����.Ԗz�����$^}�x��3Ti����8Fk퀱���h�u��>Vo�5�7�fZ� ���MԹ�}��z�0^�lt�ˠ�����v8g��5�N���5�M��f7`��U3��S�P��A�X��o@.��vFMMD�LTِ���2�t�iƊ-���|�J����w��>n�hK�O�:>���ng�{���m�x���)L����������ڗ�s"�Y�pA�8'S���=�B9��}Q��ˎm���M�(h��㽂uo���s�/(��)���է(��$�it
O:�� ���(��~M���?��?A@�"cOSp�p�y,�O����D�Aِ��t�KF�Q�b(�a9�}L'�̫�GU��Ss@B�7����l�;���0���IS��{Bj�P�ʁ�� ����55=dT7��@Gj}Rljd�NNR#Ŵj��ޙ;�9w���ja���@���d��8�nN��h��S��X�,��Π�#Q�R�x�eNQ�[\R�d�
ݙA��t��6��b0��Z�Nc5����
'��������չ\��k��u|�^h3�f�ˤ8��`E~~{]���ͽk;J�[3�]�����e����ϘV��
�C���F���L�3�-^�H.�pX��b2��G�)�H)54�*BY-U]{:'��n���s*��LΆ�9�n�m�U0t�d����{US/�N���>��蛭s7����y��w��v�����~�q�����N���.Zn�K��ך�nU�\,<�ݹ?�c_F�Ng�E�^�Yg�y�Z�j�9[���A�1I"4�r&����h("5�Dax�BYX�
�i!%9�"���D5�i�tS�ʹ��)r~�Ԕ��^Y@�6QR����o�>[��>��'cb�,15�Fc��q0���,Ο��A���ˁ�g��9x��C��/�DA�� �`p�_�0X<ލ;
�'�#랈x
+f@`"�[6ߡ�;�<�����}F�G�siYN-ݡ��Z�K��jyϥ���O�S�m����	�z�C��q�9?�g+K�=9A[SY�[w.���w^�y��@}�ܑ�M]^����p6	�.�7�����rr��T��T�,5��"e(�ir,B����gk�9ZR���/��di)Y:xw0�Qd'ڈ�V\��(u�"��A��|���ʚo�j¼�as�Sh�����t)h������Y��Q[� �t>��lxٙ)�Ȑ@vg+Aݟ�(Ё6���U��i�@�\�*iB��dyS��)�ؘi�ϴԦ��S뒴�!EYP^旔d���"�&�)/�*J��"�*�#ԍy��)����"՞�T�����X��O��/��;�ݿ���s�r����k�Z�U�R1	R
ZAC�$���Q��R�S�v�0Ϋ��T���<J�W��k�!=)l$'���Vz���f�gY�N^�W��ϯ	��ͩ$��y��=G�	gV����+�T�E��bmw���X�Q�k+0�K���!+��#�F�4�������j�&�\�?��M͢�!`SC&`�x4�ND��>� 吕�V̴�#�o�M܈���fi�Z�r�T2��ǠI+ѸИ�Q�aq/�h����y8�e&��h#�IYC�V@ �+��������54�.X�[v��
����D,,��f����ؕx�j")�D�'A��J���	��q�*+�STl��C���jU��X4�C(%*���uZ�AgV��(?��.��%��3������mږ5:ژ8�)ur[��X����]S���1Q~hw��x��X��]�G���f�`�sΝ�x�t��㝇���S�k�rv�bj�b|{���y�2���[�қ3��s�ks�
3S��݉aK�G����l7���7���7a5�* 	P�!kaSS�_45�VxK�&'���j��:<숬5Z�Nx%��g�i�Һl�A��2T�u3!s�t�2�vK����cAǾ������{䣭��÷��8�E�5��&����	�¾��{!5�������O�����W͚�jq�M���Q�ո䯻�oyo9�o�E��_���t/d��}��d�BȺ�3,x�N�߬ʿ��s�"a�Y�����'!+�`��:�;!�a�� A%~N�?#��PB"�'~��}���$�i�S��X��C4t�[���g>�?4�~����<�����h�������I��E��I�="��cp��HL�=�7��6
65w"��65� 8��65�#�3���4���ʚ�B�e��\tA)>����JN륧����K4��=m��5�����7��g����æ�Y�t/s4m^K�5�oK �	�y�F?�9�h��|�J7��GO��,i]��r�d#�bx�L��a��2<�LX��
6�G�@�8$��JB6yҩR6S�a�Yt*x<aq	q�q1� Ј���	(�3f��5�V��&i�F|l� \�A�ȫ@ �����C'&hD�d��$�R�aiɱ�X�S$�c�/O�_�Z��)���h�	�(K5 2U3ˈڙ������KwT�,�Y�&�-���6S�MMK ���ښ��)cSk��`�����Ʒ��vhf�Y�f�Ķg�ϙ������<��n������}#�G&�N�����ꞮA��-?2V8:Z86Z���cc���r��� � [qG@�̓�F� �	��FMbd@� �4O^�T��� h#�{#g;������ f;܀ɶex`Z}s]�{�j��%."�Q�S��yJ�k��B~��V��U���Z��K�P�9U�ȷ��K�@=��jqO�z@�ǁ�m �n"o�.c�t6 $1��&ڃl 5Zi[g�4&�,��V�T� ��k�����2�T�m��>Ya+5��7f(7����\���l��t����/F{����p�G����ռ�U�N{�ۍ%oT�R�z'+x+�s-��4�3j�h����9����p^��?L*x?����j;���FF񧅕_W�ʼ,�D�������� �y"t�@:�#��O��'P8�<�qn`t�SD"�?�
8�F#��$:���CD�Q2�{��>����s�G��#B�a1tPL:,%�S���G4�A5����_Iߧ��ʩ���=bh/@H�# ���p�;Y�9j�7�L�b'�S$�4��!�)�q3BB��c7b7�c�k���p� =ؕ��5�ĘRl9����a�{��.���i��:��N9�SE���65Ԣ%��m&*��Di6�[,�V;���y	���GB�v�$k���֠�#(�	��}�6��3��([�ꦠ�֯,s�s-�4�*�$B�B�ԩ�Z�^*��8b.W!�<6����BK `�\��`�iL�Z)V�ez�ڢ��4<�Dj�*]&}�Ù
�d�V�g�gՖ��^�B��R���q=�Ӧ��
�P%�Tb�Z�W�52�\H�p�,��$Ә����Ǡbc��R�_WՙUв�}��k_^�������i[o�FH�v+s�@����-WB��<m��{�4�{y��'C���r���[_n8�qݮ�27����L�r!}���K�s)�_�7�q����4�7��o����
��k7��z��u[�֙#Q�$r�H��3����Q�h�RS�SC�IA%!��'�0a�N8E���Ce��|D�@�|+9��;�NJ��^�a�x9����ֆ�k���2I^���IU�)k�C�nW��|5��-��4&.v�,E>�Q		�>6!�C=�� �+d�
��d��O`�&o�]dr��x-�'��H��g��G�|O�=a�	8 �Ǣq8���Ax��v�A�(�=�h��2�W���6Q�K��e��Nn���b�%Y)a�l&���&^���jb�� 0tK22C:Z��	�~n�&��;t�a@�[7�P�ɣ�����oݻt���[/{��ɩMIV��딐Bz���e��X��7#�g r�D@�����=�\=>�@�7L�B3��F,�n�4�B�J����6rX`��u���0�!��=��A�,hNᵤ��i �`�6r؞!td�m����#���te�9��!�Α���d+�����4iD�(��T�Y��lm��+�؞�kKW7��S�Y��t}UXY��{�k��ʠ�&,�ȷ֥��%iצ
��4���<�ܑɿ�񳅅_���?���G�.^;{���Ç���ӂ6	�.f�T�����B($�x	~al@�$��d%&E�MUÛ�g"i���m%.F��Q�c��i��J�է
��%���4aC*N$��o���H��]�J��b�`�z�L�W��-�����K-�撰,�-�.�*g�EL�̣�(��q����w_Dw<�D-	h#/�"���Z�u_�^�|��WG
h?�,�^^�De"D"���_ix�b�x�����qZ>dU0\Z���F���$�0� �(�fGF�� �Ƞ��$4Og��PA$$��x1#�'p)�,r,��cbD��OVx��MR��v!�L%�Y�ʬN���L�!Ū��.	�,f�T-� �a%4�8n�����V?��{�Q(qd8���0bpr
K��k�l��7	�����ʬ�8M��Ǘ��QS��Ґ�ۑ=Н�q xk��x���������1U�{�d���{ %{w�-��Z�ow�ι�su����W>3�s���|��{ӷ/_:�{l_�C�z��i���ضnh}Ao{v[cVkCn[cNs}nCeqcYaUvF~(ߎ2ţ�pJ�2����3
��b5�DO-�Q˴@����@]g�U��fZ�%�����7:�f����}�w�.nv���f��8؛���~�W>�U��43A�喂{k��������}�W�ɖ���g]���<�v�ɺM��B"*/x�>�Bzh!#���Ŀ��&+�C����u��A{C¿&�bR��P߰Io9����]�7ݪ���%Y���[�o!ݳ��]Hu-$Y�&�߃�?��J����U&����;!��ޟ�<��-��K�WLگYt hM��$�B�A��O�,�,�S�����.��0�J�n,����x���}<�U�e�^��x��(�}4��|���N�������h��^V6(���E�b�wp��x�]"p���E�����Pi���T�u
�*��D� �i�+t�U6�:�uC�\����+�U.�/�/�^�Hx��32�i5��Ax�,:h�v8��n�&/�Fo�ޙ{ ���2���� �5�Ӟ��H�@6Yma�  ZBl ��`"��!Bc�Y��'� a&L�1�ߘ$j�T�'�*��+7K�L������7	hFY �05\��CUq�b^�$��t����A�26]����xF�bQ1��W� $�Y	� L�l|G@Ǔ�( �L���gh1	��A.F.��P�N���!-�)+C��LS[��.,�̂�R�a��[ �Γv�{�%m���,~G��+Wzz�}�2 r����KU���5�%�g.�T���޲N���,yC�=�7��E��Z	&چ�*# >��j�P�q4��]��3�,��Y�h��5�0�-�m-����-���̡��m]�#}��v��?�����2A%�fv���
����?�ݓ�����N�=<�ijc��@��\���9<��4��?cj��eHd͓ 8�5�m��&*e�ʓ�f������\35!Z�Ә̭	2:�$JaM~E�/P�� 2�YD�̓���ͮ�V�+FeM�� �&�>KM�� �f��y���ȗE�45�SQ&י�J��։Ȧݣ�֡��l�4�4͡���>���b����]_l��z�������J_k)y�����Ozk?�����aY���7R�͡N���4�#
����@yRd8��]6�n�ï�2�d����zJֻ���%f�bt�c�ő�ĒN����ǚ
�;��O@C����l��_ �����'���$"�D:N^�:F#b���9�C\�a�tH��H��r�!�~H� ����i�Tt�^%ljvK�{��	�������faw2�;����YR�41v�����)2v��#����M��3@XӇ_݋[�Ư�"��������FL���w��R�KA�TQ;��6�YEn�QZ��v3�b� Z��v;��Ʉ:N�����u��~~K@�u&��B�Π��/���Z=�f���%�vI+"�������t�! ��1���U��x��`X,"�H�Le��m\)`��d��<���p�|>�Š�� *�F�����6G#T8���Þ�5�����^G%�ƣ	*�A�1�Ha���0�*���2�Y�U4�
2:B%@(����ccVįYM�hr����9����gOq�ь�S�[o��m��<|;iۍ�m��÷�G^��n�7_�\��	�Ϸ}s����z�׻����[�|�#��m8�8��|.��Rp��{�%��%�s�q`^�yPݺOײG]5!+� ����f+ߤNoyJ$�\�)U�H�6�@�yd6�@��*��ƀ׀�Ԩ�a56I�IѢSu�=:Ӏ�6�sM�<^�b�DMM�����R�<�_�(�L��I���i��UEP��Vd:�z!M�$���G�'��%,55��H��nS)��4����0�i��!u�5?���|ͧ�{zJ���8:�%��(�#`� "�4d<�J��!<�B�qZ&��!��T��R����L?�%����<�\7'���r�2�1�Jε���++��̶ҳ,�L+-�BM1QS��$#�#��Ĕ4�jm����6�|���?����\���{WN>�~fn�'ͩR3�}
r�����Z��VZ���o��8@���a�E��g�䛰f\��55eȮO�65�bj�v�� @�6�D���)Y؜�oN�$�ZS���T�=M�4�vG�Й!t�:2x��L~W� Н-�䈞B��'[�}Pt�I;�e��yw��'K�З�5���Y�?Gәch��7��R�`�ݔ,nN���)��L險$U%ljԩNIsE�����G���O���;n��|j�ՓL���b�K�t�)>-]�K�Q2��d9&U�N�c�p'56K���b�'X`"YH%6���?gT��AzM�՘�o���H۲%�ќ�x�S��#W֕��.P����P��T	ƵŪ�m�����\`)�3ܢ���P��r���DE	��	��,(��yjYv_#�e�����*��� ��
j"�<�����(.�M�s?K�h5k�
�G�
��DL����D�ԫ�X�"�'���T>�*"�ED��CQ�h*)S���d\��e0�\�F�1�l��c�s���N�SIl��Aѻ����uAo�ŐaФ(����]\�\@�j�Wde�tx��$��P,�#�y4+��yZ�H����,�)�r$R�Ϊs������������ܶ��ގ�-릶W�,�1U�c�t�L�����#4�8�r�X��gN��;�}�D��ѮcG����>z�ć����w�z��읋[�ZlO���ҍݍ�[k��_�����c]'Lo������ܒ��TGاK�ҝ��(���3r
��B"k(E:R��k�BK^��V�YS���p�0-6z������&|���rg@5T��K����d]�ɚ��m��k?�Y��R��R��A;�b�bs�Q��q���h�΅�!%�״ПrR�N��q��v��j�U7E���5��Ar�,��T�r�����w=���_��Or�%ɹ��^Hv��&��װ��A�ｲ�;�3(����A�����{������_�(_�I_�_�_A���H�H��a��H������w1���cP�`^�ÿ�&�����&?BA������O ��"FM�C"pO��%݅m΢�Y&k�`0w�ػx�=��x�H�C���nS�7��52�*]!C�!�E�t�
��묈��Ss�Ͼ�a ���k����{F�;�5��D���`�-����/2���Y&k�����-�~�Դ�����2��5O�)ĨO�Յi�I���ǚ&Y >5ZR���J����+4����d1�����Q ���L�� ����C��h�Pǥ�Y��A��h�M"P1((!�C��2*��N �4,���2	8.�6�g�eQ��#�֬��9 qՏ͌�\-�֯li���=9��\K[:�3wo�f�H7P��+T��K""F�D�����v�������WL�w�)���DdMhkKx�-}�#o��l��vfSǮ��M���<5�|�9>�Ț�gj���{pz�������G������S�8�'Yjg���qR��޹�l�{Wd��'���f�ÿ�;n�r7�1�[�wdI��������1��Y�2�D�,c��Y
8�4��>@��De�c��A�͓ ym�a5Q;�Y*k�i��Z;�DM��R�X�q��
+�l/1���h7&˧�̧��l��|���~:�����/�;>���Nw�[m�o����V�NS�;uE���U�s?/�F�u�e8i�S���ć�#|����X{L�;�6��Z��lw<�[�U����iH�P��x��	�?���`�ј�h4,s,������;.��b��'#�p�D �C�c�<�����)��Q�0�pX�JsDB>"��S�(���j8�氖yh1�65���#��@�E��B�.a����Df��s��(f��f����If��%�5C��M�$�15�n<lj:�;k:�Ǧ�����G�����EM��Ԑ��p@M��h��Z��6���js0a\��b�i:�Π�5(lMu�%�I��D,k����#�w����
�����3qӴ�D%ë��5n�Oĉ���Fѩ<�>Z�T��d�)42������eryL6��d� ,>�-b��L���S	��=��J���U�׈�T�l<��AcQ`"@���0��gD� �W���Z��į��c^x�zj�j��5�+W�x.f�
�H5�y��-����SzOfl��z/s��������m7C÷����n���x��{��w�p�Ζk_�{�/��ө��v��ۯ����g���&m~�=xʹ�g�y_Dи�] �6�1��tP���4�26��K�J�C�uC��Y�B��ոs���Ϋ���|��)Q9
U�$Zyx�
*������%ip�:t�&Ӏ�2baMc&�)y��<��F4����	��$�I򪰬&Yِ�uy@��Ue��A��$}��I���htBl�bL�j��4؄X:���Բ�ԏD5(`�&l���t:�qyrF�dȌ�O��� �艂��i���x\D�� D46����1	4<�M���
)#-������d;��͵=�b@T��z�^F����亨�nn�CP��8��Nv����`�8�6f���lby����nQ�'{K�=��@C�O޺�o����7�s���g�:�{l0ۧ3p�!=���2ы����> �kY�,���Z�QS�4�f��:jj@#�F��f@�����$^S2�9	f��y��F5bjM�LS����;4QGӛ�B�ʐ#�S�p O��@���ܕ���3����=�Z@o���ښM��(�\Ҧ�c����w��c�_}��;o^�{���S�.�:�o|KyZ�)�xdl��
~[�͢4��&�1P��d@���@[�,�����G�l�ĮK�4���3�JPw��ڲ%K�{
U�Q���`�t�D�[��/���t�ښ��EAY�K0��*�Y�Ԋ�R.ģ(dXЀ;���{�)�ň��-�y#�qO)�,(�J��t��ρȃ�)e�|�DD�SC"@��!��F@1	(AL��Yh-gANͧe?ijaS#UN�B'���2!O��Yl-�����"�C���IFs����6$+4I:K�ژ&Ӧ���<E"_��$������|�ޜ]�v}k�ty�ƴ�f��@g��2@?h(4)E�D��3��4�6���hd	QPL�J���J)�'g��L���Q����q�C�9����e��5�=5��nl��>��g�@���U�g���=���Ⱦ����흫��4��uj~��#;��<|дkg����3��|����s����.�t|����G��>سk�idc����-����6��o����i*�-\�PXV����OO2���YU�S�k��EFv��V�%j�B-�PM�ALM+�� #�nc��?T�
kw%j��c��&�n��Иu�6�v������6�]/Μ����Y'8�k\�-*�>�����-x���d&��8���'?�J��0�l�]W�.��IsΫy�,���jߴJ_�+^w���j?���3����oa�ߓl� ��B�?�����Q/�5zş�߉9����+`��C��E�%��s�g�W$�D�d��|N$~���' >"@����wЄ7Q��㱏bq�����0㉯%� P$���DLͣǦ�e��4�LVs��H|"wH��D�t�H�J$]!/a.	�)�+t�5&15H@�5+P�8�ż�R�e9��JpF'<n����Es���?��n����<�� �jS�ⴅ�KM"b@�;������ j&z�М�l����6�8,��֜"iJ�ևd5~I�G\nX`�&&����lӬR�]�B�ɘz>dR�~��nQA���y4�I|
�a<2�*AH#�Sb$�\	jpN�+Y�����#P�1���'��/�5/p��3��Z��3�
�ʲ8�9{��9���`�~}�n�X���ɣ���3�h��MX�f��ؙ�^S��Zm�Abj6��li���S:��avk�{Ƿ�X+O�8+�_�a5 ��Y|cj�߽ob`nk�Ć��S��G����|_�j������z<�e�&ʳLͷh�F��	`wObW��=K؛�lI ���V����Ҁ�Ec��h�(�M�7����&�k��-�U�1�d��e�f��(�$��1K5 7���fr�y�65c�D֌�����'�C)���hy���M�޵���64�jj�'Cm��T�o,|�:�nE��Ҵ{E)���yT
���M�_9.zL���i���8/�kIԇ��#2�1����|B�:��'��a���#X�q<�8�p�;���b�`Ї�(��O���5��NE|�D�'���H��dX��B��,�I6�8�6/�A���R
���zLA;����F	��2����Jx��e���[D�) ���w�pS�x�45n���i��'�1S$�	%�F	�uOpkM�����M\����t��D½\�% (h�JZ��֥�ujh�j*�E���z��	@|M����b�;Y0n6M��w]!aGXҞ$�J��$�z��!Eg@��wUM^y�S��.)u��B0�k�r2��M��$^ɢ+�4!��!$,��˒��2�X(�D�T�7�%b>�M��r�D���@�B(Q�DJ�ܨp&�2J2�ʲ<��]+��	2��%��`�ϠS�l�Ng��4�D$��X�ꄘ�V�8vŏb^|.n��WĬ\�������V�1��Lͪ�g7���.�O]>{�~�؃��$��	ELM`�&�i��rn�b_���c>8t���gso�}��{�s_.�������MG?��\ֻ�g�9��s�M��[�l��X6�4��tP6�Q5���ϩ*FU%C���M�[59]��j��X�+һ2��D��.�h�<��%�3��. �������⓵�T>݀�0b�M�3>�L*���4@���h�"7-�i�e~^y�_פ�jS�5Ɋ�TuC��:IQ��i6�_+DL�F���@LM���k!s<0y����Ɋ���LM�k>������ES�K@j5	��c�Qq 
&��F���:!�!�'މJV�^ܗi��9�E^q�OT��x����j��^���\�B'/�Ɏ�f���ee���8��)�f����ޒDW�$�-���;��'��u�����8�������s��e�;+�H/����"��L,�5��q@M��4 81�cS�T� ��5I|@��,Z��)̋�D�|���e�2M�\�,�{���zs��3��5G��ҀÁ<�`�n��ؙ���3���[7�X����@w��5K_���J3�T.YcY���[��w�����yt��Փ�O�v��ޱ�U��>�0Q+
�Ya+�*�4�K]"�S+�2���)�fP栖;���ud_'nc2��;re�y��%�bSӞ#m��eK�)��[���:�{�����"x��e��u��R[}��0 Os�|zN����I9d>��15�,��屦�G��^jj�� �x����-�,��#"j~HS�x�S<�/ �e�����		ŭb�u���i�(O�h}�U���ur�I,������U��d�#�(��+m�U��u�`�>P�	��|e2w��U"q�E{��Wa�$紷��ڰ�D���ꖉ��6or�3T�� @��t���|�/GkMH\�A��si2
���1y$��ʓ�ybG��(��T�!�7��|�9�Mu�[6�M�6on��ܳ�{���};���5���x`W��-��6�ٰ��ம����tf���M���w���<75~��˿�酏�<�ڭ��.�ua��闎O�9���\��֮��]#[��7�ml��j]�ZS\SP�\R�T\Z�����	������"*6�aS�gi)�(_�/P�(S��`�����z;g2�� �@@���������4_�t��ᡗם�N;Ӑ{����`Ã��r���5�e��\�Kd����w�m�f��ǹ����T��\�����4T}V��(9p�a����R	��D-�f�K&�U���C�K�K�K���k���!�_�օT�B��a��B��'�M>���w,k� ��^��%�����͢�����}E�~I�I����EYC$}B ~�'��oc�o�	o�����`^]�~y��5�q�G(���MM<�>�� =�S^#P���W����05pX�S�5�,psO��'\��/��W)�+T�u��y��5\�5�*��hj�k"�H@�E��^|�$��J9$���i�`��rr�ej�"{?��`�ӕ��H�5�2��\D�<��e��Y�l���SanS2�1�ٔ�4��[�"���Z��)�ư�.(��JJ��l55,%ZyX�h��2�W��k�>54 �Z�=J�KΰK�1�@,�7��t�=K|��X�p*p*�V�� �b�t��E�1|R��dC^�6�ؓ�,���9zs����%��Bso�n�H��Ը�T?X��/R""��Ğ,��?���`15�6�f��V�llڵ�w��=c[�c�'�SeMT�<�oL�����G{w�Mm�>4�qp��JL��y������ݽ���05�R�U[F�c���%�mU���D�Dj&'��*�e,�3K��Ԁ�2���� |��A�d��.Q�d8Dz���5��ˣif� �@zY��8mM�q��4Qn a5c�ֱb�\�{8C3���է�%?��x[�'C�o�W�ѳ�akɽ��[�JS_.�x�.�na��yI/��fo�xo$:���W��F�9����|\e<��S����j�A�t/���B�Q@�#��zC<B �c�0��X4`*���c�q�!�	
	p�L8D� b�R�Gi�ct�8�r�M;����1N
�'$t��D`^I?!jj�D�>T��+���H4m�dqC�Y.~���S� ������OB($�f;>~>n.f>fn�z����~��~^��"�U�՝��nz|/�����=�z�_C��Һ��N�=B�~Q�t;ـ����p�#����4���
�:�ŝ���9�'Iѕ(���򶠲�-]��:��.I�]�bd�ULF��\t���7�z[ɢJ� P5b����1�W!ˤB��'r�
�H�J�9O$�pt��!U���P�U꥾�+�,;�<Ǘ�V�!�O�KX�'��"�I�2���ׅ�6���IX�*~�JT�q�+֬^�j��=�⅕h�Ɛ�3��S��[&���d])��v�ԣ��7#�}ۯ{�����n���vӾ��y�}�I����'>�/3o���7�|����[h?�q��}_�{�q���k��/���[��3o>k�p�8xR�;��8�l�'�ߡ��QUM뫧�Ɣ��%���p�&�F�-�83զ�R�I�R�\��\���P�r�Ew����'���&\��k!�Y��L��"��A+tQkFD�p�����*IR�*�KUզ(�R��i��DY�[�i���B��e�%,���&��Ĭ��15HAfYQMfYȄp�����Ddѓ�A!��TӐ1(2&����`bh�-e�4"�E���y%�4&N����y�n~��[��仙��Z����:9�^��ȷ3aMcg�8�fJ�����������ԬK�����2��G�����?|��[�^z����7O�\�4�����add��Vz��Zl�[�"	�5�AT� 5��y2��2 ��  =��y���c@"15��4�e15O�4���o��2�����U-v79ʮ�H�M��'[� �p��,xTo�	15������CG��#�Мe�M7�T�nyCiҾ��_����/��g?}�ׯܽ~��ك���=��� -�(˰*R�ےgg�%N~��S�`Jlt𳋊6��o���z0H��	ZӅ�yr@W���5PQ��W��W9���i��U����15���E��u�_��z�\��i���b��K��b�����
nX���+�QM}[pG��<o�'
r[>Y"Ϗ����Gbj�&��g��T����
�&d�Q<jz@�S��׈ !�4dT��z��d3X��Ji���R�_�Ob�S��I�T�Vc�n1絙r�9m��FUf�.��PУ����u*2ە�M��&oV' ����i��w_e�u;s����=��vP�9��sR�5��(P��dZ�J�I���K��"!�/dpEL��Ñ��r�(=-%55911���2Ҋ���uu4��5n�\3��~t�en�cώ��;���v��yxgǡ��ûz��8�㉃�O�v�ئ����Ԏn)��۵s��+7n~�����;���>wld~���=���ݲkz��m;��N��oi�io^�TU�.��������<� ӕ6��eM�E�hj���gL�R_��8㞅�b ��X���dݮ�v�_�YMyw����?��z���pm�����l�`j���)gݦ�.
^����p�l4��A�;�i!;ma}�����覅��?n�|�2�f��G� >m�1��ȧ��V�m��U��u��]����^�o��[��l]H�/�Z�-) �Bر�/8�0�����I%��Z�W��"��
��`Q~J#~ᾄ5�+����%��L��@����!|�ÿ��yK|�Y� �ꚄWV���`^�ǿ�"��!����ф��!��+8�w��hL�=� �:s����������p��t�J�F�]g1nrX׹0�8����}Uȹ,�"��Zp�,=n�vJ��%3^�G�����bo��S��40Iߘ��t���e�&�i@;�>�)ܖTvs�%�@�.lː��˻���ڶ4ms��.(�p
���%�ƍ��PV>�%!�����PQ�r(I�J6�@;Q��i~ls<j�[�5������A�T0\J& \�6���ͯかA?��!�7�j8���Hg�UZ�d�-�m(�
}y���`��Y�?{�D=P�BDL4�f��YJ�� ,;�p�����`15���ͭ�#�e3��w��ݴ{t��ѭQ/�,��@T�<�oLͅós�:��v����<6��?%�Y��$�UO��K�i_��/�T�ej��"��A.Sg��{�Rvv&m�q̴�*�۪-����MDB]�#+�� �'Y&h��SS�cj��15O� ҳ�����2Y@L�2Y3Q�8�L�DA|bj�֙&֚&+,Q����2�x�u��<U`��2���>�����O����zo}�������O�;Ϧ��d�o�og�do�����A�����r�h9k����N�L'��Z=�N�W ����f0�3X�Y�cL�a2m?�p�D<D�#$��á�d?=O%�� �1�(�x��?�N���l�q�8�~��8)`�����2Ƽ��4 8I����9���WR��ɑP�1�i�x�n�����&h	�P`�3���8�$�0AA���#��!\�f��Ջ����á4���b��1�КJ�i�y��_((�:F��ޭ�u�i #����0;l�n'����qq�\l��Ǐ�A4MO��',�Nw�H�mj������%Yk��r8��VaPC��H"b���S��Z]ɡ����0�Db�� �)���|6����H<~[^aFnA�Ůc�!�f0��:) ���K�U�S�Z���e��E��
I�f hx0���ph"&��K�_�ju̪5(Ԋ��VŬxq�ϭ\��j4�D��݉�:YJ�X������E�N�杸������vյ��{�m��-ۖk捗�[�*��/�_�r�џ�~���ÿ��E��𦋦���Σ�-/��o��]DL�i���Ic�	cＮ�lj�v�*�T�s�����qaV?7�InЦ6H��2k����lR�^"TH2�o���2X��T�ԤH�(�B�F4�*�S����Ɋl�D�hfD�p+�d�S]��>M���ڠ$��O�}j�UL�	�b&����_�r��U�7�q4�,�e!��:S��U�(�|oY���G�A4kx�7f��J����d���P0�*F���f`e�8�N����y�y.v����b��i�.j����?N��[dg��Y���1r��=�DI5�ҌL0&��yn]Y�#˩��>xp��_������߻p����O�ޘ2�ؐ��n�ghIy&j�*�QKl�b+��d���qQS�l�ӓ5�!�2M屚����0�%Y�t�S�� �K{����Lѓ�晦������K Q3K�2e钶4IG��+[ߓ�(0�Zן����td*�r�m��cqH��6��vN�|����_��;��ݻv���C�N���__��jQ湵�6y���zz��W��;Ye�޴3��.*ڢ�,b�xͩ4�gy��2H@Mt�S_�f�T��5�(�{��=���
S�Z[K��,Y��$ل.-Ǣ`d��%���3����Ԁ���E�hp3F�O/�w�%��!M�7Ijpp��H(1���B�U/}�jA'`�-b�yNP/�>��gֻMf�Ѯ�:*�L�듥�l�5��.㇪��M��]~���_W4�����aG݄�~�R=���{���e����%�k��[�
�v�v�ͬ� ���^kV���i��q��
�|%m��:c�P��493���Xd�5�B���g)��gs�<���|I�PJr8%%)-+3� /� ?���?6ںus톁���]sS�]ho߾�={���O�]x��#;6�ѻwr�����3};�;���&�n��w��WF��:�k���'�]��uy�����-%�5[�ƶ�Ll���2>ҿiCKWGMC��ڵ9Ei%�e�����d;x��%u�Y����qL�f��SM���L뷳�y�Ӊ�!�΀���p�0��]�kÃ���y��r}���gv|�{����;%�/9����K|�k"��r��՚���_{�-�v-�ؿphn���gM�k
����ǌ�:�wL�>k��^�iz�o�5z�_���
�0�1h�[ؼ��X�p.�;`S��X9�����f�_t2������x��~��|E%|A� "��������%��9D��H� ��[jjފ,�z-x/�z�@xE|��Gh��!��K<�}�+8�L��<5w��x�-�&w=�
��e�U<�*�t�L�A��`2n���k��ᱮؗ���R�K
�y���^x�*=��sKw��S>�v��P��,�Yjj����%t��]I�Fq+HOw��Yt�
�eQ_�T� ��&Uؖ�o��f��2�b@G��#Kޛ����udj[S5�aE�O\jc��~1�#¸�h�����hia��􌥤���T���j⦘��f��[�?�e9��NY���T�e�b�HԱCZh�'�����DCqP��V�w ��������`��?�֗g��7�����H����e15����(�R��(�e�K��aj~����hL����# �XY�2O�Ss��������ݻ�7��:���JL�R;����Yx	�w���"�iS�	�(�����
�H�i���O�kO�s��Motט��Z���D� >�I�ڙ��S��"_�4O��}�vfSS�Ț��,s7KeMT� �f���S��֨����̬�L�3O�5�W���M�J�2���t�m��6�����m�d;.�f�o/}C��������p�Y%�&�~��\��b��j��z��z������x�n8k6�3[�͖S&�	�i�k�G�C�A��w�eb1�ө�h�>p�����,g�A���1�G��f����c�)!��1&�q	s^�D����((��JXրz���WJ�#�v�Ȼ��\�,�0���SQ���QR�1 cP�89a��LS��(�&�o��l��Ĭ �I!�M�MM7�4ݔ�N�NzL+�������H�*�zu@O��S�u�.=��H�2ӻ�n'����vsz�<@�����z$��#���+$�Nu'�{�%QSӕ,�L��'�[��&���)*�	
͂B��ȭ�`�k�$P�/ $��0������d4�E�r�.�/`	E��-r���i.^����0�c��}����CcR�:��`�������ʒ��`ث7j8<&�Ees�t��G� � ��!��G��DL:nM��^|���1�?^��Gϯz����?�r�1�B�i�irwAj�X��ۯe�~�=��s�X�_v_u��t��q�ݱo�m�z�3~[�vȱ�|����.}>x����O]�q���t���N�7�����h�xּ�q���I}�	C�	}�1U�Y�nqŌ�j��rFR4����%���d�j�=GlI��M"7H%*�X�	�rn@���IZ����'��,+)�J̵�
�P��\정�e.v��Y�#���ϊhx˧u�"$�15�)��de�O�c�Oz��eS�B��E"c�bW��r��7�f�Y:�B&�`�&x�%���D&zO)X4�����D�i(X;.1^@I�3���1�&���D-��L1fV���ce�;�E^��]�fF�������8%N.����"����w��pv�L#��	����4n}�V6����>xp�7_��֫��=����7O��R�d���a-�HK�CyZ��Tj� Jld�� �5��Ҁ$���uO�/@";�ؙ�v�T�  ��aq����N�D� �aj�]Y�Y��h��<�7vf�S���)}���9 �tgI�:�� p:;2�]��lmw��74��'Wݑ��)0v�[2%Ae�G�P�1���{7��O���7^�t����3.���o��&��>m�G���xeY&z����
P�d�;ie*� ��0jCldn$�f��A@�kM�_�,ӯ/7�:"k��j�ս%���1������
�l�8l85p:a�����<�I��~��8�pT�,��z� 5�z�ZpG���#O������%��Ϛ2�P��x�'>�GJ�0�>�,&�5*�_K8~�k������z�G/w�46�ɤw��.��#V��4����.����z^Z�8�[�?�*ި.٢,٬)�U�k���3��)ͺq�c+
Ԍ��F�գ�]{��-8\4x$�0�Y7l+��m����3�ԙm��nwy���Ř�V,2�t�T��.�E"�'�r���"�Ig0hr�D�R[F�������!�ף����jj��j*��*�۪��6���nl]�2��mrs��P��pߎ�����C}��F6�o��=��oj���=g^���'o�tj����ͭ���6������_T]^^WY�PSYWUVQ������������K��:���:ˣ�u*s��<���(���)��H��3
�R�ۦ�5�.8�^�����lvF�ҩ�rWP5�������z�O�m:�Q0�.��WO����_^�����w������9.��7����_*T�J$�_d�/̎.�tb�c���j�����^�X;�h>j�������e���e���W��[I-��,��ʯ�ҥ��]�{�^��ZH�-�u7�k��M����:�_��?(x�*f��}A�~FJ |	�J�����F|E%��}J�j��`��� �`�ocpo�AMxKxG|KB�D�����c�aa���c�ej��p��x<�{���J�w#u3����D�ob�A!��:��,�B4�2�uYȾ$�\�p��f�(<j��wJvy�3�XP2m
�vf��A�i�v&JWR��s�
��dYfg�d��,55߼C��=C ;�,!�#Kҙ-�̖wf+zr��Y��teK*LcXQ���	��|#�D+�2�7����ғA'��N@���g��;�NA�KX��#@�O
:��2�N0�������kゞ�Lsm��&E��dmU��!��U��X�[_�(�Z}���<�3L�����4��Yz*�R5��������М�䩙��87Գ{d㞱-�Ƿ!b�IS��n�15g�ONmn=8ٻg���L��=}�Sbj�eOY��$���/55{z�M�]����j���̙���Z��5ӑ���v��$�M�h<bjA�.�5ț<��̴xf��O��"=�����M�� q4���kp!��/55�ն�*�t%,k��f��<��5^h��lKV�&�&ª��r�#ۛb��6�A{�ڜ#ɖi�h�M:0vkNx����K��+���A�e���r�n9�p�w:/8��l���I=ljN���5��r�ash�n&io�},����a6pt9�#L�a� 8�$�s)ǅ�S�)pR�>!e��9&gU�,u4���C*�~99*k@�O�w	�����<h�C�f�&h�Qr�1v;!���LPP�T�;Aō��ۈ�qk1��0+a7�^�EX�IZ���Z�4����Nfl'�W���zuPk�=�KO�0P:M�.������:��������<\@���汩��D5�+Y���B�f���#��)*ܲb��̯+O��� �o�*�E�3I��Ĥ�*�|����Ӹb�T#��t:�N����rw�SX��}z�����s��ݻꖞFG�*T�N��er�)��Y��ጰ�f�K�$Deј<����s�����0He2h�HOFxlB|���?���_X��x���_^�_����?Z���x�Fc*ĺ�ԙ��>���T����W��w��8����]BL�g�{��s��m��k�v�l�W֝�8o�+��3'/ٺ[Y���֟so�`�t޶��u�ǶK��Sc�;a�;i�״T��U��Lps7�2�E面����g����z�Xm�*�
�V)W���T��Ԭd-15&r���k##���I)q�9!lj�ݜR7�q@+�i�-��]��⨩�IV�Ij��,3+�*�8V1�(fH�bj�c15QM�L��3(0mCL��-z��M����Q8<�4D4���b�i�X!�O���Pj6�( �f��=r����)�&zvd/�#��.�p=��"/��KG(�0�ݼr7ԥnn��(v2]�+��#�l+?M��q�2-
���j����~�ڕ�~��;���������xt����[KR�v)!���23���5�!��5�Ț���15KEL�� ��&
�[�KwK��{���ʔ <���15р���y������|cj�aw��~S3��Z_��#��zs��9����&q�Ț�Y�������\����?;����~�����7�_�ui���}��m�)Mu�����ħ*rK��\+���/��ֺ�0`<pz����	���쨩Y*h�#<!�i �%ځR��rV�i�qC���T�]��[k�di���L�8l95����r4b��/>���pV55� ^��򤩉<�Y��g���'L��5M��,	�A�p�|��I�|��h#db�������"�=:�G'u�6�ڬ3tN��%Rzx��Ȑ!v�p���P3+��M�f�I�6(�ԥ�E�d0ۥ��F%�#��!U�&sِ�x�m����C�[N�M�>h�u�L���=��Ϊ1]�FiF�(�U�٤�k�e�)�e�@�1T�sgJu~��*�yB�'fsxL6�J�Sx�AX<"s�,�Tf6��v��l+�R�Ve1�\�ǩ�� �S�6 ��gօ�T�3+��Mre'L�N�� ��y�Ȫ���l)^K�'�,�y}w�������t�ͨ2h�6��ew���fGF��ZA�ϭ�X��4�&�2Kҵ�7_�*��{?!���@.1�(S��d���?J����]��n�XP�+Q}:ɰ�*|�&�˙�����,�˳��ޱ��w�_������?�n�_�y��?�f�$��+���b���څ�}N,\?���K���Og�|6=x&/p̧�v]v�w	�#j���[y˩|١|í����ħ��*�� ��S��d�B�g!��W��on�߸�,L���d��^+��V��7��8�O(�O�񀥦�gt*����S�.�>��4ط�pp�;�=�"�=<�m�M��ܣ�h�Xb��<��Q_���刦�����b��.��^�������IX457q�k�U"�*]��I��EO���/��/I8�eܳ*�I�`�(<l�s�wz$3�xH:�(�oH�	�ejz�@O�7t'G�8��d>��	4�ғ.���@4=�z�!Cґ	;X�d�"�Fڕ� t����ut\I������[��y��L�T�-Jffff�R��,YI3ٲ���m�ٮr13cWWsWW�^�9+K�k���̜�׷��;�Δ�̈���H��%I�ǋ��#9k��0sMc��6Q�/Nz Aސ��r��W��B@�2�_%��	��E`�P���x�n~�GP��"E�TS��@��S�4.�W��@�'N�?IS��kʲt:����&е�}g��-[ג�i��4g*�rԝ���e����H���e�����8�;L�?,��w|_]�`s�XǞ��O��|LLͩɡ�-S�q15�SS�+3��3KS��'� ��Y�X-<��,�X8�����;��~D�<�5�S~Se P��`;̙�Xh@9p�hɩ��Gr�#�d��X�w��p4��6��~� ��0q r|���{
V-Ъ@����/��� P��l��?A=4���u`j~�����G}�ÌW#�4����	Pc��I?e�e&?�T�c��>Uh��6��j��CQ�A��X��D��X���[1e�L�ZΨ�=��4�fM�E�l�$_��.8�W��K^�y�uÆ(���t֬[�)7�u�b]+_U�WT�%%oQ���N
�'��\2�4�2˧�	��b����ģ/ri�l����c�
K\�2��, ���kbچ��!g6���޺���`.)�e%sI�\ѱ��c^M�9�O�ɳr2�䓒��9&���PG��iv����a�)�1r�1l�
 Cä�r�(%Џم$�A=��Ӷ��������f�?p��4Rv7QCiH(M37���&Bw��]*R���m���h�Fj��|�@:h�4��-NV�����6�9�FIL�dp2 �P�D�a(�� ��ĝ���TyC��9IY++���L��H��x�gmvtMNLj�ΡḌ"�I�5i<V��np8�6���5#-2��m�xLj�ٝ���W^�=Իtq�ޫw���w�|��7�G��s,�v�ۨq�.��k3G���bj�j���фl�T���h|�A��Il!��g�<��@
������������ߞx"<,�
#�0t"Y�W8�wqgj�bҡ���K�÷"'�������������ky�1z?r�롛ƞ���XU<��=fh�s�\�w^p�_u\5umZ�xm�9S�%}Ϧ�㬡����e�иj�_V���*�	
FY�}��f�~l�4�\����x'On˴r�Z!��$"�Z�f��0��3%�LI�"�&�F�wR
ݴb7 5M����7E�'	I'\�yyNN���e�&�^�,�(�)�dȓ?�yjM�_�%<,$|��!���15І��̶�y����cx��=�'�m��_�������)��{�
�Gc(�W!E�cws�|�n)5T�B�h��c4�d#=�� �ܙZ���cg湘p��\'��{\$�ϳ��mLh��S:�d�fۑ;�8م^Q���l��8��v�Wư�(���_�����|��W�_x����+�6���"�y�d)�@*�	2�B��
�ɷ��,8(9H%�O*��5�4���Hƾx> ��T�'C�6�j�����r�Ә"��+� ���А�H(7#�~�P�M[�О-�ȑv�ʺ�� P ��4k�Ba�v��A
۳���	x?" x��	�-�����Ç��e�۲�`ߞ�n�Ruf* ���g��ӵuƊM��Y�d<=���;w��~��k�o\]�r~��;�#}����m�&aQ��8VS-ߓ�.��Vƀa4��E�ƿz��)�P˽��(ڞX��D6�7f�����s��f'%��iȓ5�k���yH���(q�[m�T,��*�L"�����D�a�=���|�l���o����j��Ԁ��|��?�� >�!�|�w���9�U�6�!���Ph"K�`�h4	NF!롰q!Bj����J��zO:V�����t����q���[+rj$�̤��&��!�xĺ8�>Yh�`[r�*FT-;� +���"N�e��3z%������aiް$wH�;�(�P�LZ*�ԅ�����ٜÛ��S	m1Mg{�L#��C��~�my�&�Ҍzi�^qb�8�DU ue�-	"]$_n�I\��×�x|�I��x&<"��]O�䧀]O>~��7�;4�Y�d*�	zL�'�T�&�H�r��IR¨��.e�&�pT\PV9�$��`�\Zo�Od�����Q�V�e�s[}��*�J�,2
��1Eb�L*TJEj�D��)%B!�!�0$"�RL5��:9�#cī99fa����c��9Zr����#�H9Z��ej�,�&0z�E~�ԹY�v$������{DcN�Wq)�<�c~8z���wv��/n}���{w����ߜ;���{%Y�\����L�k�
�m&�%���nMo=}e��K[o����sßOt�)J��I7-��dE�Y��6M�M���q�$|;Z�^��H���z���76	2*�Yc��G�G��ON�m��L�ou�߫��	���VL���v�O����o���c|��x��D����'D����Bw��
G����b������!��!R��S��Q�Œ�ƒ����_G^E�_C?��� <��LzB�`L�
pq3"p+<��ЛO����mjи�X��*�D�F�\g������|�=��Jx^�Y���U�%=�"<ew�&�¡H�@��Ǉ8�6 �,����c�����8�쌟�d�A1а4'	[S��iRpؔ(�e (�CP���Mhܒ,��R�X18�� ��@S��� �$u��$im��@�a�����	UQ�GR��W� ձ�=q��x��	 �A����`p�_�lP�LW��zJ��n��(���@e}�
������ں�s����r4-Y��,eG�֏�{���Ŀ@#���΄�� �k@%l�0��y�l�H�⁂�_�>����Ԁr�pd�0z������ڄ�������ړÝg�N�M�B��0�������q������噮�ɦ�閥����LS3?��C�V0��&�`�FA:��	 ���C�65�������L�GBS�5�5H�`P���Q0�lXF��	��PӀ� �l/�aj �>�V��q� �iv0��Yi���qd� 5Zn��f���	65����t�}*�2�aIRE����t�%��G��X��!)m\ƘV�O�xg��%��]{)�z5�}������;����v��ߴh�~Ѭ\7�V�%�hQ'\�
fU�Y紌uJ��JY�2����$�.K9K"֢��,d��X�b����$�.�(Kb겄�"��əkJଞ���h��j֢�	XR��5�E-s^˘�l����F�壧��l�4=M�LQ�c�QR�1l���C_�@�@S3B������<Չz�5�-�?i��	��i�=р���d�4���&zh#cw37�E�h�v)�CA�T�:t�6=��@i2RM�3��For2[��H��@YM �U
�l�IO~M�/ 5q��DQG��%EV#����U8yUI�[�'޼?�[W��X�Q�ዴ�M�ۮs��6���0�<f��j�s�ά����Ȣ�袬̽���{k{:��-��{��_��w_|��O����ʉ��})���!֫��2��L	q����+u��['ߤci�`/��xF-S� ��`D)g�$T>��b�T�y*�D��]��PtxY�'��ñ�2�ґ�.hMm;�:p���}�o�~�����ȑ�������Α{���αg݀����ێ��Ǝu]㼩e��}��w��u��w���нi�l���>05��c놱i�P��=���sFQqLT0����$�q���1U��R�-�o��T6�L'��
�F!�˄�A����a�S�e#�9���P��Fs � $��&YMMY��8RX��!���O�#�\����9�l�����SO<�� ����&l�S0���w<b=n��|��<���<���q�o45���|?����5��̣��d��'����IOR���d��V�%���D-%�D�0S3��,9�N�u�,|�8��{����F/�����B'��A˳S���\;��ϰpS�ۦ�#����3���^�����_}���O��c�����Ҽ�t�8J�O������HN���L�	�5��Xx�|���.�MM��'@��djb���?A ʠf��	DӀ���&!F&�ԀC�n`�ԀC�Y�� �&�i P�@�!hВ.�F摦&Xր�m�� �A���MM{�Y�;s[�|/k�u���Q��?3����Oom���7�ܹ�|a���W�F����sbL�~A��8ZY%ٓ�*�dW��J<�2���R�UDR�|��8Ɓ$��4AS�����#���v
� %ڶBMc���P�Td<�k(MRdFI�]b�YdU��B�<N�3HL
x���ej���k~N�Q��0X	�!�#�aTT(�'EHhh-g��"5D��MM���ձ=z����4
�z�K'�i��¤�i5&��!VG
4q\]
ǘ�4��lo=7���k�ǵJS{���>YƠ"gX�?QLh
�u%S��e�!IvOr�Z��_�lB�r\�c�QS帺hP�?�*< IN�4�E�^'N��UJ|EW�����x�2+W���,���P�,<��h
�L���aHN.�����Ƈ��@��_�B �Hd��"S�"�����R�O�i\9���\�j���'3�L�QB��;���Js�nW����<�.��$R�D���4"��C3�x� �G?��W|�����++�_��!<�d�Rd�l����Ղ)����%R���h��D����F�k��s����P��{��� (k�Mr�75�f����x�CN��O5�.%�'��9}w�a��|�!���ӿ{��֛�}i�����7��K;!�]��q_S�n�97E����>�_�u~e��[/^��s��6���#�u�!/�S�
F�r�@n��U�kz�.��n�{��\�����t�/���x4���g܊5 �AEj��R~g�}k��(����G���z����s���>Ň|N�������|F�}�L�¿�E��6����� o��������@�ƒ obI/��_C����GL�
u;b[���5B�?UM���
���B"^�S���p��kB�e��NzQ#\Sr��h^�9c⟲	g��	�p$R8��F����Ѽ���恦�5�~M�7���~���r[��#]�.&����2��i����LB]��6I�]d}�P�(�M@�	����{$���[��	�A=L
���
���`��9Sٖ����w{�L Pn�V7e(��`ߒ����A��8۞�m�Q�f�;��hd�%�i��	���a��L��Gbjej�SX�i����H����3�O��[bj S
�$p!�Ssr�m�X��D��T������bjG��#��&�>;M��&��m>���\'?3��P�4x�|�45��Q۲�F�@M=�,�7y`^��f�A4��,�æ���~V�>��ɚ�&��d��^' ʚ	^�
�8���8]��,�O���ˍ�Q��w�i��<���t�i,]3��8���8F΀�}H�>�ejXCjֈ�}HB�PG��q!uRD;&g�iE�fՕX����8ϥ(�9�a�a��܌�_�.��ݺs.��C�j�.�ċɲM�d�͛�sz�V X�	�u��pY-XV�W��5])8��S�e�e9uEA[U�WT�5kU�Zӱ7L�5g�A�/�YK���qFK?���RSO�('�2" �ל��N������\�4;|�>IFM�0�D�85��" �h�H�a2
0BAQ�=�]�ا��O��~
�i��i$<	�7P�����od��"Z��2L��Х!vh��|�ר�7��VJ����f6{Y-��&/�����M����k�,MӔ nN��$I��1Q�K sRd�1�}���Q��ʎl������{���&{��O.����_Q���x������{�j�:��[����F{
�UO��-?�];6T;<�{�����^~����_���^���է�v���h��,�o/�i+�i/��*������mo�,/��f�R,��ւLcN�&=A�/�: �@l�D^��e�8l"��)����0"���l4��Ŀ�	���Ĭ�%���RN���'�o�^��;z+f��ȍȡ[��;=��y�_p��M�3��{����w3��嘡�C�͝�ݗ,�W�=MW��7t������㼮嬾yCװ�>���;+�<)/?*-�����u��rQdϜ�ӹ�J�H��+j�L�����(�0V�Iа���d#���!dZ	�����nf��U����e1� �~��=I��DYU��"VZ-)�z��nQ�U��Z$�`S����;4IR��ӄ!�jv��~24�ɿ7�>�G����5�T�S���Owo�=<no�oi���h:,J@����ۋ���4�p'�.Dy��6^�K5�2��+9�F̵�௺�M+�Ћ<�@y4:F��g�:�J��V���:X�6v������9T�V�[BIqJ�'Z�]:���_~����w�n_���qt�x_������h	�.v��q�ݠ���&V�#ضe ��@��Yx����! (�Chj�YЦ�K��!���������E��ۓ��I	65��6����	�	�	h�5����t��	�ĭ�(k@e�|�����N��zM���.?ۦ&K}0]]�a�LT'��%I��ɶ�>xfk������+kS7.,��k,ψ�Ei��Q�|�� JP�,/�d~oj~�h ��>Jum_�.�Ә!hΒ�8�	�MG���t��[��M��bCs��@��4I�%Mt�&�Q�T�"6�M#�)�!��ej��ozCB@M�
?��m�C6
�LzB#��HJǄ�I()+gb�SA��X��
,�8-����s��x"�Vb�H��^k�h,����d��X�T�>�f*d8�ّ���\_�0�E��%O�'w���9Gt��)Cь�p
�xR�{H�H�7�ڿY0~+�u)�k=�}�Yw�X=�,g元� ��~in�$�Y�R'N�#�.:�y���Ñ�X"=��dp��L���x4~�6<4�����># $2���2�L�ͣ��4P Q1XB�\%�YEkVZ��*T�f�Kb�8�C����OO�e��R�I��h�"�A�	Y![�g��$"&���
�`"ȨBĿaC���?�w�m��d��'�V��$))K��׳ru�l)�@���HC.�P5�Fz���k�i��@@M}$�!π��Hn}B�Ϗ�}��W���huq:ܼn7����q
O�EsI�&5���VF�X�/�9�^����n}��֋W}��og^�_�Z/��<�=��:_p�ɻ �=��5f�է��_�z����W�<�ݙ����݌q�7�d�3"ʚ�u^�?�a_аo���%���x�����YD���_9d_�Ŀ�����J2�5��W�;��[��;��wZ�¿��	~/e��O���k>�s
�S"�c�_ِ���qq��1�p����w	�w	�w��$�Kz�(�x�{�;D���藂x!Ṉ�5�#M��$�ƯiBCo����S�
_�@_B�/a0����e&�*�y]Ĺ.�]��.�y��5-^�>�a�4r�Y��_d�-�k�~��'F�����<�5�H4R�Դ� ;�"h�l����v�=M
�KG�~Ã8�A�L��p9�;r����{���T�>Ek�����z�]��$>�6I�v ��5;A:_>d_<�no7��X�s�Y��6�I�2���|]w���� p+��%K	� @�-Gݑ��)2�6]��|MG��=WՖ�l�V���@����	X0/� A%l�H����_bj�a15{cz$6L�מ�^�Z�>39�ð��55��{׎��;�8�tz��?;��y�`�lX�?�h��h�[	kv�f�9��;�M�̃����?Q����
�5�yH��@�2� #h������I��ng�	�|$�\S����d��Ƀwpt�0��	ʓ���0M�顩�˚�M�H�q��<Uj?Z�8Zh��1��h��}645}Zf��1�fV3�T�q-wB��1���An��瑧%�e��\��j��Z���ײ�6\�ٞI�܌�ވ�\�6]�2��Ҭ{U�^�W��]�j�]�E;�l-�e�l�,[3��M��F�9��I�i�_0).���Z���l�g��﬙�n�oX�f޲��`d�X PX0sN��SZ�I儒|\����R�uZJDj��)V�#d�:N� ���c��QlX��# ��@��TnW;��6�-r����;4M+���j�E4QmRt��У#w���:b�W�B�i�Fb����e���ޮ��i�dd� `�0��iN��&��R�`ߜ,�'
��P[��!AT/��W��N4m,ޜ�>7qi~����kO;��u�ot�o|�gf���T���Ε��kgZ�ϴ�[蹼ֶ�ؼ|�uq���L�������x������Ϸ���_=��{g_}f��b��h������ұ�����≱��ʩ���C�����;�z�;��Dܫ+���fh��LY��yT�hb�U��)�R�
��dJ!R9t��'I�*s�#eOB���ֹ���ɇ�%ߊ�;|3f���-���ȳ�c/ �B?=��o���p*u�ٌ�����F.�.����{/����k�.AS�i?�m��6�ij�U{�U�de3�)yш<�8�]�P+�*����(��*P�$
�J-3he&�ԪF��:^���CSCʴ�v��R��˫�V�� � 1�:Q��_��"VV-)�z%�6�O˷Ij.�KF��O��|
�CB�S��S�;"��ݻ�ޘ����#D�Ԁ<�����$S���A�~�;�n�!��P�A�E��<b����ᠭt���'i	�R�����8�/���$��P�y���؍�-�3�� z�I����;XfF������:�96E����:=�pum�g��{���37���?qai��p���J�scu��H~�nR�e�)ۉi(k`�a
��rCSSh';�eR`@�/`�/�����:�M�aS��$nHF�h���j��	>=��C�ґ#�j�`j�D���,E�����(Y���?��ƯiTp�SS��I2�ʓ����swk����y�ލեS���Ύ�<�R��V{T�,�$�+��p��$����v��^�A�>�~��TFѪ|��hjMc"�>�۔)l͑to'@_�㦦�X�V�k-1�����-�r�E���(Y�]�1�2��O屈,*�J��X���=���&��L�to���k�nj�IO(Bx(>d1�):&TH�(��h�P�*f���g��	F�Y�;�(�2����Q��AS��S�Dj[�T%д�tc�\�p��D����c�Ͳ�nyZ�(�S�ڣ���K&%���	uḺpT�?(���u&u��L��Ԟsq����3�=3��aE�ae���h����wKsڥM��ZqL�����&2�����\�-����w��(�ψ�ED���u2	Y��߯l�ɢ�$����8\*�E���*��F���|6���ӳ�R��6��f�&eū�
�M�щlB8%��pۉ�S��l)�.dh-�E�0јP��t�Ǧ�T>�£�9$�$�ѱ��ا�n�������D%�H�*z�������(yFj����%k)�Z����Ĩ��~M�D4�IOS�>�i������5��𰐜5z�����{x�.n��ݣ!�&�{�ԑh�P���O�}se�B�����N�z���;�����/�'_l���b�y�O��$�Y�U*�ŵu��֭+[�������Wo�������_��_�K{6�uA'�㓗��5笊��b^а�x�m��\�\����O<��\��-�o���b�[)��$��T���o��!��(��Y�e�n�V�1��0� e���������Bd	��	���B|H!�O¿G$��ǽ�ÿ�ſ�!��!��%��#���|@�~H�}@���ïD`^��@Y�|8
�\��<�B��%�Bݍ�65��Bo���En�~�����\�`6����E:�2�~EȾ&�]W����4�r��z�)���5c�N9cn��` J���i���4M`�S[���4��.A�l����)QВ,j����=�b��R@VB�I�!�3|(�S�r@G����i����Й�A{䒇d�y$�$�ޖ�/t�l (@@=x��tIk��=W�S��+1��WX��ʖ,9�/�М)��yj�7 f� �P�0�y�j��@:P ��0�S���*S����yj�ZKf�jgG���,L�O���15�?���\�Z=qx�X�����ɦ�C{��cj���t4�`�ljv�� ��;��`_�!z�4`^��-�ǚ�0�f�s���A�(���D!��η-kj����@�������w���ڡi��۪�!S��uw�Xx��Z�����h<N�<��L��K�bjF+���R�x�i��6Sa?Zb�)�Ld�'�t�Q��t�&<l��X�4Lhj��i-oR�R����aa�O�1N[e�c,�����t�G[�Nvߌ�ވ1]�5^�5��ծ�iVb��1��8�J�a9J��Q-���ŲS��P�ui�95\�K.�U�����G�&�� 6�N�Kz�-�s���+�7�fμ�sJG���N�)�U�cJ�19bj�4(��f�>��>5J�5���� ���0&�a��!"�3@� t��j�>��750����T3iW#�)dޓ_�4�#Z��V�M�i����.�WO�6���F�^���c,�V7�3���k��6E�"Y͑��H^cT>>�9NԚ��i����TyK�<t����H��4U[�a�*ac�v�g����;k'6N�.��;5>6�����64�69�y�X��\Ϲ��s�s{�O7_?�q�R�s��W֖*�N��]|���_}�������;�������VkO�Ԝ��81Srt*wz"kr,sz2��t��ugW��k�g�g����;9�93�>>��l��k��p�T��T[�ti��d��#5yrG���\&K��)�J�Ԡ�y�Q�ޜ��}�K��.'�L�7t+���衻��g�ƞ�1r�%��}��m�н�SoT�R��n��sI3ϛ���.���{/��/�������碦���i]Ӱ
M��⤴xRQ4./8"�퓦���k��|�=�g�h��F���t2�Ab׋�Z~�A���'�y�U�)fJ���fAj���wR�\��H~��W/B�G��fO�ҟTXQ#��(�*�ixd>CD�cg�3���ٍ<R킦&,���7�<��g?��x���15ඁ?�pX4&<���`�l
�KA��h��"��-�ƫ	�r���c!���E.J��T�"���b��C�x�?�C{ ���,u�J LnR�W�
���t5UOO�1sm�|�:� ��i�ڿz���W.ߺt���ӗ֧�燆��c��47ߧ� �ƈ��e��b5 ks�~�B����2��T��8S�д/�_�,>�*���Mt:�pO)"A��h�C�l�45M��PA� dN�(��F�ӝ`A��ag�e.�a +0�5�J�n�c���($|�x�ʔ�d  ��e{��1Mِ��NR%[������η_���o?}���wo�͟�v~nr��pkU�[�R�2ݢ//�êHx)�����=�,��P U�T@u�&�v �y0�ۜ�c��젭P�V�k/�w����mM%ֽن�U�Ok:|��)�QxL2�F$���<���S?��3���	|`�!2�1,�م��bj���4��K�H�Nç��؉FdE�d#3�̎6�}f��,�������,Z�^���,J�C��T�tM2]�Ͱ��L�nl-�>�A��$������~uѐ�tL]2�,V�(
��(���ݴP:y7�o ���3���ڒU�M�0(�k��}��.$aMr�$�J��g��2/Kde��L���1�<hj"�(4����л�#v���,C �qx�ņ�p�$�BA �#4	�A��t��Nۼ��zn��p����Q	� �^ƕ�L|]���ў�}�F�A���:_�WoU�����'�d4�I�Љ\�����|ȿw�-�'|�B�O�!�K��4���3��|=+�@�5P�M�\bjJ��2�{B4����ʨ�1����h7J�h�1
���LC��.a��oj��:7���i�p[]�6;�E����X�I�F#�����t�����ɢ�[�[�^�����,N�����VQ⬆�,�^�����D֦P�����S[￺���[/]C�knl�qj蛦��J��u�W��%u]��P�7T�s�9톉��S��W��O�i��S��#����7>����N��.R�K��76�wN���?[D[�_M�?i��)��Ji���%}�$|NAFF}F�~A�N'>cP>��?��?�? ��#����������G�����?��> �?$Q> Q�@a^Cc^E�_�@��B��bx���S<�	p+TboE`o��ױH"�+�E"�2�r�M�,`]�񮩄�Ԣ�Z��x^�;a�L�Yf���5M$�����;Hw� �=ꁦi�G4�%A �s��@�Pn�O}B$�߶�X	EL�T��15��҅��i@}*�.Y"
P9�
�G\[��=��ٟ�ޗ�� ԀS��Z�����"Mg�
��J�V�� ��y
p�5G��Ж+��
��,��Zr��nvR�~���Àm�cv��dj�a15)�3G�K`����ó�M'��55�6N-�t=�wi��ԑ=��150���T˩�-�&`dv ��e�h�mw\ ��s�%2X����
O�����4���	��a�"�� �^ �����`5�� �)��q<N� ��P;�ڋ$�y$���T�L}�)�M��65�妉r�T�m��v��1Sl;Zh=�g;�����Nz#6�sD�ѰGT�q{\�����Q>yBH��0�Y�9�M��Ү�����z��j���O)Z��?�]�׮&�W�����8�R�~1J��Y�jV=�u����x�g�m�k�k�c�c�k�����\�A��p!Rq�+[w��l�y3g���1�O'�~S���PS�����N�jfx�If�m�0��!�Sc�phj�1���`#�pG�������|x?.��C��`M�B	�/󴻑��o����v�M�k�c;U�n-��@�2�ڍ�=���l!5;��Q��.45�Ѭ�Q,8�i���� \�%^MM{*�i�YS*��5Cі�j�Զ��TĮ�q���瞻�pvv���#���G{M�8}�om�Х�}�/�_?_e���J����KkU���[ݷ�\ttz���⛯���/?���[�h�/����?߱���̱�͍��j/��>w�|c�xc�t�|�������Յ����������W��-�Ι;�23���77D��Ķ�z��:*��e��T�/Re6HU2��/`��,�\(��uZ�KgM2ŔEv�5����H�>�9z+u�n�𝸡;1G�F�5�\�����X�o;�&N�r��/�n}{��WE��dϽ����h>tM?pE�wIw��.�/���j�ֵ�kں��u�iiф�`X�{H��%N9(���s��D��+5X�V�0�'��e�u�x�8�(L1�S�쀩I5��SH�v45e��J��5	��D�@y�� �&I^��T�+ʢ%H^a�0�*�i�v)S'��x*.�
â1aa��	�Xa��CBCvE�<�
E"m��ՎG��m���$Aa5`�~�q�?���-�4��h&�J�p�x!�(f�l���3
p1.ZIL�S�-�<�A���R7�og�)�� v�4��=^:��p�ʜlD�8����J<�j���6�Ӎ�d-#�"*�j�ݪ�D�t���ɶ7�={���N�_[=uh��$-R�+w��r]�,3��I-vS��m�5?B�Mh�i`��r/=ؿ��קH�dS�P��@�en@`z|���%�S�8�`S�4ЭG� �c�( X�ʓw�+��6�hd:��aY��������75�yOP�@�!�S�'Y�faU����鍗�������gn�/��ua��P{_cY�G�V��<�\7�M/O��I�>jY��~ (�yO��f"#`j�����05��`Zԭ�ڎRSw�����Tb����+ӣ��6�L�[L�������_ p�X�u���C6�YH.t7!t71,��
�#,�QHq)XQn���h�&�Y�bb%�9qfa�Em�D��� S��[�Z�@�ei��t�����F�c���%�	3E�-��6E^�,�K��.����)JUeC��!Y	��dXW:*���$�$��V������w!�a>���c�Qc阡d���ae��<�_��-�j��6�����Em2S��9|��d�DL�Ja�/W����S� ?y�<���w���s<�����d2�F�18.�,�Ur�C�s�b[,����}�͗�~���_zfqm��HoVafjN�ΡWY����2�(�K����r�DcQ*�R��E��X,���cB"v��$���cw�3��E�N���B�����>��(v�S���"�F��3�
�thj��r=�{Mca�ؘ{�.6��ͪ�<�4�`�h��d45�#�<,D�x��m\�f���h2N�Z����hU�G��D��WO�p�s(5j2/�7�6�~���K7_=~䕱��۫.&�.Xu焢K4��5�e?��Ik����[�Zn����3W�|t����~����X��`M�:���Uq��̳Z���zQǺi�=����(N�Q����S���71��F+~���.��M�]��M�g��/&�_��������;�W<��L����ğ1I_0Ȉ�aR��)~YC��Lz�D|�HxK� �����!� oapo��P����Q��p��f������·P�
�n�p�m<�&�t�B�A�^�Oz�"d_��*W4�+:�e���Q|Rϙ4�ƌ�a+{�Ń�40�p{4��t� �5��B 8DӴ�E�15Y��ORp4�����S�9�\؃S�}��g?5�KI�ò�@��6���G|M��M�B$q`T�6e���2����ʦ�X�*TVn��ŶA��/k�M���h�W9?�4P���������iLl�n+��=p�H�����c��yj`��.� 15�fG&ۧ����[N��g�Ԝ���h ���ghj�=��w��C�8��5��L�;&��p�6�n?��y�g|����ޖ54�����m�aj�&`g �35^w���������<��&��� ���f��4VfxS��(�bjF*��A7�֩2�L��X��d��L��d��D�qƧsI��I�G��q� �bO�9SJ���>.��(`��D��rڔ�9#g�P���sv�9��[y֫���b�+�$�r�n%ټ�h^�7.� +1�����X�x��xۭ��ɞ��^�sI�g���$[�N�@�S��i.�(�FJ���9+甙y��8a��41OYs\�Ț�*d IX#!b����ʓC��a:��� �0�Cš��A\8�.�ڋ���tcvwbwCSӌ}�d���Vj�vaFX3�*@4M����ɭ�w��Z|���i ��mfR����f�{�H@M�=���i�f5�؍Q\0���41B�7���P�"��М*oJ�N�	��������4������ڥ��SCm������ݍ�=���M��Gg�Ϝ�_:�ou�jc�xc�`c6w�L�ŕ�sK՛{ή���YZZ|��׾��{�݇[�}����~s��{5�'KO�T�.Vo����(�X�^YN[YL_[��XM�=��<��:�:"y�x��@���ӑc���N�@_|���ٶg���ڞ�n���9�j�J��H\���ˌ*�V�P�#��Tkʁ�}��`��?~7k�^���ġ�1G���Ey&r�٘���mW�]׋�?�}n�������i��˒�O<����Zo]W�^��]{m�m�Eu�yM�Y}�Y����]͜�pB�?(�镤���	�J��L�=^n�T����hT��r�E�5	"��$�$�$z������*ZT'ړ$B�G�IV�MVCSS�绸�v�QX˵��]�&��X2C"�"�C�"v�����
م
����~d�����|� �FS�>������i��<�8��eQ�BE�!˹d�`,"�[��U��M�<;��AA4��\�!�{)��$@��� �׀'��d@*��
7���*u�J�bj�<�ʩ�q��s��'YK�4	�}��D۾\g&�_��q�������揃�S^Q��<�`�?�n%g���^F��X�dM`ԏP�ؖ5�Ԕ"+C#S��;��v�d��d1���/M��*a�h	�L�4�"R&8
S�����|�i ��|��W�(���+�2���UW��5��AxQ{6x	qG��3���+OʏBꏦ�ij�2�Ay{��1M٘e؛�I����YV�"15_����^�u���ҙ��W��ZZjr�#�^55ۋ���x�e��\7�$��{�p4�JPM�KݟȨO�4e
Z��-��Gf~$��)Bjz�8��]ͥ��,45qvD������em�"1/���/75�S�5�o�_#�`S�����&��Q�L�K�H��n�1=n��o�'[��fN���jf&[�qVQ�Um��,2�I���R������)��8�D�1��F�
�IxYE�-��6Ia���[R���kwK���U�UCҪ#Ҫa��Q͞qy^�*o@[8X<r���K92{��7/x��WOY*���c��	�m�ٽH�ev�<�]��"�? q����,��#rp�[�fJ��B'���G�ɓO���П���[H����!b�t�E�r9_.�J�t��iԋ\�Z&�y�n��j1�:y��?����?z���.߸tj�d}k}��
ObTdr�̬�Ӽ/�:/6;Γ�q'��N[̠��|S"�*�B��ˢ��P6�I�p)X6.��~��SN�Ox��,x��+�g<L����g��&���)�:B��Qa`�yO������Y�P�p�<�z�M�0��(0�i����c�u��Q����Z/��4h�䷸9MvdP��˷4��C��j�lu·�G��;z���x~�����om}���������N���P�bN�E��"�w������%�|p��/7�m�vw��綞��5�w�m��,y'�{M-��^Ҋ��C��ukUI9��^�Ѯ��:�o�ToE)�r?v>w�r�v
������m���"��,�������=��j����d�ߋY���~ɥ��K�9��%���Mͧ�'�Ț����)��yG�K� ��k�����"��ſ����AdV�����G�ij�c��{����`з�(���p�@�K�ܥ�ﰘ�y�[�1���M%��_�K.�śzњI4�g���&����So����MMo��/f��lOz��{jO�%!��MA ��AKn@������'[՟��ׁ=(wf��U-��(ܒ�h�Ⱦ'Kh��ep0�W��_�`_�&�KjS�R�����{ ��M�� ܭ>]ؐ)nΑ��:�4~��=m���P�;9(@@e �.��S�m�s�` {hj� �	Ԁ8�����7��XLM_}����������Ό�N��iX�cL��x�To��t˙�+��'�S3^�S3�4ۦfi0�x8u�P
`~ ��y#�8v��ǱC�L4A�wlg�9�����f���(S�h�$[z�-D�<���T��'@=�N8p-(l�55?��L͎���!�3�4��t�`��5#F�r��:^b�,�+���r�WEK7O�O�(G��a�`�*��&l�1=o�(8jNky�2�q���e�{��>��Ƃ�Q>����h���+vŊK��U���˱���r�i-ն�b]NB|`=Ѳ�d��d��h��켝�y:=�~��t��i�g�"�����tx:���h��=�S,�DsV�i뤁q�@;ef�22N���a5'��S
�	���t\���F�1v��$��0�'c�Ѐ�ã#�0}5t4�]�v�S��-8��4�Sj�i�0CM33���&@w�q]RB��خ!�iq-:\��j ��Im6
�t�8Mh�a#��|ld����P������iM�~�SS��9M֘"��L��'���J��=�sd_V߾�������C-}��z������<}�q�L����g*�g����.,�^^+��Zq}���f͕�{ΟϞ9V5�4��{/���/���}��������wG��̛Ϝ/\�-X[�?�ؙ�典���兤�Ŕ�3y�9KI�bg�%,�D���Z]��w�N�4���XJJ�)�(�ڡט5�B�D�j�f�Q���e��k�.M��o8��p�t�N��݌�{IGn�ލ:|�{���3�#/�[.;�����7����}��/���������+����C7�=�4��u=��ݗ��4-�t�g�����MV���c��C��NQr=P��9S���ݭ7��&�̈́h�(�(�ȋұ�ͼT'��N31SM��O&b�	15�ߛzy�ڸ/YR�d~�����2NV)�u�3��$3/J�u�F1M�!�8&Ǥ�a��Hv���]�a�v��A�����9k��5a���?d����#٣�|��o�G>P������bj3��=�~��	\��� ��( b1$,�M�
i���Q�|��O0�6!&R��W2��|�ȅ�Z*sQ�=d�PMM��y��<�5���ʃLM��R�������m�|;;��I��Ҍ��8sm���<qn�yn���\;buvhn���>�2�Y��0���'�ّ$59�}V�c�ƟB8`j�QB���iL�L���WG�*���H��&�S� �K5�H����銖%�7!_�������������&X��� P��@�15P�4P���5 j�������� �Ɵ�&��0kҭ�Ǻ�{��/�y��Wn=�������+S����dEi���\�4?�����qr��"/��Ǩ�
@��mSC�Kݗ� c����4eK�Jw��	��X�Ua�q��q7�:�d"15��x��k\��gQX42�D$�	 �H�L��� 8�P��LBc`%r�gjv��>�� S�`��A 8�JEG��/c5<�Y�p�XQ:N���l�X8�fv���|�Z��A�Mc��M�¡W��*�Z��;�z�P��%�-�"O�"�2���R/�m�v���>Ei���SQ>���T�������#����S��c�a��c�g^l_z=��\v�zz�bԞiO儫|�]1��C��.Ef�<�S�֦JmR��{J�4�,�#rpF6W�fKYL>��"H(�-G��X�G��	>Y&���R��*��2�Q)T�i:�C��R_JLU�ެ�ol���Ɵ��������{��f���#�ƛu%��W��b�zƗOd�9Ң���+�F9��g��b�To����U�TI��DȑrY<2�����	��E�������-�g3��.*MA�30򡩱ҶM���W[�{��i�9��n45#�ߛ�XA����@M��q��ku7F�Z}��(�ޥ�Qo#�f)[��y�u0R5�3�;����ે;�+�FR�ε����������s��h���=�,��l�-�j�=ϑω�b�35����m=sik����J�����|W-���2K.��*ƺ�����jh��y5�����K�[�����[���������M�3����f�o-�ߚx�y6
�j�������'�;��r�o$�_�X�0��Ѿ`Q>�>gR?󛚀��C}���� �{����¾��@_��L�
G��~)�Bhċ(�h��1�b���X�8�i,�{����`��p�[�-��v�ͺ+���o����*����A�i��3�7��E�p��<lb�[���H��`S�_�)���ŉ�j��=Yܚ�H�`��A
�75��ILXӝ���Q���������ܙl8Mښ%�!��)]�GИ�oH��Me��#��$�>�	`�N Z�2ŭ92d�R���D�U��(݄*�h��	4 ���������<F�|oj4�6,���A��HS�S��珩����s u�!�c�����C�S#ӣ�����91>��X����:=�8�Q�0R�:u0�������������ᜥ�m���o45���(|�?SiG(ͱ6o@�� ��f�>3����P�@�s�3.��(�CP	��9���j ��?�0`ʟ��o�:�	�ÉQS��-1ǚ|3���x�*(�(@3�`̟].��<� ��M��� �[�d����{$���Z����X� ˣ�-��}f��q`���0cU��Js��*�x�2Va�LVX-�MefR��I��8ňO:)�J'<��q�i�l�,�4��U�..����@�p�l|�#b���;*f�I���3&�Y5k�,{L���h۬ǰ�`YH0�M+ɖ�����+��+�����rb�+Hx�8�Ҵ�K ���&�Q��VE
����c��x�f8_*���b]uJ�؀Yo�ʟ�pN�(�L��q�pTF8���*��Z�1>a�6L�u��oݨ����C��q၉N�pa=��ݨ]����Ј����t�B�𡝄�Vb���@	k��4QC��O4�w�r�;��.!�[��W����=��Dn��Zm�vZ����ewE�;c�®QG��3Qܑ$�JUt�(���	���핞�'���-)�����dys��5E�/���q�Km���ƼȆ򔖺�=��m���j9y���}�NV�>Q6w�p�t��l��B����k�/�/;�Q�~.{�Ğ����|u��߼��߽�������g�\>�sb:qj,{�L��\��\��\��l��\��\�ʙ��	�3�Ǔ�Ϥ�/��.%Ο�;y<�䉄�G���Eww;���K5�Y�D���u*�F��<�B$��b�R�P��J�E��r{��JN���e^���=�\��3��w��O{G_t�<�h��<�|��omy��#��q潭����z�%Y���q����w��}����y��y�ܾin>go>�h�0�WMJsdY]�ԃ��R�9����.�١7���(uE�FA��c�&��)Fr���a$f�&B�ɵ��㷓\�"��ǩ��U�q�$kR����2d��i�}�
��tվTUU��"N\-�s����T;?���V)� &�'9�$��8�!����b(���>����0�����PԶ�A�*�
���.<�	��� @C�a1�8l�&0`�ǡ�z:�
EE�D��Cxv���;�� ��9��"v��B�ѻ#0! 4x��t(�Ç�	
G�� �aİPd]^t�����AH�H�J*J��yx� �#�8%�D�0Ӳl�<;��S��~���A�{)e2��M�L8��G���VG3��Y�^�$/I��� z���o!�G
K�D�JB���'��T�0�^ya����C���H.�թ͕�����E��e)�$3#Z�ʱ3+��y6"hH��#�F� h��\3&ςηb
�b'�s���m�a�O���#ABjb����,��8��x�B�C�dAC��1Mܔg<�����4>�1�hH����e��8�ȑBG�W���h`(t^���h������x:�d��LIW�!Sґ)mɔ5���(*�eyQ�����o�r���{��{���\9{��ک�G��S�c��6q�MP�zx%��2��M�)h �ۀ�3{�`t�`ޘ!�g�yA9�� x��Y��Sn��c면5k�4���$�*ri�C�$q(D�@'�)"�/h�F�m?̶���65P�<�A��wl\ ?��J��	��#��d,��E1��\2J�Ī�D���TQ�ZJ���la����fF���ia�XX�VN�������V�]+1����a��9���D�%E����ʌ	5��}�����vMa���W[�o,{p��;�|:�e�W�R5f�u8�;��7i+����  ��IDAT9���L^�d`����w��-�H>0_3��w2�f2�j�W6�):�-p�[��m�}�e�c�9�e�|�6IjH��<��#P�2:G��R1$�B�k�
�Y�u#]�H�$#E]�+�L�$�2#+J�t6�������=(u7<�������ۭ����⹷޸���s�.��o:: ~@���tz�c�T����Ku�#-'��.?n�ٸ�S���M7&DI&�Q#3��Z%_"`�,"I@��x&\N�hIa:�vƮ6U��ґr-�|;򭋬�g!�Y)Vj��V�`ԸX�<��^�(�w&����h^C�p�KI����X��>���9���]���n~@K$��A��1'��ċ{=���|��NC�+3�L��l�<k���^=vx�����¥��/�f�䗓�ϖ宨�B�-�b����}[.� %nk�w�����C[ӝi�z?J��N������Ix��=��,�p�*ʢ���$-)��jƦ�{�*�g��`�f�e��o�}�P|j�}a�|i�����U��]�G��;3�OF���?�x�(�hR�N#�F���K��C����Z�F0��ѿ�P?c�>�?$��'b?"�?&�?�a�Ǡ߉34썐�Ww�<�6x�[8����7±/�P/��_{�4�y³�Kd�D³�3���=�
�>��4�y�ż�n8�%�[J�M�dS�;�n������|�.���Zx�̌^�����k����e�{$����@�-�ז��'�:���)��T! Դ>��d^s 
�)��tQw��'[���'�;�À����2%�V�=��t.�2@����#i�6��A�>�S����W!����!l���K@/ ���\)v�2<�F�Xy�Gz��1 8%��@���C��W����vv�!���.��=��� /*a�
��P��Kt}��CU6��j����~��q �~�C�|����� D:��������>�p�!g���ء�ӣ�sン�#���� `g �����驝F&��#����3��]�#�3ݕK#W��V&k�'����-��,�U-��/��.��G
�F򖆲����2��d.N�,J]H,�#F�q�4�O	D�@S��� ��afZ�G[=��f;���45P�dt X8�}��{�5�xs�LC�TP�@@�� ����x	8lj�!45ǚ�w�'x����	Z����k�!h�p4��*8�(��7S��\�T�n<U=���S��)�c��1ʣњ�HՌG=�RN��FᐚwH��R{x����j�a���	�hJ#�)�땀S&ݢӺ�u�F١�YL4!a5)����K���Y�7s|wrc�-Hx�8�������!oVd�U��v5��<奢�gs}Ogy�ˋ��d]s��L�y�`�&,X�sʜ����-}V͘W�Լw�C���w����s/�)O��:���"D�}6�����`vY��BZ	a-�p�iZ�a���fZ(������΋�a:���_M�3P[��F+��A49hpM��HN��t'�;ɲ�T%�`��p7%��r� �)ʃ��$Es��9A�+k��w���Ɇ�}e�koyʾ������ޖ���G�N��{�bjfO-�)X[��X�X�/��Yr�\������ܣg��������?�O�pk���x�{��f����V3V�RW�W���b�fc����	�G�'-�N]YL^Z�;}:�ر������ј�Ñ��Zmi�*;͜�mj�Z�V"R��*�T�WJE�\������u&e��Tt�u�f>�=|-c�N�ؽ�������O;����lz��n���ѷ��_�����}w���Ҏ��lXR\1u]4u]��oX���:��[ϛ7l��+�=g�c��IZ3?����e�z��hי���i�{���1r�L@���f�gр,&ی�Xp��X��4��5��X�8����$�S#���ojd�Uu������$yU��8R�ie�;�	^���S-b��OR�
:��ǰ�z8����ȡ�.,�	>�� `�#С(HD�£"�#p�ᄐp��0\h�Ba�a��@��y��	G�Y�톄���D֠v��w���������`v�q���,!G
�R"�4��@E�0\<F@Ĉ)x)��c5�#e��"�WB�ɉ�jJ���cg�:Xy.�t��?f��o�2���/U>z�; � ��  �\lj*nzU$��J)�򊼂81IϬIw�U��w�\^;{f����啙��э��#�㽵���d��"e)j��V�de��35�����ɳ� �45MP˂�R�������e�qj㹀��>����U���8���k��<R��MG�����hp��O[[T�#-�ʚ^�lg~��iK7�!Y{�t5)�,7o�}a���w�}�٫����w6���v��򙱞�ũyѦ4�8�.,�J�=�/�<�]�<�� ��=1�}��?�*jL�4e��8��N��l8چ������D�W����W�ۊ��24E���$ނ���!a�y�D��T<���=�H����L�"�� @��08,�
G�Z�� ��%2�d�%�c�\�ALr()�:j���h��Z�if*�gM�l3=��ʲ�͌D;/�.��H=z�C�uN[�ݖ`���fo�#�*2�66��W�����Z
��Vt�]>��4��x&�e�����7�Xw"��xT��%���-:���7�7�*�Z(l=��g4m�xJ�H|�ᨂOngdNgt~Olɀ+��+�.�%�Y2��8�6V(s"�F�刕t����Rx\�D�2�����%���2�
wGS��`��`��p��p��D��Ԟ�5���gg�槪f'�NOTi�;~��������ֻ��ŵ�_���g_|n��F���s��7��}y�����3�+�G�^l^��9:^99��՚�ٜ�p yoejuEvuEzYqlz��zX�R��,��ǰ��v.&Z�OP`RԸL1�J�s �؈H̠�Ta#W�)�NZ�����:ŁS���.�W�o�G&kÿ05&�p�hjc�&��4G1[���Q���@4���鱳�x��/��|3;�ŉ��}c�K{�>Z����٭wn����'���Ҿ�nn����Dr�żA���˿\#ῌq}[���}����~���ĥ�@�yMAU�z��{ZϺ��]�R��9qNN����T��Y|�"yަxզzîzץ}ߩ�����*��$��"��&�/%�����w���?ٕ��4�7*~�}%�|!f�L��F�����������3>�K6�s&��c*���P��p���b�o�>��`ښ���wЄwPķ#oF�^EE��	��"6�,��
��"����,q4��h�3ϲ�����\�m�&�}C̽!\W���%�uB$��*]wʗ��Y����?a��ژ�.v����Do����Y�t$
���t�~��Ak
�%�MM{�|��3�<����qz4г�>vv;ć�@	:ʃɜ�$6�7�p�a��ؓ^�"x����-B��>"`U�a��y��x�?zLe������/�_�� �n
�I���{ga�@�����_a��ʚ�=��}n�f�e͑�7bj��L���1�{c�kb��&��g��Wh�����;96lg�y��=16�H���?�O��\�h?�_�4ְ4z`%`j~S�8R�8R�8��8��8��OO��4��45�a55�x�a����V�æ��d�/ �y��	T�?�_�����֘���G���&��4�q��؃T5�f�!�X�Nw�m@Vo����o	����w������(k ��&8�f�c����p4&��&�A��	0Yn���Ofi'2uc��T�D�z:E7����U�L2��7Ly�n�	���[5���i-j��Z��Vcw�RP�<j�zH�����)�dZ)>��/ڍgc\�qfhjV�-�i���+ّ�s|O%<[��bI�+ei�Ud�Q��fY��ՙ�w�2�(Ky�0��쨧3<w�\W�L.ŲU�b��9d`�h�-�YKƲ��b�X�+�I�f��J9S,�)l�r��k �o��?"������¹N���^LH	������75�8�� ډ�m��vrX%���Fke�"lkT�۩�u��:b���l"7�i�n&��� �6/�������J� ���])�N���aj ;َ�IS4�(��I��xiS��1FT-���TGI
<�$cEQL��̦��}3�]Ǉ���15�󧋗g��Ϯ�/_<���V��^�v.��B����󯭼�ɕ�}}���<���ի�1�C	Ǧ�/l��̥l����Ud� ~y.q�T��I@�♤Ź��Y������{h�sh����jk5ا*-Rd����^�¡S۵2�T���b�L�UIj�I�3jL&��n���eħU����[���v�J�����Q#������+Z�#���oG��{�/o�e杭���M=���i]ٸ�븨m�����m빁���s���%��}�	e�iz� n/�U�0%��b�Gm��L�E�1�|fQ��of'�YIv���a�g�0��&׊:���J<��(fU灦�I�MASS�)��P��9��;�m8���OSW����l�$�.�1p�*�]F3�Z.A�$��8�����"Cf�)�p"1CAc�h4��GD��Q��Oa��LPXBh&4yTCBn0(<C�c�y�¢A�1h�*',d[���5��GO!�&��fw*����bw�1O��Q�04�gb�,�G��81/�L��M�qH&�.��%�H9FI���R���v�E!�gU�p���*��kd�Ĳ �: n<p4��)�1J� ����^z���(V��Z���y	r���7��W�7ճ������ع����х��fGNLt���o�H�L��%�r��4#9�L�6㋝H���M(�a���UDR�;?���'pa.CP ����<�i&	�����%�B�8�M��2X���e���!��;5�jn��&0D�a+�?x�G �
#�恦�w�ߡAVIk�i�.�Lٓi��x��_��_���'����՗����K3�K�s��Q�CP%)���=��(v�	\z$��?���%��M��,IK��8>�B`�4�����Já=ցWG��6[_'����-���1�,2�F����?��ω�����v@�FAG�p��N�K	 ��h��B�Q	B:V�!�D$����Ң��83=�JO�PS-�t5ӂ����&�̈��,�x�$ڬ�t.��nt[��k�ّf��Z����5����]�e}1U���C������Ȳ�q{F���2�g5��l<�V4��1PH����3�-�TĔ��ݙ�����������?�P���m�&���*��e�jwJ]TV�=��L�w��5E��	be�L)��P�H�����
�ݪs����s[�r���zrO�쿼Y�j��k�/��=߲�޴�ڴ��ty���zÅ���K+g��V^{�í��lk�_�z�޽�����gn_�z��y���swF��nY]��<7|�f���m�V �s'�N�?>�xl���Lc��:��&%��$$zl6�J�P	]
V����g$�q�:\���k%���l�2v�vr��\��q��z�P������i�4M[��y��dadMSBc4��Ch�Vg�-�����x�|�>'��Ho�Pg��O�����''���-hq�OT�o�rm�㧷޾����ׇ��h����&\���
�0��ɸwt�ob�[e9[5��M�|a�~�㼧a��g��g?����1�R�� ��I��
ʺ�q^Ϲb�߷�_�*_u��r��u)ߵ�޵��3�>�	���)��]�+�F�/��_��9�t��hW��,��N�s�?�Rq���B����������9���S:�h����1����!	Y�=<�\��!�kp�W���(��D�$�s$�+,��,�KL�,�l��\�|���}!���GĻ%�ݐ�o(�7����%�t�*[��V����Mx��3���n�7������cE ����+n��x~w
A�����Mw��a��D��4a[*�k��5��l��t� }�#��M< �߁r�s}P�G���jJ�7�p���!���ᫀ7M_���X�W��;@� �������^�#�� �I���2�Y`{x!8�m~���o�
�x��xm�;�R��w��SH�
�3����V8
Bke�	���aj�cjjb�����f��h8=�;?1<?96;5�fv�ؘ��4������C�]+�]g��7-�[yLLM O��P�� bj�����bj�7�V% k��;<�u��Yl�P��j�\�MM�Y�;�Z�kZ�aL45�N�\� ��h�9�n� p[Py�=�x3�Z��{�npAM
;M���	Ț`e�C֌��4F�Xf��:��zސ�	P��&��f��8��GdM�q2�0�c<�m<�e>�e9�b�ͶO4�	��S	�Sq�!��d�g:�u:�w"�{آ���z�L;��/d�)�S*ɸ�?.��*V\�y�~.N��`\I��Ks\��\ˎ���{�4�Œ��KSSS��ԼQ��Vy�[io�#Ӡ^.�.�w/�};�q5�tѧ;�V�;�.`�![�
ל�U�%:�_�j.z��Ƌ�\t��&c�B�v&�$>5H�݋z��{ 
@�cB��'(k:0��,�LM'!���A
�$�wR#:��LT;+���)@wIp]J|��Х!v�H=Fr��S����#��#�I#$Iz����ҞB��#1`��:���(h:@3H��=Sߚ�mMQ�$�[dm��du[��@��<ZY�n�)M�_��y�v�����ɶSG�:����=���Δ��m,�[-8���\��j��j�ʹ��K�sk�7��C��5���gy�`�L�ә���+�Ik���K	�K�+��KK�ĥ���3I��f��9y�3}�56m?2�84��;����jkUe���Sz��mU�Z�^��+5R�V�Q"1�6�ڮ�Z�z��d5��6�͓�-nMk�-��9x1���䑻1����W�CϨZ6#������ț[�o�u��V��_��z��y	��u\�u\A�Ρ��ޛ��+��u��9m�)c�	uɸ,�G�x��-f��Z���U[�f��"m��<_%X8Iv���fa�[hYf�G�g# �����ǫ���K�K�M�O��f�j3刬�O���PCSS�����j�T%��<�<�%�7�L��n�R�B��CR1IRYD"���%�YX
�g���ǒ�X"��@Bl�a��T8:"�	E�@v����Ec��iП�ŀs.@��s(��z��&4<�!ӣ��w!��F�@�FE���1���S(�S�����4G�HQD&H�9��d�u\��O7	(v�-%D))qjDӀg�t3+��.���Ǌ*c��<D�<��d�}MMe"h����y`j<��(N��^�`滸)z���?�=�R6ճ��������顕�g�{�.�/;4�\Q��ʋ�T$�"��R��T�BV���h P���\3�g�����5P��4(#ӝr4��� �?��udoj��5xl
� 8�ׂ2<��1(}� l�?B`l�W��d#it ]�r �W�l	�Ve�%Zr���u>5�2������G�ç_���/\}���7�_]?9�V���Ѧ���Na�OZ��CSS�D��/4էa@Ms&��jk�d�_D�	���ȵ�L�_i8\c;���[�:�g*�W��Dqf!45R�OEL�@��H;Ϳ�SL�����&M��pxP��#\x8��ƀYĠ!I��5�h��\j����33-�+-�J�kZ��ȳ�s��+��I0r⌂X�ܫS�T�L�U�uZ�V����t�
s�ɛk����T��\�-�®ĊC�e�)�GJZO�7���M�����=C�l\q�+�đU�29w���+o�ͪ��m�Ĕ�\yb}2Wi���=G��ո���\�#C���(�R�K�t�Z�P+��yb9�+�r�"��eOL�+.�no��Mȟ?]{���۷�^�t��f��ٺՍ����g믞k��������+�+��_|�?��㭭W�S������[_~9~�恹�˽w��߻��f�����s�ׯ�]:�z�\Ǖ-�7���mK�}�+G�V�͵ML���W��W�NKK�:,n�����h�Ff���ӲM�<%ߎ$�B����H@M����j���8�	��C��dIs���&��i�Gh����Z���v��Z��6�P�`$A>-�s�,�c�,鳓��ru�呶��5R{w������|�wϮ�<��RǞ�9q�j�e���Dx�E�Ǡ=Ϣ�-~��k��gF��z�WZ�gZ�:Ϋ
�=	ᶂt��>/í�pk2�����U�7u���-������U����m��-��m��3��K����_y����?���6��1q~k�|�P�ѩ�ߚ%��	~���B�����5_��_	�_
(_�ɟ��۰ȀO�4?����h��Ȥw���	�7q�7��7��7h����"�_f�_b_��_�3_�^r^q_��/��ʅ��Dwe�[r�-��F|�(�j�_�+7
0x^rH��E',�ig���wqz�ܾ(~�O�+�C��D�^?���}鲞t1 1~_M�|��1�5�15�������ї�������3PʀCXeM@ӀJ�����.��PM�5� ��]8�������!G�+����q�%;�Hp���~�� x��_�o^��� @8�����@��hj`ښ������=���ytLM{UL�������}g���'����&�Q15'�G�Abj�z֎���[�����aL��� ���`4��`:�Ss���OP���eͶy�@�l��n�a�U˿gjN�0^�oӂ��ۙ`�f���kO�ŝ�H8�����s]I���d?I���7 
�fv�4���ɚ��Ԍ���d�NG�ӝ��)3�K�%��B�x�a��8Uh�)� ���N�َg[O��'��V�[���=_�8����ѷ��>:1�����^�i�[[}2���g�YCr��Z:-��Y�B�q���[u*J5�]J4m��.���dz�fE>S��La³	�$����R~"���W
�_Ώ{)/��l��������8��H�G}΅,2��3�T��e+6њS���9$��+1�[	�[	�[��u�~V.�������AB�B�!�S��O�E<鏬������<Յ~Ѝy��TnWa7���!�w�»(a��.&�����;�n9�GE��S��.#��L�R�\�i:��]>^G�+ �\o� Mo��/Mћ���Pv�e�j*0�	8��tUW�Н�����曻s�]���t8՛���2��ZZ2LҌ�y�ʄ�Y�}��O��Ov͝h���_�ݷx�zy�lm���r����͍�s��+K�+�y+ٳ���.\o�~�fm=�ĉ�c����.l�]O\�MY]NZ[N\Y$,�&.� ��fgS�g���cO�{��r�u�NۏL8����~GG��`���\��cJMR��j�Ig7��J�Vj�ˌZ�M/u�N��i�8Z�Ak3�f�>�$��p鑵��͔�̈́C�boxnD��m=5t���χ^ߚxkk��?����;�͘}��{C�vI�u��s��w�u螭熵���nIUuBY6�)E	��D��#���q�.��e�9�V�Ǭ���m�/��N�0Ҭ�t-�LͶv8�|;R� ��8�	���I��>�f�����_�(�25�Y��-�5��F+���$� ���Բ�*�]J7�i>]å)Yt�.g2�4��L�(���%�D<�%aQD��
UKXX�+!!�
�Ȭx��> x�,6��؜0DӠ��d��k$���F����P~w8aw(%��b���N�R^�X�l��B�UDvKH>91NMM�ђ�T##���u ��2151��hd�S��	��hOڈ׈�@_8U�d')�ˣ���(FU$��OU$���(�3�;��ٓ��:�_wcm������Ë'���~����pw͞���x}M��<V�n��X�>N���H15?�A4M���ԧG�Ps 4���`�  �5���cV8~@����7a�@xF�<<P��8��������ojh�lIW��[2e5���tuM��#�Hվ~oqk�˭?��O_}�����{�ޅs����Ҝ�d3/�-.��Er�<t��,
f/zP�����ԧ�,Ik��<���a�æfp�����Th-�W�8���C�Ff?�)<�E$Qp"���� v���_lj��ܐ ����M��"�� *���`���J�eHx%�����P��T;-�Nϴѳ�l3��ʷss�|� ��N2�b�,��m�p�\���3%b�Z�7py���EJ�Ҙ 1���y��Bsl�7}\^cn����ٽ�
I,l��8�J��%T�K���CU`�9�{G'VKkz�Q�rm�B��ɳЙ��f��\+�g�l�C(���6��"�e�\l�e<��Ǔ19B"��c0�J�����S�^W��ՙ��9؟1��ʥ��9�˅�+勫�+�U�kg�KϯJV�*W��N�[Z8��/��/lm����_x�Ɨ__���7n��<�_>�|�j��u�j/\��t���y@���7k7V�WW�[W��WV��[O�j��i�)��LN����zm���hf��)�fR��T`���09z��\�@4M�ԧ@4��XA ��U�#Mђ"�4'o��on��Zb�B~8�������#Im�¡hE��ߨalTe���韯L��/Iu�'W����7�>���ܡ���ۗ��R���+|�u�>�u�L|�B�J*��J�%����5�gZ�Z��R�=n�-ꮒ|]I��$]P�6���E㲁u�Ⱦ�f^Ӳo��-�l�����7킏���}���(����}��ׇ�
�)Q.ٷN�o��oܯu�o ���̯��dԯ$�/Ť/�������D�'�S��6�}�=&�]:�m*�-
�M2�u2�m�-.�?���ɯ��/(��X��8�+��)��(^R�^P
�V�(�Hn���Av͢��P]�hλUk.��]|�*8j�M�9�V�a/�/�����Fo��C���I��x1 �}�;1��?Cڗ)�͐�� ��Ag��;K�d{Y���͑?��4͏�hv�5��� }_�� ` *�=#(4M��B�uaX2_��=�Y?;:�@9X� �c����e<�����������J����ǙSs��	3
�����S�Rݽ?�Hs�t_����xL�NS�>7�t��X��ڵ��������g?����l˚���i�!��aY�#�&�ZvP3;�qy�`��5ղ�ԀC<�6@�j�:��;�_�	����L�s� &�9��j���䅞���T ( ��� �Ȅ� &�A7G\����o�!hۙ ����aj�KC%��"�H�a��8^l�*6O�ئ��36�t�u2�4�>쓟�v�l�{����u[������k���|��֝+���֡�#fu�BpHR��*�c��|�G�6�����l�v%�t6�v!�y9�u#3�z��F��f��v��^Z���Q�d��I�|:�}/�u'�q3�z-�t%�p٧� :��|�&]�J��%�`�"�p���9����H~6=�f\�9�y���â�Q!��ჸ���'��k�Ї�݋�Ճ�Ջ�ݍ��C�Rh/9��F�0P=lL/�-�v�q�ZZ���get��6j����wzYP��Y�]�H���xQ_��?U�KS �ӕ���L��LW@w���5P��di{�u}9��\��B[��?�ܛc����\�@��-�T�n��s֖��V$�����<�:۹�Ժ�P�<�we�jm�lc���J���쵥쵕����������sek6/�te����,6�/�]���8������������������
H�_M85�<��:��4�{r�3s�9~�5z�14�<2�v�8::��Q�嘓�N��j1��z�Z���Lr�^�0�]��(����mR;M�ɢr%{
:�W���<��{.��R쑛1Gn����������W�2��_F^�����5��]��{ƞ��ˆ�ց{��{��;��+��M��9E���hX�? Lk�D�][���49��f��ic��$�8��ϰq2��L-�Bd���V�����A
H'\ͮ������&��lO}�˒�g+��@��>K����D��$���fn����s��[ɶI�f��ghyl-<�p,��N��hbU� C_�"�,��ţ�p�lD8��12a(\8�#bd	B��!��ƃ�p&�E�BШL�@���	ń�a#G�C��%G�(�p
��c�d��AUs�rQ�$j�D�d�lb�CJsʨ>9^KM2��j/H&Q;+�Ł��2�W���W����ʚp*|��hd_�cUG1{ ��J/���D�rqs��T�"�<�Y=;�z�챍�C�_^>~x��Э���7N���Ƣ�������xU���-�►�n��;Ɂ�5��&ߊ��5x��g���(k$|?�)�h��P�&8��Y�		c��H8�(_�!& 1�x^8�G���!� _����d%)@w����5G��-��Ww�����'�kRԑJLi���[�[���15��?{s����Ξ�+N�I�L�<��"VQ��65�ؙ`���75ib(kZsd�Z���aj�Kս�C{���#�j.�����(Ǧdj�41�ģ��"	��Gl҇��a��bj��yx���A�i����B�;Q0(*MǢ�x,�J��i*>S���xx���V�|d�S����Z�t@���sr
��B'P��8�)f��ddc�d� �ac�t��eЉ|:YĠ�Y�@h��RM�L͓9�b�De�df7t�8�<�[��/28R��8���Z�<#K`�
�<���s��y����͚(��Tr�X`�24�]�hj>]�&+D1��gR���KX2O�e
�IaӨl
��%�0:C$���]��}�CGR���Gҗ�
/_�:{.{u�`mt��篔o^,<w6kc9se!oe�xi�hv�jye�7^��zgk���Yz���Ͽ^�����w�K����?Ww������<p�ڞK��/^ �\������Kk�o�ml\[oY]k[^m�_j?=�{�D���悪¬���8c�C�����YVz��Vh��)%�m����׸��i �ek��5U@|\Y9Q�/ �՝�t'~:c=q��XNO�7���b�Z���`�d<A[ŏ���_l��������*����ƅ�?�q�����{w��f�gBLY3��E�%�Y��y�ߪ�՚��T�R��F�������<}�qW�}ZM�����R��hW �U#p^I���_TӮj7�̧M�����w��}�Oc���*>�I?�)��+�����C�k���N�/l¯ͼ��z��:�ϵ��5̟)�_)h_ʩ��)�JIKɐOd�Od4)�=>�=>�]�]�.��m6�-�=	�]	�)����������������5��e��E�9%�i%�RpS%��]׈���,�k``��^�Ԟ���\��v�1+��rG�#Q�~��N}:/9�$;���O� zz���J��eȡ���&�G ��@S5�Sӗ�x$�Y�=Ȏ^�a`��0�Z��F&0_�K=i��.�W�B�/Af��� ���(@=h��1��эdy���㝳԰���E�F133[l[�eɒ-�̘f'����N��Nc:������q�ahg�����ֻ��R��쪞ٝ��N�7n��i߈/�wQ���U����>ߚ�����ru_�&T��IjPS؅�󞠩��15gJ.v6�v.�,��橉���v���������}ug6'��65ߌ�	eF~Z�[�iu0 ����D�h^"�

�f"�3�D��5aY�#�C���cS� (k������v6�-�$��_f�q/���Ml'ΜN���v����R�g�5��D� .
d���>��	�4�nAM��e~RL�X��`�"s	���j��"e�b�H5R�-ь�j�K�cEڱ|�h�f<O?�!��H�rW�2�8���_.������ѝ�>|���|�������_���og�V�����C0.J9�\r)��xlHF���8�v�S���n��w܆�n'E{ա�uhn8��R�w\	�ӌ�	��]�{��;N�47�������yWt\���Kj漒���r�^������n~����\�s"QgLL��C=��{����Yh��3=1��ŽЋ9��BW����;1/t`_�����$�" ���|��z���Ɏ��Ŷ	�����j���n��X�-�vRK2�B"����H�t�r��^0¡���/t�=AYw��'[ޚ)AuضfJ�x�	w4�9�\Mo���@�S��]`���v媻����U{��_��S4�����������ƁɎ�˽��m�+g7�7����˶��wVs7V��+9ۛ�;;�+W ���h�:xjlz��3o�^��˥w�ݹ�{�v����{c�}e+}m'}u;}y�[�J�]�,�f�lx��S.�ڧ-�s��Y���Z���'uC���X�=���R���F�S�,z�Eõ�X �����%%�����9A�2;��|oe{M�����Y�;�O�]��#Å]������y���������<���G��[�T�r�jW��������e��;��׵'�T'�%#��.q�9Vj9���;e	6��j4Y,	�D�<� N7�2����
^�����b����8T� �mD$m��$5�nN}:���G�>AS�Ț���/i
*N�O�h��*HM�����w����ݹ�4=;E�v��V	�$��T-����5\��E��)RID'
i>�%a�$$���������4�0�x,6:�%���x (�]P	�DŁ��أ�1G���:t,�pY󵩉>z,���cGc��u}�(��1ZL43>�G�a�,���Ѱp!G�7	V1�.�$ˈ51CKu�	!�L+�1K�X�)��NU
�*�Q�J�Ie@�5 B�T;�XX��i�f�9�L���35��J��&��,��=ZZa�r�|��l��w�V����l-��t{����+�F�t�g5�ً��F��\d=X� `d�	�`8��75`[�/�0"<_Ot��攗75��9��I}���v�%|��ϵ���Pe�����K�p@'� ��saoO�9���	��ǚ&[О- �B{���ͩK55.5� U�`{����������o��������:������y�.QQ��F(K&�%#�K�]���&/������Lιl$U͙ v�njڊ����*�@}"x�<[d,L��T���eL�����I�q�ǣ��X��	'B�@����65�
�}}�h�x�?~{�(����"r��X1���U�x=c�*J���5R|&�ψ϶Rr��\5�N˷2
l�"+����7ѳ(9��8*�}�~�'���9F<�;�;�#�P�X6���\2UD�I18nT=ˡ1�cZ~a}0�ʖ�)�[��@O��p>˦Q�F}�L���i�>]Vp"Ֆn�&��	R��K�3�l�`�1)QT�1Ca��L�K`��<!�����1l������b��D
��e(����wuM�����+�Y�n�����Ƚz���ݒ�w���ʽ~#sw;ck#o{�`}+{a�xmk��^��7��j��y��_L���w>j{鍚k�K6vʮ^�����΃�G/W�{Xr�v��[%7n�^-�q��Ƶ���j�^mعڼu�y}�i�J���陉s�j��5��W�3w�8#��i�M�<#��@(N���e	 ������d8��Ot>C A|\Pك,�|�����ڜ�v�3�Ֆȸ`"_0Q;m�a����yJEv�_i�����Ϧ;���/��j�7|t��/W�?��J}pZÚda.�b��Dy�B�-��G&�o��?�ȿ��(�����;9��-v�k��7��Wd�帇J�}%ដp[���"�P�we�m1vK�#��!��W�_�Rޱrn�}�|�~���<�����+�/-�?Z9c�����G3��F�_�Xcf���@������AE����;	�%�7J2ʯ���B�BRʗ"*�bڗ�2��r�r*���
��J��Z·Z�:�{��J�kr��b�}���ySʾ)��R�n�wL�{v��d��dņ]�d��S	�	��5je8���E����tрO�� `$x;��2P �@v�� �H|�;(D+���#�4�����3��(�o	: �2>��Ƹo�)a�p?�8�p�@�At ��<�����cj�Bbj-�]h1��8�.k"�C?�G�o��nS�l{����ځ*( ��j(k���Q.��8=ʟ�S3x�t��iv�ma�~d�)��bj"3
�ܼ�=?�9�q��fs���ԩ'���J��`�_*����W.?�Ԡ
�[=Nx{������@S���6P@c2ل��_`�(?��@PSZ^:�$��9����8*dp�)W������뢷��S�~;0��50��)15��&�ĉ�YN�AM�����@�D֔�A�X�v�D7R����F]���rEҝ��7Fj?�9����o��|~w���|����W���O��ꭇ�N�ߩ-���γ	�¸�1�#���[	Gz��niHϼh�'�VST멚�T�Z�|�&[�J�X�V�v�rס����s%�K��M�BM����������a��oE˞S0.Ii�Z�5���,�;E��Vs��`pQ�l��?�pg���G�?��ǟ�~�;��������ƼЉy�{�"�h:HG:�G�IGM��VL'7�]�"��M�����6Z���t�N<�L�ञO��;ٝ��.N�CP�8�j��,yO��'K	�Lg��0�&B���������<}W��;OMMGP��]���>IC@]��p"�|�6s��nl�u���ȵ�ޝ��������'6*�����ז
w6��d,�d,���\+�z��ƭ־�R�ÇU/�\��kzw�"�15;�k;ޕm�Җoi'ci+uf1}~-ceԤ\�b�ZL�XH��3���{F,�}��N㙳����<q���v�&�^�`��5R�Zh׉��M�LT�UT�����sY��d��hMT�R��ʺ���/�-���o����=0��8���\�u��m������>s�w���}�#����ME�}S����M�T����5M���h@��"ɬg%�4�<u�Ɛ`����&�I�ԋ�;^��4R�	���J�Y:$�0\��@MSh��'S�P�:��'h����}<hj�����t��l��l��d�М����K���d45��7��n��I�qD��	Z�������I�3	R^Bǉi8d=o
�q�8�k�x�����ɸ�-*�����! ��y���z!:(D!5Gb�"9����1��M}�p�0-�+>�O@4��Aа�:A��'��&�&"&II)
�KEMSS2u䠑�cA^� �vFY2q4���T6���ƪw�!�E*4�J�lPMߺA�'�ԔZH�Vj^	y'L���yIҡ��w���}p�����Ů͹���1��l]z����dKWCvm��cff�&J������k`| ?!.�������V�n�iN�x�n��	-����v�����чK�|	�t���a���et}2� � eh΂WA/���>�&GҖ#t�H HH|�![�䢵�+�}���|�/����ߙo��߿������o?�����v��G��}m�9iz�[^�y�.qI"bj��r)�΄����CY�15g���jj�3�LMk���D�S��K�s�+6�S4��� ��b<G���A�W)BР����_+�fO�|�Inu<6�k���M�;vs�)�(�#�
��bV�"��kb�$���a�,����r)��Dj>�a�Y�;�m �D�$�@y�{���|���O量Ҏ��`�����$\9�0��Ϣ����8���a2�P<C�K�:��ǖQI\6C,�)�,)�*`���c��S+��_�-�xs��)i	�D�bH��tF�M��PXQ$�,�XK�H|��SX"<��#����������82����eJk^~ک�y�#��)��H��\��{��g��o}7�q=�y#k�F`���ƍ��7rwo�C�Wr��z����?}u�}5��_������o������j��J��������*��R���Wo�]��{�Fp�j��n��V��V��N���ꍝ��+�sK�K�;k���Z��J�*��AkZ��g�fZ�Y&�\����-ν���h�l�M���	BSs>$k.��dMp����俲����$ZO�?]���w&s����fƴ�pJE�#=s)h��t�o�>;7���Ӻ��wO��b���~�Rvť����S�{����CϼN��|Ac��B�5��������N'����� ����eY#��Q�n��w��]eC�Y�F�r���w���J�KF���;I���������&������C��$��l�����`��M��6���{#�	�������@����������+��r�
�
�/T�_�ؿRs~���R��\��L��I����u�t�x�x�%����^S�^T�7��k���yU����^3oZe��U�]��d�Z�d�ʿhD�|72�-��Dn�����n2���+̐v�]^������5����=�V�h�yO0��;W.h���15Ow�ۄ���C�tP��&�4 ���U`\:<OMw�05p��������5І@S�(�+��������}��j= �K����W醠�汸�=)��턫�10t��bg��@��p����塧ɚ�Sij��.̏�,��[9�8P�SsPL��h��X��hΕ��6�����Z�P� @y�?s���4�]�R�;B�,u� �&ܪ������T�D ��H��h­�5 �����)P�DX���5�����K���O�J@_��^hq͇��� W�[��hdЛ��_�^�=2�	�����k����z�T��b�0�dG����N��4Z�h pTxd�^�ǔ�a��"M�@�j�ظP�z�w�%�����p�ߺ������ݯ����㗟������~�ҫ-��)�GB��	FD�>f쐈�##�j��F�E�h�!�w���$٢]�dCX���;����i��n�{ ���0s+Us5Q�e�����eͫ�rʤ�0ĉ�G��IƷ*
~y��7��}ϋ��7R��F�#���������}�5�]����u���Ң��c�n��q@/=���c�q���VL+���-����}zJ���a&��ɭI��j��v!���f�� ����Ņ��ab�������Q z��,D�t�����J�7�鱠[PF�j�Yӓ�����䪻s]���\eK��B�
���d*+34������C����L�m͍�,�,u�,�ۘ�[�)_���Z.�X.X[����\����.��-�v���ݦ�_?�����yɣG���66�֑��|�rշ��[���oy�x���=k)3���@��eS߄m`��=��ٛ���l�`��Ք�r���l�4Z�\�U\����"y�ZZ�����p�Y�VN���NT$Z���i����ʳ5]s'�nV���w�zz�'w^O黛s���N��m�k�0��W�n�}$:�+;[���E͙ۚ�7Lg������sbo� ��m�p�V�^oԫ�F�ìt[�^��ob?�4��3V�I+����81�%�ij���鼦as���5gK"d�0��L��l��t��~*w���9��l;7`�f���ƽ�����b$)�69�,�E�!�  �D����4��OVq)JYΥ�8d!��!c�8>�F�gRp\*��' �"���S1XR,��H���GE�G�w��#G��=t8��ј�E?����!���;|4 �	1Q��hR\4K���p�t\,��s��8��RJ����s�	|"��(!:ACNUS@�4��M�|�0�V��(M
�H=���Mi�F7���BA���A��U�@�Br<��k��P�H)��}�t%&�����.�徦��ξ}o���ĭ���ۗ\_���{?����w��^�k8[�,q�:B@�-O������O��y�؂�X�S�И �� {�Z(O�5��� 7���%�����7��&Z�5� �[$�[���Q��	��ǚ&Gؑ#�ݞ�8�׸�)|��Z����;��/_�ۿ����x�����|i���;���RIL�HC$��T�bZ1�)O45��{#��&�,�t ����>�G��YO����8��lL�(2M4��e�uB��E�	�7�,�v,Y�8 �x��8]66Y5)������P���AS����x<�@ ��H$4�|�C�ف��q�)D�?~����f:�4 G��a?��蘸c�w��A �����S㎱qQr��/eb�l�N@6K(vɩ$z�������*t�
��B'�4�U��.sq���B;���,N�'��L�L.Ec�Vb_F=G��Ϟ%=w��B��xG<�'�a�b0G���F={<��(�K�&�� r,IH�B�
J�B�1�6�ň��Ʋ̂�Z@uVI�-�*��XR%�/�0��^�?N��sc㹱q��x ?Ï��bq�8#�ĐI�8d�8��8l��Rj��tgc���=qν0��M���ݼ�q�v`�n�UP�]��v������ͫ��[9�R&�J�oO��o�?�m��\x�S/�U���Kw�_�[|�^���7��ݼ�}�N��M����ε����ͭ쭭­�����͒�������ʑ�����s9E�����L�*+E����O�ۨej��TiD�6"�Pk��� N�r �\\�D��5+yp��|�/��T����.�	�H�t�!�p�!dڸ�ۑ��:���v3��̞�j�6?h�w"s�khS��K�s�վ�ې��ˍ��>?��,��J����t��t�t�t�L�l��<���b�G��|�]��H�����PC���]S��H[r���!�lJ�d��Fڋ�+6���o:x����&E��D�gf�'F��K3󷉼�L��.��Wv�_Z8�62��Q?א�4P>O о�@|��������������6�̢_��Y�$�?3���O��L���o�Y�i�/k��Ի2�-)�uuSN�P��5ܫ	�kfɮ]��$�N�/[��-�i{,�1bd��Y�vߟ��I���4�a_���+����+\���'��:3������7[�ˑ�B=��s^�"�i�s%=y��|��;���˓��R����ܿ�c�.�@,ã����}.#hU�����f�=A��A/�]�=�E�d���蝄�
��r5��P�P�ӝ�
�J�`���6�W��[��]��Ok�����m����<��ry�g~dp~|8\̈́371x �v�W�/�_9�:rr��nk��bjB��h}�pc�`c$���~��bj��Y����M�f"X<(��hjPPs��@M�ÚHS�)hP�dj�$5� Mͥ��O�ԄH�q@���S�sS��&��<f��5jjPY�!P�@_3V�����55����BS325��Q�x�q _=T����]:�<_�r�������{��W������7���_���^zq�����j����6�)�_��q$�nDA�3͜	�p�)�OS-��.�b�r.I��(E|M�l5I��T�t���<	w<�{^�}�	p7=�[+Mw5Y�i����=�fL�ȓb´�6""�r㇥��T˛5�_���U���<1�����_R)��jz�g�ǻ�]��i;�n�a@/��3v��ǈ�t1���рVL7;��;����0]��Nnl��#'��Ƚ&Z���n��%RZԖj+�i��q���A���������	���\D�� q1* �	�5����i�ljԠ�ǦF~!Kv!Gq&KU�)��P6�;O��Η��ͬ_����pgc���������3��M��'6�ʮ,�.�,宮�olln�^�v���3�s����x=��-��v��.�E�ʖw}ۻ�����[��ͭ�Ϯ�/�x���V��K���%����o��=bi�os����9m�����&G��f4�F�Ԥ��\����g�h(iZ�GO����gce$r��bO�����������S���K�ûC7rG�{�����}9k�ܙ7˗ޯ�����{_T\��n�������}��[��k��Mu�EIV��}B��'J�	,Ib�>��N4�FY�Y�52͜,#=�H��&_�Z�$|mjr��MX��	�x<���o����p*�`Ss2[u&O{���RlۓٚZ���-.r����$n����3��+�kЙP̐��[e4��jW ��*�����n!�5�*�E<����8d���щ,�E"��D ����Tl<9>� �D��&/�=�(�h�HT��c ̑�أ���1:�C�����а1t\,�$Ĳ�1,�a�fb�\�YHB&:�I�b����P�Zj����!x��!�L̳�d$﯃^�d �#���&�!4��P�<��<vM���T&�i��I�W&�*��YZ\@O*Ld�E)ʩ���������K�G�^����;w�}q��k�޸�1��Z�.K�i�fjU
��F�p4�}�f�b�4�045P�D����\¨��Yi��XsY�	q0O�~45���~P5|6�O������ȕ>)��% @MMY� ��Wejg�k~�ŋ�����7o���Ϋ��]�_�h�i.(�R��,3�Og%V��v\�+RР���!��Sx��Gy���(��Vi��ܜ2ܘZT��t��c�S�LO�"�&��Ѹc1����5hMx%�5qqH\45��ᩦ4��p^vk�c�b�FcG�F������є�hzl{�O�����L�ixx��l�Q\
����H%�F-p�K\�27��E/Kc��2��L$��U��+O�~5�ɋ5�+0��1��G����gG�qv<�Oc�S�qj,�C����ƃ,c�ā-5���� \K�i<d���P�R_Ω�j@uf~�1�̕�b-�'��E1da4I� ��p�x�8+��I�� Q<���0��hl|T\|>:O��JU�'��6��|�����9���ի��ߵ[��w�;� ��w���o�J�~+c�F����R/��l����7�q�͏�_z���Uw_)��p�^��{���z�w�~���Y7�o��_���{#��5���k;��S��S��S��U�p�pv���t�p�pgu�ܺ���T�/!#Mt����|+��J/�P�L�&r����X���%�O���zg�����p�Ӆt8�	�Ԅi^W��t�x��iwrY��v;�=^��Ց@L��7KRw3�[.Ø�Y�}�����(/tK	JJ?���|'��Q±��#K��]�.�&�%��4�L��<���'b�GR�{"�B�+B��R�+*�Z�K�5ᦖrUC�Q7e�i��$l�����]閁z;����̗��S��:�_8���ϒy�%q?M��"��U� ��Dޗ6��֧&�'f�O-�gV�6��V>�K�����_&ʿ�J>5�?�>�
?�	?��?��޷�6��4r(iw��Ҏ ���_�b�p1���d�i9�	�m�x�.ݲKד�+I�y�`�ʛ4�GL�a3s��K⍤�SMMM_�����+�_�P�4p�i���ˑ<�� Z�H4M����?�O75��<Ĺ�'r�x��6���|�L�X	�K�c����{����<]�<�tH�"�g���^�[Ƭ� �9�?\Ӡ���˰e8�M�݇&<��M�d"MM_���.��>�󱩙�:9��M�S��D��D�'��~�8�0tzq�i��vc��kS��bj6�~T�@��&C�����Y|e��hg�djе�"@�L��� �΄E(̇��2� �Ȅ;����Կ Pe��j@�!T֠a5s��Z�Ԁ[W��e��Ak�M>�� �<5������!�k�Bl�S5M��ٓ5ڑJ�p�
�L=T�L�L�����s����b؎�[f�}//��k��X��kWso�ũ������.i�K;̢�`�$2pՌ�Pz��d�X���Gyɧ���-�t���E�f�!�K��'���r-U������{tw�	����/e'>X������)��$ٚE�����2g��q1~P?.'��=찚����������n��W���껝�o��*����:�u.���g:H/tӏz�Ǉxq��^Nt7;
�ɉ��Fw�c ݂X@��#�t����=r\���o����6JG"��AisR�\��%���a��9�#���:��F�t���G
@4M�
!��ԝ�l���`X��75�yʮ\EG�15ْ�l��l�I����h
h/�[��]'��ZgWG����][�؞�2ݺv�����s5ks�+sE�s��+˅WV��6�o�l~����^)�uݳ��������v�gm����]ZO�_�\Zv�,9g�SgS.-$_�s^�O�^L���7nkﵞm��<�z�tj]��$�����$�ժ���ت�$�4�GO��)�	d���a�����Hd��9C��p��3srJ�OT��T��.�z�;�0c�g�~Z�ݔ�[�����G�#/Z�$t�3w?2w<ԟ��k�Mh��W/���xiu,k����Rs�*A�hQ��2�E��n���m��&���q	1�	q�\c�P�8
���50 Ԝ�O$��8L�|�Ԝ�Q��׵�X��lm��3y��LUu��$UP��/r��y9����㷰�N�����&���v!ʆ��2�5�T'U�K�rn��cS��J�E�2��:h��Q�l��I2�:�O��iD�����yR�8q.TL49�8)�1�(!�>�096�C���L�31LB,��&�r)�<*FH����T�8-c�#�h���d�)'��f���i�T��@&=��vra�4�R�U�ЫR*S�;3�0WK��fa��A]:焛}��?���a�8�!���'��B35��(Jf$�J�4��'~����~���+��^~������>{�����^�}�ѕ[K����d��������hj��AMMD@�]�o����q@��-��|ք@G�i �m�	x?�����-JD3�'�Ԁ�n˓��ե�*�D�ʯ�<T��/��������w^�yx{��������M��L#+��̱Rr��j7�4	W롣j&���945���?#���L�W��3��Jnv5f��Vf������E$9�~�x�����G�i��5M��D�bB�6Ȳ��/hjЀ���M�i�׷75��ȲS�7�z��86�H4�H�h4)*�ǌ�gc㸸X!9NB�W�qZ.N�ǛD���PQ2�t����@���6r��^��>��-N�����LM2�(�S�T��6N���̏ӑ�(0�$�G��Q��8��8�1,=�@C ����8�1,C��)�Z,�����{.*��h��8ze��B
�K`�f�F�g&�J��M�U�y��i�.�UKR-Y ǲ$14�4���h�G��Ir�KA�`ɬh,+O�
%�����a0$S*U���֟p�=�1>��<�^[�]�M�tٻ}ݷuӿu+�};s����]������˿����[kײ�n�{糓����FŝWKo���A�������Y��Gy7�g�@4M�����W�g��BS������]��]��^��Rpi�h�b�`o�@{e����<OVr�G���&sl�B+��B)�P�͔Z��J���k�Ԉ��M��Υ�i"L��Ԓ��i�P��N7���4g�#��R8�V������'s�m�A+g�ΟN]O7��Y�l�s�r~��<��^���0{�����]�>�M8�����4)fu���)�*�M6�]>��"�R��e��e�7e�ו�75����W�������zUK�R�7�+��5i�j�+r̺
���^Qb��jܶ���F"�����'�R��i�S�:�9��?M}�"��)��!�8�����$��i�w��pJ~���}�T>O�l`|�$�(Q�A��}����5#�e����8�
�Ȋ�cFͳb���|ܚ����[��6�ɲ�DɢMx�ƿd�O�yc���5>�D�p2o8UЗ&�qzC50��':MMg@���4�����lqKh�'4=Mw��7_�$z
�y�1L��Q	m��/pt��M4a�Ԁ2�Xn���O�'����=�{����� [��@�КS����6@�oj`?��؛����<U��_Ss��ũޓs'��{j���ӓbj6�L͕��j��ojV{=��7`��AeM���W15��'/��,�� �f�}�e6e�j(J�hj�Sg3��X�i"�/kBi�S�m��u1O15h����h@M8��A�����1�ۙ��'k*�c���
5`�15pjj:��ݹ��|UW�����k�k3��S�j|k�����`�Ww���I���(��~w�&��$OMy�>�L�v6������ݼW;����"�M�_v�S�+i�+�V�aǣ��a|�m)��r��Qnҽ��v�i׭�t*Vl�y#���9���q���~�K�!�8W�\v6�~f�o��ߺ���*�G�����G_�k����ƀ�x��!���C�L�0�[�#��` =Rl|�ߥ�u)�:r��>��rpz���zG
�#�ޞFk��ۼ��tVg:����4=���4�_k�LM(Op��'W@}� l�'k65�٢�iK��lPz�'=�U��kO�X���;[*'��_��Y[\�[�h[�<�|�ii�z�b��t��l��|��b��R��j��F��F��B��t����J����+�+��k���i3�����餙�䋗'/9�.�]�O�u��9�z��\Hnhr�Թ�K��c��䴘��In5��Z^����P�P9�HO�A3��e�Y���$NN�� Y]�l�u%g�gd���
�NT]���_0�(8�0s�Q�������3F_t�w>r�������p���n3�fYS<!˼��2u�|�Ia��j�U������6���Z��fZ������35a�&�kr�>�4��R(kNš5$OMSPh�R��Ӷ��J��%hjNx�e�TA��W��ɳs�l,�緰����ƅ��cb��L���20�	\w�c��iA����p�j�YN7˘ ��e�0T��C��R6I�!C�,����Ӱ\J<��1�I�f�h�cT�QZ�q&.�zA8�X.!�G�G��&#)H
	#ebe,���5��F>�,$�ń$)�)'�(���C����4p�S����ҤP�\�J�*�V�Hc�ޙC��雉Z��bP`b�}p��儛[�Ʈu�jS���`�p0O89%6\��o`�g�O���G��k�>�z����_��ᛷ~�ዯ�Z��>���+���;s��|3��B+���kLM���S���eH��90�0G@3ԴdIB��15���x�Ϛ�A�L�P��~�S�~"N�#Wڞ+t�JH�\B�Tk��T���'�N�,�j�na��/����~��7�~u���w�/�N�M��v���B�3˷ ���A��2��L8��;�g�7��/8~טhj��`}�5v�ݜ�Ͷ�vA����dL���g����#�b�".f?��1h�4�I�1��>�f�dj��������>~�xx@����|A;�@�	�.����Ē���1�l,��ǋ�q(����7�f1�"!��d����т&:��}jq2�,�Q�ELM��\�J-I�;�EF��[�*�v��̜=Y��S��c��c�臏1��я��pԣx�1<�(�pK8��D��P�p�(�&�٨�g�c^���J�L����| �-i�d)��$3�;��Ye5�Ҽ��D�AA�2-I(ǰ��YS�
����<E�C�`�2,Y�!�1~��%Sc��,C����bqd.G�hs�T��4�G��˗27V�n^3����w3�\ϼrݿq�5��e޾�� �ƃ���_�y�������/�^y�ċo�z�������Ϲzl�!-s��˾q/�����M���;���ܺ��������*\�,\Z-�[ʿ8W<>U��]��Zu�)�<7=3������da��Qh��Y�UZM��4ٙ����4����yRL�7������1Ƀh��\��nt��;�N�IfҤ�Nь��c���[N	�������A!~XH�bD���)��\K��:0�����`�,�ތ=��!�>�2��&����������������f�M#�53羁q;�5;��.ǬJ�V$���i̒<nA{Y5+����.�b�鉷���V�+ɼ�S�o���$�7�o9��8E�J>H�~�>N�~�"�$U��K�Y��s�����t5��	���pk>O�|�R�T�o��m�g��c�a���<԰n+h�e�]	y��[�b�q���Yv��"��*�k	�e�`-Q��,[s�E��P�);o���s���;{0�;����H@��yO0��7S����h�u0��R@w@�i�s� ��D���CMP�W 4�t�G�8�ȑ�1�(k�.:���O��	�M�?(�m�
HƷ��15hW����%�� `cp��}�=%�l��(�oej�=��� �N��_S��21��x��ya��rω�ắMͷ��Y�o ��8�@S�֗��:8�)�΄[�ES��m��iK�H:Ps�����'��̄V&\ӠP�����eMh�7��15{�}�����*؅a50��~&��L���9P��4������J�X�j�B=^�+S��*���4�*:���Vy��[���Ӝ�J;rL�i��$n��Ӕ�;��/�����G2tc^u_�h Y4�Q_���]��L͸_3�]�!��f:]5�Vθ���9�rѣY��V��-��Zf��\��"�K%�`{//�v���O��V�8��6���;�g�(I�2\��#�t+�cV�fQ�[5���~:���l�z�����9��l������M*�CR���8�&�q�2̠�#�oF�Nz�n%�G�����Z��ԣ%!3����@"s��tqzSݩ��4z����at�3:��N/�˻M5Mo �4}�Hb@x4�<}���	�5���C{�&π4��t�;�y��B�!��"�eS.�g3���%'��F��\����?�R:�[72tjx���T����S]g.�6��ΎVύW.LU�\�X�/YYʾ<�13�qi�;7�67�ۥ��޵���%��gq1��k����y|�zq�65e�rLL�Mͤ�N���ںR�ϦTפ����f��&��l�&�E	:�I�2k�659YMti��Z\�LɲP�V�?ቬ�$n~"��*)�k�Ӓ�3|������@Mgq�b�е��{�������_ə|-��9�o��s����5����NB�zYW6��5pM��.3�VUb�"5I��P�d�Da��˶0sL�<1߄�+�@�L�&L��������'�����m��a@�����@�����i�C�F� ���)Nx��)| xQ)Hf�%��l����26��dXY^3�c�����:���N7�&> \z�S�JV��L;�j8vϪ�e�����B*@#���
��!I�x	3�"FH��Scy�.9�Ko8�|&$e����pr6^��)�x��B�A���$J��d)�)G�Ѹ��
~ęzt4�&B�_��x��W�j7R��z��zC:ٺ�h4�ip2���b�h�r�����x85^M2��Ŭ?�5NF��]bcd%P�UČօ����=����7>|��{/�|���/~��7����ݕW�޹�r}��TAR���g���fB��A�'h {�&<�5�4{�W:�2w���@Ys6S 	CS�<5�q3BӠϚ�A�#@�#�h������Q�?hy��<YW��;O�
=���HOf�����R�j�'N�կ��o��o�r�Gk��^�Y�[>9�RZ�S��	��<�������	�jPG>shj��g����O���3ic�='�t��xv��{��N`�	�x&*&��ޜ& �2�A5��t�0��H$�H���4���ѣ�>t��w55��BG��/�->C��Тq�XK�HRY� �Y$=�bRm2Z����$;��4=	�1�r��$z��]��9��T�3*=��Ri
��
�b'�$�S�&��(��l���,$��r\4/���p�/�č��b(�h*=�B�"R�➏�~.&����Ø�C�=���Ӓ�Ԁϑa��u��)a�YL,S�VXe�L���WT�-�4�M<����d*�H��JbY�x���p�)�Ӆ8�Cē�q$A,QK��B�O���x"�I��@��ujGq��Tm�X_��E��b����ߕ팵��ի����֍������Y���L���6��s�������O��v�ݗ�o>Ȼq?��=p�w�^���y���\��}�V��������̭m��v��f��f�+�˫��yӳy����U�]��O��ӽ6o�&��%���R+��J���km��Dfs"�)��i��NP�@Gs�+�K'���&�Դx�<�v�hB�j{���6!S WZC7�nnW*���N�M�ų�e���Cp�Ɵ�1{Ÿ.^\�7*&��c[��w���>��3Q����؟�m�H/��X���Ǟ���b̑\�2�>���M~[�}[�~K�|M�xU�|M�|��}�¿o`�1�o�i׵�m5aC�]�bV$���IܢsYwIsQ5#���Ʈi�W4�5nKK�M�ܲ2�'q9�x�����8�����tI�v��s+>�(>����+>���t�_d?��?qk>ri>HQ��(}��IϽ�a�U1n��� �Ɖ_b�-�c�(�&��&�QS��~QL[Sq��%3�&\N�,;����K��q{��@4Mw0�3��ppR�����4��NG~������;ɱ؝%9P�<���d�;��P�t�QM�$z��J�0���1�1�"�i `^^����D��'��	%�YhW C�AD4C��4h{�� ��(���p��uLMw���\�_��s4��kbj���F;�g���线ij�]L�z& \�@;�mLMxz����"dͿ���"f�5e�-lA�R(42��g��\:〲55���@����_!k.�A2Ԡ���Scj`��g�]�,�ΠL6"F�#��(n`�SbjFʴ�fo2T�~�R;Q���Ќ��ɚ�2$�0h6P���@��%��
�H�q�$a�:i�"i��ؕ����{��~��']>U`�η��ňG9��O��>�xP;�� 
�_;�����L{��骋�[9�Vͥk|����W��i��c�[�|��	�S�t;?Tnx�+.�"�l�){�@�IdOX#քS�R�x�)�橢�Ƽ�b�Y/�|55�_�P0z��ig���23��yXGP:��:R��4` ��	�>#��d�����F���oc$���Ag���s��fO:BW:����򱺼{kr��/�h�Ԡ�4{���񜦐�	�4h�3K	���>S��̗���,Q[P�◞O��uK�ܲ:��&��ϱ4%7W�O�g�:Y�|��dgC}ϩ���c�5�Fj��Vg�7��.�eN���'���Ks��9��|���ʒwmٷ���0�vy.��L��E���ej�29fK�H��LK��u�>�T]�XX��
:�n{��bT��5;A�0�iV9ICL��Z�W�Ͷ�s-�\3-�Jϳ1�YyvN��_d�Xd��J�7ן���O������~z})w�u@`╌񗲦_^|�3�(�妩iSW>����
�	^���7��iNI�StH��$YvA���c�#�o&!+:Eh.ˌ�+9Z�	N}�j`@�P�M�S�5Q�i$�ps��P���^9x?)w	�����,�oedZ�>�k����n!��3�2��L/�"��n�IV!�Ʃ�%�xI�U�1ə	R�A� $(� ����PUB�R@T�Ȱ��d\�����12FB�J�8�`A� 9�哴�NH4�I	�QJ2��V9%IAr�IN9�xr��B���h�B�	���-�B2�2�^�c�zi5��P�4�^f���4g�C�LM��W���xx�nN]��Ū?�Tf��Y�®Jf�ڙ=�)��X���wWG~�֭�����y��W�}����������w6.�vsnc��L��8YP��)Kd�%1�kLM�����:�$�I�
��@YnjspLM��&��	�n�g���'������D4CAm#�8}�\iG�Ⱪ�u�>�5��Mͩ��ޯ
Z�'�+����W�~��׿���;�m�����,�e@T�׵�:$�C�k��:��)�F@@��������A�)�x������|r�k�{�uc/8UbV�s�V��-ʯ���l����B���د���sݓ�~W���Y���T"��/��v���~#� ��9CtOu��L"����D!'�.0�5�2.8ZH��ک�	���O�:����o�OZ�Xa��"Z>��!Τ2���Ե\�K����)���"��c?G�cѱ��)�ψ��N�q�����#&�V^_�� �%�*w7�&i�eR+L-��B,�e�^�+w����S��pǨĠ��-�tF�������5�%�k��X}mP�A��?�򡿽��.����4HF��! ��X�r��[f�25��bJ�Gw��oTO��ME�l<{s<�Pt4sC֑E��A�"�?I�E{	�$Wԫ����rt+]�5�Rmg@�y��G�;�$���E�p�|g0��%I�# igڟi�6�?���U����_Y	fY	�?ۼR]��L���66����>��@�t|kx�"��z��4}q�W�L���|B�BY��?~�(q~>^�}�sf�YO
�`���`�(�iK���em���l>1��V�ɻ�<@a���y����6�dQ���l-'��|V���P�>�MERj++��H�5y��Nm�O=��ށ���nP��[��9v�|0f�|���s'���Hv:��������&
��yt�.0�4��ɷ�K5:�žȎ^��]$�V�_�Ͼ/$��h�{���PC�~s�=��4�%�ס��m�Fl7��b���k��?�%�u
�1�Yc���|G>���(��C��]鴝����(q�4т��E٠7����{lx�g��ͅ%�c~����i����)2D�r��N�x�n5�nB-�'�\���ӱ�ݞ��=N���w��ɍ#�7X�VS1֌d0Fwu]T���^�ŋ�$�6&nl�yI�WAT7�~�y�Tւj����k�UtE��!bDZ�>�x��n>L��6�ӹ_��Y�)�����L�X{cwP���@�?��_�B`����8GPS��<�h��p.b���݄<�7����.�Ӳ�}�V^�����Z�R3���J�'.������{�	��\^�Una������şs��������P~�-LҟT+8'�s����zR�մS.�l�?���I�L9I�á܁5��p,���C�!�L^Pi4\��9�J~�+���9��-����g;��K_&��8�_��fվ�u�[)���W��@6)=K�V��0�Y���@bgKs\"��ZbY���y3�#��c&A>�y�A��sn��Ng��7,AW�j��9�xI�'��ϩ!b.%_:�ɤ:1+��ϩYڱ?�i����ϻ���ק�^����իW�rhBO:ǧ�nD@%%nmp�e���u� ;1�ڮ̛ɜ�~Ű��L�������"Γ?O͂g��}I<
^�.�d9�s�*J 9�-���.4�	:Y����O�x�SR���(�������C�($֌aۘ�.�k���_8�&��n}���8���|H��=?/���c!�{H�ZEG,s7��h����\!�h�>�����;�Щ��]�'��YS�՗�"C�3���ݽS�Գ~1)@�`�F�����R��N�����4��m��^ �l��e��e�T�#���Y�<�'�/��<D����(�5���3c�{oy�(zX+i ��z�/!Jr%rR0�{�3�d�����M�{5�r1���h0	L_��xX�ǵ<���1�b��"����j��cl����uO�%�C>s_v�;�/����x=�����Ҟ/�w��{�~�+/���6���1�6^v��+c2[��Ɯ`�QI��˿L��x��+f�ա �<�!�Ia�ft���a�T߇y,\Y��)���zB�7���=���c�$A`����!<��&c MW�.F�g�u(e��st��[E���d])�K�2@uX�S���O���[@�g�L�Y�h��O�V����{�WZ�m��]#x��B�
s��N�N.$��Р���_�#��[`��y�L-9�_�B˖[@��A��2�i G��c�4\@�2���Zk���[��03���$����V����W�2���w�`�@�])w��B��9���$�i� +l< �߇>���eʜ�|ܱ��е0�:�B���^�Q5��Le�~yL,�w�)(����O��>�z�����F�٣��׫P��Ɲ-b�_�`m���&�4�J�b,��y��8�q=�p E�Y	�P;��;��y[��*����v�`Z����u*R�>���J5Y���[����g��:a��l���4�V��C��]H��{j9W�p�]�;i��-��}�ە^���k���R�߉޿��U�U���謠�(�B�ȏI��Q�*t"�s�ؔ~�Ss"������o5����Z�Z;8�s�ѡ�$�cV��B	*�I�ɂ�z��"�������j���$Lm6�qt��c0� >%%6�;��(9��o�����ã�gܖ�GY͗,Y#S�?�eP��ev��UV��,��p�^<i_�$}�)_�E�/���v����W��M2Ne.uf�s�����J�O�z�'�!�`E��m�a�298��ʾo==-��nm�98T+�2��d�L�C�>��4���RJ~mi�����i���j���&�۩-Y-�fDꫂ�s��
*,!-���.��D4�$�.5�5h��[���'w͉�H�SG"��7S.!r���P�Uc��������������dmo�q����/l�E�ޖ�����o�3�ˋ�ę�l��ٺ�˺|U����^��؛��Q4e���u��Dh�ʐ���9�QWf��j�y�s����?��&�̕ט�����v�WJ��~��˕�e�	���
j���G��c��y�������N�ò������*���/d���3u���__���OqUF"z�Tr*�#1u;�2�-�iP'�p�����_y�d���=8������ W���*ຍ)����~wɅ��eMh��]�Z�>N������9� �\%���q�G\��7%U�3�Ϧ�bw������;������k���d+TV�Vqpϙʚ���P(�kYM�g��jA"g��I�z���(�jFt���X�:v�y�L+B�ѯ5�[�5ן�)d���?�;2��*�w����t9�u@��y]Ϗ��@�I�A�_�>Z�M�'ũ�ũnc�X�P��������%���&��!�Px��w�?�����ž|?Kx^�!je��@���XKk���C��Y�a�i^j�Y��8�D�w8h���@���zk������,��w���$�i��T���v���K�Ψ'];�3�� �\{3��qު�s��P0lG������8��̻���� �r��x��"�{|nd�o����^�Sl[Gܟ,�����aVn.��U�ն��ޝ�P�#C&�&�:���2�v��5�E�р>xs�yu���sc�&/$_x� A0���ඍ����/�� ���`��	�P(�H+r�����T���S���(�)N���D��L��W�t�D/��hL�*�ھ�ʔ�x@(I{�H�^-�P����5Av�L�l`�O���i�@juNu#LO�u������Ȇs�k�G>�������n�I-��-����A�Z<	�9e�Yb�r��^�SO�>��B���JX�Zbщ%�T���D�E��G�X5�XO�徰�Y#n׼�U3�R���%j����K2u�׆�~rC�ш$��Я�`H��?�b�u)7�	O�P��Pم���(\O�2�� Si'���N&ՙ<�{wO�v1����pwkga?��p��8D�	I��	�c^L�>�=�L�КM�~��I�3r�RU��d/��.�è�%��_�5�N���N��Cr�5[I�ڮ�57ވ��|O�Vq��������ʢ�J���5�*Sc�ܮdO[N��I.��.������ՕV��DD"i��<�e�'����"�~�.6S\�$
Ε�=u�&Ջ��B���ٴ�,J�� ��ts�6�!1<A3�iB+ܢn������"�<#?\�F�
� �)�����3�_GR+�vZ�+�뀟�TĘ3+ G���Qip�c���-gM����b׬K������F��2U�L�tn�v6�����*������1(�M��Us}���� ���Ԇ�&?����Al������-~��s`֨V�F#	OQLe�,�J;����tRb��n�rj1�U�8���<ޱ��e>N��G}]�*���o���$K��}e0a����e,���=x\����]��0�p�S?�<�NV�Զ�^R�u=i�v��Ʀ���������!6z�����s����9���uj�'L�r>9a��d>��l�D̪K�*�9ߖ� `u��A�������e��9*��~"'?��U�BM���?7=+���*����R�+�QHw�Ƥ��G��)�]oW�^7��?�z�U���9K�<__�jih���������r=���vLN�܎J�t��ԣ�eN�6�u��PLf������!p�Td��O�e ;�ZH΢F��fr8�+u�N�u˫�$վ^�c���7��H��
h���,j��z�4���h]7���JZAo������ ������SW�����?U�V?�������r�F/U"K�u�Q��]�
�I��O��$Pnc�y1c;#=ʨ�УgٕKJ�sm[��dI'q��e�i�k��Ѭ�q=8;;�..�K|B$Aё=�A$2�5���Y�"�Qi�Th5 (��$ ��I�!��&>��42�?��/sFD�l�m�R\fi����џ6�c�`�C5QeX�l:a�0E�� -�~jX��E�8|q�6cs�l��恴�֧�+T�
�� H�pe��wyQ7��"*�"*uj\仭Hnf��dMj��Hb�wT;H�!�*8;��� $\��-�����}�+��?*Ws�;��sQ�OWJ���5�j��[�f�*�^V��jHi��r;U~#b�P,��BV���/R�L�`ė3>P�t��AF�\D�7eQ��O�E +i� �0Wr�ŵ����Ճ�Ӫ�ϭ��q8"�s,7q%�pE�kT���u�:1�D�DI���:i ��}3)��uґ��9jPu�-{g��~W������`x;�X�̄�u��o>�^�X-���jN�eM�f��d��l���ߢpd�9�2�j��%����gH��RW*n/�՞H��zTCy�v��K��wP�@���t�nc����ԑ�t1�4�#(>Џin?� V���g��Ol+]O u SaK�Ĺ�o=H�3�)�Ԫ=ʅ�Z����6����K���>���l��FٷJ�~F�|�����C4����j�����������I�8Q��^5Xܳ��}}��x��)��=�y�7gi��|�m�LmvW����ҽv���њ�!�����	%-�7��DY��Ko�R����~X������6*��
�p"���;�ޜ�،]s�G��s��Pn�5�<����hY���~����$������dܧ\��vN��U��k��ɿ&����t����5I4Ǖ!yx��i�Qg��إ4g�Z�`�m�x����b,-�D:��Y��cx�;��=�A��EfYJS8���N#o5��9���>$L4^����"�Eӝh��<]"��}�y.�髈�ۦT� | T����N¹J��?�+@��ɫ^T�ՔȎdJ|���?���Q/é��5C��jB�z�?F{�SG�<���I���|0;�I��`�"3��΀�;�h)}�� r��)�������S�c{t����S���o�6��3@��&6$ޅʍ(kW��z��`�l<w�<�Dk*��uT��� �VpZï�h˻�����<�I��-���j�~��g��+�Qm�9�o��-��<��nӞ6�4��!�g���T	�	�]�>�%[(x	0�|9���
huV�k�	�Dj��2����d�SSܤa�#]���q����#���I�e#�5�<�Sãy-�} �rQ uA�RR������A�X�DT	u��hɿ�V�L�����kē�����d��?<���Sхo�G�yv�ž~���c�TFV����@�.2EZ��i�!'qu�sB�(���y$?3��k�����X��Q%�5���$ō�9K�|D�C�#����^���JZ!���s��=+�?o$ӷo��8��k���b���p_���ԠN�~��|C�"�}��|tfa��R�#��h�f����q�r�.G�x\�a���e�U@���g'>G�1A�w����?�Sy���Z�\�?m�m��[@Fx�EySs��t�m+	�nJ�Ӌt��y��T�\ߙ��x�S�p↠6�~c�˵�{Fia���2K�h9<�(�S���J[���#�Ҋ���O�����fq�.o�A�<Aܦ�{�:�⩴�Q��Pd~]x�\- ܈��Aϧj�j�q��,k���������V>���#IS15�\Gm+�V�,��.|����3~Ţ��׉�'��S8�������yR�e����Q~�;�">�{���YQ�R3�i��#�8쯉K��M��ٶN�r�GY�1xa�I%���<'����*}>թ,�
�Z����bXֺ���A��VE��Nl���EG	ŅTeB�T����S=� 	AEE��:+wXRUs�� �%�ig;l��u�����s����P��N����ZY~�/�5�� #xvf��c�J�/s�4PЫ����:\Q�`n�;$ �_�#�/E]RΓ�E "�����W^ӥ�d��h����TZ7��E2*��w)U�ئ�ϓ]�o���[���Om�ƾ;[�)�����f�N#C�Wu�6��r-)����*���p�?]�	 `��	�>K��PӪO���|����?	�É��E���j3� �&D�<3
Ⱥ�R��Xs/��n��_��P�MG(נw`8����˘~��;!���E�j8p���8_���ds̝њG�d��"�g4�XS�����d���4���n7�9v�&�����ЫfJ��_>�U�pt=���-��/�v�_7��p	|�OIث�-/��%��Yr�K�j�As�5�W�JM��HBL6N<�p{8P�G����`3�'ɾ���^����h�'����#AT��ރf�������;�b�U�riU�+;����MNsM�� ڃ}�Z ���N�k��E�K��>(��]�{�`t((DB����`�咽��Q��T�i���=5|B���G���ߑ���@��|`�'#R���t�UA���w�&��!��8JeF�Q��8���Q-�).��%񳂿<)n�}O`;v�!h�F�ĉ�'�t[�S�X%d��ǆ9�G\O��Tp9�U`!�I��R0��k9����&�L�)�+�#㠊�mRע}?�kƴ��=}��,靘�ŕ5���y�p���'�%�<��VY�_LɄ8�4���Q�����ulB�����rA��%����T�)����pg��|�n/4��\�2��.��2�R��0��S���uS};�|j�~��y����z}����i?6nM�l%_m��Ky����X�?^a0��؊�_�b�szS��tYkI�}����k�;��E�v���iϸ-���d����Qu~��}�y[�z�.�>���R�V7U4����R���ʑ����В�M3T<�}���C�Ɨ��;��4�-�QmM"7L+�+��*Yd_:Ƿ����P���4���H��w$6J�-�����qzA��ݲf�1{�ST뫩�_V���`�jì%�[l8���07��Ԣ�~c<��Z�n*��Sn���B���E���}����%e��#�$���C�[��)l��l�����9��;�ցSo�wrXo6̏ʗF��j��DZ鿭�n���t��L�ǡ\3���\J��xᆶZ m.��A�N$����ڇ�LU~�%�U���DހW]���#(�������L��Vh����Δ��%���L��G�Š�`�Be�n'��Ot�gW�:�i��(`��Z���q�z�f�s��5�Kw��C�������� 	���R9�}��\b�*o�p;5��aJU@����A�;y��Z�Z�9ŬjCE��Gx�m�[�,:dz%��Z͓��G��Ag��v�"ǆ��uk�Y,m*vO���l�{� oPLR<��0b'�z�YkHЉ���R�ow�^J����K�������D�Z�pk~��QnWPG��Q��-�(�wΦ������"�K"|irO�q؀�0b� 2G�"��l`�]��\J�,zGC&�x&�I/9�`nw%�[��E湫��E6�^`���o[�6>d���!��7�DZ�W,!���t>��I��c*4�J�P�hKq�-�z;�֡�� NF�@��{A��p�M�Ҝ;�`g���+
ѵ;�V���( <8���J>�l�`�%Lq�fm��
yL�������Tٵ�J��')aO��vT��7�)��"o�w`��>3 Yƌ+X.�2�t!��ߔ��B��&xZ�$R�Q�So�8)�@��\���[���)-;bS�$(�NQ_�	Q�|+-�d6�V�HU�2r@�&���Gf3\��ڹ�0�yt�Q-�#��<�B��g+��<�t�&���sس3F23<����'vλߪ ���?���aL�Y�NZ�M��H������-o��N-�ɕ-��3��J�et&iV%�u�e��2�̵�����|�Rw�.�V�+�����2*BR������JG���q>&��1���j�8m��r=:���uZ�bIY��w��r�r��-x8�);S��
L��xc���h��ԭ�߭#�h�|��`m�Q:啨�1�����fB��W-8�= 3xP��� <h�Z�ɽ5P+�\-�-�o�<t�u0�B��M�Œ�c�^��<�0�#H�'���򻗞1e�:�e@���Ԉ\eLF�-�C�:'�����5���H�b7Rщ 9)�c���m.��s>������:*!��cW�B�9]EhjWSP=��-�s��ԯbv��V�'�n,��ભ�dh���˱3� �/���������n�a�{��|�U��\�jH%�E��|نf%��2���b�>���io[��o�&O7m��_N��gr����������7���1�^�'z�Y��U3''�Ƣd$a��6�.��F-zV=��3�	*?��A�����ׄ%ps~'���(2�Zb�vv�X�h�MxA��`�E8�Ȁ��\8<�j�,��n�+��v���8��k$B��:3��k��d�N�n!�f��G9���x�=��z��?|��zK�����}�h�p\_&3%o�]�k�m�2��Ӄ�7����vh1G<A ��̖%URk� �S��\� ����e��6{��VXnϹg�D%i����� |��
�N!�LS�" �R��@�	�L����`���b�W(Hb�@�'N$���^�6 �O;]&Ť��"ks�(Dc����b���.]0D�b��/�;��2KNP��k�E��ΰ�D�4(�b	��Q�i��bN��|I�C�MS`T�O.�`YUxt�5>���5�X�����}�%ku_6��z�Ӆ�{j8��y��\��G�*Ay{�%%D�T#W�=!��I�:Ɇm��w����,:�d���ޱ»���ܷ�ܷ�l��?71?��3���S5��8%��q��� pk���h����	��i	a�-E���X���r�)�T��@����%�ĚJF*�����^�� �\,CO`���=����o]�8���u"g��ǲ>ۆ	ǒv�c�g�j��ߝZ?}���HL*��*@���#��M�M�V��{]�J7�`��X����xeE[OvE�p'��QE�z��wK�����y�C�t�3�̬�G.�g�Jc�:����Z�L7��d���M�����	�T�C`��aU�,�i�b.��a>���L�lt0X࿠��-���}U�56۷�fS���̟mc�D�f,����/������"s�)_�t?�C�15U�����	ٷñKʜ�ˌ�7���;5�׌Bq��'k�{l����q��;a�?ş:~Xwm���{�5Ƴ�"������Kv���o�@�F�-���rZo9�'����������XÄ�*�Θ���/��rA��Ηu�����EDp�M�EW����EK���7��8�f�;#������Ɓ�"Э�A����ۆ}��x���N���ɻ��_. ��_��C��i��I��H�FH�\"NO�ddf1D%g�&qz>��`��r@(ϙ��y%A����̝PC�/
g:�cu��O��h !^C�ә�0L2�L��F����д���<\���h�7���<o\0B��{���jۿ�1eG�j��b�Jӏľ�t�êݜ�̾ع~2��Ri!�?����V��IW��CKR�U'�松�;�Tn�D���?���{	n�A�,}����K��S;�Ƿ���B�:��$�x�>B���}�����$'��~u.H�P8OB�ER���S�޿k\{	���	b(x	J��r�&}&�0c��>���0����P��&E>�[�KMY�ދ�<B�G�Jd9��9�J�]���F���<I��Y�WP�4��F^�;$�>}�_�f�xH�hJ ru:5n F	:������!!0qy�`���y�ԧ�h�:<�$���  T
��j]7g�kS_K(	����e�C����"�r�K'�	�����N�LcUj�R,K�D�OU,>)kMw�<�+^݄ͷ<�jk�x�&e$%u.���U#-6�6y�5����L�hZ��Q��q3�-.�=��1��--���"�[&�x���B�8��\�W���%�x(���X�����KL�C{	�Υ4a�=��(�/����,Ǿ@��*8��OЛ��NG[aяi��M�D�:��ƝN���i���_���52�R���F[��l�~�&��e�6Oke�ь���Ӑc;�W�Zx��1�QG~U�ޔ�oד��=��Sv��R��Ǉ�r˂3BP$C�&�%nU�`bM�6�Q{9>�G�b2]}t�`X�j_г�SNv������c�*t)�k^�������(�����-/L����<+q��`��g���s\��4�&.�6hC��ʅ�5Y��c���W+���[�L$"e�^��$�f&Wia�ܾ6=%���ظ��R_���W)IV�����b�d����#-�(����y0�K��(�w��������xt��~�'��F������԰Z��/�-��޺%J�Z2�x�*	4��
�&�����O�מ��Fj��L��`�A�3����ne.9�O�M[\���{34J�\;�n郞��Y	0B�	��s#��d/l_�':6�6dx]Lt�� ��#e=�s���}E��EE��v������A���?���i��'�Dzl|��E9c�lJ���JI����xe�xT0�x�����G,	 �a��ӡY2��<�l5��ej�J�(�m�����{h��e�B�,�e�ir�6�]X��3U9#���{� �S᪴�
��c�p�!J�(�T�8��x���DxD�cfQB7K�}�qdB��H5aAН�X@������@���{r���|�}/D
8*�b^�fC̴p�Y�B�5�|:E,A6YE7[F
6���'΋�Tl��!UZ����rw@!�y[Z�	���+k�*����~�@�C� �,�2j�|�6>f���h��]�w�@ؐy��`�_րW�������_���f�$�6}����ο'�>�o�}]�v��3�2�UX�(Z�����X��[^�G���%B�$>��NW�Чe�)�4
.��W�"�s��ҍ�m�=��h-&l�#��p����-�u�d��U�J���<�%��tpc����g琗��:�N�on5�u�����:��V诏|l����>���쳷�T�+�ӱ�U�j�4��ѱ�d�ڌ����d"4k��i}r�#�����_x׆ouTo5ZOݞ�Z���^0-�����t�f��6�����S]���ά�>�E)�6���a��K�Bl�gw���P�#+�j�r�_wk77���1�O�+�N�<Q�ʣ1���Ku-KpS�ڙ9f����~��� +�<��}�(�4�9	J��f��K����$q�o�9�̸�M��8ha���o�|���A�`r���y����x��y���xx��!�x?(��v�$:�A��m�s�o;�h���W\� ǈ˨�LTl]y�����16R����\<�`w�(^�N$4�(�ϻ+(�P�U���+W�X��q��̖�v���u����N��S��8��g$�ܸ��$�缣�?ق�;������Y�U-&/����Q~"���LAij���Ʀ��8o���s7�Q����=�����0#�6�Q���#�p+�B��BbG�%Ę��Gb���|�VTl�Xnk���z+�`�?I�+ �+y�v�sDE��-��#��T@V��g���������u�D᳥T`�m� ����.��#����b-c0�[=�z��},_�z\Q�����n@������v;_r�;�T�%��t�J2������O>Hj/����tU�Eڄ_5@#7�`�w,|@����1c�l��?=�Ѕ 6muX77�@7�j�KfN��X"\[�9��Z�h7�t�����gi��we��W���[�`>�h�3ջm`�����_(��R6��̍7~Zd<X��p�q�E"�Ɔ#\��olw�-(��1h��.���95��[���Q�I�a�<������TR����gJ�/ŏ��z��zNvTɠ(��:t8e�eh1|:U,��@s�����8��].�p,c����1\��7��6��a<��=�����������]��Z�}j$��g+��x㰹�bre=ey=ua.�X#���ņ�J2�x�������~��n�¨"�� �N��V�e���bC��U[���W�ļU���S�z$����	���>���Ie
�4��[� �t�A��s�)v[�mI�s�L����h����|�YL�£��R���V�V2f���-�C�h���a@�©� "kU$Z%���׭��}�w��<�v��	S%Zp�Gy����H���:&�ߛ��H�X�X����UG�7����LA��Q<!ך�����5DΤ{�.�,���N���
�ܰ�B�p�����VQf: I�cպ��}Y�R�*�L�����5#Jœ{6�JE"!,
��I�tG��,��@�] x$�V��� �z��ݽ���	���O$}9a1��>����Wߙ�ent��ƙ>_�E����5��M�c�d�-��o�j��V���J���+����ҪKKF�EG$�8ܿ�`\1�dO�6�(7 h��u���Y�����Q�p��Q��H��e�~�br�`�����u�{�+�/ǔ]Ϧog�՝�gzo7'��j����/�M[@��ǽ�ҾO)��V�ȬH4�����%p���Ia���	�UEB�J��vݟ-SS��5uT"�'�Z.ѩT|��.!�w��m�̑�'����Bi�p�!"qR�Z�"$a�Ե
��ﰑ0�m�����=[R��
ۤFF�||@<<rJr��c���XqpAƀҸh!�oqbrQ��rpC��s���c�ec�C�.���a6��I�,S\ϸc��Ԓ��фS�F/����eV��4Г���i՜Ҽ{K���o�������Řpu�p�&���Ҩ-���V��zH�'�̿���29��;O�y(�kg;�y��6Z�٬��m�-����� �������u�h��m�q{���x:2��'d�9�˫�ӡ��AJ�m4�M���|}�6�L!�J��|�p![w�xD�Ϙ�ΐ�Q��eJ�mZ��d��Z)��ڴ?ϕ�;E�1�R �ڐ� ��BÉ��h��A�RS9��#݋Rz� �s�x�?pR�:wnĴ�q����T�nިE���|�g��lf�v�׋���j�zsR�_��s��ߕ��C�̻��s�QY�ӵ���P+����X��-��m��л�?��L�Z���_~�*�k~2������v*k&33�I������!��m��B#b)B{V���=)��[����#qo,�ݧN�?� �V�ֵ�^��h�tz�D\+Fv�rv����!�R����y��ϴϻ2swǅ�S�w�ǰ��������D���	�����+x���a9���%�sk�n%�y0�P�N��/������l`5���:%fb ߄ �x��_���=r�P�+�w��1����i�zy*��=k��C��L��+�=�p�A����À��U��	w�8��J�y����d�1�0���17�]�"�ߡ����=���1v��?�Wu�Ӑ*b�< ���)�����(D���l���RA��0�h�����SQh�vgeG������n��
ش�������	-�`�X���H �'��V�?@��-��vr�J�9�Ƽ��_�k���� 6��h�瞉�@٘��Z�Ig1�j�3�C��scjX��&x�~+�8��9���&�F��'G�����ࠪ�YE��xmP��	����˃m���������@����e����xh���@��[��a$`�=/@>�O�䧮�`U�3�u�oq�w�j�!ݩK�>�̈́ͼ��݄�(�Lx!�S�����7���7��E��� 2%9�	_����h�'���skV�'c0�����'������G���k��������z��62�����Q?�����AAOG3X��ďJ0�!�����0��2�}���\�n�L?j!��!��H�Glris1�V���m�L�U�U2�璟�TT`�le���������m��o=ķb�6�8�i���䇱��[��+�7	�Q�@Ê�|�����hp�W�bQE�͖ �)a�g��ە�ciE�B��K�L��B����0.�i��u}�RL��[�8��Uj���T�֡�#L�v�(Y�6���Ÿ́��rfj���g�~�/�xS?�@�5���`�Wk��q��`���zj{6�T���C:�qH�Q� ���c:�Z� >k8�/��c��>����F�V��u�,���z���� J#�<t1b��yl�JD:0e �K���9aZq�Qb��d"ծ����Ic)o-O����F�j��U4ʙy?���!���˧$Z�OZB��V6�s
�P�[j���;Vھ�'^d��5?���!�rh��b�UM��;
����<�@�/���r�k|��;���<@UP}A�̄A@��<�|��އ*&ۣ�;���/O����m���[�/��q�-��U{�}m�,τ����?���	���o�ҡ��uT�e�f�yTG_QR<����-(b�� � Jߑ$�V����8r������:Ӭ!�0��������@-�̖'w�]����I�j+��Y����Sӝʸ^�����^��Z��_���׫��ۖ��X��pVGGX�/�q>9���,Z� ���gb�z�gc����*�S�l�M1��lt�ZA�
 E�KX�<#uߎ������k���kj��%J�)��s!("��I� ���5=dČ
?ˆ�R���,��) D!�ׯU�1"�#�����ka�?H-�K��=~7;`.�0��<�q���p���G�*K�JA�,b������qE�2f���ȯ3���<�	8��*���2�O!�-u(nQ9J���r{�'7�7^^�$= ��1�p�ε׉ނX�Tǵ��XʪT��h��+��C
k�����x'[�ȅm�V�o����]�KM���WF���9S���1:�L���Lמ��A�緎�X\>^�r��1����+����?Ɵ_Ϟ׫V�Y�XzƮ�;�y:��-�b�����D���f)+�����}�C*Ҕ�r�k0Ր����T�˴������W�.�����:3�Nܬ|�s�&��$��H�d±Ԯq��7ճK��� ��e�wf���#���,����iu�=`2����1��B���IN
ۤ������6�۪��^�s���qt�QQ=}FpA�Aiv�FR�Z�;�n	��ZZ`����;������=�Ɯ���yf������F1`����r$���� ��.�"�r��9���L�C���N"'<� mL��`���i�۶����C5�o?xy����餼 ��4G�ǀZmt3��V߿�cI��K�o�V�=H�q��B{~�(!���}�^� �W���tpH׽g����O�(�]}O?7*���o�G���ڑj$�����Ĵ�p��gp�[�n>:�=F_-���ͥ���i.J*��=�K�6���z�S��q��I8���JRs��r���od�>0�����]��q�������=��}��/FQY'g��٬;�nv�tw��U����Q��ũ4�,�jw[�ד�ѕ�h���q��ȍ���>����0@��%vĒ��w��|C|��%�����f҅ى�Ó�yqF>�;*Ì���<*s�Oo0�{�"�^%�SGc6(��#�����R��w#���~v<��5��g�i�ϕ�D�2���� �Lέ�
hp����Z�
V�r�<$�l1a��l 3�KΑ�i�˙���(�<#�Q���{[���x";��V���������<�oi�g�!(� '`��aǾ�t|�ڋ}�ϙ�*�1���ͲhQK_���eY�V���ќY̅N)�I�>�<
��RY"��Y��_{���:?,���E����icB������U� �.��1U�{KX�46�߁0�m�����O����5�6h�.��,�Ya�&5�?O��ߚң9^���u����%d�*��`N�dn�U"��k�`5�����Wĳ�U�Z�Ʒ0gY]�!3{/o'���N�O��OeG�l���b�ʎ�����e@&�9�\<���&�ݽ�#��GZf�B?�u'�S�m���8�Rǧb�h���>��0�l*�)ś��9��	�ẼB���XUh.!���c����8�b���08m����0
�3d�1ti��n5�q(��`�Ʒ��,����p����(4�/KycGte�2��ĕ�t�_n��w6qeM�g���kaM\�� A&�RgI}Uh��SH0"�����>z��	���Y�x�cV��wP�̂o�f�!��3�����[�si!h�1T�W�H*�	jh�o��E�cĔ�?��ƪb^d���������(=�[�T������T�i)\xA�lL*��$Na�[\��:GQ���VU��bd���؉��H��7.E�8;a>�$��4����V=�*���J�^����q�+�i����O�hLn�@�@���Y���N~F>q�#�s~M��ã�L�|~x���*��_6�>��L[B!*d�}�5K�\y��W��29C����d�5i8B��S�O��2DR���)r�\������i&���Qd����g���8wڻ5�+���/�I�:B]���=
�0���d�ܰ6s�#���Io�7Ԟ��?>�^�-Ϧ��-���wB����)^��V	a�/���e,ʗ�
|qJ�M~��-p� �R�`��W����[���LI�qE�|[%�y�-q�Ic���$�r��2�֕��b��(%=����k�H,�QC)���3��O#7�q��QVVZw�^���Z����F�CONs�5�G��!G'Iu�Oj֎5ĥQԨ�#`Z�2ъ-m�E�O��U�}X>Y8��YT\��Q1�4��V��В�7�t�s��ø���C��Q�������9R���r���j]�ß1��F�:Fh�� �X;��#����9��FKǨ*œ���"����d�b�,5t��ik��F@�jxB�>��I*�Vti�N���7�/)e6����?�����ó>�����̼����tn�O0R3�Jb��d)�`��RN�_��_��˂p�Xh�ӽ���o������:�����q�2#�Y��I�C��bil��Gй��F��@�mU�{S��@�eC��"��&��0��8��<���n���/О�ߡ{��pM���7�����@�|7��lbϨ��O�x�`�����FR;eho_Z���V�CM1"���n�·A-�Fײݡ����&!���5�m�siLT�¿+5͕'����8+gmO���?^���u���I�Z��5i����N�����Xex;�}rh����cnv;w�C����������Әq0#H�"��?�5�4K~c~>�<���X���,��s�����"1q�d���G�Y����RՓ��nᦜ4�p.I"4�l���^��1s�%ڕֳ�o�z*����v�Fo�����#�8_���ƽOF�'�[��F��Q��3=\��ۖ�������3%���v�Q�<���f��ݎ�����������ٚ�ӆ��8ܞM�Nۇ	fh�3����՛��U�����j��P��9e�S�]�;�����/����_���?�:��1>��.>��]�к>'�K����&�[y�~��v����qg��ٙ�}�詧����y��]��K���%ݟ˟��>L����X�wiL��:-�0[�ȿ�V����`sTe^$�r�{���>\E	cy��@�5C���~��A�Vyং�s��/�>������ST1���X��_�@ɍ6�d2���]�{]���%h��scTã����@���o�'_��ߢ;��1�d�z���B��i��~����E�fHBĲx����>�y��	4�	����?� ��8TZHKWî�)����Ѐ�� 3M��I�͎ (�����M�%U�����]�V������c�oub�����z҆��c�Չ\#	���o��n�z����J�>w�����6��{����J�|Mh�CȒ���a�*�!}O}*���/g�����И#�Hv
�7��l�VF�2@��<��ߗq�i+0��y_�I��GK#��|N[aG2��dBŴ�[�U��w�����L�ނeys(�?��.�0k�5�ec�8�nB�}/6�/ϥ�!]�AEZ��D��4O!o�Z\7�5�O��C���9e����F�^��O���I?0���p�_��^�J��p�<� q���z��{�Y<GH;P�@����cع�E����˚D�t�g�/8F����/~Ff��9��۞R	�Ԑ9�a�l�A�EG�[�։�"��Y�"�����\��;���C����M�\}o��7v��8��F�V��'���]���a%�
bq7O����
C��a��?�凇��0�ƁOɰ'�O7
��]��A�4�Z_����ԭ���?�S���Ʀ�����c5XG����+�AyE�Gn%B~�����H��+�o�m�r�W��K�w3f.��}M9�]n�o��H��D1�.k�]��p<��P�T�F8�Ly�U6��lW�:qA{·��L���r��ta��H�,����6�a�J�x�N���/���[�#Ux3��uF=�FL3b����Z�龸�v^������bm���
Tp�63Z�9xpE�F�l�_�Y��.��_�?���]I��%��D�2�Kѹl�u^��[��P\$ʝ����$N�F��`aj\��\V}(E6�Ƿ��d�X4or'���,�w��~�<������d���;5�rGȬd�����+��p��ꜭ����|߉v�3�xW{A���x�(����h0c+*�0�R&f�C�`�݈� q�'yY��v�@���ƒ1eM�h|��$MJA�J%�D��j[�e���Zdlty�$Fw6���=�8$��h�F�����P�:��W�����eDmnOn?�
hI���<��z]����G���С�ߏF��������u��e9����-5:c��b�fZ�@����xD"B�(�6<9#�k5lx��v�T6鄳��'�L����q�!C3���DF(+�tw;���$��^t1�0�+4Z�����}⨥V�~�Q�X)"nU�kp�Kګ�~�	�z=k�xmt��?o?�	��]�}�l�;bL�Y�,[��|b��<Vڒ��^��ʘڢ��#���j�D�%o��n��j��Tr�g�ϳOν}4�qW��Ko��7pD]�LY�Zb��2�fFa�c
�`K;){$7vZծf�!��OC鴧Sm��nU}f,�:g���>�x�:8e��Aԕtr�r9��Ӿt;���~1�o'����L-3�p"��Ӹ����e��:���`�cƩo�$*���o��k���i�����c���5c��ʲ;��f�Dð��h���S�/���DXV�/`QN�����>�g���nXyfP��zF�g�x�ۛ�kE�b��U_�K
�^�}5�a���Uo#v;��L=�<�&��C�����l�WZܖ�]�Lm�h-��O�nG��"C&�${􈉼~o���f�x2873B:x�0{���vx2��O�8�4}����)����o��x��{���U�T���)��J\���}��/�u�e{�'z��&�Uck
;�D�Zt���5R[��:��]K�Z���a�Ss~�l��+f�N#��O��%���B(F����m;B"��Ƀ���-}�7�M:�	�k���)�����Yx
?*T�%������������(.@ Rmeة��^[�fM��3�SUEd}H�g6ޡ����ï?�;�'P���غ�-?��.�v~|��5�D&�>����>��!�w�W���ؔ�q�M�~�;>�z.����v�w��wЧ�]�l���ۧҒJ�v��F�c�䓗�
�q��) sk�'XaG���P�����ƍ�n���8��B��nVn7c�}1{ۓ���A%<co�W��W��.&��1D��!����B*;�`��j���0���$��\(�OP�F>�N<e(N�d���A3��jC�Ǹ��Y���F*��i�����pSH��T�8��� mʒ�\�/�dv�g*LSFy��������qJ�Ƞ
a�]���,�����X*-��4��dR�����2��{z� �ݡۺ+&� ԗg#��
l+�x�R��%��K:
�� j���v�޽w�7��\{�dy�9�Όkl�g6�N�Tq^��x�[�� �f�6)oG��b�����.Vp����їjy���[󵽍Z3d8ǎ�H^�f��l%g��a�.��L�f�Y��z��u��Kw!�H��H�r�Ȕ���R�S�NR]܂(��L�`���ȶ{@Z�,�ٴ��Qˌ�\:9l�2([�,�
|%����l`/�J�n�-���@k�+c-t���2��@�w~W�NN�̰(�6�Ȥ�S��9�b��,d�T�%d�ߒj���k�n�wmG�#�f�д^7�j��(-�R�~���Ư@z�d��z~MbC_v�L��n�hy�3��&�Np9|NcY����]�Mb��x`y^p�	��2��iCf��Rf�iM�'�m^IL:�'뜞��9���3v#���`h`��P�U�y�ʔ��t!F+��Q��ƴrT�wnvr�#ĝ��v��P�v?�}?�}���u�x���a�h�u���E	���o�%�K�2۸��D���0�,������	���}Ȝ%��W '��+P� Ҙg@"��O6
X^�*��
f���j�x���u�� ��%Ì[jVzr�����5���o@�x0��cG����L���r�׎��K��k�3ؚ���1�׽�N!u7reG��%'vܮ�G��J�����V�W�����b�í��PQK�J�
�*k&)��$w�������^  j#G�U�C��ZEN.*m��9��3��?<���Q{M��������#�ǌ�'q�g䁊j]�,~r/�kp�]~�*HX�A�sV�c^gxIkp�ϸ�VsM��+�f��:S��(�Q��:��Ʒ�3��al0xO'����Ć��P�g7~$E|�_e�w��\�A�%����UE��R͏�U�^+W�t��$7x7*u?�t��H�ޠ�f�
]�#.�SR�R�@qj��f4}��fڗ�8l?9��ŝ���ה��r��C�.�SЫ����f��V��K��mԙ��ɭŰVɹ����@tx��Q?z�ouhd�݈�J��~�ă���
�XԤ�C?�z�B,h�9|�|}+C�g�L�1&;��'��j�Tq��of���l]��py�{��ev�>�m��8�o� ��'����ծz���'��5`g��ѕi�6YN�ޔ��4�t�8f1wL���CT�V��%��b� �N�m1cY�}����>*�09e�x�vS�&�9Wh� ��BE(�L��.y��ʒ�4�(|�g����9L�Y(E�9����t��A�\��Z���ogyO6?����yth٦K�U�a!�P���AX����o���յU��UL�u�/�W5C�ߐ����9�8�:vf[F7���V�ꨯ��3l�q�[����A�����m,k�ʑ��Q��CBE�p�B^�Q!�Tt�-dIK�He3�dn��,�붪�b�r����Ϟ&����Z��縯jfX%���^���J�e�U�9#�i�+`����kLS�'�D	=�&�~A���2��ı_�ꮹjI<\������`f�ܾ�m�-gc���ynǅęB����W��B߭�ծ���|�j˺���/�4u��ǷKu����v�^�&K�-�m�oo���SA�'��aB?m�e����(ݝlV����k���sG�к�@ ����7?���Cn��҃��KI�r��,�a�������#�w#�?Fi̶�_JYxI���ӄ[0[�Gڍp�=����ZS� 4���`w���%�^͍QM�H/�xK*a�%�)����^F���	8�'���Ŗq�MÚO��U���"㘇�W|䋘YIM긜1�
�hr>m��v�)���n��''EcI���������r�Ӏ��%r�96��q7�ZVh\V�(�)z3���)���P+y]�6�u�X�ɪs!]�������S�� mD�0��WV9v�& ��)��pԌ�W��1�tKA'l��
�m�{�{(��������5�$?�j���z�	5�v1��`��t诼��xơ�K��s����9�5���gZ�B?x�OG:p�uޙoO��(,��XR����5��"۫�����C��G�(�伇-/�衺y^e�S��
��:���@֦�@�T���R�A�y���P�%m�B��Dq�9D=Ν<M�>Bo���f�;�������`�Ѷ�A��k�`�PUc��^g��<�c}RM�)�0��;����>p������b=�%K��Ȧx��D[쮚��L6��!��w0�/Xj���Y+]y�êoo��ڵ�����FC�11n~k�`��n�<���7
��w�%���I�㊤qfS��c���؀֖qMB��0r�V�)�N��/h0�EW��U�ԇ�yS3���rTރb��Ҍ3SI�E���[f���}�hv��K��Z�ӾܧYY|knF�y��[��O?��v��aI�c�H2��v��o��j�|(,���
5�,�m�7�S�q���(s�.�M���!'9JmӴ�n]3�q2�$���O6�Az^���x�(�������6%u�
m|�qS��m��_��;p~W��Z����K�%(�D���\8�\�"B��E����=��t:�C!!��U��)g���* �_�8%5K�h���sX[9��+��,��y˲��" ���Ks�f1o�Yꀞ��,�\�Ֆ��,�7�\��Z�"���4h�PPy��]�U��~;��]�)۶G��V<Oz��K�j݋�&���B]���.�X��|���y�x��i�a3փ'�D��!�$vhCkÑwt�@k6d���fàAj�j�yV�^GD!%)��sT%Ũ�N�hI?쨌��i,��Iش�q���� �B	:x2D�)Y�Ѡ���2

�q2��˸�kr"�^O�--j���0�"wx"s]��
晆�tP��1ُ������T��ػ����������.��Rk�$��G�Ϟh�:P�l�Q:!YԚ1��S���'��=�ӱ�C�CVP�x�˗���D^�rhјM�݌5S�VX��x.^qZ�.�hM��jm��<:��4�<�E'�ң���v��G���[3>�{Z��������:�י�W����2����c�3��.dc_`����0��c	_A�T�D^�\�~��9j�o�k����ϡ�5���#+Z�o��/3�D�I�^��,�^Ԃ0U���M��z�T�eU�����4.����� �{����:o�����X�/��j�͔�d�Ly\J\N�Ny�㬐�8)F��Y������7��;�R�}Z�,�R�12�Ŵ�B&��E!���<��ۣ�<4�O�X�5u5}�'#�]�t*��(�qQH�������
��&.5#����}�Qu1$�����wEZ�Y�)<R���x��܌}�Wa�K�/	z�]��ZnMf�Ԭ!������jl��P��,��F�.���2��T�i0�kU��V�&b��o4�/I�C�j�a�p�7 {����SW�fEl}���3��Ih��o�<;�j*1��ȃ-�M5��晎��\��<�	lħ8N����+n,�Nu�J#�Fџ�����Ֆ;\kގ$T�$~�K�z�%�f�{`ey����UquZ{��3[�Y�5*S4~�^�F�k%��Fb=+R">*ր�_Ube��Ơ�Hh`3t�y�G�i�
�m�t�Ả�`���i��N��7�aO-����(N���`'>1�i����1�b�ؐ�,2� q��o�إ��|v>@�b|��Tٳ�F������W��H��G�b�'��f��"7h���e-����4�>#�Za���E�ʱ@)����0��1�ΖT �-�����[Ǝrnk���3�j�*r��E���vE��ɗ������j�]���[؃Y^�����]���T�C����)���}�mu�wyl)�4�З>�"���.Cl�
�����O�( ���W�2("&���8��ޯk�_F�A��
ߑI�g5����%��yo��׽(�6Q��C��;S���x=ݼ/H��;�@5��*q� �Ca@йE�KK���2��	���*|�a�3��o�GĎ>��Ћu�tNB�6jn����(���ɒ }��gߣO?��e	�y]Z�_)���_G���z�-��Bb�+��f��HX��I�5^YP�����բo^��������?�ݛ����!ף�vk����b�	�:�X�&��|���<���H7�*_�
�@eU��w�� ��!�1���J�mJ�a&"9�fʩʘa=� ��ZbK�����f�᥎��l�a�iw͢RE�������n�9�ckP��?�Z4��@��R?K&��"�S07��b�T��O��y�c_>��L��_pC2��˺���j�5��ߠ7�4`��Y8�ƶ+%���]�.$	ߣղ�X_UҞ�P.ו$0���u��"5?�Sk|ǉ/���vy���a���TP�T�r��b���������ЦC�=��@]��B�qUz�/Ц�3eIմ<p��,0mh�g��� b�`��]:�ll��YK��l���=�sf��FJ���b��(��LY���YE�
Cy#k�0�0N�g�@Ι��J�Vz�A&-�{�P\1"�=Y�h��ꦂ���L"��iM�a	��;�4R�3Iv*���Y�)N��^����C�]̈#��ck����QH�~���Z~�/��"µ�����GU� +�eJ���T��yqg�A8-d2:�WU����YQ��Pnn1fRFVc\�&�|K@�m�W���K#h���Ϩe�QTD�<��@��h+��C��O$i�M�S��$��V(����XP!�^�޾k���8��%��(����8�	C�&E�u Ե��A��@M%�Ui��`H�A�\������A�Ú�K�K4@�Mޝ �]����y�ӧ<j5.Z~�������
h/���:��8�~B�r�#�=�:k�,�4�O�L�JK�X�ػ�>
�̎��6>�1�H��������:�9������E�p�P kT�p�w��sz�2?��;E59+�X�;��m�l��m���a&ib���
]W<Be�?l�>�y$P��(G-��5'7��3Z�S���J�N�JΕu�ϛh��\�^v���hf�!T��o���E�UV���Rz1�8ȝ�����-��B�4c�5���g�ଙ�-�y��	7��I'5+n����B���G��3w�͕��~׺���[M�K�kE�&����}r\i���kJ��6*��O���d6�!��5E��F� _�Lh��Y�U;l�*���\8���9���Ө����V��0����XY@i�` Zrm�|Z���A!��UU}jXoZ�W��U}�ąVbe�o��rl�	
q ���r@h��)NS���o�'A,��?��,��5U������(��?�:�u:`������C*[c���D9*��~���9ʭ��Wt^30y��x�ypz��v
���L���2[,��V}Jse&{�	gH�D��bi�;pՙ�B���a�|z�
I��t�JD���D�5F��V�0F�-�b�"��_T��;<��T�i�n�.��k'�Xc2XC�P�4Ld����(���A��4xM�n�'����n|����{w�CLr��X��I_]��o�
d��g����������3����y�����c
)�辂��.<�d���>e��0�q���m������KnG2}�an/L��`_���˕|��W�-�a�ф��T��+�K޶�{[!Os�{��ޔ\��e�|�E7�%�D�W��F\]�p=���Kd����Ix9��Nt��"1���Vo��H�xx�����ѻ�������`"|b�` >�Xdd�<nI-���+���v��f�ɤ�9�Wɫ'$��dx�zdk#@�M�8�nV�\l�����:	��c΀T�	�)=[�6]�nʦ�=x�pZZ�����m
��m茻\��|�^"��CS�r@�w��w��.J�mրˠP�37r/����:WQ�9���S��4DSv�r��bsy��7��|�y8=k��P��6ύ�KO��G?����{ϜG���*$%�L+@�KC=�t"���5��^i
_a*襊^��+Z�5���k����������F^�d.�l�����'x��R�	@�nс\���uG��!�A���j��ߓă����CԿo��@�q�Z(u��PO������`�޿xh]�K@�Q�hM�?��w7Pļ^}�f%����|O�;9>�NEp�'1:�-�@��`�Ä�ޜO}�(x����Z����)��e4H>rr�1��2�`�p�3��}1������
������U�?�~J�#�! ���#��F8�89��#����+�[�i�����m�|n8�z���P���~�Z|�Yu*��?�ӛ|��o�V���A�wf��+O]��W��gKQ������1��ds�RS*ח�������X��e&�7�%LTE�
0��|�ڸnDwBsj��.����B34�p�m���$��`�����]�}��z���S�_쾗flҍF��ͪ`R��Q�d�t#��dz����`S�6 j~������E����S�ض?x�L�<���{�ͧ����h�3YU��̧	/�eBTS�-waA�(�e�A���<Dע"r�a2/��2�a#�'��u��ߠ���M� �eE+��h�Ae���|��,i�w���U�|��O^�MEs&ƱPG���`�6x��I��/�� 7v/9P�c¡ AɒR�H���<��W�>S2�ǘ�e̾`aKy�+	������o�?�)L�iL�8,::�j�r����c��C$���U鑡�o^���L�҉&�h��	ɚ�DƷ���3k�k�
j��M�`;�]|��s>+���ENG���)c��BA��oc�+��ܜslu�H�/+��9#��duK�[t�r�%zh�P}�͚�N���˿|�;����ڎv����F��5]ڡ1Vg�n9���E1�	b��h�*��"�&z�&>�j��Dϋ:�S������	��TD�sen��7S�2E7v��e�e@����Px^Ә��~9}��vj^�t����<�&i������l�}��"G1�ͿOydj��ڻ-?joώ�]�N���ϗ^���q�>��g�m����}�w�#3V��Ӵ�M���C��ߓ<F�#�G�x��{��!��AJ������ܽ�Gm�N�89p����넌9K�U_=�J�8L̂�K�ReԹ�UG�#��w ����qp�:�������j�'˯����4J�3jA�U�rRz���6S|yJ.�Ɣn����X��A!<�F�)W�ƦB���p�9��q��ze��aZ��?�(��0�=,�3"pϟWDD�'������%C�XFK�-�L~[��Σ#~���;a�5HFQ����G���%��P`~������:)��s�U���|���]9=�Q1:et��nÜ����sy��r�	/ĥu�by@�Q���F�|�`F��"Ɋm�w�=��D�ET�/{�]���i��;���u����Uh�b&����U<�_@����.�r1HE5+�c#Y�"�b/A�K���+���'��1H���~4�h�^X��0�D�@��'2�d�=��u*<S�>ڪ�V�a*��b%�+�](>g�oA#��isB</�ݼ�m{<k��[�7���s	�!�2򛸭�
y�`��O�S�C��~�4�hU�X�E�(���B
)>��J���5�O��p���d�O �zB���q����U\f��hQ�����I�����bg�=D�>DǮ��M�c7�r�r�Q(/n:!up��B{8+M=�R��v
���H&B���(�"���S���QH7�qL#]7߅��R}g��d�T�.I$�5trk"Y޾D�v��LdX��A��T{�o�*pc���2;�,l���6��F���x^��$�]��/�%����`M���6W���^��R��M��.�<��J;{aE�������"�ڒ�:'���Z�t��߅sv������J����p>�A�(dR��-Y1Jo��F-��F�r����b��z7ӊ8�Z��衔ZS�Eb�0~ ,���-!1�
U3�qYX3C�NlC?�0��N{���r'Vᩦ\Y/���;h"\�չ ����piG��e�'�/���B�\��1V�"Vl�*ӂ���0�����q��Š��V�m�
v�0��+p�� ���=m�M����>�n�o���8��k{�r��H�d ����bi�9tջ��S�TZH�3���6��n�P��4
�z�e��R���
��kLZ3V:)��j��n�G��w�*��;�<��iw�+����b�g��wO�K�^��Qާ��mOO��jףWN� ��,��)��bG��3-���NZ�������M;c�2~3�<H�2G��\Ѭ���n:�&�N������XŻ�T�(-`��mz��F��*�X�/��7�d����h�N��}
��QA"	�!��1S�C�ʳ�������Mz����{#�1�rSg����O��/����������$�c�piP4�K��n����2/A"�G�5|]�YW6�cQN�|#�7�5/cՇ-��*&�=4eM�u���r{UB�����:�e�@=V汄-KԻ�O�lA�wU���Б��c�i$�
��C��Y|9¬USj���L�T7R�6Ue$�ύ���~�/s��4�o����ug��{,�sr�sؒ=6���Y�X�X}���h���v���«<�uAq�'�fm����b/�ݪ�3д_�p'hGʔ7|y�y�;��wQs����L�q��ouA0��rۭB�eY�^*�hS�p$�q����g�ut5Rk���L̴���3��
�_a k��,0��-p��u������>r1ܕ�`k��c�E+�$H7�c�0�$�װ+�^�3��(6XZ:�6&�B��!F�C�	f]�e՟��٥�tj[_��[9�'��b��!d�'0n/�����z��eh�S����r�mx���jR�r;n�K�����F�%ק��M����lG"\"�n����o?l�H��IT��qnT( ҭ"�lop�D�|Wlp]R�}0�
��)���� T���6�f7^{����B�g��@����!Fy��{�U+m4џZ���
��pt�g�;����ٌ�m]�C:�I�Ȍ�J6P��b�G���p�!?��f� � D����Q���׬0j���i/Ҡ{��t�}�����M*��)���h�1;��Ğ�>$_�����07��΁CvM�$�g� �RG-�_��ʆO��X72ek��~I�9�p�HlV��ݗ��K)]��Y�4�NÁ'#>�5d=��k�38l7_��M�zw,������A��q�����VV�X�i�gG̦ W	�|�:ӟ��FP�!�5��I�b�W)~M����w�g��}�"9"-h:֞v��r���wD�_SvB,�~�����w�e�/�4�ޒA��`s�����-�д}���ny���Z���:iBM�}��"�"��yWh�Ƌ*�������{c��.4���Y9"`87ȚW�����o<�[�����a���%w��&/2�۹u��EmR�޽�|��"4��C�( ��V�*��K(LS���F��q⒐]����x�RbFb��zA�k��0�<�h�)��u ���	������i*j'�[I�E(´V~��1gy�Nߥ����:|��:����SⓨOߑ�²D�|�ay�|98��{0Jq
,�������!t>�@�FLO%UO�L���4����G�mí~���:Rf���|������E
�f�Q�T庻͢�Vmb��z��q�A��N���ȣm��5�	�]�d�l�P<s�EK�G]�������b:�i|����"�|�Q��>�GX�M~�M����v&��j�%�V�����R!{>.[!C6�e`d2F��Q�U<w��@�����hF�hTJl���w���<�U���4;7��^}3�oA����a�,�cܾ���PN0K��9���Mvʆ��#�>B�W�ߎ��|��=�~.R	���Q��+�������A��p��b�m���Y3Z��,�jk�kM���� �'�����9�h�5�l�-�����!D\�I�|Y���:�T#��Կ����!��!����L	�������v���[`z,�ӯ&��u��߼�BN���JZ"d���UW�g�G��|���zU��)+.".�T,�߽)��ms:Z�o�����|�;i���z��9�o�:NOݙ�f���������|m���Hk�
S�E��k��r(�tW���ً"�`QqT�0�(�O�+��7�N�ϩ�	��B���2X�o����W��ϻ:�p1��7/���� �n9�����U�Fй�g�����v�hF5N��l����Æ/l۟����-�G��~��">[�$�js�x�I�����2��+J�؛�i�`H�}�
�F	C[(3�ٵ�����r���`���[n����͸�ʇ�I'u	�NRt�&H��3mWpL���8���}ں��Jm���t�������`_'ڠ�2�[��\f!q���1�|ƥ�Q���mUʍ>��의��>�T�Y�)Y�ǫ8��FϨFO"��٭����yԆb�;c�O��d���.��qS[�W?nzx]���i|����k�T��VFO	�f���&��_�a�/�C�U��Gl'c�ϋ��=KXfdf���#�}#��#�,�2��nX�8=[?���=�=5��q9�cd�����O��ͤ�I��n�N��=�U)�S�(�/��0O��
�;�����lK�\�$���0�G�ܟ;�#�.L�<t��A;ƾ���j66%*��Z�WبiU��aI|�$����O#c+����1�9���|����YZ�ּhT�b�0��[˩�e�<t[�3Sv��<����<0L��6���i3���С�R����r��t�5�˱��%��\����|�N�ݑ �Oy�;t�Y��R��k`v�m�X1xW�����2��׻_�ؚT��8�F�I�� c�j"a君.���Ѝ�u��D��� ʶ,(t�����K��\Z8xN����]�#�����8�����T�YA�	M�K2�6UtF->S�ܟ�0T&��Q��aQ}��?
!��")��J��1t#! )�1�Cw�H3t���ޟ��{�����\����u��kg����W��c5��s�p�&���6�kQ�s���&�*��l�eG�C/+��a��dѶ�s�1����� ��[k+t�R&`Fh�,^��UϷ�xJ@�MR�o��3_�vm.�+&�^�V�:���h����c�b��8�1��ݶ4�M��^��dce��o��֜o�H�=Dd�+~�X���e���+�`���҇�@��;�����p��S���Ջ��S���d�Z���p�C�)���`H�5��r�L���!?.~�u���Ղ��S;�A�[��3���f�h�[
��^D"��Laft��k�һ}���8��[��^57s�ag�H�v_sx
�Rz2'���g�D���_9�����B7��.F�D���Ly��k���֘Q�{��Y���<�FU���5JL��%�C�q̩!����^��\�~�4��A:���K�V)��!)������Y��t�&��3I��5z�;8��hO��--ba�;���&����^��<]�V���|]B:��;���?yI<��!f8|Hu���A��::U�6>0BN��4��$d�bL�n�zپrѭ�Q�Պ�v���)��c�˾\�-�����$�o�tV�r��|���U.�k��^�
F4����9��(�5�V��V��|�i���G�b���Ex�JsaT�t�C�\f��~�E[�huB�a��е*'��74y4^����5(ߨT�h믟��e7k2��(�����"�FT;�j�f�{����?�?E��L�L�u�?Z�y��71�ƾ|d-ה=�{��֘ٳ��ܕ��w���,�!R+�b��lrG�N� iXPV,���q���R�4y��FL�(5f̇�;~�e�$��{�:������e�s�nȮr�x!<W��Vu�h�)��Ċ��y�Qr`��^�/�Ƈq���Y�	�D40�L�Ř�`��^�A��cL���o��<p�W� ����m���o�γ���+�Y��N	$��t^�E�T�Ht�zر�����2���ԗ�Bfb�ߥ m
�_�^�Ki���ʜܧ�R���*gcϬ,`�Ȩ
�Q�Z �/	;������cgTHL���5��f�}��a��H&Ә�e�k$U��c�=�\ǆ����Y�����o�V�OL>�]u�J��X���Yi�+pwD�#M�&��!�n�&_zVM��>-l�����+똘��C�M�=:����f�*����]����s��W%=p{lX��ǹ���[Z+��G��vڧ4>�Sm���m���p����rһ�(i���E�?u�
��l/f�� ��V��Ğ��l�w�6N���g��T��I6)�ӡ�5�Y�/F��QbiQs�b��c0oϴ2ߦb��./.C^��O,hx���Yz֯�����)/p"�}��=��lb8��wyspzh�|�'�lΠF<kF�o:~���j����".������������� �����W��v��$�Z��V�k&v$�ڦ���Us`���v��ev`��dy���av�aa���mE|S��mom��+��2P�1Qw����{ N����ɯ��-ߵ�ܭ)�y$M��r�7��w�~�T�5�����ƛ����USj)�
�'�V�u�?�n�k�!y˹n���S��X�)�W���{�m����]:����0�t�<O'
�^���n�LlbS7UɎg�QI,�ܿ����Y�	����A����c_�]ʽ\ʈ˞p�{.is4A�m�q]!wS����2�cթ|���6#c%`���X����mir����U�:�ng�T�Y</��xU��r)�g0nDx�0:ZC�H/�^-�|�?Ó�"N��-�"��M$/5�쇋��\V�ߥzp���4}�hG�����12����ؘm��d\,�͒�CJ}ˣY8;1whoL={�C_'ȟ��XZ�n�K3�!d8h���x;8P�ZOJ�<e!_�b�����h�ɟ�=�I�­����;�bd��i��2�v�z�ϓ�z�ߵ��A�ؤ"��-�ډD�pP
d�Iu���� �ܞW�2<��P��Pê�D�oc�n��Kb�/���D����`�O�k�o5:�N��f��u���[�갃�Xaͯ&��@�7"w�9d9�B	b����4����V֏vg����3-!��!5� C�#Ѯ�<;㉙���.��'s������qZ�`�管�C���}������O��w/`�G��)8O��U��ߗlCa��+I��1������]���\���>��0sm��%�}h�3�Fݔ�������3�&#�$X�:����3��?{T��&��Ʉ$��᳹ȼ��"$��;�V�A���_�*���8���A�'A�F  �rk�Բ܍S�/�6<�m�]��G��E�\�4�pň�����w}��i	��o�����I��n�,�d3)G'�o%�N�Us�TU���}�����:O�i�*��Oڼ��*O�|����rԖ��z�)�U�(žOLM��F)sc��Ii�S�e���E��`p��~����mz����,��";����1m��}��}��c�G\	�Ʈ��\���"%U�mx$�ͮ[}z+�Qt*2����?�D'.)?��dvx��$�Ǎ���*��kȻ���ֹ��x�4�Y����e�#��>K�,A�?���7<�`x�*��\8L`���%o]�,��optg{
�MR��p�Wjb�QVh��9�8v���f����E~&��xy;�@?�N<��+���[���&����L=�{�������ʦ�3$�Y���>�^߻������Yg9
�C��R��=�s��>�Hן����Y&���C}�<�0��^ϾDx�6���bQ0�f�}9q1{��h����2;ug�B0TN8:� c�}�`�����(�;��!T!4	~�?ِ�N/�.���Ű�=||,z`���G"6�N����W'�_�ɟ��ofEV��;LD}My'w*��(b�?4�/eNŲ��ſV*^NY6ۯ�1;a6�5bdU������N�a.��%���{|��^#�F��6��������|�E�N~p��p׳����)<o�����پ��6��)�}�^�Ύ�nm=S��)��VTƮ���b��C�so)i��;���
��'S�޿1�.�wȹ6"����|�M'�o�N����TA�fZ�eD�c@+y;��j���6[KĿV�ފv|R��<��"���i~|�����z�)K7myD�+�cEʚ�@%� ҎCt�[���[4�mzS�H���?[�����̕0w��]��݃����Eg� Һ�nǉźr��R3��s�����|*�n�����O�E�����3O��f�V�T母!ʤ}��J=U�w�Á����T�bQ9#���r��r�5MՁ�a�n�s��l��@�R9�5JP��]>��i&E��?+f?�T�
�nx��ږ��oh�����V��
��]�S��%�V�S�m+�Sn�3C�u�Y*�'�nf;Gi��{��W��oN�O)��*덄�%�_��^vG5���hf��6��;�Օ	)˺�v�M��=��S�c��*w{7_��0zs�ԯ���|��;��D�A�a��Dq��#J`���;�H��U��S�q�Ď��]����aT/�dg�/��:���uE�Is�����m�gԨ�"�9�wz��+}_�՟�����s<Ԕ�(��(5�T�'��IM�Zѷ��N	g�8ªq2�`�`L��&�?�a��M��)�=1�hl����[�pi��ӛ�6����o�.�ˤ�/aI������'!�ļ��ZZ@�3d��LI�͂K̦�B1h���G���K7��iK���R��َ�2��)S"����'��wzd�!�������� L� �C�����+�b�#�UJ�M<��"�9%ҐiݥАQ����"3�'�(�Q|��5������Pkm�ȶ�|�v�;1:����(SL&<V����Y�k%ԟL�ݼ?a����oCƃ��'f>�5��_Ij��:*���̶8r��="e������dg�0aDj҇xo>��q�i�^A����kL��/r~�%�����ߘ#�M��sT�MBX�C�Y}�Gym.��I�|[=M,7}�Hk�E�ql_)�Q��GX��;�rz��0�p�i�旦&Yì{�܉�x!��A!8*��=A �����?*�u��j�,����J�:��Y'�nXbɏ��X�4���ӑسyxs,*-�m/16��F����c��J���͊��Ug�������of�h�a�3(��VWC˲�����c�A�oK���s���&K�J�yp�� G.�c�Z��v�T�7f���F^�G�V"���P�k�&7���3KnG�O&~�^�ٿ�RvfM������-��M�hP]�%�K�()#�B��g�_�	�G�B΍�@Q��]+X$BJ�/�d��6�`�ϙ4���
Z�T&���'���F�,��G�\�n�����!�1�~)%��nBa2��
�q������������խ�7�b_+�c?��;EN����а��N�%�*%��C&�o������M���Hd��
���hOwd���#ذ����f�N:�+V��C���i�K�wr@%�������ݺ���÷O�m�]ws!��q\TF ��Ær@�B�P{\����E��
�J�@��&VɄk*��9��� Σ}߿)��7��~Z8�qoXƴf$d����d�~q�`:�'C��=�?G�B� M��7z|�;��<z���Ӓ8w� ��GkmݻS��uiT���a�y�����m�Ϋ�o���'W!ΝwW�Ϋ]՟���ٶOPκZ,n�.�d�-$P�?�G��'�����GaV��n~�X2�?�� :���rRڞ��gm�?�:?iZr�T�}�7�n�P?��YssU
=�Zz �,zf��E�E�G�+���<�X����E{K#��#Bo��W�+jL!�>�)jv%����y!߳AgN�C4���M2�?�ȏ��n�
��EBA��!)x��Ţ�{_/'׏0��]6RY5�b��(U���m�xفݡI#�������M�8u�.��ʅ�@	%G�ĕ�d���蔚�<���Ȝ����|��T����X�Y��!�O焼�S�nR1�P2�7�]VE�Q��Svh
|��q�ط�����N9���<���q-�^%�a�2'�.����K�׳�m=�a��jCl�55��$�\Ȅ׿�r��������A�Ui�]��$�$hi���M=�K�jnv0��W7����m�hLA"�P�øY��֤u��K��Ř��
�t6�S5_vȕ�鰢pZdȿe��W�l%VG 8��?����
p��?Qo���v��ס�L`"��n��/��MU�y��޷�C�A�5��-�5V)1��,x���sO(�T��$���tx����"V09꯮~8����h�O��E���P@o������S���7H�c�Pc"��_����ɝ�΍
�}]Д�M����� `6�\O�!H�����8�l]�~����	�B��ې��Yڼe�)��?J��R���0�#�2v��8�i�W	�aDLKw!=�T5��K����2ͺ#N�Q�"%j>d�_eovN�O�W���8o�}T�[kR��e�L�7��7*�E������}�"��l$��;:�΢G�ň������JP��
����dmvb�5!�;��8j5l��ݻ���uÔR@ߨ}��Iluy��9}m���Λ�YZ�8ʟtZ�:�?�^AQ6QHy/�$���G�"�R[�2G��ϮH���:�������3G"��NLS�E�ߗx�n��7y���'-W���j�_��؋6-�|z�� �<-�\G�<��8�}�3l�p�X�80	�rvX�B��BT���tS�6�ƕ�U��!|����h��Z=W)��ٞ+��s֘;Uq���
ݗO��G|a�5&�+�{\M�꫟�MH�M_Mф/�,h�5�)Q?�s	����x}�0s������q%�x=7�9b)�����sSq4�=f���I���ޗSϷ��R1+ԣv�b��,Y�:Ixh/ş[&u�5{����N���בU�hۗJO���0[sRW�IĔ#���y{��2�]=�C���u=�J����KC$|10Ku��{W�����!1����/�zf4���gS9���
��e�;p��[��|��^W� G0��|���n}t�p?��v�;��E+�^)��q���/���x�8dyyɴ��hRg�U����J1����a\����J�������j"��6`������mˎ�i����֬��	�W��ۊ�R�m4q@�-���Ȋ��v�P�g؛�/lr`.�ئXN']���)�R����)�sv��+��jJ���SB���ds���%.
����l�h,�=]������J��X�Ke���V��iκ��y	a�"ф#`��.�	�4���엔'ցRl���'i�a�\����!��6Ft�=D��y�����ϟ<�3�jKn��*�;Y1q��r���$e5L�AQ��!Y�*6�D���&}� o[:̣i�r�ހ%e��4�4Q��t#��ԄLK���OK���
�Q���v�8���v}&�Ur]�g x<,]ש6�+�ϣ�t���)5Ϳ�[�P��N�^6iX�D�ﳌ�]�O����`+�>*Y�oMJ�=J`-�Z�E�e;���c��6L�^��;X�?�6	<�?���=O�K����ĽHs3T6A]��������,��c���Z�&��[�)���4<Y�M_Ӫ��)������OO��Uܠ'��"M0���`kȖQfIˈ��G|�`�ۍ��P�����e�z��N��8��RGO�M��z$�xdY@��P�H����&�n-z�NEs�ɀ�&�Ҏ��_3f�1�~���|s���ݮ��`^ЕI����{l�_���[�� ��f,��al�d9�wwt��9n��Ӄ:G�g��n������Q� ξo�[/Uڵ:~|�̧�rg�y�^��/x�֭m��=+�5(����?�Mf.��=V�yu�R>������P�%7�r�GRԐ+t$�W!vc���;�+����hh8��"���$�8$
nή9�|8J��L�D���F.�6��.X��)����<�*�i`�C㥩n� ���UFt���̶��pI��*j<w��jP�<*�I?�Om�d���j������w�v
�:6uԆͱ��r�L$��N6E��G�������}�=O�s5��|W��!���U����,��d������` ]\�p8��C �m���f7���nN���Sڷ�P�s��I�g�Ȳ�r�t�!��g���l��c��o�ֽ�+��~t�m��]z����<��F�C��I�o��o7���=����lU���`O�`���.�H�� ԭ�*\93Y7�`s���PtQ�^됤DUެ�rm`����p̒55�!8��L9�i�Pr�Up���nt��[g��U��_�狼���W�J���^���qC��v�����z�%�T�pt�a�U$.&`n٤߂���7����22��c���uǦjGg��ps�x��;���!����9�c�l�s.4��+�V>�h74]�:wE<:�"�S���@�p`�)�O�M~��C�Cd��y�~���)�j)�N�zX*V0�U �u\��k!�$fD�<�==�8#�tRߔy�e<�����C(���Poc��v�O٧��h�8��M�Boqp�7���`,��+��2|��y���yn�mlb<���jI�e��cw_�`_aʋ��rZ&Eٙ�(���|N��UD���Ao�N�l�?
����Z�t��R�H��=���T�7nN)�&!�_�x���f��C�?��Pz�k�N�g})�>x�"���k5
�p�-�%�}�A��j��88n�-n0��f�WB��W�z�=��J8���ڟɢ�����<�k�s�l�*,��xk�0�߀�_�I�����g�qBBH�}�00��'�V��G��?c�ϊ̥�dr�KT��p6G�6M���0Ӥ��nx�3�J@�m߹#r0�����Ş.�s�ͼB�Z�i������
H�r����3�L+�A`�黆B)ęr����z����%ʭ������	:�F�!��b ~Y��~�$�y&� ��y{ _�Jq���@3�΍\x�i�e�$��W�3�n� �=1*�����c���MQ�0INQ�[w�jp�}Bxz�1}s��0�|���l����c�g�6����rћ�\(���Y��)J�-,K?�᯶�Ntzo�����;z-"�y^㹙zA/�,�����U��S�	�볲�
�[�D�u�v���E��4����#ggσ�s�5mk�+<E�4�M�G{sb:����'�\[M�5�V^˭vW���a��p���ʠE$o�W�����7�r�F� ����m�:���_*C(=�%7�[.��괆7�׫�b�T�&K<�3�[��
���/����N>�>ݛ}��K�bW��WIL��v�x���c��q���� �/�9����ļ����������vn��v��ԛ�.�3Q��9,j���i,j�i�/F%�;���~c�}a/3��	��s��yyg�q���N.��>(z�CH��[���}�އ7Ev��";Vx4r��ɫ������|t�:"	c��t���欩��\������<�r�۱mE�k���l�b�--\D��j�?*9����Pk�d_o�3X�/3�l��$Դj,�e���/"����LŒ�?	��U���e���|���5A�\���h�I:�P�C,��u�\O6���`�[(��|ӈ��IW'5�7���ݗ��6A��KI���bS��8�ӫ,+Gn�T�ů>w��~���,Z�ο{_"��OhO�*�Z`Y�Ir���B�FR�Y��;?�����hP��}
N�Љ7)��Տ���!L+ �BMt.8������>��+~k.����x;f�C����a	��5�(p���S�F20[�z�n@����M׃7K��6�=Uɛq��ؖĦLP��\'�}�݈B� �p.�x2�hV�΃��j�愈$�Vqή(�X�6���!X�c[��j�ڶ��P�������=����I�K�����j@�)��bdq��bMdS�KI3l1�L.��P�-+YP��0��	�J�Q�U-�b)<"�{����7���7�3��}��W��e��e��� �=�V�]a�!���.��t.��-��+��S��I̴i�)q�AV}[��3�K�J�Kϳ��[���Ev�6���}�6���iM�Uv����������Hk��ac��i��+�N�~�!
|�Ć�A�dZ�P�!i�
6]����6�7�4Y��&oI�ct#H�p�
�S����\�g	)�rgVk�:F%�������sReK4N����	S)7�jM�����n�)Jt5}���r����yw��q\��C3@x�����~e���` ��x�1�8b�Ŕ,��7���zI�t�e����N���,WAX��;��A*A���c�[�[PP��idfB�揀�5ڢ_�����jv6��ۙ����Ik|���4g�c7�t����;���6��,�֟�&�-?�G����Q��O@���5��.�# N�ϗ'�J�&Z$_O�$�J.��A��Ά��a;��:��}�^Ͷ��(�yJaa'1�~�Pg�������F^��j_G+�)L�ן���!��l����z'���Z�
���X�ȖzPg�KIw�}_Vw�E�bV�T�+��1��F�mFz=�0����q��3lAk����e����63�4A�9�\����tEM��X�kj�ĸ�|�Ik��e�S_,���S�?Ah;k�,��Ҫ�\��ez2ez�o8����C*����V�K�KZ�Ͷ�A'�R��y e�C����*LD�/Z����Bs��}_	{̇������H��.����7����1��Q��5E!��PTs��O�)'b���V��º߳��wW�������iZ�x{}�V@y���`1��w�LH�Ux���>�������خ��X��əw[zO��!�R�4TS��?����c�z����v-0���=H�o���^��pܘ+*���&����=<�k?�����\bi`�K�%R��9�e*�|�^��Y��̓��v��	�����C�-�p)�鶅VF+�Ⱥ���������ƚ"�u����r� �3.���&���&�k��KL�%��T.��>�������_��� Ya�4��_�9�%��C8�� V�z����s���H��$Px�6���0T�hgIY�Sq���,��sB�:R*j�O��o�:7��c�U�o�����/w�A������������D�2��WNu���#}t=��<�@ǿ��	��������w\O�~i��oO����pY��.k�jL�`�������GL�ORA�[��l������D���~���`ߐ8�x2UȞ4FR.����\Dz!�pN���"�F0D�h��5�6����^c�4t T����n���^"��� X�X�yAx��Gc���s��N����2i>�6��x�kxSWp�)�u�����K���',��±�Ƴ��uR�崛�~i2��`p���J�X
�?Yd,������!��Rt7O�c很��#7���IW3�#pd�9�poh^8��$p��J&&�g&P��9Т��S���Mk�o��p�Z�݉�.��|�>�i�e�ljt��50I�(-*�ձ4`s/�j�>�z�lc"p���ȁ;�,�![��=<�'�)������u?�)*w�a.�=�Q�8{4^��_=�ӶvK�P�ek�Av���uz��.9>`8�DF�*pb�ߋ��o�3������ϋ���΅�n�-���e�`��7'?	ڷ/����P���mVM��M#�ǚJ+�:�[4���,Z}�ٜoE�O��nbr��l6�iʎ�G���^���[xQ�7��,>En�,N�f6w�����{*y%�U�j�m�)����͞h����V�{�ռ��P[m��o,k�N������ӭ�џ�'��ϯ��n�zWu�\�r���ޮ��J�6�o�XXZ=��8�-.�gu��"�r��H:��q�y�b%�TU��S�ep�╙V��bWF�Gء��w��۫�^'�<R~�F֭o7l����U���O�R��{T��|�kM9�b�3LA���c���T�k�㤈������@��%GD��F�Ѥ���S�mf5W�$��^B���$4��N�=pC"���٥?3��
O'Be��Ai�OX��|%R	�Q�H��Θ���M���g�㕿�g{�y'jc��Ř�u(���@�}�'�p��J�f(\��cf���Wb�u�� �ya���O��4]s>�����P�r9h2/$�:�p�]a�A���ѩL�.$� #5��5���;�s8�7���N�jn�2R�!�B�j�vT���ɬ��^� ~j�`5��e(� Oi�.���|y��v)���
�%�.V7T���
A�����'��Ū]H�1t��zuS��pd�|��,��+D�k�N�`��n]��V�L�/�����@~��5����G}!���5�gU|r�\r�ExD<	>�ȅ����d�Ǒ�S��.����]��u�/]�G�[ːj\Y�E6����&�ĝ���V����H+v���9�O��������J��C��SqĦ2��V�bϿ���پX_�Ú�Y����Ed::,����P���D�@,kOY��ۆ:�)�p���1-�Ow6�?Y�-���\v�X��~Ҷ��r�_�]I�Ӹ�����]�?��Q�G�0�y�v����Џl?I�s@�]�p[I�iE������T�N����%c�[<����O��EI5|F�(�8��ڪ�� �J�,K4)2u~�-��4ד�E<^T�NN,���rs�p����=�h��>6s��&j)5rA3)����2x�BD�����yǡ�5d����k$� �ޗ��Ѵ��N�F3m�>��X�(Rw�q'�5N��}����.�����Rn��	fl<u~p/i���	s�|��p�z؛Kn�?6w?9ȴ��s4��W��y�6��a��>���c懖�<���܂<��'҄y{S�NL� +U7�`p�,�X	�T�RN��n����[���C�Q�Įg�j��a`��������sky�Gc<}�
��+|�a�2h׸s9w�n�D���y�Rˬ����vFi���X`%���,���*���f6�1TfŖ3� Ԍ�m�u����#N#!;b�$$�M�<#Z,�	�5����g�e�e'~�U��Jr�pRS�7��R�}}��l�=�1圢s�0Ix��\�rS�bY�77��"����ܰ`U!CEf���\J�n�M阀�nA����8�aq��F�� -��.+���u])�d�k��3q��u��0LN��q��9m�;ӂ�h�}-D��&���F���h6��5��]\�3�aZB��o���I.��NoiBPP����ee������)ƛ)��w��%�{r�Lݼ煷R��^�q�q�����L�ږɾ��E���/ߘNm�SQK�J�/UV�M�	���_e�z~c�T[�j���պ��2�<�O���V��E-�B%9_̾`�4�%�̼�2�V[m�G1��ϕ�u�q� 3��R4E1�Ռ������V�jS���q)�p*�Q�w<1�޷}<��wz���L�qRd��b� -U�����E����A�n��J��Z��Ø��e-н���?���I�=sk����cx
=�ċf�8k��ۺ4�Ӟ�Eȯ��_�f�t�����쀝L�ٺ�U7��������$r@R'���W�>n��+V2:^��|Q<�Z"�6cD}�b\rҔ��{8Q�C����������#U�R�w]�3��<���Y���c���}�!��
E����@���������l�+ߨ��Ә߷�æ���͑��G{bTD�����r�����'����r�xr4H���t�[�G����7~�o�B2�,	��J1>���U�sP(�� ����XĖ���XP`���F� ��\�a�Vq&��`�fOR�q�L�[�j<8ѳ������Q���7^N�zgs��R�̥����4|/�<�=+!�޽������Mb��x��C*�*���@91IGARk-���2I;&(�M򶊷��0'��	�i)j,U<�g�j�OD)�_��A�\؃�����S3t�0����=L��ñ��kŝe�:�{��+�Dh�$��V��e�t�/{w=��^�z�t���~�ဃ�?�J6���Ӯ���'���Rt��2@�ߗ2��r�����g�N�g���1�H���N ��E���i�FgOo���)Kk,�	��1/���y��^��]���p�7��&��X�{cp���}�~R������oYn)|���)D�Q�~���q[�/���r���Q�JD��NX	�6%,��ӄ��$����űb�1�<�/S��z$a�u�� ��`���~�%ae@ �9�S������'�F�P����X �LM<��f\/w{+����K�x=`�j`�C2ɽ�?�4P��CX��"�FO�&,���zTp�=79�f|���-�6����������B�~-�%��#1>X/>���G��u|�F z�?���n �$��?��>��J�b)m:�fъ�<E�6l_M7q���ɉҵa:ϗrtz��![�r�50V�:��@�T��b~�0�M<��iJ�}���rs�0��k��Q
���[EC�Kȥ�j5k�]��ɾ������?m�	� ���&3��\i��Xا�*��
c�1lE��n]Ogf��Ԇ�3
.��Zm���<K��xܠlk��8����N,i����Q
�o1�C�E��dqg:�9������΅�l�Kn��~dp?Oc*_?-������=f���P���q��s�q�{���ը�۪��^	|tR�Y�����X��m'c�*� l9�x�i�-�!i��Ū/�m�yL�kh� �_��,y�|Ψ`�Y��~%Y;�YX�e�0�l�����Ӭk����W(X�ћ�򕍺f�/��	���eZ�T����z~y&]���M���R������C�]�%Ɠ��K�	#T�L�6��(V��m=�]���I(��u:˱;�1;�b�j���D�b�N`�C��uᜢ,Β�k$�X�#�09�8��s�'�����������䩸�튈"6���lLP�-Ѡ������=�OU���S�|02 �«��FBK��vBAqS`��/�?�BGd�ʠ3���+� �2��Xna�5��� 7���;�����.�k��6���&��>��!X���gc(s{�1Ǉ��/�cV�����Y�x��i�7pUn������ZJ�E��ӭ��O+��-u��2��/�sh0�7&{�r�qf��=�a �^iXQHYfݝ�)��":�稧hk�L�~�aym�"�i�APn2Ci�/@���)0�x'O��;���cf��?\�%P3�Wd<���HdOEf8c��"[Ps	�Bk��r�Af�\T�B��Gb����?�y��*�QSB5�a�>h����1`ը����6U����#�궨������2�O|kO���i���P���̡4��V��� �昆����g�H!+AG�!!Mxy��q��ԅ���0�xRH<_j]:��r(�2��?ZH�R7�������'�
��Ż����Ed�I�Q����E�@�)�Sy�Ɠ^�@D`^C7,�q�Hz���ƞ=K�4�TF	���_1����w�E����j"Ot��N�9����;^&� is4������VEfF�֬�,X��'��D��Ό��o�<�th9ƹ�Pp9	z;��OW�Vu�ɦ�tUx��p�+����omj٠x���p�h��x�4����T.�D���$�̑]��R��avX�֧x�M�'!�'��V6k�Yr"�F~M�H��
����i�>�y��fE�j��o~��h���a���^�E���������ʒ�h�wdjZ3f+>X��V��g��ŀ�:v�I��t2F��r�k$��C9�)�ӱ�¾�v%�e$�&�iQ䢌X ]!�G>\^Z](@g��"K�Hlr1Lj>���r�}%�+Ѧ�:q���jQ*�s�wČ��"��&m��ҋe�q=�C1�[8��ʾ�2�*�Χ�Fl(��0��j�G��`~Kt��������:W?�>��'4An��N|lͦ���+�?o�Y�����I�/��#\W�<9�ox�)��0<���>˷z����m%�f�B�ɤ��l&�b ��?VC�Z�9���{�'I5
-�'ՙ.B_��rݫsyn�v�2{��Ƀ��	nL���-�Wơ'�j��H{�?���"r����B�f��a(W��d9!ɧ͸g��C<F�<��R@?�!C�b�A�Az���Τ�t���A����
��s�ǣ�\C�ǝL��8#��)�Z��+X�����+z-���I� %�,����<��p�X>��YB�� ��'���XS�6;����6�>b���IB��[�1
h�Jk�^������"D܁����|�d�����(�ٰ�a�n�D�qH�.ۅC��2�t�9�2#��آt7#ڒ'Ɋ0LZ�وS�jh��	����nP�{������#�^	���^ل��f!m�VlB $x�k��n�����	?�d����i��ߋ~W�������	v;������h�u�]�ܑiZ.kB]̳e��ҴDm��.//f�g�����W�s�
�v���m�iҠ���("Lȡˤ��$qƤ&l��&+����>�=��Z�Z60�7xx��]��� �z5��y�	T�$=�̒	e��s�Rl9�,y>��NY9�_���ޙ-�h�&\j�Xm�	��[�ԉ���=۽��'��~��\�N>A3᫏�&�&��$n�7�V�/����i����,��3����zI��ԏ��ĨՉ�� ����F\��&�1�`{Z�u�*�й'���W[ɛ�&<&�8�� Ï);�o��x{�����j����c�b���!w��eS>�r�ׂ����øs��Q������c�"byzNlX���ǁ&'̢��MgU��m)��sH)ia�������A���n�n$%��n���|���5���u�����羗��t,��Ò��VVZ�__�6t�8_^����3^+t�$�ɡ
���N��Є(�o�#����?Nz�eq����=�_��My���L3τ�U��b��������X��j�[�S��RC�9��؛+�!P$�I��ߺ=>����Iۗ�;� �ƅ��)��xw��AC����(b�Đ�J�w�%]l�j�)�1�<�ք��b"���(�f0��^�E�L�:�Fi
��N"$')����PO@�,�ff#Xql�՜�N 7!�W  �a_�Þ:��J��n[x�@m*1�U��iɝs�+�`��pQ҅y%O![���rg
B|��`У@-��	�p�.�cZ�x�Z�:����rQ���T��[�M-L̻��tAZ�m����z�]`�p�p�T���v��~wzp3���x�xDBϞ�#P��̠<���1��{m�V;�ފ\�<b\��ؒj�_@XK�Ϊ�{ �0.����>�,.ay�ݚ�he��$5S�6�N�H��0g0��P�AOYrT��j���x6� �˓�f�� �ˑW3噢"�+�n4I
j̿Omz�����c�yK'�k1��H�SaG
����U�t8`NuR9I��e����41���k5�-��-z�g;���H��C�X�HwӚ���c����i������@�^b�k_�9�73���|��6�������t<,�.��ߪƽr<�i�q�%�e��}��7���p;_KƮX����D��x����nH����礍�×�L�6\��Q5�t�pe1jU#k�TU\P-"6�?�inY��5�aPRR۫��9�."%��t�>��z�������.V��m�����t r�����ܦ�-�[��Q�P|��?��i��]�"
$O߇���%���)MeŤE��ߡ+$0򂁼Z�f#��R�\*�j��?�S�EVlslp )�,�E#&I�O�P�<�hRm8;���4�
�I�55�/�1�-�8i��D�a�J�_�m.n����O��
�+��O�.��d�^n�ʖ��{Ry�N������~Gp�B��/`{����3�������9_���(���A}n���|j[In�S;�=�Z=ZyV�ʞ��l�8}0�@��*����l�b� ���MbNҌ��=���z���Fr��
)_�	����B�l�g��λPcW�Y*�4��`u��D�Z�ާ��g�ٍ"��^TF���vo�퐂*dG��%��ZS%��Z)���E�s�&|a&�?�����ʍ�ia_��L��^�=s�����rF��5���v����Vp�)�i�,�5�j]mm_a�ś�ca���q��SX,�\�&6%�������UgjmgG���������΋̶�̮��Ih'������s��Z.`K��.���ݨj�鬓 �ꧬ�A�}9*�X��9%1E�*�٠�^;np/���TМI>U�*�����.��e���/E�����1&���0�����{�}e|'o_����������p.��/�_I��Z|��Z�J��u߀�=�tS:u9�BЬ+�/��b���c.k�#t1t|g�	��*���>��.��e���[�Y�9���VV俽Cc����6 ,>��!T��v6 >��^��l��h�a�F���(��՘��t>U
�������3�]�	V�Z��(�h/To
Fl�t�kh%'W���@(.'�b�V���5�c�y9�N	So�-���tf�n?����A�[��;��sQʹo��h�yFv��hF���e�6q�������B����r��-Fe�kۙ���M���TQ��	�~�����!�J�|���Ҕ7���_��{Ϻ�u)�N�6��K����|$NFդ[�E�g�F[����[@3s��s���%�!��69(���Y[+��{T�� $�+.�=!�.�0�fDn�[�0�81�2�V"R�$�����S�� ��(ZT7���U&13`�Ti��Zz ]���\���γc]!�/m��XQ�`��ϡ���;�������g�X3Y�1��ǯ��鬧0���Wu~\�o�"��I��o�y���r����ٸL������Rsב��3�t2���Y��xepڰr7������"ె��r�������ճ<����r�so4a�bɜu�p��O���G��u�L���<���S�x�E�d�h^Ӱ#�y5>2��@��OiǇ	RV���&# ��5%�z�WK܎+B׻�{�Y�^�]��ʎ]+���j.f-���_��@ۛ��DE[딺�~��*,_��#��o!�y�L,yg�$�����_a�1�k#��@��m5�J��]�UB��Ҿ����i�`��>��/{�����Z�w���re�+���/�Z̻!M!�U�����uT�9w������א��*�6�q�VH��]������		2�;�?���`Ӕ���8x{-��������'�x��+ [�L��O�}!H�$�vq�Ę�Ä���6�:t3?�7B�z3Hһ�`4�rs�9:�!)���1���1�[�VM�wc���~�N3�}��'2�,��>`�M��!�v�K�b�}[�w���<#��J<�8����0��ͽn���������..Xr��#�kj+<q�kσ��o<��zX�[%�r������;֑�OɵT��{Ak��0)�yx�ø�Q�]l�PC�k�E�����<������,��������久�Kz�������NH�:��
kR��r��������tܵ�-DT>}��!�d��z�]d��#q��C��c�f;$c����u��f$9��b"9� l�L�t�\�����i���Ƭ$�[r�I8�HXhc���<ջ��vK#���i�pCc?R���_�Q[J���U:��-ҽ2fq��n�ν�h��#��{'�WF���2"#�>Yq�`��+ͯ�N��?|��tiE�M(�����M^M�#U���\�����ME?O��w*�u{<�x*��Oq1�o����=�Qy��~���|�����a�_���7�{�R}��DpM<w<M��*|[n�B�G��wYb.s���=��:�US�~���jZ�J��t���Rtb˼��g��X�"Z)e����gnVtj��*=
G�0B�.t~�\��V���h9�r���?��([����6��v�����^9�����l�_j:#8���ذ��s<���<̈́�{Xe�(�w���������~�6���vs�2x^W�!#zb�$�c=N_)aB��T��.Qx*H���D�i]����������
y��?c��v�3��ݫi��"�9N=�Ɯ�6D���ֆ�!F�:Ra)��{���"k�u��\��m�M��^8V6�(�T@�	Q�H��Xe����sÍ��4�/���$ī��u~ϻu������81�q�Z�Oz�݇,�����A;���oo��B]i쓏uwpJ=����Xݳ���V��K�F��ǳ ��PW�@�^AB�j,S����ؓ�s���C�����%d�
�9qm���G��o���_� �ˡ�0��֌��ek\q	��<'�t�E��b���<�/��r�(l��,UTB��=�6��rR_�$����RqL��Q�v�R�p���.zә}]�y����+"��J�:Ge����\۶��˸�� #?2�s�r7��I���	�� �&'#;����u�m�?��5���s��q���Hs,��S�;��s5�)�o�ȱ�3� �K��X����&����ɇ�3-���_�V}$��Y��� ��*r�K��W�{�Yif*��R��|
�u΀��RI�@fl:ܫl�5?p$�JL���w��:3����>�;�ޝ�y��]��WZiz\=��������f]4eh˲�S6x�q�XCx�N�z�����^�
Gغ ����'����^~A�`�i ��z��kQ�9������Y@����G�m���^����&6�NZ�G���|q��Nf��n58|l�?r\i���ge��jv�7Xg�(��l��S�պYi�w�L��u2�II ��ϡB�D��RHy��.��g���m(b?�o?�E�Z��`Q�� �B��d���b�N_ˍ^Khe�z2���FdW�*�o s��!��X��ca�zar��̆���k�eW�:�y��;{����k�8ffr�F��y���
_���~�V�oh��z�/�j�+ϴ�.�\X�u�P�M��Fou ��������5�\����ӑe%k ��W���߇u���`>6��Ny/�e����"�iq5�l3��7N
[ N��.�,d,�n'Y��{4��[]�iXn
�ڰe��/ �v/ߗ��2������� �"�ŴWIj-�Z���kȋ6)ߍ�R: ���o[>�j���u1������������)wp!9;�D9��?�H�QS���80Tr6˘��r:Q�� (���r�7�2~����v�>�a�(�)�+\H-�q�Q��O�e�RP�l��xaGc%�|P��{���p����R4���݃�&�b���oЕ����~ 򷤓o�q�Q�_��>ǎ����i�k� �Ӈ��!5��^��Z�zL�iV����e�+�����j��B���UyWXzqI�x�U���h�Ab�9�����HK(�ͦ4;4�Q��[Sv�
�+$Q�\<�j���L��\4>�Xy+m���a������+��:�J���h�P6��\����ژ�R"�3y��mTG�˰�l�(Ю-�����A8N�؋��(�+k1��2���l}����/(�${F���B5$���Le[���� !ms���T5Zk�}J�>.��
��N6^ѽ��+��/�*���%q|aj�?1M���L�u/�Bޒ\]��@�CW�In�M+qVs�姍A�L8�HA�؏����L�m�FE�6��@��B:m�)NAl)��u|�ªw�� jZ[޻���%�����{oќ6i\�e�cg�ii�<��J�{4�x̤xy��uu��e��j��݂�c�5������%��X��m]4�̓��	���F�Oy<BIS�Cnbe���^�N�.�h�yy�:����8�sj�s��4?&z�L6~��s�Bq��u�Z�I�E�����=OHϡ(��~EYH����4H|)��(D��-�_�E}ґ���4�LKc�c��
U���hܩ��.�����0�eZ���)�����i!�\��́{�ܰP�:���W����0;~���@%�^iF�u�]�	�E�(����g_�?p�����䠘wcP^^Z|
-�갤8Z:�,�-�jb�T
H�.M����3@d:j�~熸ի��f����+�]B������Y:R��b�ƕW<�q�k����u��43@]���sx6�7��Jj,�g�����W�������9@�y0�@*�h`�)�/2�z
@���2
�_r�.�$/��h��D�q�x�z��`���){�;}M3bUؐ�	��=��H�{u~J�(Ȼ�z�W;�wn:�%��~����wz�{�L��=R�G�ҧR��=��*a:o��1/x��U*H!O���v�euz�K�������{z�WʓFZ@t�n�Y��w��Yp:��dߢ���b�ZPj�t썭���#�ּ��h؏�}O���OG+��OцO��+��#|�+���W[�)���zd��3�|!g�C�Ty#���4�я�ׂ�(U0��9��Ѕ��
^�ǵ�͇,93#�'��H/ ��q����j�ͯ��&�^����oO��������m�OK��Mg��׎s|S$�s��6P�*hC���\���u�[z��t�HI�B�#ޭ������`�S��S��ԎbIt(�`p9w�ϽHec0�p[KV��+)+��=��A	f��ts���K^�}=߈�U_���m���?Q
�����s��.2v��'�h&@*������J������pp���ŧZK�9?W���O}�ۀ�5��ƐF
@�f<(Z��2t<�� �f$W��f"���D��r(N��ҹ[� j�}��>⮣!��:d��10ig���?�=�{.{?�u��8d�:�";�:���+je߈lh���e�?h����A'���,��m8�M�q�X��3���N�{�<Pg̯�ciGa�=�
m���9o68xyv�i�覃��&r���뜹�4�Yf08��8��&!��o�����@�Ark�:_�����[�.O��9�\�=����Tp��O�r}��J�x�����[�@�q���M�M�n���+3ڋ�(���J{��W��W��'��}p҂|�[n�w��>f3���������`���B�X�rm��*<|���0�&1`�𑌕S[�@��?(��P���EHy�8����k0H��h�iFf]u���04o�ha���{�a�HgU}���d�S/�M��5)f�A?�{�n�z�3u6cq�;$�0��AV(~�_���7�0����8�v�H��D�O(��]@LđKGd\�{�~T�U�p���8(9<��<[�S���7�r�)�<y���\	l�t�.�,L��f�*�	~���A/���1��EE�Zz��`�`Y	&L�f�H��bw�{oXf���/���c[ٷ�v ��1\���)��Z��n�T�8͊���Ix��*��-�� ��l�9����|W��0L��<4|T�`O˚��j����2�u�w�[^�pש�x}�������ˆ����@����tr���ſ�_L2)�k��{�������؝��M��"kȭ?��?[��c�M�CgBt{b���I��_B.:'�f�JUT�5糹E�rkp+Y����qkh��e���IÏ�+UF�O�WS�ЎOF��5��-�Ysu�X���.���e;@]A�pǹ9P��n�KM��9pN���,p�bT��'��^B>�m��0��MϏ"W�� �m��7.q��<�wܓZ�%	ikV	nP�r�].Z�R�%p�=Qa���g2Ck�skq�gޝH��{>_l�G�c#?��(�o�6�A������4I�op��S\���c�@W�Ԕy�jHB��#�ۧ��eD�$���|5�7K�E��1���J���,mU����K#�70=��bru��`�B��h*��ޛ�i����>�.��E����/�,�.Wz�/����~ �1���ًW�T�	?,A�Z�?;�0�g\�S��d�N>Vƛ,�,z36>��$k���i�����'����_�/a�0��O�Kn����gj�}Y�W��'+��"���ُK��Jm���7}�$��zG������;A����&�bF�����ئ�[�
���t���v!��עH�����*uΘu��pcs����=�o������u!B���k!��0	���f��
р�kQ�2+^�$���d������8}l{��஧���j�+�t4ᐞ��)f�8t3�	N�����+tb�-��!qt�I\��=���UBF��P��8RР��o9=�kA���t&�&�7� CiLO�%�kC_33�]�/����e(ei	T�y;�(,<��
��TfK=��ɪ�a��|�X�`N?`Υ}���dVͫl�m�:ê��Z^P_�k��YE(J����ր�	V����1�$���F�ŨG�l�|�[EkeC!nM�ƶ9��H�$�;����M�騟.;�#M�K�_p{��I��s�y9��⳽[���BZp�ԡ�c8��}�w���Dr*&���<���2���U&��I�Wu�-���lK��hqT]��M�� ][��uEr%5��U�L��Z�����$8����U=�Ζ#�6��!ޝqVH"����Ò��}�Wsy4��LSŇ�����1�7͓�o��������M_���CF����م��eb�]݋�`�1,:�.*�T�WhS��Bbup�w_Ұ�s��~�iM��w0J}�8�Hk���4.8��.o� �߱^�̢M�gE�Ӹ�g`����BM���il�Ϧ1�>�p�It��Q)7�:vQq��iyV���*n�,5�i�Z�!��u��ʹQ�jg��E������Xw���=uD��&��s@d�ϡqᢘߜ܍W�]da֏N�Q��(�N�W;�3�d6�t�TE
��0�]V����_E�l/����tP�����o��d�
�ж�-s�������T���Yl\��->�ڸ����'�Q�:�Q?3�]�ػ@����<����Ykܹ�|C�~#�#�E]I���r�w�������;�\����V��
	5/�ͥ��YZ��ԛ�iXng��0R�p��P�����F�e�*7�T�i8}�&,��+t��0�����x�����/4[�a�U��X�z�Ց0?���%�z���x�O�Ee����;~T:e|��Hb�m �<Z��s7O){�O4��ȈI��R�F�؃��*Y�f��~K;
,����r���^�����}͠z�'C ?M��<2R��������x�Ӯ��������������V
詈,��Wo7���1���Ҟo{U�y�H'�X��[�w	�Nx�Xe�/ ib��`�*�ٽ��\%5�F"? <�����0Nv=���ⓄS=^+��VkK@}F â�iQ���u���t���u�+/[�4��3�87�]����p�
�Z	��*nC�݃�@tV�~s�Ԛ�����8�q��<.� C�n����>��=�Q/���T��;K1v�)��G%�b��ԤWJqnt#�@�7�{K�A��g����p6����ð�B�n`�v�%���୶�F�*{U�|���TEqe�*�hc���|�|�a�¾��J���H��.p��NWC'G��̅u�1{D��.	��
r,E��>�Ъ��� 3�P����J���o��-�i\���OO]Fln�8������)ᔚ8/�pg
Ll�HLf��пR��~�`V<Jʿ�\����T;�ѻz���q��'�o�z�92�)�pk�t&3S�������ox/�[A���>�}/��8Z���ǯ7ܲ��M�Y�	�Ӈ߈�T��s�>�'�zxd�и�ךC�tl��K�`�r����e�,�<����Sw�����+��#D��.�g�����S�U�鵆䈵�t�D����;&8�g^���;��{���#� ���	;��a�
��+|�
�o�H|��\�V/��'O9�D��G���N	P�^Z��kNߕ��xm?l�[�6�B��-	cܘ���9��N̓L�S;��aK)�OK�;	�?.2�e�"4��n�%��6�7N���͟�J����2��� )ૢ�Y6���B��A��~W�!�U�R��b�S���'�Q5">�CS?ڱ�_��E-U�h�y\���	�x�mAm�S,5,��ꤕ4UA�`��ۭW�.h������p�B�M|�K��(%x>�p������k��N F}�V���R��U[��pN�O������l����Q�鼲�mCx�|�Xp�M+�*u�F��M��)C�DiE�����.2��13�o@ˆ��#�2����]�%)���Y��5�m�L��#j�ً���22<D��U��V�|�*o{(�'���әp�ٓd��Z!O<�`��Ob!I�-���X��Ƅ�Y/�d�|����b�IT��o���]��s<]���Zc��ǼmRu��������P:����F�/�MDN7=�,R]S�d����^�1�wPﯺ}>��K�|j_?���fb����[��a��� �
ɧQ��f�\a����GqMe�q�}�>�(HۦӔC(!g VsE��a�Wh������l�f����X�α��E��_��E�.����B��T�r��W`�?[��r�n=�[�gxa�q5rɗ�K�xSf�孆��槠s��ׯ�����i�~vQO�h�|�����g��P������#I���~��v),:�z��R&�`y�ˏ��[��R�h��u�S7�i�����/TD�Z�K17U��[BS���hs��Q����ڋ���� -��Ը��a��o�T�d�O������7�b: ^��L�"�%��M@���C84}P���A/$<Ț�h�:�ȁx��b!1�m��M�j\l�����`"�����:g(܂-���C��PV���y^��3D�3�����Dq����f��,R��BC.����X.�.�r�wmUʪ�UC�f�$8��]�ߒNh�������`6)� 0�tH��͇A��$�?��q����gr�7�/Or8�x����"cD�h��;�{!���C�w@G#���e[Az�O����R�$`3	y��PBGpH���2(Jƾ��ΦF�?7��˛,sz��Î�B�����{5�����m.&����I���&C՗��@M���������o5cޱJ@{�Ŝ�U1F���wp�j�BN0z5��g>��"4U���/�$��K��$����6�b��X���Gɽ;�Y�<?��]�h�+�Ma$�)��&Z��N����*
�N*I�~
8�;HOw�wh;��^�h�۰M����Y�=|�Eo'��=ߩ�J��w�Z��_��U�d��Rԅ/�
'�z��AX�%��=�Sx?�6�3�KcD�Қ��K�瘲�o��Y5<k�T搲�_�=���[ʉ�BG���K��W�ѻ����OG+~�Ev�E���]]�Y�y��1(mӒS����s8�����3�FJ�.���"r@. �zK	^㧚G�\U@��U�����'oc�q�Qh���j����CA޹z.��i��_��M�3��o�d�y� ��a*&[��Q-��m�݆�Q+�e�Bs>�V�2�&���dl���	7WHm�G��6�?F!"8��C����ғ��=���V�:QT�8S����n�	6�U�&	���%�֕��P��B���8�X�>zxl\^���NQ*�Ԃd|���h��_�θ;�1
(j���NB1 ���Z�ߨn�E�D���P�Xë��y!�:~�Y���5p�xCH��!�\m��Q���1c`�o���XL��3L9���C���n���a�#�� y�U>�mn�^��# �:h��/�V\�u�'�n����.Xێ$���ح�ΐ	�����	���>�N��y�D���B����z;Gi�{�6a�O]z�'��+���!�ғr��dNsL% �%\�$���3E�|Y����kF"�O�������I����o>�������p�*���]������<�C��z�3=���mHa]UE��cM�q9'����i񾕔y~�*�� ���u���O�F���[��w��Ye4�.a�i�W��m9�8 �Q1I���|-o�즅�);���Sd	y�K��M��B���?e@2^/�]�K$J0���|MF�fڒ�,���������9��bQ���WV����˦�˷�>mf�G�?��́�ڼW���:����h)�K��>�B�����,3=E���M��umWiWT���N<q�jQ>� 6�嫁���3YyH�7,�|��.U�)ɲz2s�x)�<�x���j#n��H��]�d:D6[a���1�Ʃ̕t��9<SK?�xK6�[�7���|"�� ����v!���I�L��D]��y7w�Wx��yF8q���_��툋/����!7"�V�5Q! D*<ۇ�UL��/����0H�H:ym��$�@��¥� S��������>���^r��'��S34E�;�	UA�rT�b!�Ē$�z9)��$/=���s3�g+�@�qkjV��� �@a2�D�w1wש�u�[jp ��_�� ��C:���[w�������n�?p���Uu3�/ĸ�c�ȓ�,��;t�{r��y�qc����w?eG"���jx�uHU��[��Ӑ����8'�Mw�@	��ǰ����
Ͻ��-�lٮI�`p%�uPrt�j%�����ԥAT�5i	nb@���J߸�B_�u�}*67NA�PYX�$;!(B�b��6�lb������M{H�L�1��B'8���J���$�+���CBp	>I�%��&臲��o+f9v�%��*^�c�~27�9|�yv��/:��݌�uj�̪D���m��q�{��A�>�4��_�_��n��/�ߧ^��Eh*| �*�]'�\.T�����eҜ���H+�{�E4Y�i�� �`k1�t�*��z�nt0��21F��%\������ۏ����ev������Nf�6]�Yȳ��\��J_H�k��S;�i����1R�I�XZ�� �r!K�)^ɻj{���8YBr�`c���%>��j��E��6m��_9�GF
��MM�P1�0ʭok:�:�c�o��!��Z,(����(߯��8�5+����Ҙ�+�g|�wt_ز{Oz7�<t,��GB����w�f��;�J|�XT��k���ܲ,��HYF�ʈ�������b���u�Ԇ�4�J����"5� ����bȓ
�AVyR��K����8H=+����U"����<Kk9�D�������v���X��2E9S)�ºyx�-�
x�O����+��Wk/�U|34����bU�����N�����B��N�-�i-�������e����`?�T�s�c�P���[<�uW��T�d��'�u��$�R��{H������\-��ܻ�}�=֭���t����
�ͦ���
��������?+�]S�:�z|���4�������<��Iѐм��� K�FE����&n�����ҳx�,��S���E�\&��B��nq*J�(�tY�
_�c*z��&ᜯ��N�@�R��E�MY`�p���zӄ}�(��eT�Y���[�>)��H<��TG�^u���ǀ��b��Ţ���ꑎa-��>����Z�y��ֳ����/�������0{�U�L��L�S�:�#��1Eޙ�����C��^�N�cά�ʻ`e�������srs?Q2��*��W��: ��+m��
.���Ʒ�\i͍.���m���R��e�	�^H��K�����M5��֥�a �{�q}k�Ypr�A{;^�� ���@-��_ʂ5uN���W,+��N��)�[l���BX�z3�:�cp���F߻I�1�v��õ���T~�J^V��g���N]Ѷ&�h���B��M��!�,�tR�_:ux��㢘q�Ou��u,L|���j-ě��n	0��׼��Z����s� ��̹��)����GuxO��8,k#�:U�-k���s6,<�Vޭ���F�M���P����"�=��)�(�r%�ĝ�h������d��;?��<�&_"�C�qu#��8d��R�������b�a�sKa!�+�x�ۃ��H)����!ᲱL��i�u�_0��&���}t��m��\P[s"���9#b.�����G�'�:�uc"������a"����z��8yC���U��Hg�VA����w��� ����rYA�/�R-�f���ZofM�K_��Kc���20lA�H�d���Q�?4�?#����7řWHE\�Lz?g���!�4IF 0��M4"�L	�wW��jH#:�:�f>w�{��C.�g&��'ᯱ�h�V1]~T�){OApT�߯Ź�okڡ�!�:e�P��p0��C�v1�+d��jz��`~��h�M@ͯ[�Pp�����h+�������\��*�Ñ���9��(� ���|�53?���Q"Ā�X�9��v���G�h����J�)���( cJa%�ҙ�`^�H����R��|���c��$z����l��������v�u���L��̽�7�X�//�;J)̍��[�ĂH��W=��~�G�ƍ��E���o .s��Y�W(�ƦB@+ʌ���D̾��.��ܔ-�SQA��ߣ@JO�����R+�RZ�� ՟Z��H���7Mo��N�M{����戾t/
n��	�[E$�ұj))��v�:7�D xAƱ�/��Pu���v�ڑt�+�a$���V�R�E[���@��z��x �<���ݨ��ͪ��Ir�)4�q�+���ij^mk:��tݺ����d���٠v �;����y�|\][�0V	}֏TW���b0_�X���a�g�6_�;���,�a¯'���"�5۪K� ds��ψ�l�Gϡ'����
q�/��5d�؋�.Z�@t~�/Rb���Hb�J�X�6�+)H��I._K�Eu/��J:��.!�`IM5��H��
-�KL��5F&�V�D�=����X�ĕ�d/��5̸�����s��޾�=�2�3�k�[�ڗ���TD�!pj� ]�&eXR��җ�tV a�ٗJ�nĞf7�|��Fv�P�)#RD0Xי��VɅ��=�n%���d�	;���Cgwb�Vz�^U<����LWw~EUt�n����6�y���������4YB�nB1W���CDO��]�S֮F���:ʦ_����&�e��;�%�����_i���.�@m�7 0��ܷ�UW����O�
T2����}���D��u�����x��7`��}���k#/�t�t�gh���lz|>�6.�/��H`���'�̪�[6��zF�UE|/2�q�8P�]S�|����/��ڐM����7j���^��B�-�-uB3LjI�ܳEYk�F!5����b��J����{j.ݢ�qy$�L�zo����JL<k��n>|S���(�n�ϹR�7��a�h�����P�^�wQn��B&=�E�YH�w׹�~߫Ԓ߷�0�J�'/�TŤ�dZ��8�ֻ�Iú֒���|�&��U�m��)�V�_��>8��'�&6��[��a����GȞ1��8� zO�YIC~�i0r���tY��Z�n�M/b�D`G����[D�YO5�����fg
�a��nƛ�C�F�tD6��M�Ǆ��#���#$d�L�S���?H$�ʚ)��F��}-;D}&t��D
P�'�%S��p�T�\������33�tͪ3��R^9[��Ar� �ҥU��@u�o�Sdܘ����I�ߞ�/�imw)�0�k�P�Φ�q�,�x�3Mg�V�n�[�ǖ����Y�%~4��J�j1��2ѭ]��	tV��*�셆P�s1\9�؞��9Q�D*����c��R�!ny�{�SJ�q�4
}���� B<.���OU���(�U�� V�)?����I�7�� ��xq���*��+�r�$��	��U�f�]�6L���
���u�w@�z0��2�r���}_�xl�/�m�~w�w���tNW����|��l��M��x��
Q����~"��C�w�� d*3��~R�`m]u]�/��Hs�H����ްxS,�c{����������Ǎ!Ǉq�����W�
��CJ2�v��%��9�-�4�#"�\LG
���ث��#n�86�R�~_�m�^t�2�B�ǲ@�"q�L��(C�=[t��H��Y�	'��(?��R]^$��[B��@����dr�ϋ��ĳ��G�͡���DQ���F�$k��_�?�8��
^�^�B�la!�Ѿ�u���O]ޱ��Ds��~�<�-�)��_�#��J\�Km�M�x���.^��$��	i�eSȨu�6�ȣ�_�&_F��"�M�[�%�5�X33QY㮚t.Z�K�V:�JcK~c���% ��<��>�5L���r��o���g�����	�TCz�~��l��χ������ɯՇ�6^�H���q��+��-aJ�pQ�M�w���.3��&I��Pĳ�����T��(P��c���;䇳]��O��R
:,�o� ����U�U����"&���a����78�v�
oWfig�\D�+grno�UM������Y��1�M��I�qL��I�WP"��|bĢ�V��_���rR��\�jHuYK	+b�|]\�p�Y��XZO&�_̿X�'Ή2R�s��!�H��n�2m\.V>m����Rp�~&�+�U�3��yӟp*��Hp�2#��I�dl�
d����g�����b��c�����7�]��P:�`��1:��z��1�G�>7��*݃o�����AH�ȽdɅ$QE�.�!)T%�]��W�8�wE!�+;&���Ɲ�#�as�@�"�qx_Sќ&���#x�!��6ow�����HJ� 5"����ؙ�3Q�� ��4/�ړ��[����^��4��0����rhdho?��W��v�PI��g9E�GB��׮�R�AQ-�>�������&ty�R��3.8x�8M1��������	�np]\'A��Bp������}� !8�,Npw	�Y<�!hp���޺�Uu���������6CI
�N��1�m�
�vg��7=�fW$�T���#�WkJ?����E�Xo��(_��~��E��~�����5�D�Aǽ2����B�U	��ՀY�)8�R:��V`�n�	��W�'�im��Fx֐��"����� �o�p�E�����a���'v�}<�����E�^�F�J/?҂`�,��x8���.�.�`�E���2�<6��(+)�*R�	,s ,�Ck�E�$�>��"��TOZ�*��z�yV=���B��d�i�q�x�D���@wJ����O'K�Z�j����U�)%+�����`�c�T���t7 ��� :�H�7kɄ]q��;��\���^�?
O��6��a͹'���Tb���\7�#��*���&\�@�w+$;ΕA�PZHTo61) >����,�6 �cΙ���E:ST=]^$w���h��;k&8�s@H����4�4��.9�O�4���[T�oٸ�p��c,�V��Z��"�]�@��3�l�f��N7�V�Y8�h�أ?�hTޭ (J8.�G��Fͳ����`�g#?Q9KA:�d��&Q�T���i�����"zf$`(�dxh#�m
5����*U��FNG���"��-ف�����{;��T5�5�+kN�@�3F�� ���gR0�?���N�D ��]D	�|X
��n��	\����Jh]Äu���!�Of�W���2|�׹�����w>��O;*T��+ߚ��.ʢ���� H4_�oG/�%Z%z��qX��_�D�vb�l��9��]������2��2ş$BA�������/
-��e]=���L�~J=��9#[H;�����{9��A�m�����{�&�AOѷ�ϛ�*���z�ή�w�cW+WԾ�U?>|6�̺n�!�n/�֟P�'�TМ��%S��sj�i,�?��`�fjW�k+'��.:��V���쉅��*��y��
��;}8)�X�ܒ����B<�F�>~/�"�9���D5��hy��j��t���\�٩A)��&tZ�N��re��q�}�Bw�=qk�_�[��Ա�Z`�L' �mf��j|�g|u�S@�m���|�g�'Vi�=�E��O|��)G(��3�~��å�G�/<��qXM�����A�ww1:.��ֳ�%�-{��W��-���1BXIT�B+��(�i����f��$��\��_���4�y���λ:�z՟z�B^~}�.�����a�Щd\��O���7�`�U��YBY�$�"�0���k�(p�2��iA��;���F�1Θ��D-�3v��]�~%H��.�$�����@R.���H��=�T����0KF"�7���]���3��N��XZ��-9�,^��L���>�@�_,I�G=���Q��I�5�� ��o��!W�YZ"Duh��^�u ������-�E��r�J?�_������`�����vJ����x�T��r�=���1n	�N)K�f�z�<a&J��VM�W3HJ���1�z�n�j&@�4�>���eK�0�o<�'2�G9����%��ل��fKaq����\�HV�Qm�{��,]�4�a ��F�"D�쥖�@�X�Dj�vErI��+�k���嗒�&��_i���cp���B�%�6���н�������͞�}��;T`Y�]��Ҁ����c'i�h��&�<�﷞n����bg�O!��P{pFCk���{x���v*�����%>Ö��Xقb.x�+� ܵ{=����#<z��T})yz��"�p�\�ja������%�RH`�ӎ������� B@�O��D[Q*'��_��#�8;�-Ɣƿ:1i�\��z?��]��g z��˅�9�z�̨̔�(�,�I#��e��]8�;��������&��Y�����)�0Νh(q���v�����ۥ���i�/�쯦�s�|�O��L��}��k'*�>�W���P=��#�K���BU`�3�V�H��²[��ý�
��6s�h��][���FWt���G]s�F+2��`��d31�FSC���5�N=
�����(�����o�!���t�}|$�OV�p�1���8�jQr�5̈A4�X�y�$^�Ua	��C�N���#����1s1�Y�%˥j�8I���ܪ6��^�������N���wؘ�\�N}�Y�`\��@��]|U��\5Jri^�����7���%��Gd	G�u�lmt�(U@o����y�L$�.����:'{D`�j8���`?��!V:���+w���i3j������Jn��jwȌ�G01��L�&�oV:V+����yJ0(����!�K��'>��V��$f�U�c)r5��l4�H|���$�&���!<�	m����ZYn�<���4�P)F����� ��o�܇�z�BtRR�o�L�2��3�yK$�ܴ�4�` c����>#�e����f���~��Z��7Z?x�fQlu�I$4qut��iSk�槔l5#t�`X�æZ3�V��(�Z�����X�������xq�5�	������� �*:v����c_o&T�DF�{�m�T#]4�����<ơm���U��!>L�&P?���pG�v����� `W�TF�~�#z����x����8��u�L��a��J�i���K,5H�Y���<a�d�I�/�\�R
в/��?z	���H�v�~�Z ���]� ����N v?�k��7��ۋ�)�x���t���86�׎~b[Vb`T�6��#��^�����s�(_,��O�=����w�۝�7-H$�CUZs8�x����.�oS�О?,���Y����c:�F{�4� <��ȵI����$�?���v�Z.�}N�Aya�Y-����1�8��l��=;�H�ɉ�]���2	�~�Z�3JLi�/���Z�RX���[_��vn@���=�g��dT� U��(�J2ҀZ�P�fQ��P��*�#X	�еT�7���f�I)�A�=�z�f���ԹOTY��V&�U�:T�=��ouI8���Q�[��`��De���R7s~���	�:�}��CA=�Z� 6�l��O���qbE�ESqNQz�!h�Լ�����Ĕ
�l����I��R�2O���z�����܊q�!�B�bw�I�?���.��z�9Z2�X'���@]QM3I�*��'E�M�a�_T�4�t�=�_��e6I��W1kk�a$��G���Gq^��	�32��&sf��o����'懪$?���z�t
���fsh�Ə]/�|�S���GGy�q�Z<K��� Wڮs^�"�]��X�+��.?��v����Z�7���&ת=��3��NI�̥��i�α��7g����3(^��Z���o*�Wx�(,r;7�&�4B%s���Ա��3a�t�tO��������\�
!�_����1ȇ�qܗh�8��	�1	|"���t�R]Te	x�e�������R���?�0y��G�:�զ݋Z}�8n|v������EҖ�y��~��j*}O���m!+���i��xE멕���`;�r�_#��m�Z�ϥ�:K���7����K�왱-Q�=�-��������nle�K��ev����PG�}�Q�������xu<N�6��.p�0���^/��ͦ�{�;���2���З(i�����~-SL�#^V\#9�������$G��2�I��h/iQ�W�`�\�����eC�(���'@�J's����oA]J8�B�Zb�%��DN�5��A�[��5PC��9p�M���>��bUE4o݉a����o�r�1�L�T��&I-�H���.��M#�z~¤J��ؗ�iL�j:�%"���֡��g����#�T������ �`KL�iv:%�^����y	�?d�d�Ev�Rw���+/�i[��T�=q�(�����+O���{��3O������88��n��]t�����Jv�~Z�"C﨤�������渍#F��!� �f��-��꯱3e�%�Ar�8w������� ��ꇶ�~�>"��+�v�����ڬ�8nfЂ�N�؄��f����}�.��
�5Cf�B^���$Z��1���9�G�%2<��yF���1Zǡ�����[>g�,�˹d��ӓ�m�Zv����SO���5���9����	����B�AZ���E£����&u��ϙ?�&5�*�y��A�_��FdM��'��Z�����V'�Mw��_�>�,3�_�r����$xϚ��.�W�3�Գ���~#+���P����zw�a��TX/��Q���E�k�u�k�:��&�vr��VK�[j�Oo����H��0�e)�I[3����1���Y���c�P�7��8�g��n����T�컦f��\F&߫�cx�n�Xe(�dA���'�/���-/�<�ɵ=g��M���)|�FK���;Y:�S��OkR�ϐH�d��y���+���˙���Xp7O�� 3�b���Dn����Uء�^
�'�-56���������c��F.K˝�F�5�])/%��?�5�'�]Ӿ���Ե_�f�G���Ⅰ�6`}v��P��9���[�{ #ɶJ�ǸP1P�6��jҤt���n5iE�'JM�c��lZ��
)/'f��߅ޝ�Hc� b��b�f���V|n�;jXHM��D<g���d������xc/�<�3Q&Y��yK�U&�u�D�8��A�m�9�x��&6��RC7]�~������Vieq�0}?���d��H��^������v��< �X��7yV|�I9�ЅX���3�u�Ĭ�ig���s�Ch'��7���=Py,g�B_�[o+�P^�J�����a~���X�jV����UP��|����Zzʇ��Ӣ�_DR���?[	'�??������� t��;�޿�i/b���6��p�Z��V:C��Eb��N����@T��������v���+er$��ɦ�>�L_�ZЉ�ѷըmto.�o����$��f���p��g��]�I�6*���9O���T�C��ݯ���܀qs�t0vք�=ِ�H��Y|�lo�	�vT�}�(�~�h�/�}	u4��f�7��Pl�_\�����j��.�[�D��y��N��2��]��|^g�jKkt��7�H�|���w�"������$� ��蔡:�9;xzqn�?[j�	"�2!�����6���}���-p4p�ȼW/�iw�"������m-�h�.\��6uvoi�ȝ�����!5ם��{��E�b5�ٕ�M�:�#ě�5DTC�I��U�Ì�@Ќ ;�?F� V��
�������d��8oO�"B�KK�T���(��9 �U@�K��͚]��9��i?���FL��a�E��NʣK�"��=������"L��A�q��}Y�,i�E@1�Ӧ	���K��:.y4�%�ђ�g[GX˞pT�|'0�����_�[���k����[�p.o��{ؽ�|��o'�D%�6�7�,�@��� ��a�Z��	#��`��pmi�HGS����]���aeF����Ųb�W�2�F!e��2�"��T��3F�%�;�1W�_XE��lBR�(� �p��w��]7��U13,�$�`����(VW7�7�0X�$�U|����u�.隩�q�#���Fc�N M�,U<J�wr��7��7�����}���Ξ��|ؽ���_k�PR��>K�]ˊ^�t��ǖo�J�ZW*�	RIyi�In��>���E]�hXF4	,�:�%s�lE|�;��:4}t�p�T�)�(sv
zI~m��<x�?�)��R/�)��(�D��m�9ڦ���s��J�f��)͈��������'�^<�����f���K���#c�˽�������J�ˌ��L(�BJ%I��f��?����KN�7`�%�u�p��k��c��V��O^3|���1)���J�g�3*��j����@Hin鎟e~��R��Rܵ����Nzޟ���t���>�j�:Ǽ������I�>�j}^���e;i��N8Wj��c��l�J~j��t� ��$���8u�Rڪ�ۧ P��1☫�>�����$����,�W{���9<T母ͯ���rM����J����GqOh4��F��<����������P��T%s�Ģ���Q��
�i��̈�wq�rLM�����{����0sb>��r��� N�l�����4��Wr�ĘmZ�i�H#Q���'�L�F&�5K']�S��~���������I�R���s��L!���������N��v]]�aE3R�y�)���d��é�ü_�L9%ΏҬ�3@�iS8Rj��O�ӗ�������V����"N�5�	�>Σ�&�ؙlp�v河�)��QI�޻z�.����2n��ɳ�[�z��A��L�:���LD��>�`�_���{�.�nВU��T���C������M]خ: �6G�+/����`4�X\1p,�J۝g(�^���$wU�͑�s�L?Q�<-*�`k�����Z���SW���Jm�3���P@�b��4����8Xq'����й���]��i��U*�X���Ӗ�]֯�\��/�G�]i܋'�F���뷅lF���
����9�v�L�,)>{��/�/���m`w��Ҟt�c�8����~~��'?��x��I<e$��0.�ly<��]�Yl qN)�T�&pF�n�}�Wq��9w�n.���]�Ň��?�K@������i��G��H�Ը�H�@��y��_��>��,ܿT#`�\�WO�Fq.�m4��G���]�K2牱ř ki�9�Je�����(+G9J��*-:Lm] o�R��J#��c1�����X�G�k�<\���|� �13��]��[|'�:��^u��&9��94@=Y%e.T�)�[z�D�����������,�f�f��7�?)����o�BN�w@�+5��p�v�E��=1�]Y��+{.��]��yR, �������JQ�����יo�G`%.��o:,��C�*LT�JJ�	��ꕷ7��S�y�I����y.g]�	#T܂ B�8Ԫ	@�)��f��� ew�$��GU@�&�Cz'>깵;c/�Ib+',��/�G��?p9�FT����IE��i�8Ő��Qf� ��;���,b(�$'G�+��N"xכ��5�2���I�+�PCh����l�d�ܓ�%��D�Z�@òү�kt}�X�^暼��{{���)�dT�/F٪'ر������ء3��n؟�nmб��e�a�*Y��)�	�ފ�,y$�D��C�uq�*QoR�9�9!P�_��m�������?��*��wwߟ�Š���L�$�6A�c��YXՐ��=	�R��;S�欫d�q7Ҟ*y�߅jc�f{��"Г#�)=���_��s�n��"�px�p�Ō�M����Ԡ��^�/-�ݲi<��-5Yދ�^|U���,���O{���=eH��d�T��/�9�ĿHkj�Ƚ�����������S���L">�קG���O�ǻ�2�$_��Y�����գ?��ۥ�����'��	�G1$�p�H6�7�'8�Z���Z�[(�H4^f�R����2`ŊT[>��5�
F�<�	���gX�����(<+YP\)����1�%9���)����W��*x];|�T�Yk�=s�5n�0e��ȝ*���L�mr�ڈy�JU�7 ��3!Ǟ0�w\A� �~\�+g���7g���$��٨�-19����w����[~�_�_7S�5�r�������ݒ/�7\�
��Krՙ[Iw���s/%�:��j����O(1�`OaSsT?��O�-}���`��Wz�vy��M�^c��ܘgs�O�������_QX�y��%�U� �錢���
l��+&b���8k�� ����X�eE���,��:a=�&a��&J�eᱸ �������%/��Hߐ���*$XY�[|�y
��>�32�Jh+�r�c�e|i�FE�Z{�B��'�<,��xK�N1�$�ȟ�M��;#� ���Hc��ӝU�s��n�H>[Ȃ#KS��
�y�&�sk$�lJ�_wm�<��,����4�}�-j��V\/J���;����-ݒ����>��t�ɲ��qN,[�������*i��.��eF��E�醰�+>VP�uJ�nW,�j�/	F]���nhY��B����5�*��_W�{��WW!{*0�������)c�z���c.,������19y�\����Es�4���=!Wu,M��Rri��^��9��T���>W�3��r�|(ruӡ�N G�Ə@�]��'֜����2_�K�DK;p��5#�O�]���JW����ࡒ�j2��@3&f�:�R�b���W��g�]�;e�����7y&�D
�� X�g���"?{�t*ax���ǉ���i�a#!v�^q)V]�ض�M���&�Z����;�f}���">o������l��÷}���,I��7�N+YVj��B�K~z؉�a9&}��#� �z+NBE~ټeA�ʙ�x��O���X�g�uw���d���3��E����� �������h�t�<�	9�hHЉ�3��@1&�x�N�'���T1L$�w\��<�������8s���>���W��`	�7�I-������X�"`!ԡ��tq�K����#�;⊍zT��S8�w��"'-�Vvkљ�����q(��ssrf@;��쬛l]��6��5;��WaB�؝�=��|k�����w��=vVV�u�� �2}j�N�,�=��i�6�\�ƞ���U��b�@~X Ty@(�(��keus���U$�T${��H�m9�s��x:��?}ً��~�jR��yP��}��s�U�ޮ��Ƭ�1|J�Wv,��#�FC�\Ӝ%~�}��U��ه� Ӱ���&�B"�p'S�-����!��?��%΂i�CZG�p����ŧT�w�\>�	��J}
�O�ɩ�Z�#B���n���S���{��⋽,�D޿M+���c��w܋?w��xA�맏_1$����������1�'E<����Ls_t��g�W�����1Zؾ�z �Y���ƒd�-]���["m.�H�R����!�O��X�CʼWڅiN��w�rr�4�Rp�Jg��O�f�ۡ���'�R�.���\Y�}��2�b�F>�Q��4��e8ṿ*|�Ю���^�'5�%��4I��b-��b�ɱt��s��s�4�F��վڡ
O�i���\�L%�ι3��:g�8�^C�3���$�h�ͬ� J�Z�.�j���wZ<��+�/$<���V��kdye�U�����K����nSb�;r��32�du�pR���ם����]�F�:���)�Zi�����H�#$�xJnU�uƫ8?�0�|P��c�>	���w]
�a�ŠVѼ�[9��R��\�{r�d�U�T�l��k_��F�� :|e��cW@�,	,�rҒnh�SҞef�}ى��~��zz��,z|���\!Le�Wح���ouh�TCv��s�#�c�A�F���� ��E����Ϛ�)Mq(+���rQ>q����y?S�&�U�]��x$�cю�ZiM}A�m����kԕ佊����z�˥'S�GS��5B���9�<ʖ�n���x������˘�4wP��הR�U�p�5e&��F`�Ql���� ��6l�R��l����^+��O�oa-p{��Ep5������$�u6��ld��R*�C� 2<�� �%�ꗎdR� �Ƚ�J�^����Ms*M�<�.��d*"'�2sQ�B[��Fǫ�V�\�g���1��W��b���X��(�r���Hŏ�!���I�u��!q>���L�J�K!�N��d �;e�m�c�#2p���쥤j���J���ߎ#�8�X�r��x>19��<�����H$�jB�`�z�$�C�R�6 8�'z6���l:F,�^Y����8���0����wwś��z@p���߻ u%ѵ3^u��{�t�l��P����� �T�-K�{�<�Cլom���<͢ۯ�(48��aJ����D�8A"�v���x�07$��X=8���)FV����W��W8@�oŹ�z��C+�TH��9C�bd�Ja�`L	ǨK�Z���_�F^�a��EȔx�0ED�!�����]R7\֛yԔ�2>��]�	1������@ns��cb�ҁ���ç�<��[Ǩ=9�+5ʦ�a��|D��*1h��ݭ�d������0ka僑�CK�{��}�����U��zp88;y�~{y~�C��ߺ��[U�D��;Y�o��Z�gqG��G�q�c鵁����	$l'$���<��gB��ENIó�^`\�KG��W-{��7H��FC+�HM�/���C=_����h�M���������^ݍϪZ;�-�����eLZ}��N(m�:S�U:f�䒻bުy8������O���P,���``4ߗ���$E��hX#O��Q��Z�l���}���y�/֥J�Ă���	���ϒɈA ����#��	�G���{�ۿ2�)��3�
���٢|��~���nz��Rm(��:`���si��dB	���?@'<g�녋 r T6lᐓ��H�����k�մ,QՓ'�Q4p��ת�}#G)�ī�"�h��E*b,ޯW�q�zDAq�lzZ��yʎ�gYی�R���曕+�j3dۥ^�֏�����r8h�`]���ЂT/��܏T��8A' 8���VJ�c�A�!

%�9%o�w1����#���$R-=�Op4$� a$��Ә�o.cE��
�.�垽;����ud�qb*�M�k��0m��K�V/�L�ü�ߵ�Ҭ�V�/UC/_�eŇ� �T�S͸�t5�3�'�잂[�s�f�D��J;�R#HDu���_Q���Az���/֋����ߐ�6 ��/�H��L�6���������
?�,P��剝FRi�a�[zm�����x{J{���[��'V�l:���x�k��kh;s���Y
�+I�뺔���˽���@�](��j^�F{�B��� ��M�uD�d�� "��Al�g�$�����a?Y;�"@6��_EʹS�����Cª �+b�۲�����b��\�?t��CL��s�Z�ۮc�%�
�n�O����?cu�N�M��M2�E�L�+�_�N5���k����;����%ZH[[>�j��_��� �oy�E�H-$�5@W��C�bF�d�t��L�(MJ�֞�_uXQIw�|G��G��[vg��#:���E�N$�k1�f�$q~�߷�R��VbZK�Nl ;6�-�o��!�{��s�(�J����p�y=X��w�V�=<2�G�)1%�9 �)}K��2�y/�J�;x������j�qı�6F����-N�G�y�K&���U�
�a@ؑD�ҝ���*��)�ٸu���4f�8�g��GG��{�ʀ�+"�l�芩
0��a�@��g�2�VV��~��QX��ۤŁǛ��$1 f��@PN������ ��S���u��_D�"��G?rb���S�T��jÁ8X�C��y��ܸZ�/�>�����g��`�mTØ .��X�Ю��[���q�Axw����#��W�A='.�Se�u%��3�d��K��E/���sݡN���,�A�_B~�1��O�ec!�M]���O��ݰ�AC�� ���9*�����K�eC��LF��C����� &'IOb�.�~l�2�G���P�A;iA��[:?!����+�W��0�C�ӕ���ʷ�t�[�
�w��A�w�ׂ.�.��m�m�5���
�)���=�٪����H[l�x�/���C����]uQ�T���LL��AZ�t��lT�,(׸�xW��T�S�|���EՔ=U-��λ%�h��N�h����q^�}�Brn�	��pC�Po��,�5Z��Dâ&��"�"���O.��G�Pŵ�迳����Z��R���P��{�`Q�9C�0H�$�c�k��Q���e�y|���q��	>�c�o�����*O�=�xw�U1�{#A|�k9����ؠ3*t�SnͲ�fԅ(Ew����	Q������^�����W�/�v��H:8����}�%ī�脊��pg����A��.��C�Y��k%\F���l����7c"�9�~!Q�bj%�s���)����k�[�Z�T⋳��L�>�z�<RFxUۈ��X�p��`S���A�ﾞ����-���_	���k�T@������t*�d$+�%v����Q?��I]�'��xWP����ḽ$�M�{��;�
�?}*P��>O8�֔1BĪ⼴��ct���^��-��Oi�����ʲo���<�ݲ�����u(�*5b ��߽�'�c#���I��&tJ� )yT9qL+v���o��a���l��V0���QY��lx@���c�M���}z�V���T�K4`�E
��A�BX��� �-��^���!g{��H!����G����y��	�ջw����R�G����90U6����N8���5�#8����Y0$���br�S7���c��[�X��*��*O�I�)l���8�i�э��V��g˼x2���ԫ�I�P�e�؅�O���"��&�����S�@Y��d����>&�k՜2V�0���7�rQ�w)[�4�d���_�j��n�h��63Ji��}m��|���q)ȍ�ʥeA5��8��������o!U��`p�4���з+�v�?/5��O�9��O<�\�8w�F���z��O���<�OX���,ġb�/��9�aߠ�y+�W;̳@�'�����⿐�-���*��Y�}�vչn ���}�K�^���(����~1�$�����X#�68OrJ:G�W�L�ڼd���S(π�ʌ�� W�;�P�gߋ��j��Z��ǁ��z�-�8�[;R�Ǉ]�� �t�cl/y^�#��1��hm#�b�G� �b���n4���%̥ps)�)�FYW�H�3�Y��ͳf�&�m�ʵ�n�N@Ӧx޸xKA�eO���k+�@�³y���͞\�hHV3V�j[z3_��V��75n]��ڨ"�] ���;��o�\ ���|X��}���c%��2-�l��U������D0�l�g���@%���`A��)�#o'��4#�۴����@���ܪ��8s���(}T��b���>��㺦i-��<��=��DF����e��iN��08}s\�N�F8q:]2J�o	{j����X��P��(tӨ���;jd|\�(TN3���� �X�.{W��nc	 �Ay������&�l!��|� �0l�L$�(��+��!�8�P���܀�qM�ȲJ��O<�阺(����L ��G�otL^~������?ʬ^���.-��:�L�w�wcl��^�\�$P�����'+�m'�(��Km�^�ј.e9;ƬN����}q��jC��{�ЊY)_�-���o������fך���x��o�	z�RR8�f\Y���w��;�wsl��H�*���0�*�9z؏PVM,*��;�� �Aą�	��UWE�C�ɪ�"�G��IM�W���uv�Xb$J�\���I����!�3�;ֈA+@M�x�:�5j��#�ќ���ʠ�%��<�4R��`���7V%�����vZv�\9�����-3��8��� m�s��v���K}^i?Zq]�(��m�*z��X5&�k@<P���an��_7-�>�߼��D5�S�O?��������S�Z�n��s�w�Xk,��W�/R�@6�pT��^{!�gu]M�:�#��ۉM�Q�����Q�VI�V> �f��&�L8�1��iZQW��������n�yp�]]�\�n3z���R�'��p��������⩛�>Y�/�w�����i�J*�Mp���4G��4�'�h�G�r!��B��J��Y�Լ��;[��5U'��Q��T2ٌ�浗����<��Z��|h�W_*��an癯�����zُ~�~��wz��~�
)��f��b!���DEⅵ4K�Z����=� ��]�P}�~G8IWMuH7��8,j=�'y�Oat�:"39�szn�R>�2�{-������ί�����w�O姡��=:�w�j��n�݄�����&T/{�O�w���Oe/q�y;H�mtܩ�H:u �n�!��, yh/i��i�J�7S����Dc��ufuJ��Z�s<�� �%'k�\�&��C\��s|E�|��{q���\��ʉ���t`��v����q�����Ka�/zAR�^��9��_2.�/�>���������m�y���0��z,钛��;� i��HH�i$h%0W�"��(��H���:� ��tt����vŐ�.>�B9@���o��a���OW��&���~��PnK�/��93a;o!�h�xIt .j��I��K���Xv�h��K�̭Ih?�KfSj��)nw2 �h�2(6?���ߔ#���0-�S�w��n��괻��Fa���R�����9_�a��W���j+�L��Q�cϙ��r��*YQ�K91�x3Ty��ҿz$ ��az+�oKmX6l݁�gJZ��`�O�\��"Ņ�5؈)����&}�<��'
ָ+�E�_���	�7 E�ԽK������z5�=�=CW�#�,��³���f�� ���|o�� z��P��d�u�>�i���,ދ=*��]ɣ�yU�4وBC�Ћ�Jt���UR@V�7��Zc\�¿�?�E�z���:�V1�LTO��+1`%'vy��ɽA�KD�9�œP�G���c���|F�� 0�)ggMX��j@n�9��m�TLTQo8�Y��@x��~�D��v��A����o0[F�o�uP��l�oC"aA&E��K���x,���'�iAr�b_1����������
�rLs�������m��$�J��PO��C���ƫ�bx��������*z�"�$g4����W���@�4&ޒJ/�#�1�R�|�*���"d�^}.�K}n�$U�1gL8�O��8XJ�|�y��]��9��~��O���2�Ezs����#�հ2%�)G3�g�H�D&�0����>k̝J��߭���1�d�	�"��4�Y{$�u"v�H�������?�"6��Ҭ�L|�`SA.���*=��ksڛ9D�\���E�ٻ�]y`�d������oFG��<2+F@�µ�ݾGT��{F��	B� ������v�JHyms�S��Ю�cK����e�l=�ո)��u��͵36c��]�daw&j)��� �b�P�[��m�I*�]+kǽ��7��|N���7C~�ݛP@至/Tʃ1�K�����
 ��<o�!�	�uc#3 �!8ә^�B��f��
yqҕǹ�JG�:܁3.�_�\��c;ֲn:���5���A�S4��V&�jR�E�}_X�j~X��Hnm�ʺieRLf,,-r�д��W�Ʌỵ�'~'J��}��{��[����
�A���hL�P&�8��Fn���Å��1�3DUu����d����)��uJ����%�pX8����u�*�-�E��w3g�1 $xa0�mw6�y7��u���d'�:Z��̏�]�$�5%��\g�/����k`��o��o��?if�Lº܊J|T��?L��~��Ȑ�:� ��ڑ\��j�Gx�I���|��Z���ƔtPG�xh�����3t�4���5,�M�����z*z�w�Nw�1�[�q��ҝ�s�o~����4�N't���B��[�M������m]�^�d�8Q�z�SlU�4U-��C����H߾1��{�'O/�u����;T��Q$:���䊁d�=��y�a�.�m�H[!�ci��}�)�'C��RZ�.^��+�u8/\�C�8�yH:�_�d�LZ6i���y�l�-����� �U���)�' �����f��+�q�X�B�Y�L�#H"��h2pL+?�]�im�_�+��;`���rd�̹�1:3����s�{�C�1F�0��s�^��c=�i��Ř�P;�!��`8�VB����ipU��b���15�v$.�&1�$�E
����.�w���,��9'��IOOP����A5�N���]������.���j�jf=�j��;�AK[�G�y����c�-��h����w	N)�� ��=P��	R�ݥx��$H	^��'�{�+P�?�9�]������5s�ﺮ�s��f�x�+��[!��,�k�z-��=��$9
�
�ؼI�J���E�cnɡS���NN��EF�S9��iI(�"4�����?a������)(e���A�4��=Np���4 �@���w��/ࡳ�k�;=�%�<f��Fwd
�Lh+�����˂3X�A�.�f`ή�"E����b�($����R�D"��o�_a��&�Ys+�����{�U3�W�C��"���kWƅO�ӋW�O2C���܌㫏7h����$8R�|HP-kA�ȏ7���38q�$�	w���O3`����0?�*�ΐ�K��H�?#�Xl���^~�Z4����: ���˿6cEOU���M����?�%�[��8M�__�8??z=ܻ�RT�OR_�V�k=�ƴX��c�ǰ^��{��v_����7.�鉖	�C#!�a���(bb�S%滯�9d���2��T��B9?N��|�s>��p��^��rܾ�=dp��s�t6<b��]���w}��b̩A��D2 ��I�Ć	r/n�uq��	%wގ:REy���^�@�X(;{� �G �W��Rj�@�;����QH� Q��J��p������w�y�C,$�M��=�7#'�8��3�m�5�l�#w֮�h�Ҽz�`�p�_���`O��'���&�5/%۞GfO�hlm���}��� ,D��o"?�.���Z$�6�Ŧ)\<b"n����:�TX��/��N'ʃ�d��U�)��|1{B:�uڀԾ"q^_ޞ�W`�l����������?����I;aKM2|e����H�jtq݋,+l���~x�����a��a
<��f�ױh�Yi�8lG/=��$�A������Bľ+�2�����Y~�5:�W�^��x��?PS�w)�z�$�ܰ���zz�8��J>Ӓ>7������o,?8�㙃-�+���vy�GCZ�i��D�j��N�MX�]���-]���4W,�&I�h�4��ʇ�'K��]B8���J���%��U.*$F"���9�B�Fe��c��<
��6����Y�n>һ�[�n�O������g�Yٮ�ۚ7�f	��^�b<�I�g���A5z�S6�]m���q{c�A�bs��t����r�����C�%���F:(�ZN2����Vs�oB�4�C����4��w$V&e���3Az&�dT,��0��[Pz4݀yZQ�T�'��O�!:�c��##�jU\_�I����<zH�l��_���/W�> 3��)�R�P5/�Kz�p
��.��)��H���ua|3��҅x��2���,t?�$��;��������@�����9�u�ƯCY��t�!j� �1�"5�F�'.%\8
�n*��l���p��B^��G����% �l�>��=H ��8>�^m�AwhX�^�wdaҬ�m�d��M
w�n���(�r�j?�������T=Tz�R��ӫ�.޼��9�Ka�}vm ��Sk���f^/��(��xK�8�L_J�{Ee&���0�����N�Ν~�ca�A�=_�I��g� hX�%�1�j��l�R��`ǟf����cqD�{�k]~rH�_��Rg�dr��N���[�t�| �J���O����!g��k�}�pa��9)���V8�J`L��5�Qf30R�0��"��.���JJ��;��7��
��D���L�K!C՜< ��l��	�E�Ag�-� AP�/C���%���d���v�EƇ�)�(D���t7'�>��3OZP�Ʒ����ı�0��}���sk��oF�:Wi� �FD����$#y�3�t�9�@����m�s8�}���ɖ�F�(u�8���x@�1�D1�$H�f?P��Ef��ϽM�<#���[�J��s���O�qsE3��Bf3��ͥI�B�Q�]|)����b�".���\O{i	Pڐ��������2j��+گ<+;b�8a	��ʹ�Pr�:���3��;9�K*��]���`���zyP����;��:�śe�'Peq�	lmrE;�7�o-�1�yp��!Q��Y����b�� $��ng��h:�T���q�'4��q��hg�:�2y�i�D���/��\��<���N��o�jEh��=���_��>3c����t�%���+W��Ҹw�8�4���j���SR�Wn�<�ظ��U���E��?D�WZ�����=g��@���37T��Yl2ݔ��h_�*� *0�"�}��}
$�'�ws�q��h(�U���V'L�G���6�C2��a��{��qnټKۦ�������<}͞#���Qn��+0� Hdy�!����?
�0�7����vI����df�������vi�x�G�~��g��ů8g�;V*�&Q�YL��k#�M�b��� ��D���׭�j�8:�?�FܕCt����p>�_L�T��ѕM�0~��y��}y��S�P�ݟg�onZ_�ặ��Y����6�����^��ˇx'�|Cl�G$r}�ȓ̩ ���"�7s�ww�W$�O'���Z?.���C�E�v�
���4��D���d �{�N_�bS��x�ㅆ�F��֗�ځ����Ӈ�B�'���g�2'�<�O{������]_�O����h�7GA�b��\��z���_�3�<)����T��yQ�%x������
��>[ J�	w�K��'���Y�=����ԭ,�e-E%��&����_�sp�V�^Eq�筋���f8jq�+���&��2A K�����d��z�6$�*%�o��S���;I��cG���s
�ᷢi��mL@�uriM��$��nA.B������w���B��7MT9�}�]��.�?\��,0���w�bMB۶��kH$�����FΊX�����Hex���,ɛ1���)	�_�b.L�P2�ר��Wz��J0������H�.��u�^e���-��,k|Q���Ci��A�T�*��G��J�s�Dż>���㥂�I��Y;F{A�ң(�ذ�c���L����qB�*�2v��NfN�1e�E�
"����+�(�H�b4>Ӽ^ݕg�ݯƴ.� �����}����C�l�ʸ>kn��6�~׳�^��p�<�{���m�N�)T��#��]��T���k����}P|q��"�S�#�;ח�	�	���|@��x�?�����K�~�ޒk�j�U8���� ����(���3���Z�	�8�[鏱Fi£����g�41��_��K����_���N�ף�+l�i�oJ��1��C��ǲ
;&��{x��pC�!D���4y�����}p��S��%�8��\O掻(�Wǃ(���م%ܓO:����H�oNA�G@���t
G�,q�kP�<>����G߃���+1`.���e^�����ee�Z�v�ಘ�g���p���lUI��˽�Z������z��V���S
tf�}�e��tܶ��2� �X����c��~4G�P��X�=t��j�"�/6�N��	!�����gD��!e��k����ћ�����=��[��&����c�c���X�I���@���?���m��s徙B�N}77�`𢋥����{������ѦW���n�S*��j&�����	���^2?vk���/�1��������nd��\1�E �ܾ$8�4�J.�b�&G�c��#_g�~yٽk��Ԅ	;�z�}����L�6��?�YfH�R�4_y�k洀��?�����@;8��ӠuW��>! �#M}�Ꮣ�R��%� ��0>���^>Lǩ���`�q[�01G�Q��_`Q�W��y4*j'(x�sqGXD��I���b��??n}~:�x�?�Ls����*����Ii�����&1���I�
aq?�� �i7c_� 7%�ve^Cz�!�?�pm�Gs���R?�p�=�k����b(��C��M�nt��e��E�I.�F-[=5֐�v��Fs�g�p�L>h���u
���G������甏�G�B��f��O��y��&�at��V��}�OW�~���Q�F�7���{R�|PZ�L3%�.��r���C�����G���A`�x��/p�!�{ԮWPvzAi�D�Χ����
#�Hu�����@���4�_乿�<���ۙE���>���+Kt�ijeCX���u~}�W��5���Þ͈#�������#�/�K^���<&.��������}N�g�;t �oR!��ӿ���swl��\��}�Ga� eswCy9�O© �#=�T��?�W�Ĕ�����rC�攰^���sBڇ2N�3�k��r)��N6𻱕�����u��if���O����m#�y5��B�?L��9|횩��]�v�QdmcƢ�^sı��J�B�eo39����;���&��)V�-�������]��=n��ħf�i�E����
<J�O�����B�(
�"Tu���R����2t�\N�c���ͅ?�ʢ�OX�e�23����β��Zv�$��l:�|�>��K��U�ɇ,��jo籿�p΄%}�6��������ң� �z��`�}���l�w۬�f#i��~/�4/�Tz�oo�;�>F�*{ ��e�B�r�̶�!�˒␈�F�g�(�4��ܵT��A�ĥ�M�eg����w���\��[�T@0?�đo�����6i뫗�y- i�i�L���:̀���_j~��NuF�;��������.Y\�EQ���I���+<��0��a~��]�q�������%�Cq�9���}�IM��(�~�hE��-��9]R˚��xH����C�w�ٷ�?�f���=���"��^W�ӧf�A�;����̂-$̨�:}T�D>�HsP$=E<,�0]���m^uW։�w.�މPi5����/����Ѩ֖�Dj�a�w����畣/u��i�s1�s�qa[�:_ٵ�A�����?��a^Q�#7�P^���*�I
n�	CMZ`�pr)[pKM��Z�������j�I�}zsL	��O!��y��>���/�
l���&�-�W�)�*/�\hKD'I�o�'�TY\#XT2��q�'ZڧV�ٌ�T�'��Z�@�b����5��I��a�u��r�:��_9#���S��H�+�.r>��]���H� �^MS(}�#*-�Hٮo4ꞃ3��gz�»)�U��{�� ��,�N8��(:,+\��k���u��<���'[4�Q�%*��[l~c�<��o����گ�@��g��*�X|�������.���Gӟ~�{�-��vQ�棍�l�}��zY�9{n�%��x�!x0Ku?{א���~�?/�|�1I�����CL�">-�(�:���N%��"���kג��7����y}V�ܐ� �Hk�e���p��t�7\!r.�:����ϣtg�z���0��9�z����C|��kap\ ����`~<�&l���YȂ||�G�9��4ǅ��T��<�k�:6���5��5X�������f!y��u�x."}����KF҃���D�b���Ý�ݜ�E��Y�v{�v�TvfD��{�*��Y8Y5�+ȍ����'%E<�+Ͽ8�����9���>�d�cG�E&���gҳ��	|��OU�i?�F��5��^QH^�@s#e�{ �~
������:�(q<��۲���e�8Km�ܬlt\�Z��hj�?X�I*R Q|A����O޿�ڿ0�V����Xڒ{�(qQf顭)g��l{�!��Axw�k)#|��A$�%�+��r~pǿ����g��v�Z�B��Mֽ@l`��B�b�N� �!PLe�`�2Ǥ)U�1kWT	�.6C�O	�jF|�Lk~Ԍ�ڲ��#T$�s	��갻,���Ɍ\�_�
@`�j�ą[�d���H�G��I~.Շ �4Z	���ˍ�����d\<�,������:(�u�LR1etd�E����YE�/��Mq���Q_�ڳ���l����Il��GN�ߎ���+�ز��s����#�_�d%ҷF�>�v�N��2.�6��<�woF̨"ѷ��2��8��l8 �b����71�D%�G��P`V4��GEm7��G6�C�b!̊3%����\֔#�xo��qZ����e:�<�#��p��]8����e\�

r)9�M@r��m�c�d�K\,�G�h���8�}@�hNn�Mxh��%Y��M�d>}��BPa9���hMSh����e����I�F���hod�v<�M$=�¡����	m-kw(dpXԎ]��@)+��NK]���o>
�q��߆����?Bu�+.=�i�0�3�$����=�g��]J�V��s�/��1E�3e�+����`�J�2Ц�Ύ�M����P��d��.�v�.�����Ewd���GӇB�E$�U�#L	�$�uU}�ZK�p-��~mA_�L��dV�AQ\6<�����\I����<��$uv�I0ݒ�����g	�R�W�k8~cF��@�|��~���aW]�]K_�Q��j}�U�RoG$�nf�B��h�#𸽅����V�@M$�\�x�N��� B�[)�C��:S`�+�-��">�-�O��t��(-��5e���7n�6UO�]]�6ַ��d��m�i�hֱy��Z���
R�9�/^g�-8˥V�����L晣�� �2�P!|�,W�1�(��L;�c�١E
#��bIR"
�X(�b8��?�BV���c:uN�T����]�Z��mG�(�]�"Q�9���YE����v��kx���5S}���7W:o��=��P�EN?��N�r᫆g�m�hޖu��H������׻ُ/Zqh���7�M{+7�櫨��;HD~=$;��	L�ua	 �һ\��o���V�|�g���㥯���2)Y��Pz��o,*��1{�ͭEr ��^�Au���!��w�s���(�(�`��d)?�w˷���YG���Z�i����'��i�K�_ێ��L:M���P�ϲ��XV&�z�o�`(�]���hI�0�.�/� V2�����:���ω"(I+��E�����C��\��ͧë9ydך���u|:Q!����o�Н�>U��
?C�F��m�����U��;��8*�~��O���FJv�Ӏ$
ρ��@,U�bh���G�V��Zh��x�>$��������x����������ڠ��*fM�?߼�����N;ʏ�8x຀�H`������/���IMN	�B@�e1�Wr�M��O�:�w�c*l\&^;d�����⃨J�hA����f�	Y:�)M%�ï���+��t�Ӵ�aF�]풋
�%�4�c�b/z��z�tj�ϝ��R8�4'ǶKȳ?p��gn����_�\�s-m�kҾ���"�e��JD��f+�����Z���ǔĵ�N�`9D�'zu��������J�'��U_5\f�ua��^n2�k�s��l�V2���~�IR�M��s�jG�Le{�g\k?�]��ۍ�VJ���AXއ���)�;/�~L�gg�?�4>j��o�y���[���"��3" ̈́�`�Rn� ����,�a�G/dȾ����V��'.L����(^t���S�1l5�
�Ŗ6Ĭ�9�$x���DfC�{�:���&+-�ʀ���������e*��{�z����ʸ1��v���!K_ߧQܐP�]Ӡ��~��gDw��1��ӓ�X4�h�J䴸�0,0���4{�Gz�.4��7�9  *��
�`��{�+�,�y_�>��zX���7�Ngt��~����yviE�@N�d &*t4��OE��aY�s���P��iakn1�~�ysu��ӻ�40?C�2C�0��Mr��M�Uv���x�����;�*���|C�N�;���������������i�R���許�wUK\���RQ��EL~3��-H*VͽZ�V<�ԉ��rAB�3��i='8�L�1a�.��~I�u�V���&�Z��o�iC=�NJ�G�m#4�*y�2�{�j���-zj�U�~T�;͕H�#ɭ֫�4N�'s{���m�м�~2m�*�6�9��c��pQ��Ϫ`�h��k[Hq0�%��J1ȀO|����?�������~��&�)%�������k3��;�I���(�w� �k�ge�y?S�r�����Ȝځ<�_c�>��,����ޅ�[4���#�.�ĩ �n�g�<�r�\$�L(R4U�Ë@N��J�)�g���<�>�R�<u�}uk-�-�>�l1R�R��庎�l����Ng�j��PBbD2c+�:.���"�.�
75�gդ�ʒ`7ˬ�dU�+�t�vz���\�]޹��q�!?�$���_�T��� )^V��y��t*����N�rxM�5���[oY�Qe�ƐLj��c?(�Za
1��i�_׺cCC�z�)�$E���fߔ�������o�`�J�LԽV�#ȃ��e�3<��M}��ϳc˭�˧N13�^�xLwH[�p�?���M���q�h}������KSd.;�r��I�� -�j�(�v5M��r� ���	}�l�!��Ty���c@j6���q*��G���}�5o��A��\�9=O�9c��������r�+B߁�JX�{K�rn�:����l��_��Ҡ�r�͸���e������^�5��;ح�����k6���(��9;�b�ߟ� L@L��c50�H���U'�[�#������;��CB�w�	��:(FS��OG��~�G�LM	���Y?R�|&Mud�1E7ɑ�/qb��:6xt��VE͂��/�7�˖ġH�hb�.�)�HŴ��CP�|:�w�5"�-��ZQ��'	��--7���K��G�����8%&`��V�F}fc�#��b[5@�z���<#�e �&ȫy.Po�����؜�H�䪊��a~�\�4�CA��}|卖
���Ăi㈑e����K"_���(.���q���}e�<�77G� ��a��b�O}vI�G'�x�d\Π����a�^��xe��'�L�.��hߋ
|�]�#�O�y��29s�~/�x*�k��_QE;��2\�>,6ZX�4�P�q��gb��
�Z&����$);�W_�dܳg殒�|��S�����4�����)�,G4�E(�)�Zp�"�JO�����#�Ƶ D�>$�.��ﲡ�j2�ag�1���=���>���|�L��Pw��+���,�{���nH�wE}��EDz�}�:G���8�@sI�c����Q�d�)6�6�����x�0�69wGkv&�`Qk�ڹ1��=�N�i����%	��^��!�->�iJ�#)*K{��gRТ��#l�zL⴩Q����:ZJ(��#I"�0s'-sE�S��� �1�etl�=l^�RI{�7�C2����=���nRA[��s�S�s�u��ܜB�D�]Z�2qx�E����IЧ'	�uӍ����M�JL�J��h#�l�7P���2iF��m.Ϻ�#�@��r���2���U���;xo��7�hW���U��|QuM�WR7PɌ,�63�6*�W�4���H\Ʌ�Ez���}&o�C_OʤR쟴����:�OA���a�a� N�Aa���5��?�)4W�B�z���5��5��|�CB�^��62"���ʙ��E�{�L�Q�ē�����z��w#E��j���)��XC+*RV5%\�0QG�W��C\�}ec�)������J#�9�zY�u�*s���lo�a���)��n��r�oUk�_oV\T�0�uBQ=p*����;�+�o�*���&3�M�b$��Mؿ*H��'�,]�H��3;��B-��š!�I����v��� 5���8�D�P�w7�y7%*���_��%��E��+�[{�
3���t��B=;-��vLG^�럩Z�!�:"z��~��V��lS���e�~C�[w����qP����������ئS;U\���6��C$�a�k�UA�]ە&n��^�C9�vl�-b�h�a�3Q��}-Zɧl��O���d�A4�<|Β�"�=-�[+?�;%����P��?��Ƶ�/��U_����E+�:������rC;�m"�>G�G�Y&�7��u�u\����?jZ�����i�Hx�I�n��ڡJ��RV���/o��v�6�BNgJ�j�obR3=V)37��A.�ٴ�6+��h��k�G��br��h����(s~ZZYE�^A�V��&>mai��֜ͼ��兟�������d�D�1�'�������j[�ѭc~*��lggYW�@iGY��&5C�-+V�i=-�L�/����ݵ�(~�X�3슭��"��)Μ	���p�[�D4Ud���H-\�[+9uЦ.��y\NU�q;�HR��p���u�~;W�.Q��_� �1�⏺�ΐh;\��*��o���.��}����-xuØ����k���XE�3��kƎ�<8ړՙ��]��X��K3��tnP�����k͏�Q�ʁqYA��i��Ӵ��]Ȩ�8=�dT�$?m�,!cc��NF����R^�@��,!_1�8��+�f9E�g4��ȢD��1�LE7)s)9%��$�\��s��M��xoL����Oؿ�P�5��(%�*�u|>�����[�7	V����R�t��R���-y�M;�k���r;y3��nn{�׊Ď�KoϭS ��;�� Y�q/5��̃��&�?q̮ߵ�g�5����n��֭�X�:=Ft_j��fa���Xf��tk'��s���,�b�S��i���[�`���ClZ[���nM-nK�� c�,.�L[���h�͓'�q��t�
�J�@�u�a�#�?q#I#�CrG� (��"x�̱�Q��SìQ-9�=T�(�?i�������@��x���a�V$�8[����˛�}���^zF0\�S�в�`~��D����ĳ�%E-��q�Dסyh@6��Z��W�`.�7�
��9���S������������s���N���K�t�[q%�IO٢-��S:�ӿK���II�IZ�7�KG)�O��'�l[��b�l�EU/�I������{~T�+5�����l��J��J_�L�@�h�\�7F���:7{KD]�� پFm����_������ˈ����X�&C��%={H(��n�}<� ��~8�ٗۧM�N�#��X��ZA�M��o�*=�?���Y�j�B���N�Lx�ݝ����W#�9��ڇɦ�~(��=cq,b7�,m��(��>0Xf��;����@>A�ˍ����f��6.��N�_By������R��R�]�[���L�M�9#���\����ކ�|v���3V@��g�c�(Fh�yx+�����k�
�x�6dq��}��+�P#����2�TRpbz���D>N�0g�`:Li�2.���ٓ@��Z)Z�՚�duڎ������%D�D�uχs�<<?��~�t6�y�),S��L��4��#�b�ۖs�J��,GR�^P��h8R���L0p����ѥ7������Tݯ��0�fq�T ��(����L��"�#��}�˅|jRcC��)�X��O�����?���&"�n�%��aG�a�3��>K �Y��/��R�v٥
���9}�������4 ���;�[SP�<X��/�#+�U#!3�_6�7�CPT�Q=��*q�K����8���8��_��t�~п���������GV���ty�Tt�߇�)e��z�sBm׎0b,������"���bJ �
nQ��c�E��U��o�"y�
�!�#55�H�?��
8M�y�|������y����x�|sVc�xy��S�%���GD��V4�r�-�Ǐ�TY��R�ŏ���d�ç�E� ~f�k��B:ܨ��E��motP���GIE��do��dmWH�*���n��_����Ô!�|�l�� �I�eHҸ7l�JB�_>����c�9�R��{����ɥ��(N	�1F����Q+Q�کe��w&C�]i�yL��âD��C�Y���{�5�_5<�@i;3����G�x��Lÿ��[��v�3"-f��]6�a�A.67J��R�|c��~qsZ�a2E�����{w�@�D���T䅙�n]䳗��>h��Z�)B�b4��o���?6��~���Z�7���7�9.eA��`Nȹ��tqMV2`Xq���J'"A�>͠�C���G��}�%���@pve��������dd�E)k'�³�F
����$ߏׄn����<"P$\ps�8eX�cJk�y�zt���b����~py@���)�W�ԭ�qwft�'����i����e58H�<���V�+N����:�ϑ*Ϧ+�Ǉ�ѐ�շ,�+�%�ˢ4�ݱ��`1�]Z�wL�JE���z�~�9q�S`u+�)�#I�o1d���9��]u�W��W5�܅���N?K����dC�a�Q���o��{"�����nS�_�8&qgө�I�1zH�Xó�Y��v���Pi}�@��x� E��H9f!C�� �F{����������H� Ů��0ׄl�M�7;�ڑ�W�t9/��V ��^�N�kj i���̟I���ۿ;`U�ŋ�;��6ûy��E�4����Ԯm�k���>���b�������6���\��Y�H��94��by��C,(����F[��;5)��9zSi`MG߫r��fq����!�h{ǰG�;���\9��q��:�lTI���������Z�'<B��tW#�����,Lć����|?jۮ��L�K1��@)[��x�[g��4C�6��R���&Zg`ī�����v�wF�J��<1Q&�8v�R-3qF����/R,�����
~*~�ݙ���yK���~�V���S߷O���W��`O�61c��/�q��D_����UA����]SCd`�<�
K"U2�0��ܚ#�fkk �2�G�iB���
7��փS{��gi��c���8"���c-�ځխ�YYݥ�iڀ��V]g��'�Z�E]�8����9�����'������Z����8ݔ~��0�j�:������r��vEe#�sa���8������ݖ(Uq���g"�>T�׽�H����Cz���f�
v���_��3�c8^�A��	�A=�>��6}>�꺝��cg�
�NE�����Y#��Bї�8KBÛ�f�7>�Sht0���*�M�OɆ��H~��ni���
_ٜ��	,� w���Z����E�b���R��n{�y=6���ks#���c^H�P�C���7�x�-���fLRy\�Ҥ:����7�osQ�c6G_�M��۬{��ed�0�T�S�zs|�������fc;
�������&Y�%ڧ�Rp�;]����{������º�N�9���m؜�b�]&z�ͣ��\�%q'�|X�|��`�}o��И�W�h���ݏ�Or�L�~ 螽�fĤ�m����|�Ѝ�%�c�O���`7h��XI�
Q"ld	�����k�ґ%����I����h��#"+q�8=z>mȀ_-l��c�%u=���nH6LH��1����ܜ�<��?iI�͙�H���$3�g��2K��W�S�QKN���|����s6A��-j�E�:����I5��Xsss��v%�����<^Gf����q��q�ZB�]`,����z���vN[C�o�GQƆ'C�%-�f�4�~$�,5:4��=��6t�?c�7�uU��`��m�+S5���XA]��a�����a�w��ܑ��r31߇Ň^Pfm�G�f�]O�ֹVh�"#V1��'�upJS$��������%���;eZ��(�P��'�� )��%�,.�l�Ph�#�c{N�0��<�2/XxW�!7�TR)R\)U*2�I^{R�X���/�`:�	(�}%)C2�Pt�,)�E�G6>#h�AX��d���#[�'l�.?�f ��������(�1<c�#�ϻ
�%].��+0����=��3ʸ��1W��s8C���GA�|����x/���v#��Pq!g(� ��A�%*��_g�Ջ	;A�o����K֍yg߭���t�̀�"w�}K2��$p-p1g�I~Tm�{+C�G&�^/Fn|=�	��}`��X���0��o+:�3�T���r�*����A({��У&d��ǸH�騦��]��3x������3�5�-���vh��!ߧn�f�_XJ��ۋ�ڎ]LAZ*5��r%s�uZ<�0����3��Y�������Z�F�4=�~�8��/�Qd���1O�kU�0(�<(G;�p��z"���݅�s�e������M�?�D����Ý����<��5��
�����5��ڟ�#�|^lg'�muf�����!2���;W5پnG9�_��*��BP=X�g
������N�!k"4�ҡ���w��o������I���.�6�f���W�|��q�Q��G�O���x|��P�9]TR����Wϗ�rҺ~(�
����%�Fq�x�vő�uk�����EM��٫�C�q��FFA���D�<9�� ��a*,$��EW�İC?����!L��۟��ŕT�ð�.y�Qە�
W#o� N�����(�^�=9�:(A�m��ӫ��C��5�4G�mIK���x��@Y� [;ɇ^2A��/d_�러�x�ǰ��.����u�,�m��Ϡm'��W4����Fn�,�5�bi��6"�{�[zJ,�^/�{������z��v3��������z[:����v��x���h�����=*�?���L5<*�kXA	4}��;��DPK��#��K�B�(��c�#2���.�����7$8�C9�_amg��� �����|@4�DIK���!A��jc�)���K�Y|�>
ny�a.H>)OǏ�x�ˬ�_���ߔ�(����5���4����"Ҟ �ܖ౎
S�غ�N���|:I׻[����!��-+I����D��:#:?5,�\&Q��)*-�QI��%�?��ېJs�x�Q�*}	03��@N�P��^S��8��x��3=��FǗ��**~ٟIf"���#;���AW��Fi�N��%=�,�ο��C�+])g����\LOא��W�L���%<�#��;z�{�#�A�-Db�C�<���(�)��/�u�����F�Z��6�;�0���R�H���:�#�"�r��85X_��T��>3�^�#����x��C��Jo�$3~k"+�����	�Ԗn�H)����-_�4�������ߦ�,�m��:l��%M\���~L��+�a!��3!MJ����,�1��#��0PWC�� ���XYy� ��=�;�hu���D�N��iв�h�V��{�f�s�$�5#;�EZ�M10UJ?]�^�l���	��OA�>c ��]��W|���>�5�[��1\Ɇ8GD�L׬c0t�]�ը_��T�u�{������lN��8�?z*ރ���v&�JN�^�j�we�	���B��&I$���9�N��D�*w@�	%pdiMڤa��t7��W��ȭ�Q.��t��.�xg�.��2�gBx��=b���ߌ'(�I�ur�g�ꀲܜO�[�`�;;�T�=��gᚂB>k��É~99��T8��CJ�/��L|�q���?��1��R��c9T�}���w�"Y�l0tPl�aC�H�8���^M!�{ª7߷7w)/�:QxA���[$�f邞<\�?���l��H����������Q	�f�M]�����Sg�����i��>M�{D��C-~б���:����^�U�}(Ι$���&��b��a�q �N���ѮJ��XF�^�D�^6���LL=�/#>��XF�N���ڰ�4���%f �F�-Ͳ�O�l8G<$*&�*�K܍��Ǜ�nms{�gm��"�1�@��n�o1�ؘ�[�:4?t���[c�8R�g
�?E$�52�7�&�LY���ď�����a�v�$���O�V��W�%��y5z��ʣ
)�^@�Q�(1�$�W�V�*}{Q����5��m�'M�0�	��������O/�w�,�� �ݟ@|�w�v1�g��1gX9��Du��ޱH���B��r�:�>�$�&���$�7�۰��L��"�Y�VQ�+�1��=�}*/^ݸ�js�z�/����A��I$J$��-]�9�ߓҁ�s�n�(�����=7Cɑ����gT}��%W\!�|�����F�yă�04M|����]���;i���e��R糚�R�o�f��mS�h�")���܃K��R\Cq�Kq/�w	ܡ���b��)������3�~�L�%;�{��<��v����}��<����/��H�]�J���5\��3�>T�zZ]�p��^,ҡ�;�Ba,�p�!�71�@(�B�w���P���"z4G��J��Q�'Q��ýiֲq#��(���V�6��� {#}�0�Q<��I� ̬�!����Z�ֱRD.şP���g}b�S^c���y_�����b"��Fٳ���H1��=xsw�*H�5:��7sϰ��S[��珢��tPj���ny�.Vc*f3.ÕW����� K~����`��bc^��;:��5�>�l�i�0��Dv0���0L���� *_.Y����|L}|	�Qvm!q"qp��0�Bv,#,}���Hn�Z���0%�2Zz�g�o"��1�aHoˤ�F�a(����*$؅_��C�{|3$D^cҁ��뢞�L�#<n�@u#%�ka�	��Dx�<�j��8�sWt*�A@�2w�|�DUl�p9�۶��X�o!Щ�β6B`�$�]+����a��q"��j�L������v����`Q�R�T�Jm�WvX�fm�a*�A&�o��rP��zf���
s0����}�w�c�چW8*�+�l�Da?��f�6)V�3��&"���O���s�ǽ^�́���&�w��6j�BK��)��t`�?k��)4�ᢋZ4�R,)�����~�tD�tD�����O`��<7�K0��m��EP�p{C ����G&�W��mg=$���ԲZ�Ey6��`����
��(�3K�K�o���(o��Ca����߲e!�4���h?� z�\��-����hy/Bm ����D��!�1b��_�(M�>-�s�ת�x��� ��-	0{�h��ԗM�ܩ���GHQ��W�ԅ�ٽ�Hv���4�i�	�&b�K�l��XM�G3�:͉��O�7� �c��.�}���'�!�+������w\9��$A}��H���v����cƩ���r:n`�G{y�5
��auY���4��Q֬��DVǜ��� I��
	��f�%6f�m�K�?Z@&����S�?��g�O����(���-Z�I~-��w.�����)KT�����)D)�3%?[c��Ϡ���	�j��!y�w�X�	�������r����2Q�����i��
nn��F�u��%�M�G
�'T#�E���L$ۅ���	�WN�0�O�b%�a$�����N?�0��;�o`>��E���~b��,�7%>Ln���ycn����td_�9�O��buJ]�(�����eU�N���5c�&������aX��
��4d�2�{��Fg7�K�}�[�����)qϔ��Sմ��c���J�����M�:x�Գ�WKYx�����~��\����eIx��f��nq�b�n�m����N<��]5i;��B&Wz��1/�E9��W2G\Hv
E�z��Fc�vߚĽn�������O��b���p�7+�Ҽ�h�$�ڊL
�f�/Bv�eQq\�9(Y\VUV'��I/|��Q�F�[9��M_QI�2}l���+T�����6���t�В��R�,�'�������%�1���0y7���:hO��XDpw�<dX��z�%��ga�)9�����q���p��-v�R�b�!�óŉDۆB����s��A��J�N�������nߓ��8��,^'��X	(�u����eq-���M9^�]���G#sxr:A|-�l^�NmV�f-�Cjڷo�Y>�C@
��՚��(I��K?��YĿ?�����?�(X>E��Ð��f��0��\|7��2����;���]��=��	�/\s_��̦��&|u��L�W�iE%{�si�7a�Э�غ���G��vJܥ=(��l�y*^�x��иt�_#f﷖u�QA�Z_���3�u�.�5Wa�C�^��a���/N����3��4�/*��n7Z$�>��p����n+d݀���m��@���]�q{��)7x�t�*�p�4�x;xwJ`�wU7���mm{�[�gy��v�����˾g�9פ��g	�E�-�k5���X�yIa�� ��U�$B(ݎ��i���զ?xڜ������'K�8��Z%�~cd�����p��_Q���g>��O}���ZZ����C)U��c�Vh�;*B�uK����@T񏉰�Ǭ��c��|ᬽKc�@^�):Z&��oz�vC9��H�M�( ��:`G�`R.�Q])�r@�8)\���W�d���k��$у�*p�݄�v��b]9Y)�F��]�~�83�4��n4ut]��H�4�rx��x�L���!�b���h&�=7����YS]&�X֋�n7!W�k�����z�0�^hr���N��O�bU�:��<F����A-��`f�������O�p��zLpI�~i��s����2�Ofm!�����u� 9�R�/�"�����?�,F�v,y���Q4��鎵�(ր����ɡM�c��t�q)��N�=�K�P�s��W�	��?��8$��_q~i���~�1�W�Sϴ�:���ܲ�LP��&����oފ"��^yؠЂRkP����/�N٦�D�w\k��ú�7���JO�
�q�g1�H����}�&�tl/q�����o+��l�I���X�zo�a"ޠ�e�q���� �9�H|-�������Y��^���k0��5�v�-E� S0�)�<����%|�?��\}P���7�����L�J�N5�?nv��}~�w\̜s��;L��cX�����왷]F�7�=ť�Q�Ë��ͼ����̗˲M�R�Ogz�(��S���H�K�U���.Ef�Ϭ
�#Y%�g^Q��|/u�ˉ��:��,K��7u��`�U(uq9g�xd�P!,�6���"_�D��0?:y�J�6{sv]	/ۨ�B��^�|=��X���B�`�,q��Z����7�KՏ�tM�FUꪚ�9�C2׵���T2�d��<̰��:���Vq<��꺖��ى�K�/�P�����$����w{f��~�gM8W䦝��+N��Չ��)ѱ�\�U�`�}��
�},�������g�f����j3:3~"~p��	���K&�J�*��.-�O���
�L�����5�!�/|{-ϵ��"8Wf�K���k��K�K3�Xo����R�,Ǖ�{�0	���u/�^�4�~-%�Ps�G�_Q<i~R�ys�7��(��j6�i��x�~�$����Pg��?_�v�����A��	㽉�g��8 �y�Ƒ���؍�����W������4z:��,��.%��t�b�@yx��T%��($ޮ�����X��|��n�|A+����}2�z�y{ش�?�}�n�����I{AR�s�xuEWF�4s1A��\��X0��CFw%S�8hro5Gn���<Ìp��$��n1[=q�cNm��*�U����Q�f��Jv�G(��mlK"�@5`��%��zn�i^E ��=!+�C!�Ƕ�Q:!��������.ƫ�"�\b���:�wA���r��4Ұ�p�b�H��ɯ u��M�;��R��\zx'��&�b�2�F�|��$�$����zzF�s6Eۇ����r�Ұ5�����P�ͥ�G�?,�v�y����v���hNդh��۵̸�6傟)��.Lo�!���I������/H��hC�-��0�pYy*��u5�|k�v��R�*�4t�G�(�Q@��\i*�B�"C���F��L�oؙ�1�ݿJ���V��+��J�'!3\�.h�Yp�+{�,C�?Y�RF��4a�Zq���n̪�t]� �N2�a1�=y��;&�Ko�$9��M�x:5q��i���qk��uP���g3�q�i0h��8NIh���)B�C�/�k쯭�����ܫ|.�d'��?[��9��'�o$�6�Nڞ�	�}��+.������֋�bs��q�u�N0���NAt!ս/�uꡅ1�G1�q
ؘg��=�����������9p9�mYN�8��X�4i����@��߸s�N��Z(
��Qd���~��s��������_w9�1.=U�[è+���B���Uufy��Uu������/ݠ-�����!�G���g��Cgua�<Ŵ�$� ��ٵGE� f��ܟeZ�[�|B���aH�t�%������2��A�4Wv^�a�dX��LBˀp�V�� K�&(�4�Kiz��%H�Z��rW��+���M��c��uZ�2�pp�R�yV�Y��{\�@��
{熢p�G���8_����dU���}��ʄr��]<T�4.�^9 ��w!Gro��ʃ�k�}٣��:%д��`2�V'�:��7ؗ�����xE&gJ�~V�;�^��%��_20OE���`��v��[W=cdj�4�Η���UV}�8_�Hc�xc��L���f(P���t�P�^)�����.�0�|�%��(2�/C~W�|��ؠԮV�8�V��|�p �͍���\����:��`__/�R'�ԺZ�����?�<"?�׭���9�7�U�����H4ۓ9@f�V��t��o�B����b�з;��idY�-��?� kI5���8	�1˂#�#JAL�&D
B���`ȪH	��4�C�.K��xǮ22J]9F���9;|O�~�;����Jx���^i9?V�� .kM�$O�'OM�!>&�g�w+�{�������f���X����A�/�v���e\ID���09����<�*�P%��5Q;��q��B��P=S�Ņ�7D�&��f������y������}�b�vO�}0w�k	qyn�fLф�������N��rIQ�U�����o�N�f�˄���i�`j�k-��1��DJ	�N�rW��N�^��r�3�@{���ѡ4��C��иϏ�ƾ:�����D�1⮻�.��
�Ѽ�I_c�������,L@�p&� 9�E*^���;�'����o7���ۼ������qcH��I�)�:�� ~.�xt&1�&���e��Y���RL�=��k�2��-JH��+Ң�ܴ�?(s�&9��D*��Ya�if񅖌E�f-�5c���cs`�K!A#2?V�L�x���8�Pi���7�������ܔGM�u��r�\�P�K�&�ڗ�_�����&���MH_g�ѴJ�������ߗ��I��!��@�c&�GO"8$	�r�M���͜���eG�h�8�5�8-�]� v
C��\��2���B���:��;��7����o~�ܮޞ���q��d@�'kz�$�{�L�갌/C���d;R?��n�UY�o��e}PZ3�Ȳ��I�����>�߬	,���.��Vx{����kk�+kJ?���6���~�C���}f���ٌx����Dω1�c߶2IH����X5�[��>��I<�D>�w9�aX;�M�>��y����5h���0,����3|�}��j49C֗��� �b��s���h�;/�8DK(kZ��zv�ŽR\�Z\(Ӵ$mPimE|3
�e,����{�$Y�%��}�ċJ�~}�F?@�[�iZ��UQ9#��8������99�ZoN��+8��j�~�!5�Bg��e!��'�f���=�����H����v�Hyz�]+�X���<)�կgJo����G�)�xĒ����q�N�D�iX��7�.6��:犏�P�$�N?�<��"��7����x�e�&�tG��T;~��nD�!��Up�BᏙXޫ��o嚪��nz�S�����.�Ҩ�����q�%6�� �]R].�6�R��P�����4�*���J����ǔ��ߕہ����8ݜ��_�奖����*[v�#6�}��`��&+������ޛ�p���UǢ_�s7�� �j�?�7_a=�r2IE�)���x�lW?Q!o��n1�׻a#������0�H�/����4,S)��PM��ۣ�}WH���D�3o�J�t�՞�T씸�^f!*�H0�)����_����VdJ,���D���P}%	�NU�+��(����b�����q�5 ���׹��u9�}���>)�|�n1�ήr�������Q>��<)jb�`���i�"�v]_��hB�T��Ͽ͞B6J��D��������k]R9�(�-�f��i��� ��nsJvB۾?|����&`D^�0��^b-��(i�����@�&�� C8�;��G �10~�]�Pus�|�NV�A~A�NVSNV�F�r��;O"e�1���m����$
�<��a��A���2���`P�@���9YE��P=tX��Im�\�������)�y�����j����ӣ��$�v���g{`˻�W�����/���x��"���F�_���rP	�$\y�+ؔ�wC�����i�i��$�YPJ���GO�g�)˙[��q�zs�q�|��uR��1oՔ�r�����wM����LՐ��>tZ��V�x��'u��N��Ũ���%@:j{د���@�����m�g�����Qf��n�U��i��Uam���P��=�Б��Bi�cizER��4�[�3�j6ַ�/r��8	6� 7����� 'vW*���� ���ӆ�BeK�x,���JZF��lӒ���T�H����0]@7*�k��Z{�j�Ei8Q���KԻ���z�h���MLH��@���3:lՁ]�@F*��N��sH�G�[��v���hu���f� 3菱�!�	���yȽ;L�&�������<����·������7��L@������F~�z�A�)�$�q�JUaf`�w��pV>b�1��ؚ��$U�Xe�����W9�T��o�����~$�����У0<�o����V�v�B���fS�浳�4[Ł�]�L�g�hM�h[[IY���a��[��~����Eto�t}z��� ��ho�o|�;E��5��J�wG7"�2���7�=7z[hx���5�Qt�gy_��N[�����j���i*�>��QrҤ�*�	������Qz�`�}�K�W�(ԍ�A�N�Cq�F����n�y���9�:e�r�ä&Զ�2���+��6�0ɠ���e��,�C����Y;��9�g}nn6m��l� }�
�a2�)O􎯢�G�ǮKǄ�w;_�t �bѼ,��W�͙�@3�J�]���Y �?���.I��.?�K0`�Jc�	HC�1��Ȃ�W���1�4��v1q���?���#��V:��R!�{@M��ǖ'X�.��A�	�z�~Jxs�\�����U}�����z�]>�����Fq��f>��
�<��e�kJ���W?#c�R�!��C\eM��Έ�o,��v߰.9uV�>e<�n�J�<��_	|ڳNI�ع/_�F�-��]#�G��gq���g����v7K�o*�F���o=����%���j\;��bk��o���w��UN��k�h;�}i;�N��EV��{�ֈ4���8ĸWݍcM2u�md����
\PӖ"�M�]���ĚLi!S#���5?.�,��8�������o�ڷ���t/V���e�"�_�������[��|����ind��P-Kgf�r�Gׁ�{�V�{7��i��x�'�&-��>3�׵������;���кP��&�%�nm��� �B��CRJ�����/�b�*����j?�/[� Ƣ^/g�y��7S����qoʓ X�~u:V/i͗ɢ<e�n�Lr�|��=rC����B�w-�}�N�l�������ܝ�n2�������A��M3Q�J�%�ĥ���m�DbH����Y��׻���V���iڶ�;7]�r����IO���?>�M��1�k�͠)�������N��+�<�Pl������-y_OC��W���<�7~����J<o�=鼛r����3p�t���>@���:�]�N���]W%��tN#*��?�p�����ߊ�c_5��сj�b2޽����T�6V��=��;9?_�a�W��|�c[:q��P��|P��}d�S�] �Ί^vS�B�[澻�K�_9�v�A����X ����K!2W�
d*6}p�&O�e}	��,�3�PɁ���EF8��h�ԅ �յ��e�������S
�ǥoȏD��[��r7�',�BFˆ�2s�?��,��JHHx;Z������eI��ѱ����ޱ��1$�8H����H�12(i5�ui�q+���7�VD����jYy�u�����r����+g��O�{&l�_�a������k�+�4��i���?�A�K�䥛�D����E@��d�8.����dP�����q�~!���P`�ĉVjE�J����e���O�Лu&A�_<)�C�!y=�h�1J�SFp���e��+��5�����}��£+V��ݽ�r�_H�خ�,}�,^�Uꩬ��O�G����9Ί_n��h�be-�}lKh�._ }J}���#3���LQH�A|�)�oj-ij�hkv�lh=a�ڏ�zh09��2 �*�Y3 �c���N������5q��#��˧_+�c�k�9��Z�4�|�����}�uQ��q(c&���M�9�6��/;�%|2(��wa��H�N��%ˎw��m�E��Ke�E�$%��J-�*��\֔|�C����(<�>���~���xs������m_��q@7�����O|���n�lU��I��v����̪?�tC��k@�Λv2����Z뙒H�:�ъh�Rؽ�����E��ڇ����Y�� �:��$��U6��Q����{����Dі���&�[���f���H�K�2��%Z�CC�$m ���%�}t^z�������|�f�P><х*��L(CU\�����!|١i�gf?��Ј�-���L��Ӕ�������%ݜv����-�:*Dg�7f\�]���+�*_�5.�+��Rl�d		/��{�cSA��zUf6R�g����e�5�4�,:�,,�V�W��m$��:��j��47�m6�yVU-�Qf9����}<��=�|�d؛�m_���Z�����Žǘul��X�ު�����'�� V�,��%�N����{?Q\�P��j(����9Q���\�e��D�5���S�}��Nc��i�J,����7�umuwV�'�V�Or��/���NR��s���$�|���2�����W�+9b����IM;��=R�����lz���H��c_~$TЄ�0�M�w����2�h����`�V5_��.�kb��[����Z,,�,s��ק��*�썽���n�݀)֥��Ve���wi�eu>��5�qDK۩�gz%c��'A�*u�	�
��o��29K����i��s<��~|���$��&�����1�=� ���XZd3h���BV��)zt��a�m.��|*!�ތ�Y�9WI��w�Tբ<��xF�Z��KM�?����XI1呿Pa!m�^ыAt_0�ԕ�����x�k�Zp�[�u��&��4��.��y���M�6�ʺι��~�w$�fb���_÷k[6�Ȣ
�xV+�>�S=�دME����L�
ԳO�"Ry���Т�gSӉ��o�[�K����}̔����z.:γ�o�t>��<ܴ���g4�_2V,L�F�!H�2��Ŵ�F���lW
�����R�N#�뤻��7`��n+)�ef]�8Ro���?[��E�n��B�ƙ�����&��ۈ������qM0��P�f���E)�%p5��Rk��ȸ7#\H�ę��@������S��ևP����3�g.�9��%e����C�����}y㬟�+g\lӑN��P��R�j��~:@�9A���B�aj7E���H�th�{�����롏^��nc*�G�Ӕ-Y�M��޻��m�^�V��1��]��G%b$ݎ��	���	�I�F�Dj�'�6�,|����.�'ķ����T���%�v�lj�x�������^gͿ+~{�Nϲ���Cև���v�����ߣ��7�;�2�F�ŋ? ��7J�65���K�����-)N�S{����]�-e$b/��[�ݿ�(�V�gr��Rr:o7Gqg9�W���F�����<)}�]}˦Z�zk���>�»�`�(Cg%֤>L~��>��ۈ���AL��Ї#)&�Њ�#���A��S�x�dH��f"U҆{��b��hX� ^�O+?���j�h�lUBAB��qN>���h?\x������D'�CJT�d��a�d�m?%^�h�y,L�xv�a��S�H�?˄2H�	tS%TMe4C$���.~�6uG�?PNc��j��ƳP#.�������p����V��
@5��iX-'Ӈ�g9�f�q�5h46��ܦ(ke��h_��c��/>�������&T�*�}Q��7Ԃp\جf- S^$4g�GlN3�s,�\�7��)N+G|���a�Z�^11;d�UсȤYpf����I�]3~�_�zI�c������1ʢ&��l��h�hN��P��*i��s-r?��%I'��B�+��-�
��}��f$����RZ�[�\PhF+���I��=���>F����̩WH��d���Ӝ&�·�hB�F��ّ�n=��1�	��(����'C5q���0����w8��Ct������*G^F��g� �lR}٤�t~� �쯘u Lwl��TU�s�tc��d�ҳZD�w�/iK�F?H�-�w�w�W�?���h���:?|Ϥxn��y؝���l���E��������u��io�0eZ�wD�W�
���;<�ӯE0�H��!��M]���Blq)e񥃤a����_=���0�
0o �j�"񅯂�� ��Ά?	%��1���_�_!W��g�0TKh�j��YLO��9˲���'���t ١�P@�s�����εvM���	��Uy�?��J�����G�E����j/��z�C���O�94���pa�����"J�]�b�cd*l�=�G�-4uw����<���X��!�$��{�8!��J?�����$OP��ꮑ1zc��!"��1��;�~1.�ґ�X�W��ޞ!�'DO��m?�|8��~z���m�|8FblS��h��}|��<����ح�=���j�U�fQ1p��<�YޘO>X�ޙ.:�X	mtu�;ُ�i|�7��
k�'<�v%��_��7��8��ʾ��0?�eW����_&X	�
i��=K�O7�pۘz8�b��Q�W�R��W�L�
Y�i3t����D"Ϫ��p;��� �5��#�{�_S�6g��{�D�����;�	�
� c�}��L��kd���T;�2YY�z�u�x$|�!|�9F�$��PD�'!����A�~0>E�}`M-.����a�uQ�yDل{�!$I�R�x�	M��L���_�����������2��W%�k;;~��"�0�z�ĦZ>ǡ��e�e<����l���$���{���[�\[��ʏ��O���2`�e�����Uc����ׯ9:�_����r� �	��}/q�2��b���$��*(����˩�)8�@�^}]�Zd���d5�� S)|V�{I40��?f��ወx��ç�N	Q)y=�C�FW�SG�I(2|����C��'�CB��RL�b%�v��,q�"�{�)����"�.'�6��?B�T�{��l2�u�7"����\�e(�\"������^dO��	����܁#!����-��6 &t���/�pll��{���Z�:��p��`�}X�>T ��)iA��im�
u��m�X`���\v1'�@]3����g�i���s��$��45���&d�x�y͕��"�}��V��7$nO�ϲ�;�tM��Xv�j�n!ccՌG��wI���-R��K#}���cZ3���64�:����+oHs[{
�_�.�>��W^;�������[� ���<���|��+Gj~g�&gxkB�P�l_��@mJ�_�DH�F���<[�~4����ۺ.DH�qcDT����y�BLeՏS��	�� K���RȺe��E�p�d�wh���L[j��9K�J��o)qn_�-Bw����Q.)�%��x �LGՇ��z�t2�>��ǜ�%a~Q���A��=�T�pkt�Y�0�uKQwt.�N��
(�׀�R��F����M�����av�Ҟ�D1f`$��_���-�`�sd8��4�gAX� �1�8�85��4��������맛2���?N�G6�w��Ǐ{)���&�>�w��a{E�@���5�aQ�aA�J���8�����O��m�ſ�(��P�V�_|I��>�H����f�u�Ҳ;�i2i����&���hn�'9��y��
��\�fr�}�����#�͵V=�⊤w�/�@���g{�凯f�Y�Cj���Cy	�����x ��@��ͳ�7�'��c.G����Z�7:Th�I9�SXΊ�)��A*��y@�l��6C��T�(EԚ�]�)w^��[�=�,\HY)��H�����4
��(�VR}���_9JS^�&2�޲R���^�����J���e!���@$HA)� �1�R%MO�w�)㈛���B�� ]X��Q���������;X8!2��du ��?��v/�&V���k�����U4!�e�|��ޥ�SZ�I�+�Q����ZVͻ�����ST���]�|mP�Iۻ)l�ȼгH��B"s��r�g������..�fE]ĭ��uz�!(��AE�DZ���n01ǟ@�<f�e"nf)����u>#.hp"�PGq��ř$d.�v��2�(�Gzy��>~���}_���"����>N��p�������������H#H����L�5j�빑��~�_�7�-5i��������7�~8p3�T���7�Ƶ���j�����,���T�v�hMշ�!�X��pe��rm���8�ox�&uV�`�����+>�q��>��q)�ꈛ�7j���T���a.V.ܥM����v�K7�0RW��j��g��8[F�a��J���x�*v���{;X�=��Bv�Bu����(��h��_q{��~ �~��� $��r+�&��W�^9�ޑ\�J%4p5���E��%f���U?g��������:_
|��]y�ݨ�%oI?|-�S#�Fь�����_�=��1Y~����kL���ّY��z��_0��?�&�}	O�B��ש ��`Sx����2���s�u���œ��`CW|���~o�<xr��|F�y}]L��+%��b2�/�!!�`�g2�˪�mŧ�!!�{Z�*���@]i=��T����-�>�3Pr%�{o���IP��аu/���-dPT����h�P0Z:%�R'j�&�HRi����BeQ\뫃2L��^��H塷�:J��_�]�&1-up�~}�#��w`�C�0��ƥG&$�����g<�W���IUBL
�r�i�1��%�<���k7ť';�S�V�U�<��ꃤ�$�=>*4�)������3�[g���G�;�A��c^���	W7�@So�h�7&���D�N�r��v� }#�wJ�$]����=4��c�n��q�r��J?��/u��w���@rO�P�B�5��vx����D��o����im:���O���%^���^��g/R��B ��8���ٍ#���|�i��t�I�+}{��w1���B�G)���Ǭ)�C�X��妊����� �"�GKyYw�/���N?�2��O/Hu��9�>�9������yŶlـlV�lI�jL<e X("���vd�*�\��Lj��j�
�Y��u��lhG�Q9�����FT�E`(��4�kW�.�ӓ�ܛA�[昌}�_�Gm��� ]���f�����{OL6M �;^Lc�A̦��Kg�c��5Q��R�U^.c���]�G7Y@��O�����Q�CqQL��F����5����%�zr'��O�����B���Όвf�T���\�ۂ}^�v����_�X����غ����=t��Xİ[����h�%c�y(U��� (�EH��1���5��톚��5���!���0����.2���I��y$w�+��z͡�EW���Ò��Ò�C��+���]�,J�4�,�O9����.��S�镅b�Eڢ`p >^*�(��nq:Y�A�/HSrE
�l�.��.Y��y�pݗk�k�u-XR�>���H��mqn��,=�
�Q
��"Y��-:�4�>!^3�����G�a0���]"S�Y���ӗ�A��_��O�������~��>��:������f���S�˒����u��n6�q����]x6ÿ"t��
�=��;!QI;a�ee���urv=�:[�F2c�(�t!���o�^���0d�\��\̭��vШ�n�"��%��⅌��z����7���2h�<~.��7�E g��<��jq��|�S��yCk�_<���@O2��=yJJ_�	ۿ�/]�0�q����1���P���ppABQ�Y��]�CB�3�'-B��h���y��t5�����/�[Q� [ҹ_~��p�J�yv@�y�}-񰻿mmS��'�(����K�^�#�t1���+��Del����sUZ���O�/��S�u����`���{�����-�{BB,U����*�ߘ��A4��d�\I��%2�EC�?��B������+�FW��N0q�����,N����ƝJ*����TP��hjA^
۠8�߱DV��-A@�:D=aL�}1�\I�厱���n���^��'Ҧ�}��+������ZF�F�f%1�0W�2h_i�����`�������!���;|��� ��~ �10���ݶ S8�j;��K8A�K����kcj�����m�ʡ)�G�^r�����Q��ӿ���;w�9����������N؁��������ޣ�kW���3���lʎ�&�9r
]�o%����hCvI���~��]�>N/���<6pa,*��r����Xɖ)"���px�����Vǎ�����V
�k��i���Ɉ o�j��X��S�1J�_R� ��Y��>5�}�-�Ky<d^"��r���,ѿi9��$�F�4]iM|��}Ix���t�,BD��F�pG��	��1v{9{Ц2~��PUl�,��u.�N�+���ń̓�ڥ �F?��a�Z
�E.E4ye���4�{��Ȟ`��7}�*���0챺��"b�F��w,���,V����pÉ�0������U� 
�U�X["b�z��D��Be����E��j�';��ڄ�|���q�!��EA`�S��Emȶ�a���pA+�eJ
99���Ϩ�[��j¬�ko�R�ar�3L�L���ȆeK�B�~t{>�P�|Y#P5So��X�$3J�m�i+��H��	�q�Y�u���e�A�6�p��jH�?Sl-8TO	ݦa�M+~\�-`N9�A��u��3�L�A�WF��Uxzt��RNo����h�]�c$��8�q�[u%�a>P�2z_�w��5��I|�>V�hb���'<�I��2���԰�I^����"����L����ϬI�ՀrӲ���]���vN�cq��8~�{�P���X�&��Ō�����&�(#~~H?Sk$�vd�7����{?z���%����@�Ev�W����Y�� &=ƫ6�x\{�k?�����J���X=��7�:/��W|�.�W�GYS|2ް(�𒠊�(�	&����/Sşj����d�?�.�"��c9�.�{Å	xն�s��~�%���T�-!�vt��:�k�u��8�j0��U�����ӵ�ԵT[�l�N�ȭ���\��&��|����R]&e;>�8e� !����c�3�?!�r�����̒z�B�ݺ'���nGl��آ��VwH��(�L�g�߸��g3�2b������h��³��,�/+���jO����KZ{�m�7��>�����kg�үW0�Z&�3�i6_}��G��8����,��^L�\0p@��u-��ox/`-�#?Rp�pu�[�'q���3Zn�Td��CI�[8JT7�M�đ�
��؟6��T��nD︛��}�4��8�?"��bp�A6����a���i�����M��h@�z�C�Pb����`�6��i�P���7WFOl�T"��mhk����^�t���p�<A���4�5�'���C� 9j�%�q�/������B��<�f$��9;޻�ݎ�%%�bd���!7ѻtB��o9r�?N��: b�#�Z���10�����n��#$�����DU�͒d���\6v��՛y�����/��%B��U_����/]��h-1@Pj�F�tnt))ݩI1`t�tJ� AB)QD��9�w�������<�^u��u���&3�㙹��]�o�̵k��.�{�s��7�#�!/�2	!�Yρ �BMl�M��ܷ� �E�ͷ�=�m�ǘ�;�lv8)��r�V�U�ɘ���^?�Ho5�b�8�R����R����p3	��/@��M�
&d����0%�5zL�#s*���֏��>�P<�@ �[)7.����V���w�Y�e�fSp�v��9�@���&��K4�X+S��E����՝}�d�>��#��?T�C�B�+^S^Q'9����z~#?$��©�λ�@n}��e��Z��]��6��Y߁/���f�`��6v�^�Iު�?\��i����L���~�m���ݡ6��C7�i��F��E�)�������i��l��S�A��à6��Ov�����z5nh�*+���ߺ���~z�%{���+x����"���TU^*4q!���E�g��R�$��ss�S� �ߊ�υZm��D���z
S���Ӥ���Y 	E�E1t>�HDv�|��L8�Yq�R��n��'��h#M�きw8}�������y�Ԓ�{������/�fʧ;!�Ֆ��L�����@A"M�H!�>����uWw~k��{A���(�Y��8� ��9".g��~���
=a�{��0��@�G��/�-.]�W-��%%wR۞�^%a�#|���S�J�I:�L�5٧���ĉ� U\���]���ɲ�Or���I}��!w�m�{Z��ϵ\��O"ị��˒�������4+�2>g����Уo��A'bV�S��ᡛ�w�A�c��� A[,iv2��QXָ���{�ܖ�ܠ��;'))��؁Y�_혁_(�*k�o]�e�@��b�0Rƺ�ƞQ7I��<:�V(�����(7����o/�|ͮ�'`�j��7���w�/��@�%�fVT���6���z��2����[��.Ya��oH<5��&�i��d��a��/kYaq!/�̀�*�@{D>�1��v;0���IdcRY����T���j��}ڟ5�Ϩ����V�iWf���>,+��,�_�hјd�%�A���Q"�N>u�Λ}~ʅ��_�Ot՝5�M���j��Ҩ)��0�}E�U���KV��l�3B��X�s��g;)���ud�-�4pb�#���������9�e%��=ϩO�S܊ܽw��K��J�}o���:� �Xfh"�|L�X�b���f�P8}�RBh=S&R.;�$DL&�D��D������q����}����{0�}�Pk���u�����f����^1C�N�U]g�iy]���2�F%�B1��Y�Bo_�/��Z�'�^Ԗ���o~?=h��	./i���@���4��qax(BQM'y��P:4(�,��ݠ(=y�Le�"�V��OS�3����?d_�N>��(^k��yO���}��s����=�3�,k�l��)�)��]:�h���5��׎��2��xX1��T�����b�h�ӓ���%O3��������R�xL~�v�#��vũD-K|d����X4n���D�I&�{�1LxƩ�TJ�p!�1���w��L�5�����n��M �����W9�*ۄSwҫ�k�v���7;1{��XE�����m\����@�������џb�����'�B��Wǹ���Fd@�^D�-M+z��Yz��ۢ1=�~�1�8go���M��z����2:��0�G�����ֺ���ۘ3e|,�+=�h2�Bp�=�&vkc�I����g��p�Qa��$���jO,E�,Ix��T����Ef7�O|dn���B�Y���ѿ���M-��3��e������3�U�uŃiP�WQ�٬M�M�-���rH�<j�^�񺶂x@��A8��(��K�j��kL�n�p��~�e!'�m�bȁ��G�t7�4/B૬.���g�H���i���
̽J#�Bu:�M�w��j�s&!]x(PK�i����2*;����F�$L��i0���y鏤:w�5ɮ4K�Ո>o������|��mbT̹G�9��,�V�E+��H߈�ݒ�ʶ��@�?V�z粲�m&^��t*�ᾈ�����*|���IR��KT
NWU6E��#����VL��t/d�s��	��_üU� �#�t	#�Ԣ$_j�p���O�p��=����a�E�/H(�&�%�Y��{��Ȁ����g<]p�{s���d�#ɀ�y��'^�y2�K�¤�`d�l?��q*�p��kQe���X�/�����)sr�D��&(��r�X�h�ӫk:����|�M��u�5*�y�^�D]�Εݟ�+���*�>u�;�����m{v�AT?�~��`3]lN�6�{��p��D�)yyԼ`��@�L�~)4�P�?8p�ٟ?mv��̔4s���&8��4�q`��C�G_>�}[��w`;�Yջ ��ђ��N3�jgha��W��ݚb?MrPֲ6ʞW-B�X0�sٶab[���܀�>Q��f<���,�j�/���a�.�S�
�D�Q�0K��}����m��~��ֶ�<7Ҩo�����B�^x����}r
s.�6֐5�Q�u��]q�Bw�!B����<J�TՄ�j�2���������$�|`��g����/� m�LAqe\�A�U�g˱��Q��嘳�+�t?>��jfүj��B���^��rA���^���}��lE�������zʷ�Zk���������x��V1�_g��z?����s��cN>�+�Ú���o���1��j�	�GsI#������ek=km��X��eƻK�+�*��������Սm՝��z��u���gn�����g����e~vߩ2qL9wk8#����Ͳ����!�a��6&�?��m�C�iF��j�H z���ΛR����i�'"@����1iHw���A$X��p=�-�Pi�Z
- �<���
��1���a��w�����O�[c]1g����R)G�#x��2��z:a�/�D�%�<D��;�c��	���̀��l���ŉ����:^~��VŮ^���| ���<�U�t��H�yy�N?@���J�O4�2�]l�?V�2f���T56�*e{���r����3���Ն	Q��A�ˎI��摞�."9�3QE	-�h�dd�!n�"Q%�C��#���;CQ�5��J!��D|�4��a��zy�r����ٛj�����!(�=P{T��l/m�Wǧ@a0�56!��6�[f>��c�$cL5�5�~n+�2c���/�}r<xӯkh�c��d�h���*��[Ρ�+�"B[B����K��d��P,Aq�M��U��E�/U��_ӽ���w���>��j�d���f���������w���?c����@���ˊ�x�����l�ɉ����fs�?sm��e}z�߭h�gc������x��ņ[$�Ϛ}V�X1�9��\�3�f�1��Z>�i�&�<p���%1��=��O2��fF1��4Ȍ���{��l�1���њ��pT�>�i���]�:�I�p~g��m�sf4��ft�YՁ��aH�!n9Ӕ��ڙ�7�8ZŪ*���OK[�yS�)��хC��۬���	���ǀ���j�����z�?CdqEj2pD�pG�J��ј�.���A��:�-O���H��h�6�&<�T����V��|���8槐���w^���k�����%|S���F�!��p�K��r���ɼ��<n
�~i�k�#_�n��W�2/f�9V���I��%�z���݃,V>�{?�(�Dg�uv�����2L� �-�0Pj8o����f�����g���U��A�&o�
�����7�ev�U�8��R�=��i�g�Y-����h���������� �H��J��d��Օn�.�o;���!Öi6�h��I�j��u
�k4�G�
S�K�����9��lE/cO����1뇽<�a��	�Iw4�qd2��EQ�zJ�P��A�=�ӝtK�F����y}��g=ޝ�5�~"����X7������C�����~�L��F��GxT�'�jiD=�IŸd�hv#��}l��'#)S'+���_:��XH�e��`lӂ5��Ǳ��{�R��m�M��;��ς(_�z�bpQ�։-�^j�zFP�L����m�S�΅�G�̛j��P]|)�ƺn�z��D�*Lno�6�H�6���C�Q���$,�B�����Ȓ ��!�a+�<�	�5�k�J~cn���=�F$���D��Y<�a��R�2�V���/���!��fثT|u���{k�#d�#�7��t`ĞP�.�o�+Ƈ�!�/��VP����6�����6^�%&~l���d;�R
0p�w�f!���7�Y0��(��Kw���u�*�;0]�F��/%���
h��K8?���/�(���L�w�q�L�Qb`V�U����������� \�\��s���D��C�7���	�W�5c��(W�Co��]h���h�a�f�/� .:$5ɸFJ1���u���}�x/J)�Ą��"l���m,h�����Py]�j�GC�#��ǃ����Q���m��t����������4o�!�k�����F{��D���G��M����v}���8�ȏ!9�P��`W���G0�D>x�HCҐ��@	�y<�n1�[-E����$��(����ca�}�5�h�M��6��;���R��k�	Xfm��+�p��e��U'�hRq�<g^��ŋq6&pQ�	߷�:/W�ׂo��V���T�ns�f.�rt<��j�֗9�.����d�v;�uD'}n�'�T|���] .����*:��d"?he;�e@!�'V�nzk�1s����פ�J������p盶���RY��9�k�N�I�GJ��`�P��<��Y=��Q� Ж+�&DL���]�s�I��BY@mA�GQ��������3`�j0/����i���l+&Ͻ$��N]�X-m��|�S�7E���=������B�@�*@1.4S�&6  ��mуuJ�aE�(b! g�n��������|fB8Q%�������,���5��a~&��F|�M��'YI_Oo���(� � ��B�����{|�,�AY���n�H�V=������� x��/�Ł�3�6�ㅵ'YY��o���┸�4)N5�OVg:�;sL��Ϳ����+mU�t���^�ҘiZXV}�����f�r0-�ycC^z��t4Hg��E�ڽN�:?�ke�.�ߤ��gn#�����E�#p���ᣌs9Kct�s�1�j$��.��e��tΚ�\XF�,��E���|�!	��xIY�TN��}/��^%�K.���	��
�̻�j����_3L�0z��k�OĽ��l)�TH���sT< 5�!y�i������t�[_�Zl���c� e+���o�T����s/�B�)Y�k�x��X�J�W��k�򧆛ߺX֩]\�q�W�$�+���=ϥ?��@����Դ[6�Ӱ;i�@�l)����/�9��~l��F������(L5��g�E��C�)����v鑯w7��M�Q���hl?x5�k��k$jKC�-zg%,w~�$�b?�;}c��p0������B���$��|��������>��p�����sP9J�w�x?�5�ڴ汷��Q�8�@�o9�
q�j`ᱤ��g��Jv���G�u��C�4��T�Sސ��ķ˟�3=�_�c��֏����<�T�а%�$�է#3�o�1�̵Y�6ۺ�^�nB��O�,��Z9��<ns!&F�!�8���Y5ݡ}Z��Oi�-v�
*����H�%�n��:04�ګ�Q��9.IFN�
�,�]�Ԉ^� 9l'Pr]3�ss��M1�:t9��ǣ�B�J���V,ݤ�D�+#0%_�ábi4;��)"�����{x�}?FO6��F����N���nU6�w^��}��٪��Zy�g�Ʒ[t�d>"F�ϝS�_S��*{z���oNW����y�!^vH�����<٫�_�%�H�kH�jJ'����_9BҴ`��~n��x0?x���t�tb�+�j�jū�;z↉4"w!P ��1�>�`������9O��b�N~3��
�Q\u0Z��b�%�-����s��gR���_���燐���f�~�#&\�j��A�A�c@q�&��l����^D���kԲ-��]��N����F)G��r�j�O���j7�
��?�!i b�i$B���e6$NI�CEN���^Fj��o�()Vh������M��R���jQ0R��\��%V�����$_��~�~r ~r@շj�8,�OE��oZ���N��i���M�E-�,�g;Vǈ}���W����?65r6����釸1sj;��z6Y�nй�s�Q�����J���a�eZV9����b�tR*�.��׷���R�>�O/������u�`���;b��=��Z(��7�����;����ʕ���j��q|��wd��[�U��P�7J�u���V�:Q鿽���g�h��,p��+q�H|��*ǐ"G��+��g�~��T��V�<EDl*�u�����y�Lk��c��{�f T�^'O?�A&�o��=דB���>�~�{�m�R6�ɳ�}w���7�t����|���&�l΁��y�w�J���O5үP��P�%����߿i�E�y=#֜���zn��Wݹ�K0*���j+R��Ԫ#6���q~-P�E����T���Ƽ�"�У
�� W�@�6���㘏THP�^����RG�U!�b���M�`�3v�������xS����N��H5�ٛ�z�������8�񮎩�'��R[,0�;U����)�:K��?|Ū���L�������$�aW�OzY��;�-$���K��D4�$0[C>f��3�Ҵ� ��OW��y�\�Mwg��S�3vq!~����&��}��[����Ht���{�F�B��V�ݾ���fc��y��/]I��O���K�#{յk&3�)v|�嚧O����?:��R�T�y7;��\�$+�:�
��׮o�
�t�껽tS?���~4��h�C�8��ٻ����J�+����/�$n$��ތ]�c��h��,�8��^�$6H]��曯�w�#��Uv��9�Q��L��pS˱�-��`��	9���u]p���v�E���3�Ryл��gi ��6JH���>Y���߮�>AB�;��IY�� ´_,B�E_���+�_*���x��3# :=S���I����j&a42��c@�%��XG%��+.�҅���Tմ���A�W}5��r3��3�ݳ�f3�d2��}&�&�"<pl��ߘ-x��s~{�oۇR>��?�̔��B| ��V'��C��yPQRkyqG��O�jO���Q衷��G�(��;�Ѣ�I;��A��$#^��у|�k[@�O(	�GE����c�����ўh?i�E d#4�ˈ���pnБ�Z�����,Pp�?Q�Vq�7�P
K�AaO��1?�#�_V����l�m�s�](T�`�i��m++��p��wx6�+_]cW'��;�w�.�z46�y�e��~ϧmZ�� k%p<
�@o�!,�Z^��������ɝg��Iт9�S)�z��ԏ���o�4_3���.�2{�vg~�����U֡�XI?�=w����md����ʼ*_��(, ��
�5��8g꺍��u�pͰ⤈��B4[������zy���/*�d���3j�8ES�99��%�F��	ٷ�o��^��͆��$�q����l;LH�o��S��UlFZ�֍R�P~��Qo�<7P-&�F�����$�kM��}��0Nyǌp(��P���չcfo�x[������k�֟b�K�}�okwA��V�bc�D�͊%�  � D��f�z��:)7�s�n��ZL׏	F�Mɉ��C2_��#D��7
��w���W��|e��N�+�M����$@�!�Y�q�'�w���q�[�yrټ����EbO��KeR�/��%��8��P(��qg�6�/0r�'I���	�>�q�����2V��U�1�]0>뻴:�Ww��۹�s�Ӂ��:��9e�-�RَS�O>˂�'�q�s7��O�t�&>�ٞ ���)CCȅH ���W�lB�lOD
`=�e��j�o����ҽ����3Cb���}���G%���&�O�������i{���*J��w��6��e���&�!N|bp҂�\��Gp���>Lg �Vp��we%Z���m�⦑�O'Ŷ�(A�"���SpЙS�l��z��� _� �B�� Z��Hw�A�{���ޠ����zJJ�QW3��_��77��n<����9� ,�|\y��i�|Ϗ�i�q�N���$D�@CG�\��)3��YbYn�=� � ��r���k����}����)��?��	��!����J�܌e�(��P�"|6��tsC�1+T��]M�t�U9-ϟ�_J�.���v��[E:�~ڭڀ�mk�~4p��y�ɐ���/�WMt�@p$�W������Y�����3d�����H+�r5���5V�c;�v�V��a������|��/%�L2�rzh����
�a��ᮎ�f�I�㙂SǑ�6�6��ݟ$F�$$�Ͳf��nU�:���]���W+F��k��̸����G ��I���gC�R:T�-�~komҧh��`a_��gt�=���؇��H|��#��w�^�Ɱjş�&Jx����o!a�q��o�z����R�!�)m��<���M�Ґ7�{�#ƽ��7�[2�NرT�Gg��7:�ő6���>��P9��=T� �c����?`�\�]bh�<F9�˸Z{[#�ũ{�I&ҶiV�yR�N"�� �Ǖb�1[����u��1y?`�B�[9�	9�6B��L#U��cĠ���`��h�QLz�5�K滨�������p��>��k D������r')w��d��t�|��4�P�����'_W/�n�i�lukM���{��:��f*0��:硹7'��g������j���;eL��_��N*V&FN�jX���K_0ZN�6���v>���:��ֳ !�U�Ǔ)�4��y�K�u�v���&�]4$�Ȉ�~��՟4*����o�+^���+U.�8g�Dp�y��Kjg1�ne%��dj�.Ų�-��朗������~ �f��"0��KU"#�t}H"B���INng���%c�5�'T�l���!����/�#x� rv�\F՜�	Xx���%�	�i��i9��v,��&�a|�hv9�ç�Aĭ�s�׫������_�5�w�n�^�Xȩ�v6�wP����BrYζ/V��:�wP�rM�ɼ;�Ꝓ�or>P���8��V���7GR��%I����C�~겈����NB����s�0�Y�Ċ$BB����{T��A�'Su�%C������)|w���X`�s��B��"Cu=����=�[�9��Ԅ��<��x�,�]$�#�Agmm��������R�'A��?PP����:��F]2?�s��p�nU��q�H�\���w�HS<�c����f~=����¯�s�\b�Y���,���vP
�^g�QS�$�ke�����ŇʲG2��F*f�n��~�*\Mo�|>�N>2Ec�~"-��m�4�+�ڎ�hȯ^�=*]��>�E�С����j!j3�����~�
�*����p�O$�JEh����8�Xҫ[���t�Q��n�,�/U=��yi�!4�Q����������ۺ�X~�@�},`u[��]�"�@�:'L �Śi��G"J�� ؝Wh��*���=��#<���"5A2JYB����֭��Q�{���(������
b"��#��z����bqh��J���R���!ZT�G��({�i���.O�������Eת�O��}�:P
���+)�Vc��{�����Ó�����(@�X�>_���	�@>�k����1����t�ʳ���<�5x����%}�w�и�>���g��ڙ�y�ҕ��e���oY&@"~�qu�s��*�Cey$�WXN<�+W��IN��1>&at �V|�7[/��o�&;]K�正�j�
x�F��af,r�.'�Q!N�����'�����|j�Y��h�rY�%g�K+?�r\�7��O��N��m՚K�ă��,������pzr�5Xʇ�H[l��Gt����R��~�%����u�6�s*^ΖX�k�Ƈ�S'뻸���~�u'���^�.Á>� ���ǧ(lz���w���&ΓOl'�a��@�
􎌖�����;��:�L����J��pQ� ��x0Q�lXݲ�s�b��:3"DJ�z�D�B0����?��z���"� �I�8ݩ��Cz�P���IM��4��|K�b�GcU�_��~/��k,�=D�J��@|�qR�yѮ���uc-��'�!�F��H�g>��7�D�&�z��~���XD�8{a����:��A�LK����ai���
+��W7�};�՝���:��! qY!������+|<^"+�)�ru�Qkx�(n���̂�g��奷��X�V�ҵ��Ֆr �R�P��������>�i����4���ܑ&��K��CZ1*�E��
�go�OGr�l��R�s5}���	W�&F� ���|qG�������P�=Y=��E�ylJ,�IG��j�m{�?���5rF��h�I������8�&�װ�a*}��y8��P�9]���"�%���!�s+�˃�&4�5��S�k*�Z�Ts
��"��O��	O9>�$��5����~K8j|r��	Re����8d���}��F�PmeSG7 ��ъ����\.\�F\7�]��&�~-���)���������n�T���128&�������ՖW�|��|�LlO��x��K��̲p�0�;�����و�"�_������ˮ��d�yA��^^>�~Dd#�q�3�Ӿ�I\�3�b2�]�m*&t�yK�����'#|w����%�-�ٔ$�ä?������Q��);�@�0�߈�� ��Tr���8i�@�����1�ֳ�����8^�QK�ʧ1&G���o�C�?i�k��jT����Jt���*��?>�f=��_��kP�PQ�,5�[x]kD�0�3g�Я�w���T��{���S'������n�<�2���]�^�d���xE.#-NK����S�f��!�9Ő��{i(�2���rUf�' ��^cu�D#�r~��FN���Rߩ��?B�OSQ4��<vB ʢ'�
0�B��|��h���:`d�^�RI����q�
�&��^_" �iFx�(l��C�j��9Y�x3�;b}�Y�o*?�_�}����@�I+/��T�f�T�!t��
���iY,�ټ��|��^�I�YRo_����r;2�/I��6j�cɐ8�>,����M ����8��Us���j�)߸"���ILqNՋӲI��t�7�'�p֨��>�DO
jy7f�ŉ�r���u���*"-xFʕ��Η,mF�I������
,��-��`O� 5hA��D�tE��q�rS�|���v��D�w�8�JI��$
	�ue�o���τ��W�o�\�0�M�� �K]����@�Z�z�K�_&}�{
j�����P-<q�H��t! �t�ik�8/���`�Һs;@w���Ĭ�o�U-�Y�(yܡ�,���@��Ӧ����n�Q�zBz���r3�A,6F�0��j̙�m�A����;r�͋�����é��?2n��6���]g���8��4n|phs�x�er��Y��*D9[��vk��E�q��3��r���E��9*_7�������W{���_�y����h����$��� ��-S]]�����8��[,g]E[~�(J��|�Ke0/_��n��`I=�*$��͒�?���t#�Y=��m<?��½�c3<꭬q��S8�O�Q���#=��㌊o�>���j��_��CE���'���<�:��L~ej����	,?�����k2�f��*����12X���K[��Y��)�"�����61}Q��W�D���p���~�a���1KXhIH0��zɵ�K��)c�S
��+����"*�|����Q���I����+B����@ ��ϼ}��[AQϚ�F�ˁ �n9~��{Rkr>�ԥcA[���9 R%|��32��RXF��`��~J��$4K�ƺjY�νK�?���9�*�I�<��:�i�X�
�$��}�������i؜�Q�w.)���A4C�0W+�0RE�
���o��G���m��kA筆yw���Y��맗��ܰ���Sy��߸�ٌ�}�a��	�Ї��#�"T������
h'A���{��P�Z�$ܔ)����Ӳ���ֽ���&���,���v� ?����b�#�g��u��r�>��5�:ƈT6�&>�^��.�W��7V��Ac��W�������~W�O��s�Ȭ)�
z�]LP�R�أ ��.uZ*��>��^^ԥ  ���t`eAQ�@U؝����l .	�C�̑�,Fy���2�P�;q�ԽM�e�-��l;�Rh���Op��=��4c�?�)�S�MN�A˰k��Q��1�2�iB`�S����<���4�]R���l�7�>�f[r�����h�t+���s���}2+l����zdT���b@b8
S�Q�410�ɭS�ؠyIc	`l���r��(=_�*�x�CŠ)�W�����Z���K��c�@�K����J��{����_'e�*��Um���w�k��߄�-3���27
zi	.n~:
T�l�l��l�g��j[b)F;L��,�iHL��d�����VU��}�u5M)����sYL˹JX�[�z��8raK��3�2��v$���|��T��x�����y��2�������e-�d�grZ�څ'/���ěf�U���S1];�ՐpQ)<���s+(9�2�r����"�W���M��<%���r��9/����	a^���.8/��O��t�I���"5L�I��@P��1�jI���FsG�{�TΕ�,Blt�=����:@�g�S?`
,����c�����8�ߨ�=D���Os����KΪ�ڏ
�H�ikz�l�4f�]g&���4xxZy^�u�e
^%h�ٯZ�{n��}P2��e�Xd�y4j����?� ��ڝ{i$Z/��0�|��㼃K*������E*|��r@~H I����"�c�2�C괂��G���ρ��d��d}�.$��{�>:�73<!_��'$
�	�]��#�76­lP���Ge8~K!���Ze;xΥJv���7�L�8	�?�F �#�8i�y�:�Xyڄ�$��jB)p�n);� {�r]����N���Ź��w�U����H��������� С���qy}y�Ⱥ�p����� %C�.x]��F�$��K������p�j���emS'W3�Il�Z�7�3�v����ɈϬ�jRP��E���>����,.ㆫ6��⭟M~%���������&���X6/�o!v���	�t��?39�������l��8qY���֒3���~[ӡ�u�`n��x�j�����{�v�0�c�Bx4i"�b"�Y�Q�}��g��_lj?�m����.�T��\M�ʐ��Ӏ���x�f�g��r&/,8�k�0`���̢� ���_I�^Z����R�Y����΋m��,�误�/_.o�m+�)i����7��o�g1�1
�L:š,bv���� ��S�0�o�HQ|w��o7��r|ؗ��R��4�K,W��a,���~SՐ�y	��z�jY0o���g}�S1m�x���GJ��Ϭ�q;fڏ�6E�wO�bWZs~������e���,�x�1� -i%^d>�V���"pF`
��:|aS�Ēb,}@�#Wؒ����.\�d�>�C���w��g�G$��r\�Gx��-��/�����:��q`h����<�܍2����Ȗ<�;��&b��G -,IM��m��&�@��PFq�� ��,�v �D�,� S!?{ j�U2�\r�j/CĹH��������o���+��ʖdk4�gR���HX
M�>9���q�!�U���5W�\�U��:LbgP�����g[�[��S�#����2�~ˍ�Z��f<�k��;O��^�>�ہ��r�r"�BvN������D����j��� ��VT�`��~>=à��e�\�.T9W�������C�5��o}�?��[ݨ��S�d�[7�^G�#ŷq`���燂�{�y߅�*�wD
�LHųb�?�^?tw��'�$㽙�'�/�.-K���?2�	~�����TʬO?!�@u�
��' 
:T9��W�_�[z�]���cPJE'Z�����5����l�����?���C��I.ۺ�3� BB����f]�V�Q��,4B� �B���.�+z���v��QZ��STR��C!y�'���T���e���;,SR�w��ܦ~��c�O	�ކ�!�$Ɋ�ri��`T���A�U90��(Le�����I��_ܛޠ��o��]<^�:�5�ظ���{�ؿ�v��S����1���Q���q�g��N��*N���:��j��\��mi�EC�|�SӲ�u��������I��uܒ��Mbӽdʝ$d�QQ�&̹L�i}P�qn�p��sF�����9�mFE�j��W��;�/Y޳�ݏ*-�2�[+����p� �fr���]�;L����w<G���Ǚ+p�(Ne�m��!����B�cZ�K3SJ��*/
�ۚю�]_oA�@��5*Z�Kϡ,���Ҫz�;�m3��P��}�-V"�/��d��R2���l�m��aP�'�o���d�a����J~�����܏(�#��ӰIڱ��_:����N<_-�Y5.P��Q�GCgMw�,�yxA�9��i}s�f���O�u<t����0�ov��x�b�|�q��-N�?�(ګe��2���#���̍��rm����ȟ�!�������h=��ϲ"��p�>jG�f^�f����z�����@��ҿ���~0��#��W�J�l�%��i&�2�{�
S��FQLh؃����,G�i�i��	��Ș���e e�G@��>�}=ʛ���n��{��Љ��Ċ�u �:V�����C�)!��̈/�͊Ⱦ
����S��j�6�D�*�� �!��<n"l=jY�"����'�>ӥ&�L�X��b��n5;�(e�=�qj��Q#:�- 0uNx%}-�̒7=�VM9�\y���b�yM���O�ǘڹf���K43
�S�}�:��c����{���.eb��DPu�Q�S���H+<{��!���&���\��{g?WgeW?5�N��S�C������Q�y=�esw�;]����U�`��&�P���kR5��Q��?g�$Uܑ_�\�|l~�c��~4{����9|W���`^�����0g��d�#���Iĺ�$����ݭ���i�Y ��d�t��E��I@�^0�q_�����!Z�_��*�d�?e�#^TdQ9L���"{�{h9]9��t�K�"�{�G��ٖ[�V]�HK��>=��U�~�v�4��<r�AXA_�a���T���)�"P�'o�������䘻�p_"����̽�$ҹ�|2V���BY�!zF\H�a\�)�ǐ�k����0��r�n�2�^��ʾ��+�N�h#>�*�'�Cw��i����FV���"�e��p����:s��˦|�p��k���A1{�r@�eR��z-�N�brC���S��V��Jl�k�/�៥��.�qj���J���L 	���.�E; � ���d8�b�5t ��|�\��á��������%�ЖT�~��2��������b�2�͛�B��c.,_��Zn�3P|��o�P~��J�$��v?�I7`�+1˪{�3T��]�~`��N̿H)�~ ��<��Y}�¡�>�GB��c7J��S^���q��z	zDn\�e.��� ��#���Ӎs����}=C��N���o�k���~qo���"��<|�I���D5����Er��V)$ѡ��V}5�`���C�>�3M�<8I�=�/[Ŀ�tG�F��f�����IY�t�&J6�2�A�\>�
M^�J�κ8��y5�4)�s�=�6��R�l�֪r�o}f�{���G-��!io(N�g�đ{Р�l㿺� \I�HR��"0�ˉ���'�0��8�!b�,n�Eˬ��m�v:]t_u��ޓH���v���&��g��4�F��乐�p���Hp־p�	a4k�yȇkc��'L��U-�e>��c�,���n]�@qk���"��]\K�P�xqwi	Z܃��/�)P���~������uF�9s=s��&���5�Fi	C�B�NZ�����`���}��C1�u�z#�����~�5���!�����m���/�D��-�	�� �F5���֙D��3�y��=���e��#%�|b����N�}_)"b�q��m��f>ǂS�i#l.����$��U�,�s�v�#�0�"K	d[�d�&�ƀ��ɿ~����fPfP���%��O��߭�a咲�A$��Ԋ���<�w�=+��'�O�~�%�_��**:�8.�w��Ά�'o�ξ��<F��y/�bbl"e-{��t��jw�l�=�*�z/��Z���v3!��8��R�B�/��N���s�c�gJ�X�
���Z�9������Q���Qǐ���{݊8iޟ$��	xG[=r��/�����	�q]�rAA$֟F�z|��TP����*Jc<���~Vs|�_lU�FK�T�fL�n��{����r��D�u>�;��������� ��"*F�Q�X�Ȁ�>&���Iǈ̃Z���uq��K�,�B�\Q=�U&>�}0��X �f�_v@H�X:}��MyK��m����`k1U�k��1
��[H��*hB*�g�F5Y^��{� �t���?ӽ)G@+���ھ�X$˳q��"��3
2�y�[$ЭYq�t�Q�����l�'U�;A�y��Z���]�"�Or:����.�%T����J��w����6_�Q���HO� �[�Jb6Ť���C�D�:�
�Qѿ��*s'�LW;�a��![�,�~�r=ۇ�C��W�(4<�@��+N��l{��}����[�}�P�{�ѨKv�7�7�^��0EQ�T�E"۪x���52&��g��
��k؟��rj���r�a9��EpMȡg�]s�@QYs�X3EL*#i�*_"r�X�ev �c��n��,�nԅ4�����X! l�7N6)�F�"�<�[�3N(�]γS}��71"���Ke��+��.�z+}� ��p�x����^�����;�f�.c�E|=�=G5 )�)Ͼ��!J(����G{�gZż�JL����˸j�u��V]@6O�&�QP�m�: �a>	Y_Nm7�u#�Αآ������k�_�`��	E�Ȍ����P��r�b�*�&a�^��"�U7�������[��3H�(J�P@J7��?_����p}��},��K�v�B��qW��ю}^Ҩ�����Z� E��D�`�k��,�<�Nk:E&dH�jB��S�9~��pND6���?�{R�7��T>{F����v�<n��򇃨�������%=�Se)�U%���mU��>�)���pڎ;Y�x^N2�u�-�>�m}�kW����Aw�.�������f���Z?V��Zr�q��Y�[O:|�wb��*:�.�T��z��ÇM�Ui�&Riq�kiGcg�w<n�<����F�І��X�BY�eYD�J��J����7"r?\..��N^E�����j�`zU����~�^_aV8�_~ϑ���G�.��s�(6r�j,�$:}�$M�U%�w������
�e��|T{6m�b�T���B�����^C������L}�^[LT���@y�K3oHp����\�������/�M��c=}�����?tG��&�9s�[1���Z��~���3Ju�I��l�q�k�P���]Lc{�}���K}dM� P:m}l�:�מĮ��1-�52�rL��Y/�s�q�e�W1i�wIu�w���q%�t2����m����M�WxpYW��f& �v6z���D�͝:J�,��.AP�V#l�q����f��Djʟ٧���4�Ԭ������9��qډC�=�J��D�!�?����i &���O~����*�j;�~��L���9��.�� #�I,�r�|y�r���鲴ԧ��͞$��$�%@�B���ά9ϻ�������Z8�)��珃�K�3��]Аs΍� �q+]Ѐ<S�>፫����l�:�˽�ܱ����a ����o�pc��v�<`�k��0�=
u��7�)�Rq�"�=@(���(NP���!N����B��������B>lFZ�l��[#�k ��Aso�\��@l��4���ouN�7���_D@��;#���]@(�UϚ��3��ͩ�4K��
:��Y�H�������y�+�i{�	��eX��5�1Q@���yj�c|t�l���d}0��w����83!��ٝ4ME�ME4�y4-��m�m�4��������<�՞<Nǉ=��dz��g�Hֶ�#ò�n�ے�]r������si:��t�2$z�`������:i���i��"�Ȏ�1]ڰ���Dk��$�2�`���[-���[�X�����s0#�vɛʝ	��6+ᢅ�H��
�o[=�������'��JB��|�
6���� ����$�W�[�e��
;�W�T����XN���u2��M�_�����/I������t0S���U���Xjh��(�bު?4���'�o_G��`?����G8����y�Ck�@0�P�{zvK�G�9x���[
{�˵%4����
	�ʆ�g`��乽j�2Նű�K�g$�fc�FR��������j/Dm� �/��M����Oy��_�E)�FsS�2�_2�\v�I��5��5�R���Eo<L����U7��ȃ�?q���|:O9���5���S�Ce��ߖ�rG���^}�v`A������c����_������|�'�ZH !Qʢ�t_&�;�� ����q��	3�
��a�(�(o��5$5��p� ��S�cS�}��2O[�4��Wk�5k��8�XE�X��_�IQe3b1�w���Qs��2��
Ƞ�l��*0�V�๩�7�����KjB��r{����j��Q�����z6�y(ϒ��[���ךmʁM�q�m��Xܹ<��w��p`*^X-M��y(��+��V]�//τ5�k�����EM�C�<�b����i c�a�،j̫�BT�����K$�����R�vg���\ԜD�����nϚ>�v�P��/�B��Q�C$���P�(j"�FΠ�`���~��;&�G!�q��zg��#O5�?��>�I���j����_���}S\�zj0+���J����3�YXY[��MHI�$A���[ل���$��V�!��y�u���]>�S��E͎�ז=������K�&�����
K����-g6�{�[��`�Y�7�W�>w���F�+>-84���Ͽ+���+�������eL5���JC]����"si�d���˿�����l�n��C��w �C?�����i�"V�Ad�E�%�\��P���)c���U��s�-^�Jj"�3o�
��s��Su��e��u�.~J����]IG'�X֬�lZ�ė��쫷p �-*K�%؃F���J�n�eY�:��M�Ru�n�,ˡ��)�!����B�� �^�jɢ#H�~NH��+$g��x�#����P3+v����!D�ӆLp�.6��F�����i���,���ט������
��u}����V�Z�66�m!T�Mwӫs�1�3�����j$0d\��#n�L&ъ��n�/��p5}��p{�P�b�6����>}�=�X ^����$ξ9��6e�z������������g�Q=ؐ�A>̱W.�	L�.	�Tó���H��%�d��ϤU���Z���|��D�����*�IT\K��!��z/�k!Q1�-��(a����&��`��>�_F�
�:K���C��͟�[����(�f�Z�)l>oω�E��(�sp����t�]�^���-o�.��N*ə]L��5���ڗU��x��W�.5.����T�We8��m�2����pɌ�т	�$�a(��v�o�Ҏ�џqhc.����8L��h��qw�������<q#(4X�vG���\���*ʘ6��oV&k�0��7"7&�{G��ɶb����(�?���kđȉ� ���-u`�wϦ��0u�x�J�PŎ��Cy�L|�2���E��	,��.�۝B�����cc_w�-)��
��lE��R�2�g7{������V�ω9���\eN�)ʊ2�W��I��K�R���q�"
xU�M�l�l]f������Sw_��h��|�(h��	��9jAW�٥���t�A�^ճ^F��9�+R?sE8����C����:��.A��1RW��`e�fV6�:
�F.Jw���: ���bZ1��3�3��#�AP;_0�=��b�q7 ������Hc��a.��.��quI���,Q�ᨩ�����~z�r_��[`��vv�j��_�1��x�}�\�Xᔪ�=��r�\6�C��(2��t�Ҏ��%3M|�Z�%X�V�'�O�^�"��A���ܫ�6[@�\���[rw0��L-2i?�Nn��c�2	��ֈ����������1�,HP1�kXJ��1g�uI�"�����U����!O/��r0�+*a���o���V�u�*5� ف���!�5�s�	l�F��sO��XA�������-�N#`��z#�t�"�Χ�պ��#�y��Y�l�?̜��r���C7��]M`xf�h�Գ�>��!�6	��L\����>-����<,�#c�~`���>KJ��7�/
F���cQ��e}�@��1��b�ajyWy�#:�؎�F����ز.{��~V(oL�m9�&�Qb��TV�����O�gPq��Ȅ�k��(I40]��R�P:9G��������!������u�t��Rl��|�)��z$fM��bXq0�O�)��m��sX
�' (��!c�2Y�_L��QP�|�f�.��i~�sӘ�ژ,�:�p�c���Ũ0�BiHZ�L��b_V�S�"��3�Ⱥ�.��-w���3��I���a��gx(N0v#�"�kG�BO��15����q�L��rEͨ?S� Ԛ�ʎ�f�s���{����3D˻�M�9�m����D/��m\�j�,r�jT��I�+��i�����-�V�h��NZ�ܽLu�*�鱐�QW����n/�m0�!��rI� 6�E��.(e��q��� :e�����?��5�����J�I���x��iOQ%��.���H��.��]F� +�ú3����&u<�~��%��xq}�p���X����C�>���\�}�Q���q�F�N��%����ɲ�$4L7��E�K����ԑ�$\v	��tY&��qS���8�9�+>�����3��^a��mz����,;5�ʏzƒʯ1��8�Ĵ�̖��ۋ���Ҏ2��)���N��Փ���'��K�Y-��w<�`��j�s���9��]��Ҩ���}� ��pԬa�@�%������Rt�o2K���I�w%c�s��g"��%����ʔ�e��{�όY9{�+W�g����*�0ɿ)��<����G�� �����}|��i��`,�S,H�V�ڪ��>ˤ��)a��C_���9���~}#H6���P�$5nZ���V�nbl4��.US�����g�qP�����L�î��r
է�SF!�ɛ�?�eH�;@?�Y�{��~�e�΁���L��a���"z� ��ގ�>��6�`XoK.�#�'?���B�@4�/��b~�fW��*�Ш�Ĵ��[G��@����]Z�9��A��+mˢ�`���z��"��rfeU�p;����ꡂ���I�D�0U��G��F�R����S���N�ϵfwQ: i����3=����;y����*��Ȉ��q��
hZ{�!%�>�|�AB43���v߭�e���SyTK2�n��y�(M2&�!h�-o�T8�<.4d�\����6H��&���ô��?�S(�K���A-��%�JQxA~�AR�(I��_�#œ� L"?��8_���d���OJ�Mg��g�wQ��RzZӽF�K�;�z91�w���'H��
kt����]E��L�v���9K{�K�Kf��_�����R����KG+�&�e"�E
�/ �?]WQˌ�v��V��5�	��G���|;|3�B,��[i�����.a��0���F��b��
hk��UP|R��v�<�z�.�ݐ�`�pb1�F�d��Bg�ԡ�o���p�KSy%ɲ-㲋��(/(�����{V�����W)mw#Y9�/`��R��
���U��rgy�$�tL�H�x��c�z)������N���23�E�2�����,�ȴ`��:�;�jF۞L&�k�ͯ2$�
���_��a8���S~�)�z�INo�.���x��e��)�-���n-u�d�0�AxϜ	2�Rb�;�yź�rzB���K�O����Ё�t�pE���^�#�h]S	Z?

�z
�m~��8dd�	j��Uf�%	(}RE�hS�����os`62y�*0x���*���= �Fժ^I���B�ʩ�V����h[��j���i����^AHp*�@�^�OX���"��;Er��o�t{�Q�v�إ���瞝�Qz�i������C&h�M�g7��}��'w��m�9��ߚ�o���Lt��?�_�75�^�8���'���/~�=Hj@���$w�,FQ�]ς�w~~U��L����Z�𚣤|y �O�U��_�uH.e�)��F���T�~�)�nQ�Z�0U[����@?s9���!|$����>
���ԏp~�>������!V]�t=;��ٶ:�	N��u�+�i]�]��rU�����|7M���v��`~��?��X2�9�DԏVʯ��c��wq�9�����G�!�؅k�����Ω�ԑx�P���ؼ�#�y �Fz�ճ'T_�8�>��I�F� B0��F��K��?M�|_��\F��K��;�/Ȟ��{�?�����A�!�֔fJ��V���n� �DZB��阕�Ai����@٢��b�����Å0)��IŐ�KƓ��SI
UI���B�[N�I��
Y&l�O�:Q�2j�6Nh6�W�+4#�z-$`��T/���O^*8�O[uP�F�@��Բ?5l.~y&~J;yJ?�w��ɷ��lj��9��f��:�-1ՉX���_���WXL��'Ƙft���Iy�8l!���8ic��[�������w���Ţk�l�l���Y��jդ���&�	8�W��-����}{, �
��l~�t/e�VB�De�A��!��X����J���g�������R7�if�@�W�Ä�X��1 ű��@@9�D� �SJ��5@�,�d��gº�HP�r��]�j �6"8�&�����% 6k��`$�?v��6���1�b-�WI��~�r���h�).����2�c�5�i�4�%�|�����re 7V��1���(�3����.�G,#R'���R��;�s���a>���^��s��I��n�k��� ���i������b�K#�B�R�,��%�w�fh6<�j�e*6���9�j��f� '1d��P�`�@I}��ƾ�W�z���Kvj�^�~!�X��0q����~����@���
n�=����h���C�����&��{�Cb^Eq���}|�MhE��:��~�
iF���0�pB|�2{m��ʂ�0$�)�����T ?��9:/ҁL8���|�����-��sg����'L�Ƞ��~���rf`�U��OBQ\��V��2��,2�s���|[a
�M�^e���8K�1�v���5��-&�6����d��Z�	���8ո�w7~TJ������������%B��Q3����	M��nN�����
d3����P�����+�	~i�Q탍�\_*j����l&���.66gC����b>v��+��F�t}�8�J���*��V1��Af�k��VV����r�	h����Ę?É���̽R�B\�L�_8h�(��M�*��� ��l�'8N���2�� ?~e����o��	}�� `��I�Q����NLMF�i#��|v�$Aߊ�6,����Y����?1�CȌ�U����ܱ~L�N�/
����+�o��'OX��
�9�al�f}	���o�P� 0Ù^y��n�&���J��D��[ff���&꠳��xN���嵔h pL�9�=�tzE'�'�,���_��*T�~��󕆿�Ŭe����q*x�J��Js�Mƻ:�kD�VR?�����O���6#�= �[���;�Rٙ} �%eD6NW�����x��0�C�u��$��:��8�/�.������&~��Q�֊�2:&�J��� ���ϯ2WI`��P�����D}��!�!c{��yZ�ߍ��@�C7}�eM���}Ǒ���2�˄�*C3��rs��.��������&�_Cv�1�����X���\J �o�Tږ�IHJ�&k���n�ma$p�����K�RDj| 
x �.M���!�-�-���������ZN��zM��z�&�߅z�N-Rg壼��E��aVR�?����7� w�+� 9�j�J�;(��9 �
.�e��Hz�RԂ�G�E�,)=<�LKb��L�qZ��pJR���S1�X_
�n�8ӣ����V�:n'�|6�r2�\��0���+�G)㪳��&)�D��R㳺��u_X��n�q!T4��M����T1�Vw��b��g}�ҧC�Pq���st��ޮ�t6�*L�c���h�uaN�B(�y��O򴔼 	���;t��z�g�2�D�GM��:B�l`$v�ͻ&3msJ�{P�هy&T���g���@�"���D=o1�q
P-����Ϝ��IA���-��㪃��ը#����T�0i�g'��`=��:`&����.�3� ���5XfT���g�Eݯ�& <�aG�xq����r�t��t�*�eu�|�^�@�Vˢn�St�͐��O�m�,6�u0�	^!�ז�7��[=����7;�/!&�*�ɟP��D��T�װ��6y�D�ZJ;Ώ?ad?���޳��Թ�9_.���I��r�з��5qUf[̍�1|��W2�J7�+�Ա��sZf�u���T�_(���erY�ʪ����V�F�j�t�%�τre���>���O^��jDLF^�e���A ����������8�8z�#�֞D��� 
�N�JT��uͮ��'�/��� &Ѧx
��A�fE��W�?,��k"E1�ե�:>l���BTyfC�#�D.�7N�)�+��S���r<��]u�|Ԙ��Эؖ��}i9�)�˝�'3�1!�0�~�*%��g���ƅE������rdM�k%n����rdQyI��#;��g߷_����~�u�`�HL�龈�MM���W�b�3qU8��La2��V���ōj��E�G���x(P�[��^"@P&K��X3$D�[68ޒiC��H��j�����Q�5h��H12dP�1%�[]�\I�+���!��.��|���}KiA�7���Z�z����X�� �jČ$L�>��I�<U��8��O� �=����8�  |�����I^�[�L<8S,k7L&h�����9&����P��Z�H�`Y{�B^H?�%��F�_����Ӽ�शȪ��tv�n�p����7��N������$r�%J"f�(��n�RKQH��>�%W�'�����C����Dд�f��`�\�d�l��v����b槛�L]R�Bd��M ւ�k�q���X&�B��_�/�Z��x�=���a5H�*�7�z�~ɔWD>���M���<�o�Y�r�وЃ^%l���t�l��H���|;�+6��L��z�d��y�x������c�a:����YUG�7=!Ԍm2��8�����+F�C�����5h��۫�XA=o�U)�w$$�{"�b��l©x��ˤ�K�f�Ht[\uʺ�`� @�#�&fF�GX�ԄI�MQWh���?o: �\���Q�j����՘�A�-��̔�!o8{C�u���o5���v2�v�4-@�����ם�'j~��'��|k��^�H�d�@���=��h}�����"��k�|�����U� �og�agkH��@���pE��3�����60������Zڤ�o�i��3~�vTq����5�MӇB-��4�C�1��<5����|r�]�[���(P�D�+�9(��IL���L1���Me�~*��9Ҍ���4���kq�2�ǥ6�z|��S����= Y��C�R�S��f�֮@cf�7N<��U;Ҁ��"&�S�H��$M�"�3���W6�Vg/��;;ͪ�2m�ބ���H0s�;E�2�\~ IP,��ib�y�AR�O1��/�L��K�4;L�7����J��p�s�e��d�!`\���\��h��w���8�X�����_,.��n.�x���ef��R�/�LypCӢ��-*`:?ϩg�ax�B���r�乫,�w����ó/;�d�Qr�k�c���
B�i� �
з���ŵ��Z�q&��lP_$�?I_���mĳ/6C��| $k���x-�j���Da�p{YOF�f#X G�͞� 
����d�c�0.�m�/����@u�����A�9 ��aV����E�ķ��W��� �jT��ԁou�	uv������8ntU��Z>wΖ�M�LU'�-�썧��}͵j$����*�O"�+]:���������Se��5IQ�� �[Kƻ+����+��2EKjgi �2�t F�,-���9�w���Ae��͹���	^��'un�p��d�k+he�HR�I��2�]T���t��aCw�g��LҮ�~aޠ=�G=�1fa8��5]�%��Ϗ__G�C�1�DR�>Z�g8��#�G�r�����Q���[k܂���0	C��y�b2,�V�9Eu�:"����Ia�!����2P�Y7B�b�\CD�]�o�L�o	=�a� �@m1Y����l0�&j8��idZÀ��oƱj8�뙁h��"}L�[[��:c��,
;��9@�L��J��}��ӝ���h�Z��>�I����� ���������1�.��� �4\�Y�}�_�he4$�j�fp.�8xҤ��4���8�jKhh��x~�{��X�������V�̂�s�H����3�VK�&���Y#��Ӣ?z),W��u��8�T��n��3{-S�S�U���L��E:i�g�j�����h��l�T<�y$� �dU'F׌�5��7�?7�v��u��kr�m}�$��bCkӿ(a�q��Q�Qw'u!�_��6װl�?�?3���si�m����i�<5���-�؋�&�m���_��u�/�GE'v,@�����N��}6BH6�Vφ�hAY��B�3$�@�	�^���x�m�E)���s�ede��CI�!�3c�{�Ҷ/��,M�S�������ט�
u�s��{�/'e=;�[���j�9����ʵ#�j߫z��L�%��[���gd5(>�9���/S�&p�߱�_�J�I�6�=� �U���Q��p����ұ�W0M��h?� ��I�ӾׯIa��YL2�op�5E�&�^�8�����$����DΒ(���@��UX��FaNU������I
���Y)�g ��L��%d�Ό�&e�چ+�mA�!S�"�oQ�e5 _TIA�s���ʂ�{?�#�KH�΍\}b<�zRBGקR��|M��>��g?����u�Y�H��S���~ܾ$��nlYQ��ܻ
���_��D�> {��i��>�l��0�" �(�^���S2��MG9�H�0���H>�H�!�D��ϸ59�%WH��=�,��~~�����e�����T�OX-�x�(��Uo�m_��M���p�k����g1e�#�5<Ni��z����9&�~��xN���HJ��Y3�}+������\��!��ޠ䈅��j1�x(Z��)��T,�E�m��IK*>/����.����M2H�����\$`�B嘁�=����.�����\����mVX�Zӧ��I�ZH����S_JݼV��iϜ�g����ǯu����e�������?^fٯ�|�n.Z�x�!=�_HM�4-x������4W�dŐ�n�z��0�,b9&j1&b7,h:��7qw���!�.��ot�����5�m�Owm��}L���L����~�d���k���_���'�KÉ衅hZ�(:V��?�6j���7ΰ�<j��=O38yo��WFC��5��#����$y#@�D��X}=Y�㗟� ��	� #���Κ�N
ά�FEǍz%���D�̿�m��F�4�=]���F�r�fN�HzF
sq*�"�F�6�fK��{��5������Ϥ�Ϳ���uR�h�W����7<۽�x峩p������}6�%y�g�wqm�Z
Q�?�Y�mɛ]����V�f�+�kO�邝ϗ�u�;ˇ<������t�h󫂙��~���ཀྵ����~$\q�?��.�PMô��E˱d�#���샗�c�̳�V��y�0E{����!c+�#�S<̅�Z+�f�kI��RW��ؤZ^nmZ�Bb~FM��^��k@��\��!t��El��	�BHO�4�{�~��A����*��� n��t'�P�E��4��j1��*�����i����<���]�k��}������vw�o�j�J.(����NA�s7	#�?��lހ5���\2�?򈔫B����U`ی��ӕI?�͟����xH�A7ʷ��r4ǡ\�{�f�;�6���,4��i6F�F�n v�6~���k���z��z�K0��>[ȩ_4a�`�g��6��=�唄ǂ�r���K�_��a�oI7�G$GO"�{-��~S�*�f:F3ň�/�8.&�i��_����~�d����������O�������$L�r9���^��"�m����M�_ܗ����'z�Ѱ��T�]�>�,&ٸA����r��̬p<^y�Q�a.9T�m#qLu,ގ�(D-j��@�*��2� �v ��V�\s�4����يX-�((�����T�vv}(���Vz��6*)�]4K_�$\�6g�~�*���NrǷ5d慪ߦ�QIK$�b*�,�<(�6:b��i��wq�M}��H����͛�}(���c��y��H���f�h�/���xq�����aSx�(��^l9]A)�YC�yG����������-�$2�2�	���c&b���%FI�s�[���ź����Í´�Ό�����Q����鉶�Y�F"l�XF������_���L'�Zٝ߮_.�%-��խ�pڽIdw�Q�FJ������vW��a��)��VH��糚I�&�RcP��nt@�5��7A`�Z���?�*���b�wRY�t�*sU�;�:]�njwqD-���a����G���;G�`�_�P@�����T����!M��h��"�9ȧ1ћ.�I�da���8�D[Ԫ�iĉ�p �ly��oE�����gv|�i��m�C^�����AƲ!YZ�es�e���A]a�����~4�~/����f[�^�,9[(��e�r��.��.4=z���k1F�P��!�^G��fI�Z�����I��~�+�8a�����6���u#]��$q��{��ܒR̖х�{_�\
Z�oNf��V��J�5*�¦Ŋ�Gq��{��T��3�z�zS�N��0սM��_A�KA�����|R��M�h�S� )��n@�uT�,/T�F��'&�$��D �����6��NaESW"цƊ���N���� �o�o�-�ZMX#��I�@�Ǥ���mc/a��sc����!l��"ġ�]=E�uʐ���̺��a��=������♰�pг�4i��敟���]-)$vi�����j�����Z|fu����]_�:iwK�Qx�7n�7N q�c�_Ϟ��SzQ6�� �|�9�A/zB��q{���W��Q���������ɂ�S����-4!�������Y�Ի��4�\�n�q�ewW�b̥���;P��Wk�_J����$����?H����A���=e�����OA.E\�g;�&�e�c��Xd�?�ަ��3p�/��B��&*�\�Q����\.�*ᧁiϐR���D��\�)\���Zկg,�1����m��IUX/E��{~���2�`�sbv贚�Z���h���]t��&��O����%�Ρ?FT��~�g�11�_4|��e} �N��ތd=n���Ɖݛ;�\��Z���ط4ԉ'��:EJ@B���2�6۝�_�~�I�6���r���Q+�B��ƕG�9R��C��i�KF�'�mم�f�-,ͥ�K��m�+3�""�Bw7��W����gh~�$7�~"��d�s�"\5,���hحn�8k�m[^3��]{{4l��Mt?��.�9�QF�IL�ۜ�[��f6��%[��E�H����J?�PJ?l��j����>�f�aVKd�XdrN8������U�$Z3�0�w�пe�L��R�q&��Qt����iF�U���Ӫ�y�P��jtj�AP"39�բ��:/:m_L��I��0������c�v��>��#����\�6�
�4��/�Yy���E>(J!��)bP�����r��]ʠ|C!"���VO*k��wX��z�uL�r䔣�����u��G�>���ގ��vOF�~�'Ȯ����3���gl�39���$m�D75i��%y��^Y�=\0�:����	��y��)���CD�;X��M�������Zm���ԍ˅ɰ�߬	y�`3L3Z��G�/�}1�$!��B0��<s]M��|
M�:�74��6�o�k�~L[�1*Q��+���yj�SO>d����,������f�|X1V�Sc�n8��^գ�xp<���Dk
��v�Y`k�0�<���w�;ʿ��޳�֕�X'�� Ǩ��ġ7���mw�(�_�wps4A�� ���~�7��/!֫��nf�n����[\�L��O�{�����7:ޒR'Lg5ٵ-ǩ-�Q>�����d����0�v��.|�B�J�70A�{кv����a#�"�#�O�_/��Ǩ��-���`)�]D=���Z���Q+��F��t��������6�`|��0v&��;�{����ߝIg������c17m{��Ǒ�f�m~�;嘌o�f�o[���̜��nq�iBoU������kr�+E:�l~	�֨�Ԩ�����M��W�sⱑ�qBa���:���w�7����+7�vzx7ɫ�M��^�&�	��C&���;+��+
�疇:�(�z�:��vO۟�4��?A.����)u<�}���w|T��RIY��Z�8>��k��A��9�}Ͷ������<J$@|<�H^KR$�j���4�4��y=�=%�S,#�tS[����S唟5�'�C�&�:��sټэgx(}U!�:�Lks�  �E���D����,�a��{�����(��.�t)��&�m�cU��֯��C���{�nӀ j<�:�:�8(�N��x
"a�^/R˿-󮎸�#14S�������L߿�A
��.cw�H"��F7U/9�3R�Ҍ�|�ɳ�Cf��t�2�����c�U�%�������J�%\�?�����[�\��5Tl1�G�Fdq��nw��P�ַ���i����-Г2�^w9��:�B1�!��Ns�2{׆�����������Χ�λ!��?��u�(����[���?+wg(��,p?�?�����Z�k�=
#��x�%0��Z���<w�u���cCPTx��6)�+��>V?ch���[����:YM��qiy
3���2�hYn��N��Mi%���O�
O�;����l+;S�����﫷�7v�J�5�ܭ����N�v�5��Ή�V�"uh�4pjh���u�+��}7��Z���7R%ʩ�0�Ԡ��\�:w�N$�A>"Ȕ	(R���m�CD�ܨa�A���ԕ�A�do"��)U����w,�c�8`�.�1œ�Nx4j��#��?!�d�_�
��o��{Cpi�0�QM-��i#LА���媘�ڃ�y��#��(�s�/B�/�+���<��ly�ށ7X@l���O]��5&N�����ފ����=�t&�����[���,�E��rC7���1($�3��F��8��G�*~a��]�W�.S�)S�6�Ky�R3��xG =\)'�!��P��g�-��)���%�h�e����d�.��[#�[�ؑ�2� ��V���!!Ʋ<X�j_c��4�2T���C�U�{��`K�������V,��z�ٗ�{=Rf�Akd�Qc͚2�L%o����dTj����ӰIh ��b&�9����2C)�R��$a���f�T���E�:�;] ���\`�5
2�RjZNOxNnWmG���x�Wf"*c�F�޿onv�0�� `��C�Y�E�{DI�鎡Ci�n:�CA��a���;���c�9����5����?~��k&#������v��=R���R�������T�:v����K,��\�6���߮��i�"�m�[�N1m
�S	��>%T�$̫V\h(�7B�N�z�|�-M����{u\Sm���~(�����Y���~#���_|_��kv;��h�v�q?�	��I<����o7p"��N���C3��=�ϳ��d�q\�f|�ׂ���6�Y�!o��VpvU3��َ�p@9jb́t9\��Nڤ�
�5ٌx��L��
Ĭ�'����Y�����K�s�Z�� >�N ��9h�*[Pj���ӂ���I��i�,�G�xt٧�Cmy��g���R�CF
D1y�G�A�}��f�ky�D��pnmJ^`9z�� �Q���?�2���П��&5K���W�,�1������O�W)���D�E&�%&5��_�x�ˑ��Cl�>G����`��u	EK��7��:ʅ���\��ް�Svı>��k��ɶ�fD�Q$<82Uv
:��N�k�Zɛ�V���VY�p-^����nS�'NE��;v��Ҧ*��m����i,�q��qP\h�G�!� �o���#��1�_�����%��Nd�{�iJ]��[�o�|������u����a	ڭ����!��Llj��I���5�Lv��(b~B4�*��ȮPA�I����%��Ȭ�����M�I�9���u�,�e�I���a�R��Z�0�����6�:�}U�m�3cPu^rKW��|Xp�k_�~�[��ĄDB߳y�k��)�ljI�o+DTg1`�m�*E\.�^��� I�bm�l��v�k;�G��|c|���-���<��c�Tq�\�p�b�OgjjR .(b��C����C3���Ǡ�ɲ��#��(#K�g#�<�����U{B�i����Q�����K�t��s�ι^#Ku�K�l�}�Q�
��ǺHP(QKL�=��>j�uT��q�È��;�x�&�й�	�?C���F����l��3:	�a��%��gK��(c&��kI����ڟan�?s)N5���e�Y����^�"�}#�|�۳e�I����p��?��V_� 6a�|x��.r.����Z�W����=�ߖ��?,D�	��yoz�������?���� O���W�m�I'-��/瑶���꼓�\!���2#(��|���>.���%�i.���'�gj;���>�J����������%��0,(���
��?gm�����|0?���&��--����4�=6qg��\ܞ0�d>����A`� ��L|�d1 
��0n(g÷��i2E��?h��/�߲0��
���-�|��.�X�>��GA��̵��j7U�������.�:k:d�q�d3)x�>�|�ȵ(�%��Ţ���f��#+�b��D��s!2�~%���?�'��.q=�N��l�O���$�L1Da[�����PB�C� ��BmFfq�-&�1q1u�%��Z��F���,�w�*�|' �u��{�A�M��W�G�'V�Fꆺ:RImS#����5
�![΀[\1�����}*����Ŀ����s�m�_�)���b��b�%�

-G� }@��-�"ʞ�A�͔S�V�3��g�fW|[xu	�x ���:@�R�P�N�w�ؾ���W%�VׄD�ۡ@�h�S�I[�L����Q�zN��0t?�Yl��8�!��A���aN�{����~o������Ph��Qz�S` 3�,Hr��'����\���\�E�3���.���g2��j�<(?����`�'���vq�l`���,\t�3��;a��e�5z�8�y��,1@I,��}��&�p$@��7��2�����6��Cմ�9��uD�P���Q	}�:�Q�ɼ��T�Pi�yD��H��B<鋟��)��di�a؉�g�Ed�ET�8�Ҳ�P&��]d�
�拘�����2��׃�8�@�;��(X�Y�r���^�Ha�c
�I����(�ݜSޡ]C�$����j�X�g[� ��l�I�\}�1T!<���Ԝ�ǻ�*�/���ѻ�&6�a�W�ڜ��:V��FMƂ����I��B���4w�ڕ�qg����Rh����M�ص̠�>~��r��D�`�g�^[�X�{����� U)f�S��B����/L,n��������Y2���>�������^������~=Z��ueەh'��V�_�;��y�>�]��!���jZ?���W��A f�����v�,1�ū�������B> �k��#��S0B,� Q(���R
�]�*���#�-�Sti0$��$���C�*�[�!D�����y ��ֽ�~B^��%ew�/eJ&�t'|�<WP���R�"���	R)�� zz|�7�< �T�$
�̲~VD� >��xŢ� �zԣ�:�k����e����.�7ʪ��5����|�"L��p����_�O�������a98�m��z,w��dwv�͏���Z�K_��KD�,K\|�\
�׭o�3������E�4�N)�m� ��$W ��3���1T0%x�Ӫ����ݩ\��n/U���f�T�6D��D��Ww�L�F�Ú������3���z���+��]���
,2[����8iOz�D�����P��j���bi������)8�Z��$��7�}�,uh	:y�%���+rߺz�p
?���}�B6���;�@��|��[��W��'�4S�D�j	gE7�38M��=�zE�!"��Z�~��/�L	����+z�aՙu;S�sp�>����ۙ�-�P��<2���zS�;=�� �����X��J�y7�EID��!	��������'��/`
�A����M��F��[��2i������sά=UA��ӑU)����A~0�ԪtH�W2#�[��O3��ZH��K�L��j�Z��ߟNq����Y^v��n�u�"E���o�"N��8F%�:O�����#`�,/R���1~�ߥ��ҟ����JT��Ȭ��zT2~ZHxl��X�8-4�|��RZ�w�Uu
W�Q:�D���3�N��4������)7�'��4u-�B����5M�5{TZ����a��G�����~��~#����G ^��~[��D��N�򼬏�C�@��)�8SŮ1�7ۿ���b�쀫���g�Ȃ��>Ks�ÊꔾDϡN���!���jh�t��7�b���X�A����D���X���Σ��9ж��_���t)zU���>fq5g��������Sdy *=�J?�۾�_S�&��7���L�Q�p�m>���)��/�-+��:�9����y�*����66og�iQ�;#-�^���:v���
$��:�����{�i���q|E:�S�?+y2�f9���X�e[�P�s����I����;�~h��~��|��,
*��0����q`�+��m�SU��g^qh0�z=������Xy��e!x���0+V���S��U��(k�a���(�8�F����Nm��Y�V2a��u��c��J�I���+b�K�:�_u���s_����3^AE|S�����O�N	�n�8������/�_���G��I�<܄\gS����F`t���z���fjN��@ �h�By�ƒ�I�{�zq�q�lR��oSܠ����pòW<�qR�EVBcù_"g�Ѩ����C6��	������)�����M�}�~w�4�{�0����wб��ѯ|(���G6��-5ځ��(�o*�o	�/_��O���H���v�@n�
�k��;�$�N'����ʋSS�z��c����%r�6��a��èʜL��7�V1������Hx�� l��������ǠcܺwE�q���;{��h���'D����`��36t���0<-��T>`W�H_o8ӓ.ʕ�$����@K�j�á�� 1mKd�X=��"���nD��>��
4з��OG�2������G���!`�F�>��'r,�պ�����I�-o����� ,z�E�T�Y�d����ы�������%�N�����E�l_�Iq��-�  �9�Y��bSÏ����es3�ֿ�z��ʑ�er���hZ��@vA���l!��z�X9���k_8�B�ӿ��S��@j�ƫ��]d��Մ-?h�y� �$�v
s��0�m��u?"�Ϊ&?�z����o�>USF����,�kO���f���K�
f�?��̐�)�?)NŻ6�zJ�>F�&�O#a/o�Ƴ�d�����0o`��nE�v���_��clGX��-#������<kO���;��63]�n`���
�{o�(N�ʛ�k`'�ԩ.>i���-y���&�B�N�?��8�6lNW}ļ?���K>�ۻ��8r�ţ1�R���.*���ƅ4՞�|;��c��Dǝ����)�B�O�eK��!l~�*��6�
�7#�M�)-���͊�*ڣg�[Fs5x򋐾� ��'M��F������I5v;`�.����M☂5�O��Xu3g�C�txy/�7{�,e3�M{�6��j���MI�	��N,����?��'�V��� ������F�H~�ݛVO�rjJ>�S��9���TԜ"�`��m����r�q�]n������*�Luw#����d'q��>����ތG��&��[Y��5�BcDx��]ߐ��<<�`�LG?P�.�sh����f���X�a�uP>/��M�]��Vc }�/�E-*����i�Y}h̪�{~�%�4I`�ߒHq�=w�s��v&-�)\)<�u�A�>����y�0���,�<��u0���P�Wb�Ц [3�jcLA�-�gAF�/�,2�+zў�QF������qqboU�*Dd��Q+�-�����4.�E���6u�Sh���o�q:7x}=N�b��H��P��f��]zy@^pO6E�2��8��`�^#��z�VS޿+����%]�%�}B"�0�l���h�{�J�w�>�Qj��&��;����I{ő�=jZH��q!��v�Ps�o��[���E�́�* [�r=����2�kd�2I^�o��L��G������`� ���G1�J-���0A�7��o?\=K�Y�a���@��oZ� �5Y��0�w~_���ܹ
IJa���	:�̒_s�M�$��Ё/��O���Q�b�S���,s�/��j�rJ/���G�yl|�n�?�Jf@���9�ɬ���*N7��+����_̓</�܌X�f�������m�eK{�%�����'{�BS�n�����? ��I��ԗ-��I��S�����y}�U����?�U��t�����7Ӌܾ�W��yo[��ns(��b���(ઐ�æ�t�q�,n��{����=^$`El�~�b���.�YR�M:��<h�۝:�rz�pѻJ��j����5ӂ��l��U�'yf&%iG �a
z�� k).T�uV�d��K|>?���Ssi�f,���3���<o8�)�e��_b�1���F�`�\2��ǡ�?_�|�4����5��B$<l�/h�	�.K��.�i�v�9��řov�ݽ�ƫVOgeo��O4�B��4rHw�׺X�-��O�O*l��G�/	!��r�gw����i@c4L���@����	��iU�q��E�t���yʐ�6���=����G��=q�VߍI�=�G%����I�O>H�V]/|�4��f\�?:�7����W1L�^m*Ʃ&g��������i?���gkN���2��3z�1�IF�h� T�kYChJ�{�ϔ�Os㭇�I@����h+�Ӊ]���l�c
B���wo[W�>ؼ�vUt�㵼��^<�UT�mҚ������B����B�?G��x��DW2|�2�'m���)�hc���XĐ�<��Y=*�T��a<��8�4h������J*[�O
�g�G3b}�<��SԢ;$�������,�����k�誀�$u^m6�`�*xu�k�s�	K���(UZ9�R���%�rIܼOk|��������6�o�������!�%t��	�	�z�8k��o=
�*�Ơ��7%��dM����D��n�~��e�?Gg�*DXP ՞��:�jL&�_�i�4�%q3�A�]�:���\�t�qnh�Q��  %��3�,�t���Ҁ PKA/U�@���Ǩ�O@�����x7&E=�8��9]�!��Λ��q����)�1�aR~k+v�����Ӟ�cK��?Q�&��Cc�g���c�����7ֿ�b�����*8b g�� 
���Qxb�k5:��jݭ�L9o�?skF�����JA!4��W���'������xS�m�?NF��N՗��3&�=&}�ࣃ��r�6�\������X]~at����V�bU�?��*p�'ѧ�%G�8˵R�
}���������G\۶8
w;#����o�!�Ҭ˨.&��$-�u�Zu�s��n����~�'�,�����ԍd���1� &�6�ߑL���H�#4{��ۘ�I�Z���R�]��=ΛS�EԆ������m2"p\�G�7]�UB�J� ���KM�s�w08C��~���8��V?�ChG���]mL/9�\GhAǣ6_��\�9oCIra��s��e�	�����~�#���n&��+��|N���׎�C�O�K<��|�I�'7�]:�MD�0�Հ|Q�/<D����ę�[�s�$
08/���
π�uԿ����c�'��K���/����n60˼��<�pP�]ގ�X�pP�(�8����f�~���Q|��q��k�x�r���g}kQ�fr�l��_	�v����}��'p�<�g��L�����	
����~����gƠ������U�W�&��?� ��C�uw���������
�r�ߵ��yź���l�Hï?��Tz�%6�|�z�	����c��F�Y ��*��&-��K	/��.�:$=;��P*�޲��s� y�1�o�T%MK@�Ɯ[#�ƃ�����������ꈨ]P��~:�*�|��p��b�Y}ƛ��l��TjՀ�G�z�ih8��˛��n�i��h��_e��Kv�����m�B��T�w*ƝO`׽�ok?�b���}lH+�����&E!�ݚ
�/�\�\�>�tf�8������Z�!���r$���� d�*
8�V����z����ZYj~�e��׏(_V���dz�/]��_g��;�2��P��8"�X�s�,#�&:7����
���II��K\V<����AS�sg�W����x�Co�v�N���(�E4c�j����'�-(�S b�n2uta��G�B��m�b����c(,d��~{�^u3s#����I��lfj�R�hK�h��ILRz���^_x,q�
k۹��A�;i�����^��#�7
��9mǶ�[ke/�o�S��W4T��Ǐ}j��t7��y�Vr"��>5BO���J�e��q <�u�pw�#�&���*sͣ�O�E+��nQS�s*0	y�BY�x^ƺ���Pu���Zqcy͠n��)K�Ӌ�������G�}�C����3�/ *��Nc?�N��R�@3c�ə���Y�8K��!C1E�,�į���*z݋"��	�H/���/K����![	��R�4�9a��d-�S��C�-���]밎1m�����s���g�T:�:�l���>y������lqK�G���C/�?�Br[��uqU>&�c��_��K������8��6���+f^ 6L�ӵ�����i�Tc����Ԙ�����a;�w�~�TG��uU���)q�r:���G��E��I�w֣f�i\vft���m�]�q�	3	�F�L�����ω0��YOH�I�;F�lQkS6<��"N���6���8���D���Z�O�qm,�)�~���٠	 ����"FZ}x��������(�~;s��S��C�p�2�5�ԋ_�N<Nd�Ǫ�^G���������r�.tS���CZ���%NUY��tKe}�U�p�a���?��(��cS�L�������[*W2�=�u<��h��ԏ%�P����G�k���;���﹵��\���ʫ�o~S)N��u����6�}(*V��)���ٔDl�P��N��*řRT����R�漝v2u�J�B7��c�h����t0R���R�3?t�م(�ƗG�9(�,`�饼�M��MK����k����%>Ӑ�`;��[@���¢	>�pu���g}W}����M�4���	����� $4�<U(��w(��;�����v�KR��Q)�ٿC4�������gl]��=P{u��-�􏆕��5�R%�Yܕy!<tl*5X��=�z<�5�0�P4.�hә¬L�ט��J��xkG�H�j�lA
j��dܚ��/��q�?�I�?c�g!`(�1;��I�k��tpj�Y���qݑo �G�'Iy{��g_�*��Ӕ*S�ɟp��Fَ	/�jL��ħ�K��-���{�)�ˬ��3�@�� ��L�jS��YC8B�Y"mǢ,�U�wU�#\��ڴ=���)Ore�I�������q�/��m!La�`�����-��8��GA|Ǖ.�򉤗˾�:I���t!�؏Q��i�]:-`�d+:�ϕ�qGU�ք�������k�SY2�  ���/����T��<��[��Ws2��.4�w]" �W���׽���}=��>J�a�K�ahZ��I�v�Ԅ�=�,����Z�F�N��.�}�f3��z�͂l¿�X:����A��L��h/�[��+��|��4�%��}����H��T��ft�t�=-�:�I�HVO�nk:s��M��7W�2<���V��vH��N���b��4�O�����DV�}w�iyM�]��6�(���f>�}�!e8�]�B5��Z����i�<l����1{Wz##-��ғ�<1����'�����n1�ڡ#��n_�������^e����x���H_�j_�U@�aB�S[��%)ނxj������e�5½���!Ǭ��������Bn�g��>��4Gh��)�`�L�
C%��%�=�N�}�b�ql�k�E>�1p`�_h���D6�M�f _2W���Ne���� �C�G�v�/o+;��uhdGȑ��a�"�@����I9�kŦ��֐���i�S
5Ț�mt+�
���@����7��tӉ���������x>�}�
�	�N8B�j%�V��ƶ��59��8 B:+�tH_��D��z+buWm��F	(1+��7��@��͠��M�`�fĔH@Wf�����Y��ĨL���&��^5�9]�����'��:r��	�8�~̽(��tAt�zfW�@�*ZW��%���ɋ�����Ֆ��Ƞ���,���M�h�CuU���XV[���2�f���`��P���!ɧG�?u��rOGoj�:��J����	��@%�k	
͖��c%L ���vI�sp��R����y򹝮܃V��F)�qH_�>�nzby5��$3~?��\A���h�����][��L��$����YA/ܒ�+��/�5^OD�M��k���
���)����d�16�Z<.}��S6��,%@[k�}�g?�ɛh@��ijK9h�O����<�;/�s���)2�=S���;~��4	Aմ���-&�,3��]�I��p��*drю�nP����UXPE�c�DU��(�DY� �����t��]a�ף�B>n:'CL�/�:�H��B>�*6@���r�����b<5+g�-ҽӎ��=o�z�*�`+�y�� ����W�*d��\�$|V�=''�8�hG������=�5^M|v�Y�����D�H��S�e��t�$gK��]�e��j�ٷJF��w&�*�'aq�o����:Μ']��+
^�[�>W�2ĵA�Q�m�ӈ�մ���_��=�md��e�ŧd0���B���夬:��O���i?r7�2��;K9���;�@�՛XҶ��m��%�0۴���ѧ���O���_#��"�Z���?)�n&�����
�<DL�߹&*!>�t9*��8ծ�۸s�V���uqj���1$��������D�m^�.��� ��3�8�tQ����E E��������&���Hi4|��J9Z����-���cӃ�Z虝�����
����}A4���N�?�թQ���.��B�f���z�(�*���/�3��cM�~]e�$�݇�����V�3�є���'O}���c��j�֊.�6�w�'����#wY��V����>����ұ��>*��{�����Ms7n*7�-���rߩ���>�J�R��+ڽ ���*r��@IW��e+�h�z �@�q�1?v��C��<�m�����ֵ@D��p>`������C����K�Pa^X ݐ�PbBm0/m���
��5Z+uaV�� QS��m��k�U|~�"�f��c�����
R#L�I����bBLj�D
����
c�gK;�#��Ο�f�ul4�M2(�z�xn7&���N�$�Q��5�g�����'k̨��O*�	���%�pn��wŋ͒�Ҿi��nz�QM����%[��S��L��x������:yt� ��a%���!2�B_)�X�4�(Dx�b�-o��WV�qk�5br�kQ��Lݴ�b�,4�Peǌ/{�����|ݡ;��.)5����`K���97��=�O�m�]�|Z��äp��ɇ�O+���躋"��[�y2C��m��+�_�]��6Z�~���jIl�\��H���d�6&�HW>�Geϡ���8@�3���}
PFE@��Ek2�s�h��ӱe��'=��79��4��>���Y\y��k���恻.�^	�H-�;>�4ތ�y��ѿ�wPzږ!D��V}�W�x�>���/������;����a��;���@MU��R�����x���w]Q5O�
J? �=&z^�{���龀 �j5¶�nS�4jU��ViR����C^\��Fp1C��+ F�0iI*r�h|�t.��{X��9P��ao��������t
�����@qS���|Kh'q��=��|�O�<�����b���r��=*\�
�� ��M��8���$��)_���@�� i��n�\RT��0>OXz�a���³����%([t��-�:���t�c�2 �&crt��$���ȿ52Wx!GT<v�q�.2L?`_����-��BgZ����{��8��	�J�ҥ�I؅'�;�Z�+h�p5k���8�9n._>=�T�y��Q��i뗯`Dz�v+0����%�$�&��~7V�O���$U��8ߎn։(�U}3���-�;���G��LV{V~"�� �.����p<�,�F�����b�;���q�
� �������7�2�2�b��"�)&�.�mZmv~�P ZJy�C"uv��%<o�Ń�3�񼌰c��y��6���;�Q� hu�&GY _3�ʬ�IL${bwۿ���>��`��hH���˰��Y��	Ky�I!�=�2V�&2%[yP�O�Z�!|.�n��؍��}�\�)T�ʍF�U�tTi��ʉ��PB�;�n�����ʤ��C�\��b�Y.e��)D`�F	���W�@��U��$����f��e-ψ�}�j��5�+XR�7.2ǔ�V�g@/�H��&lA��*2\z��D:"��)]�b觃�%A�Ϸ��)���k�tImj�8�-Ϧ+���מs�GlU�>���f��A��?�*�l����gX�������%��t�q�y��Y	l�Q�v8u#�&��'QTO��^��7�F�7�툂���&����zƿ��$zd��{�>o����uG9��'	-�6g'�@+�k�A�۝�j��~����ҹ�]��4��f"�1���˓҆���ɫ=�t	�i$\o�>��N<��C\�U\��@�F����o�zh\[�\VU��PO�9�B$Fm~ B 8���_P�
Y?΍��hm�g�!�Ŭd��\�Uq�|�M�D��Mn��@�}Df*=�b	�}��Gō'S�������8���6.���߳�Z�á�)X�e>��T^��A�މ���8�%���������[�ynY����_���������~k�yMO�JQa�6Vw�n0y��H��g�31��x<@��]b讼�D]�Me����n[��+[)�<?��B��d��l �F�(����z�^���O�wM�ݷ�o}Db��2��ʇG�U���m�9�B�طiu��BK�<˹L+a<�д�`�Jq���=41�߬�nB����)���Gh8�-!4��.�,�� �\�[C���Ȕ��sjM%��*Άe�\ZX�[�e����p���nG{���拄F��Pی�$�Q�(Ѓ�2� 0����6Ed+A��@r����r4�y�;T�M����eKݒĺuv�S��1ڇ�Nw��k�[H��,Ύh������� �%鋺����L��k���U�v�H���K�!���G��G�������|#懋�� :))w�NO��t�gr���ҁ�r��t��*�K� +fI���ɦ��oѾ�Q~Qg�|�fC��M�!��ج�kT�۴� %yr��+d�#���_�~��R��U�7)8�7L��Yx�8�����	�RK�TDElir�L	�!e�&}?K̐h�k�#�||,g𡇝��
�0�#\}�KO����i�j�v%.�0�ѝoX�#��"�Ҩ"N{KL�~q�v@�E��ڴ��{����ɯT�<n�OĲFV���sf��z��W��:�l�Z���*��I>.i��<Σ8So�S�������2c����79�.��t�xRQ��f�����+&i%;��1�X�pՋ$���$>���&��"��ۏ�,H�[:�:^���F�ݎS$�Mġ� .�HI�{R�
�r�����uK�����v��)K��4����e�n��
"t^���ٟ���XvhL[D��)�a��}���ߪ�����q��ls`
Jї�M[6�V�R�S�Ľ;`HbQ9- �ҖW���~�Y�mr�=� ����<2�uv�3е�֕dl����}��6Q�l��nZ}t+���XF�e"x�5t�Z%l�g�}�H���ALq��ö@��3��	K�@�S͖S�K���'(%�l����}�1V+��1)(^T�[�T��)Fp{f/����M��F���K� a�݅F\ǈa
Bq�T�@�����#�m���I��ӜIB���N~gow��c�]�&	@�R~�l7�<����|)%����=Yf�R�z�15c��\�	��ίh71���� ӌy{h�?����l@��v٢z��8
I����G23�A����_=�U�}��$���ǰf��>�q�!����,^̌N�.&����q��_���N>������֡ɵs	�T��m�Մ��P�>6�F��9N&8�\�L<�!VGxTdI�%è{m�^����Ʋؚ�v�\iad���IM/(�¶T1��Gc��c�������Z�۹�D��8�1��o\��������F�}�,�1+~�=Kߎ��Ә�p�y�^jYݭt�E�T���#�`#��i�`�Qa+��o������OC�����f����!�7Ώ#ȼ�Yh�V�0j|e�,�܉�^�`iUw�a:=RQ:W��ƕ�q������^�I;"6��V=�2�m�lA�+y����m��=�sd-va����藶r���j9���s=��\�:����``�D�SzW����	���C�h	�A��r�5���d5\��f2�V@K�y��;���<aT�0�|s7l��:��i�\ 
C�d���z�[����mV.�>��TP?�rH����/*D͘��x
����p���B��X(���t�+�9�={u�YܧeM�
n F���(1�n��^	��ZM���ү\p7��X�z���U��HqF��p?,���w�y�d�}�I���w,Z�Z�C��#�at�Qf���6P�Yvpd�u92v��~�w�B�t�n��P����}�L�q��6���5Β��m��*{@]�z��.���\�~a�������,`ܵ�F�:{v/��֮ _�&s+�c��SA�8�)c`�ec�2�Y_���5�e��}R޺��������Mt��V]��C4�U�T�1�x%F�;/�3T�3�v�j=���]o˂B��Y?�"V�?�z�X!�K�<=B��',��4���d�)�ɀÛ�Mĳ���<���v���U�4�+���c����~u��p�gz$�xAh&8�!5[���fFqj^H���[-aY!�K�����z�*�0�8�ܟ�G�f�y�G���(���%���]�X?�6���T}���b���ԡg�U�C�^��yZ���6�P�g�\�\� �:�P�W<���:�8͛���`L&�����o�̵OR*m@}5�B���b�会�":��^.���Y����O-��˾z36��'�/���=-k�Su���,=����|���E����0�۷v�º�׋]o�_��2s��b�J�v%�`Ap�Hp�D�����)Q�������<�"g��#���$���`��x�L\ä��E�0�Ӱ��(���{9;��ȡv�܍�䙖��hY�U�]
��/V�M�0�����t�q�ѯ�<ߓE5)u����Wǌw!_Vb�
�&��!�+��$u��������uPK�z)B`�ϑ�BDU�`�퉦�M�#�u���o�HYO��n�+{��4x�����O֔��s=�I	����{�g��߱)��k�usQ�~�3��{F���y6C���%����C�b��%�jOu_?�ڨ�)6*���U�J�xF�%��ݣez���¶ɰ��Ǳ�]}��rO�}�*�s7[��F�^������J܍M�l�
{A�S�ưڱ�������ɬ�`v���s�٠����#���r�#�����PCl)ȅ�#��5�k�&��!|D*��^���ƥ��n�����f�_�>iq���8$�z�2M�Tg��$S���rvDZ8���jYF�V9������f{CK�7�3�gmab�2�5��W{�y-��5�\^Jz���.�u�G�Gn�P�
Ի>�)W���ٔT�)�̫Q�1��ٗb�g��w�c�ŭ�+9S����D��ɳU�T��`��pi�r�E�e���~!l����+��x��xS�cS/F�)�P�R��!�q8�v��k&�e�
S_�v�D���n�� n��3�x~��~_" q6�_���S���~���b�Ls�A���CWzB�!�UN贒_�TtE������Ns��	5j����c;˴�(F�;�D3��ç�ᛳ�xO4;��/-�:6s��w�W��4�`��4c���)8DľF�R�|>=�-DI;�������ۑ�*ZLvS�_ll2�W^�8�p�cb��^�vBg��G,�>�6��!��6?W�C��� 
������Q��q}���7�&h�%�����	��8�ݙɜ�ʥq�8������7��a����S�b&v��4��ސ�Zr�?���o�m`a�L�{�^[�/��^�[�BA5#9 ��A��ݜ��Z1Eѓm��!�Յ����V�����bfP�l�LB�óLo�3��W��Mp�L$�}�))�i��]4�>��F]ٵ��G�}��3T�ǰ�⑛w�ɧs���鶚~����p76s�3������C�6�����b3�k�&�$�m�*W�wCv��'�-�������=�XL7f�o�d7��0�ۚ�*���(�J����g��<Os�㊽g��EQpn��]r_ zտ��z�����׎0;��Z��Xٻ���TOJ��<��-C��8�����~:3|�#�L�"�8jBt$��$׍{W�lhN7�e���IP���%�|v�G��op�����p����I�K�^�����fM/�4ͫ5pHb5�ٷ2��L�ι�x��;�{����a6�Z9oS'��;��>\����:��j:��S�;�`|�Q�[�}�~��g�>7��O�}��wyt.YM�d^�ݺ�$�Y�Y�n_��D��>����>vR���s��عxT���K5 s���Φ��w!�����M�г+@`�)V1�8~�W�`��O�9K3�L�ߩ�ӧI��%F�K�i����.��e�m� 骪������P�:8���}���c�������oo�J��rޮ�<�sB�K��1[����yQ����Yw�!�1�y?мo����LP��ӊ��y�=��I�I��U���ב)�)(ѝ�"<���Q-��1]��8��\`$�p����3(..t�s�}E!���SaR�
H���;������H�E��H�H/b"������H�i!)"]�t"ґH�MPD:7<�;�{��7��Ʉ���k{�������<4�{�P��;��a����\%9{�d�B���S����Ϳ�Ūl�-on��Ntǐ�8pn��%�O��`�?�[���-g4W�@U�x��'�g�e�(����v�I�9�O/B�O>N��+v��A��
�o�i1�O,�҅�]0�#�:�G��e�yK���3��c�?�]����	���T7]��dv��5谗��������Q�K�V&�B9��T̖�\.G�~�1�Q4�k��S��21BMJ�0�0��i�j�(��zŉ�z_�x� ������a�y�XlB�n�r�_�]s�P%����F�b���+���o'#��_<��WP�\ۈ���j�%���z��J{,�/�<��^~�ZG˼z(B�)L������#ͯ���q��	u�"��<;X���M�xPy���-�2���7�g��'��.W������P��ܚ�<�ּ:���|�dܮ ?�����9���ùǲ ��
U͇�͠w�	�1�o¡RpRe{n�x�섰&oQ_Gi�����R" ���Q�^�.��������H���9�+�gO{U�l�T=y���5E2�N��\���WlA�m�͡��'��>��+F9�0_Γ��p��d�t�B�~��0#y����j�v�ZcJ�,i'b:����t��b��s<�ÿi�4��<	���ۗ��<�(��B���5��DUI}�d�p�
em|��ᴻ�ʍ��ý��!ʚ��2{j��<,>R�����U�>}���q���s����3�:�,�w\����ũ��cE0�B��f�2$�a4j��k������	������h�ǈ��m˩]��Ů,�"��9�tӍX�$͜�q�ε�>e�gW�hM���e��jK+NnA��bKYs~��!/����?��� z����I�e�U��؀ P =�����;��_��sb��@�<Vglu\&Q�#��X�>"'�&���I�$f�=�U�[ɍ�/�1�P��'�q�j�����4u����ԟ: ^����l�,�8��Xp�+�	_~	�5x)��F��$^��D5�@�O��b(Ai#az(�J��� 1.>��s�|e[֡%��֌�1�L�jWѫ��#`�Ƒg���)z�뉍�-��8be���������	:��L�3+��!I�G�_��75,��R���MR4|٠��A߃]0�(Dsr�>��^+��{���B�w��c��z�$���/?3%�`��-���]�٭}��O�㎈��hWsH/d�K�).��u�����>���R���"h��9��~=?���_ԯ���^!�VD���?n���4��Q
�l�-���?@�a~�"�K=�����j��jD��~[p���"}�g;'	�fm��)�A2
z�KE�K���C�6<b��}a���	���>G���C�X�?�`�)�Mz^Vբ��ų�w����>Id���k�WW��3p�j��hMg.A	���3q��u�e��;i�I%f�v�2e����'����h�xv�zl��B��Nf�f��s������'�g�����'#g�_�e�f*����6�K�����f�K���]��='��'j�(�
�|��<�T���l���Yx8����*<��B�<���W�/�V�o���%bj>�Z�y�A� Hv<PВ�y����ݞ<8�M��4�.̲��v���.������;Ѥ� ��B�	�.��Lm2�����7~���J�X纗*��F��Ţ	��bP}s%�{��M��e�K�1�Dk�[O˰�|���]����9�UVЈ`��^�=�+���疭�ď>e~G+�����j�p!4�/f������J2��m�BL�~E9<�
���"�o\:ci� �b�`���S2`T'���nn9>9%�Ё���6�T���y/2¼�����ɷ^�X���C�4W�Ta�����maڨ~a���e���u͘hJ��2%'�� :��ItZ�2m�&-��j� V�#�u�\S2a�E�ڜ�4��=���ݵt(_�w&�S�:���}Wi%�nu�{j-c2Ypk�%����Bqw��S&vK|�<�s�H>��LN1��.J���������6lȻDG�?3K��oj>>�R記�A�]��|�&���l��&g	ӳ����_��]��PЦ��%��Xr�����HI�y*��=ES^v�)T�X��G��un�|?�̙ɸ���'˭dL�B����npt����3db�n���� n��w�� �-{���`�V�/��S��E\�1��td�_���J]I�/m+#�Շ.��w�r3��>���Qy�7"���1�}�z�/�O7�V��K�u�qz�]^�ă���?�Lֆ��}���pn��OÒ�.��6��&�I��ڡ���JJD6n�zV�ДF��Pu�폥���!����N�UJ�����X� �� 0�C8��Ɣ*�/)%��~a�6[~����~ �L��B"�M�@+"��w����]�������,x�M��v���J�T�h���7�� �d��k�D�;om��<��\Y�I�W�
��&&R�~4��s����v��B���t27�+�ד��V��1_�I��J�H�V�IP�*q��[(X4&5�Uv4f�\f��B��S����o���"4
@�S�B"��X��2D:
�uǌBEViz�n.At��N��F����{>UC�:�6+�����o=2z�����S(dje���t���6}�y�T(����e���j~d68�?��bp!& Z����G?��_J�����D?�&ʹ8�(��ݏ`Fn���V2#���b����ު{|���f&]9�Ω"�}�J\[�>K*�~~�G�b���z�bAgIw��l0"+0��������`�Eh-UJ�½�<W���LN������vwJ��#�����"�Q�Q
�U�U&\���P�FИ�ف���lU�oO��9��������:�G�W��?��`�D�h@���*"*s���R�ͳ��]���n����xy���?B&��J����׾u_G����t_!Ь����7�����9X�^|!Ş�Wa[�����`/$4� U�ᘒ�40���5�?4y�)�$;W�c�Ə ���?nk�)!+6^mP6>��Lm�5A���䨠�&����n��S�?��PV�.v&�ߟ����Zc@pL��J;���f�u�ìht�%T����N 21�f���Kݔ�{c,b��d��St��@̚3�m1�,�ai��~����8(�`�2'�kq>b�f�Σ��-��s��vp�D9\Dw�Z%[��h��	�o�à
�^o�0��/��;-˙sX�RH֍�t�����A� V1O�:��>� q�[�`�=97������}��W �� V[ӭr�7����n�Ha� K_i�$�;Sx*V�[Ո.�P�@G�I�s����0~N��q�{����JU�A���$��F�2�5V5�A�X�	��d��!$t�:˶#\�#3F� us7
���Z]�������C����8!%(�`�D�rm�,�/ג���������Ja0�)��B>7ß�qۣQ�-u7D}�a�W�i[�ʺ�B�qh\Q�+�EQ�wLo��4�w5.=��m��<]Z�s��	��=��F�'K�љn��#H3���ՉЀ�-���ߚ�+�	����r|3�J���!�1�{s�l�s4��:�i>W���o�P��l��Z�s�<6h�n�"�b�l\���}��w� �E�����~X�*�[�d�BӔ�p�������6���T�����?���w	bҤ�Pc�D���h�����h�Gj�8��ZVk���>𾋺���A����pR��]���|�����k٭����ܥ�5��ԩh�8� |�H�F��F� �Xp�\CӺ��Du3��}�v�!��z@��%�B:�����`"(�O�W�3]��|� �R\ĩ�\�M�3d(�U��(�*R-ҽ�83	�z9�ԧq�C��dr��B�@�:7fr]|K��0WaҰ.(�����N�����~(�2�4��ޗ=p�������q?�#�u�2�1����amN�M�G�h��/>��{�������R_o��Q뢀�������j���\g��Y�[fHv@�ءtr> l����f�=ie�
ꠀ�\�Y�5��̈́�}��9<Q��1_��7��Qc,�;��5S&�m��k�i��J�� ����gU��PXE�����%��C��h%���)���_�bM:����Q��k<M ���2�E�dֵ������/f�oڱ����W�����7�?�V�t���!&�d��vwV�,A�~l��o�Nߨ{Xk>�3���n���k5wܪ����%���P>�E���;	=��A��M9t�oϢ.mpE�����.��}�5�a�t��yߍ�J�~����ٮ��u�/{�ix�D��,�3��ͥI����
����{�B��U�-�f�e�]��Z%m1)��=��;�Ccw7h�F�q ��ܬ�LÒ32*f�!s[�;��ن���0-6(`ʧlI��*��0jq����*?��V�NI���v��KvS�������ÃD=��e9�6��$����.7�m|��l�C���׸���	�����~/�}M,u�Y���4W���YcW�iȲ~,�fm��=d�|[��� �P6�T/��E��`�Ph��+�-	마'�GK�� h�E2P�� �n����;U����4����=)\�����4,ܲp��h�#Jl�U~L�l�ŋ��m1�Ν�vq�B�7פm,�7��o���s�4�ɜG3���� dz�k!�wQEz��lYP�DGH#��)�\7���DYB2���]�"L���J9��t�h��2���AT`D���}���O�+I����.�͂u�8����-��m����dF�ݚ;���cr�}���[���qD��Z���aT�o�F�W/=H��z�>_a�Dn������o�_~i#�H�rF�j��pK���V�t+��b�<ؐ�-��y(1��Ƒe���
	���i񠰧xj�/����cgn.&�;Z��a{�C���ԫ-����A�;-4<�:v�KMKIӗ���*�>�ī��ǦO�aP$"ﱴX��������0���\E��J�����XH=
����\���ٸ�n�Dv��v~���`ύ���h9X���<6���������6X~��`z�`UM�nƢ�����dk�1�$n�}��*�mI��p6�Jx&�u_�$���CI0Wdb�w�m$mO�����%����O9ҧ�� ���ߓj/(��
��;J���͛II)���2��qniFh+�r���Ab�����r��ه�Ц�O��h���u|�n�����~��ֻ���2�25�_�k�)/4�n��U�\�3IW��b�f?&��Yт�\������săU��C��G��I��i��T�#v[au.�k���'R<�������D"�+����R	���.�R�t�twr,�#����Xd�%�Y1|�3��|���֭��GzM(d�PU�+������ ��]�©�$�����nœ�<���
�j
\�ͫ�YE��~��c�% 8s[R7�ru���~a5o&� � �}�f�G'o���8Ұ�f�|5��Nc(�V�����zu�/�� un\,�_Z��Xf��oS���)}���Xp棛�����v������^�.K�E���Кs���e�g/�� ��zVf�n���G"g�l���cUDyX�:��
rg�#7��$�_�`QdCiD��&v ���o,?�\��Y����Gu�h뙊��i�P�Mx��f��ɸ���|���c�� ������;��j�Nn���P�����=�ܮ3+oy;?���Q�ΰ�̖U��Yz�p$G^�C��v�i���ݥ5B�k��-�Z,\���F?)Pƞ��1�3s�6���遐H&�3�6H����[QOt�L(���4����tQ���/]
A�U�[ڪ<O�'�M�1Q���e�0,�8�.#K�a�R���4�,��v��B\�qfr4>2�r���z�QE:�c�J�R��ȫ_�	�/N�/NL��(�Ԯ�ڗ�S��D='M�yp�5���F�>!Jl�u�aqw� Qо�>M_�y�n����&Tlz|��\����$��?�Z���s�Z��c���ա�]�0����:��ܮ���W�]/����E[*�%1����A~������&��OKs�BU�mL}
Q�~�Z���Mt�F�5��$�����q�J�z]�|[�-"����4�¿�0*��I);�]��G&7���G>O$O%^K�ܘ�ޮ4ڕ�4f�~�Ҡ�O���,$�b��_��e���t]��������ܯL�o��?�YN��H�@�k�]��W�3��t�:�!�«⬣���q�M��n��xX>�����Q��×���'QVb�K.ż���#�=��8q=����|U.��m)��G�c�e5���l"�d������t,�p r3��Ƭ������3���w���!�	��X+���狊���������9��/��j/�TXO@�yq��#L�����D�t�t��a�>N#�0���(�v��=u�B5-��:��]��suy��@�&���|;1�wO6��!�3���7g`�����Y�r?Z�Xd$�D㎱qA�H��݋�sR�WG�"�w�Җ?&_��k)x��]�������z�����-' ��=��;�a�-�qҵ�������)�nɎ=��*����ԦO���/��pE�]�&���%d��3}�3ן{A�� �c"]Jk(��\ڟ"��JeU�w	?�GK�.��T�����\d	g����i��Y�i������DF�{��ȨV�|��y��ڝO.��[%e�d�}�a��W���2�i�;�-��3~>�=���\W�N~v']�+)3��iP@��8d��K�w��^=W|O<����/'%�*�ؚ�+.F(����NӢ�P����#�
�Z+���'�G��)l���)Ya��z��!�4��{;G�
��0q@E��BD��C�|���(9i��a��X�1�뺋�k,�<\g�z���t����0�D���#��KVz�Nh��Zr�lM���s�ՓR~�M)���\�5��@�yB�f��A�����;O��:���d�9Y�+̥Zl��a���H�9	�!\�G��_G��(ȧ<�C%�/�%�<�G��9�ԥ(�LZY[ye�� p�h�f�Θ���(z��Y�\�+ƏHB(�3�(s E����^�g�տ��{�`��g��B�b=f�Zp26�Oy� :>;����˸ʊ�̗���&��;^�	\U���;����NH&(E�����:�m��GD
B��<�B��_8��yƭU��>6,�X�����O�*5�|�[���ɘʌ���h/S����,��.�{\-�� "6���}�p�&-�5�r�3���#���LVer�����x��.7C�VH+�?�'s�����\�Oҝt�pv"{����v(�^Ր��*��.t�!3+��h��V��+��Od��<�hʧ�V<�sz�;286ǳ;�`	�s2���l�8:�
/ΩBgʤ{����dDn��-���m������i��A�������̞uN��"S���9���N"#�o_0�f�p��X�߭�n��l�o$!�/��M�������%��^��y��/܏2�E�Rvt[�)��^�w��ah~ELy&�f�3Y��+ŕ0��y�+2����a�@��s��H(y���z@����&%ɨ2�X7H�'
�P����]�}+W ^��%g���4�/�|�ћ�{�%@��zϭ�Rj�=��r/�z��2�uq�(W���#V��X��oy����^8�,���Y揋�M�t��z��,�T�#')(�,����ĝ��!��C}"=�:q|%q�5W�*3�^��3�v��_��!��3���x�t5{���\�g�#>Z�|�i6m@�}�|x���̆�z!���_!����Ԛ�R(O,7`�M�P�$H�3i`SA��$��p�ǣ�7' ����D~�U6�������y�5C���v�tl}�l}\h�l��c�Ʀn�6�M��>�<�=>�����qo�Q]�������MY�s��"� +�h՛�qFB���S��M~}uZx��&�bI��ʧ#��R�����^�Jr����gciܧ �D�Y �k�@tW�����\���f���J�={��"zɟn,��F6wl��� ����CU���ߛ�(� �Y�x�x����c8����Oڕ�
%�u�����
�����\˳\���җk���'��Ȕ�9����fX/�2NwY�ל�x���/��JeA-�4�00���5"�瑾H x���=�"uz���N`��WT�~4�t������T����\�"�yȣMw��V<���wQ\�An�Z�d-�ȗK�/�ʛ�K�H�e&Q/1����BT-lxq��.^�ʀ��b�����t��l�_���^�m9GIN���(8}�|��L+�^�BQ�
HWG��Ѓy�����rح�1�'4�1�Љ�U���Q�.����La�=��dE�Y%�J\�D������:c�M[_{L�R��F���,� SL�r�u�iʹ�%�G�Q����~\|C)�Ƅ$#�f���ݼ��Đ�Z�w��7��Mn7hv�ؗ=��{�_�hu��:��^5���0_��vii��J&�կ鼦Ofw��hz�Kqb5"�.~R��<�o�X�J�s��~P��	@��笨��|y͝њD�4,�Ok�2Tg�e�=>r3�Ҕ7C��|I�^��a�����@�CD.;N���0��%�EƩiUg*M%Q�t��׀ ��82 8����M	�����a�!�?׭�;��(^w��[;���J-��6B�Tר9�;�2oW_�j�(�ܺ�}ݺ/��7�,	1O�u=�j�L�\j�5�R�U����s=x���?m��Zi�Mmk��-c1�n0X9�]̳�6y8x���-C/w+��IE�@���OW�P�O���
ծΑk��9�&&"����1�@��V��P|j��k�%*G(p>IV�_y�\Z���W����(Ta��R��h_v�=/�W�[�e�y=5n1ϻ��n������ZOVVD�hB����-���빉J\/@��QІ�R@���*��D�GӨ����.�ko"}*��I�dj�����:��ޒ㦫����w��,�� �/Q���Ǭ��";��= pCD�s yL"A����dyTE�گ��k�N#�����������Qg�(����AH��'n�AX� ��V��k*m���
��o_��^d jǒ�]��y�$q�$�4\K����L�r�%`*�	��j�N��RNn�@D/���9kuVljI{���v��Z��d(��)���m؛ 7�'"�މ�!�v�-k�S���b�⯊[�����1v6g��Z�T�����˭# 8��5��UU�	�V<�?{�h���kIo�5߾ku��L�gW>�C�=ț6�7Ϛ�|=k��Y�w���trs�����s&,�h�?��8�$e?wO���%O^a~*��,��Ҵ,���w��Ek�+]:qB��j
Al��z�g��U��ʥ#�8P�LT�)��&�]0��bIJi��*�_W_�d�8x���#�w��"�~����L�i
�Yc8֬	u-5gԦs�����w:�� A����a��	1�<�Z�-�6a\�gO�W����	ۋ�I���v��^ĖA��Xxrڂ�@}���^F޲X�F�1��d_&0Ԟףdrf@�2b�z�bML ^S9Gt'�VR�������SA���5ȅ8�T���I��ϖ�����v��qߐ�SVc��z�U�OA���(N@Z�3n˕�k��;�!�H�{w�|W�����ދ��2�i&�G���#}�� ���Psu�˜��<�WJ��K��S*�����w��>� M١�BhW�8c�������k��Q�d9�������B�����>�oJ�����u�����[}���m��}������x��!5^����h�9K���B�)n�&C�;�9sew���8C��R�w�LrC���Be��� �X���(�&��O�?�f��2�]d��G�+wz�M:��Η�_��'����/	�9�u�j�8 �D<�BH5T�Ђ��O_�:��е����U�����I�)�����a�7f�`���d5�m�E �ޖw����ɦ�������S묺��E��7w�-�=d���7;��v�qc�c��?�P@�OgU4r\�J���xO�k�}rFq �I�	�K5����������������&�y[��<���������<L�t���_G<�D�zC���m^���욜j�i�Aa��\�:S 7��A���z|�2*�p���CG4WTp��G�+!����ڷ��j_��Y?��L��⬟��ab��)�ąщ/l���M���Z�2�Bd�.��p+��!�B��S�����?�+�L��'e/J)G�ѕ,��0�&UEb���
��I<Ȑ,�֎��n�Q<���h8��A��S�̯� !Y�j�H�-��\qD��knzӠ�3�p5����g�?(���\�7�p%v��&G�Q�W��Vo�ڏc#�Ӊ�� tm�]�� ���\��'�7"&�j?�*�	IgD4��rZ/�Z9��sl��FR��u�������L��"�A��% TSx�hE�?v��#>?�eN8��xE>�|���w��g:��(����T�p�^��-C�rg�D�0�ʿ��X!r�Q��i�f���4�qa؛\��wj����u�-��Jo�7����A�I�~�f�k#��ʕ#�����λ���9]�w�C��fwz�n�Z��G^�\�"gN�^L���I=|��a�g��v�J�t�|�;�ˎhz��V̛/t�|&BMh�ŏ�q��J
�O���o6�-�F��xt�=�h���Y%Vu�1+�5FD�-��0�vO�ǝ�J0�Mw��O��L: �N�� �R��a�OԇH+�����n~���ßp,�v�7|�q�&�w*�(�&.uy��I�R�D�ƅ;�9}o8�oߒ�*�� �t�\�l�"��ͤ�L���.32�����ҷ���{џ%�_:�5A�އ�?@u���ߢ�G=�y�)YjuP��O4�Y�|��¾*��!"�-vQ�(��ƓXԂ���B�űR�7#�ڝ;�j �4�hh��'�x�������r̥"�T4�
��G�=�Wt?��Jow���cY���sg������o�a_�!߭7� GU���]�UnV���O��,�H -�T��0�����P���T.�]C��QPgϘC��z��bb} ��
�2(u�Lt&�P�`�<b�{o���Α�D0"���\��C�ޫf6,��W	9���b��BD7��$�GeN�V�o+�E�xBs��q:'׺�'�Kl�P���.�&���<��V��(��C����C��2993�+�<l�IA��/�m~��K�OY���H�V>��� ���:v(�.[<K$�Mu���&�p�XrJ�M��\dq|��� �"�7�8�j� s�t�^�k��d�M0�"�'e��$������A�ism���Bg��R��χ���7�~Q��R蓘5����6��
E�J�ޤ�J{jtw�h2�>��0�,��/�v���",90� ��y-��5*"(J���[iA��X�M�?#���U��E
J��
i����8Q}�<��ٔH"/ۑJڕ���y��UX�9Dx?Ex�|[h�~�����8�o�R��%s��t�A'-jv�l��N�=@pn�Gv�Y�������a������r�>|�N���$��4��b(�u#�z!|8<��u�#�<�r��d�@���>Tp�J��������ZT��[��	(����
(�V�%&.���t��,эCN	�=
,�ʎ�@�����\2�╹\Av�/�w�>��(�s��매(s^�v�"�]ɠk�=y��(I�NTΈ>��rJy+�n�s���H��d�)��Pd]�T�Qc��m�"H�7�4q��?A�Qd�q
��-pP�)�����¿,_,�x��
��̦������
qdr�Dw���?h��+��^IO�c��! �Y�;c�M:p]߄ER�}���)�%k�J��2`������NJFdh����x�?ͥr�!���r엝��D��D�pS?ܧ�J�c�}&��;]V�4�^ʵo�g��qkW>�G]1�S)�q�rp����+�7�}��(�8�-G�>�%��To��!�,~A�1�z�"�0�>�"��qf��`�%��X5 �w�~zc�#�y2�N�U����so�zxIw̑ɟ����7:�r��*��֒�>��}3�+���V(j�rg��z��#�5��{��1K��dr}���[ā�I'�*�Ċރ�}�y~�������`Ϥ�q!����\oA�Ѯ��oh���ױ�����uc���Cg	� A7'uf���VNaQ�G�����]��l�s��LLܳ? p�I�{!X��{.b,wz;V�X�ϥ���#�P/Ag��;�i�2����ϟ���$������kWSF�Xwi��Į�����M[ |����WuXlw��V-�@Am�Ck��g�Q�(KI��?i._}͉��x3�p��K��}Oi����!�������������P7iW���Ċ��'�-4b9�'sT*ɒ�Sr
<U8#m���[�:�܃�U��D�D{Yn�?�_�zy���f�N�{!��I`�.5D��N����x�NH�ڱ��PRWn�t1��Z����$��{Hޥ�`����+`>�:,�x^4!Ё+����*����3ň7ƻ���7P'�nBfjY�����YR�u�}w6&���rv�a�[I�`H�z �+i�BM�y���Ţ��8,k�7��^��4��`�ᬜ(���S����t'�7|HJ6�O��m�ê0ի>��FM�R/�X�h��E��B6Xg��M�j�bR��!���3��T5w�+»��{�K��{&�ފ�I�L�7ݭf\�*�o}��-�c؉�IJ=���Ôɏ�/�A�n�zn�+�e���nք�M+�n����r,���Q��	t��~�gk�3���(/��:h~���~�v;xpS恦�T���&��g'�W��#R�5�æ�NZ�\�?�������1�$�\~���_G~
����W+c��b�{*i�B�5�m�� ��lU�����i�z��U�����W��?������3���р�"�>�妮)����|�]�ң����&�kB��o�n��� M�S2�?�\�����[��ҿ&�.\k�Q�Y�썧��TTw�wbM��h�43���Nr"(��j2@�Vh~�q`��2q�)���
�Q0���T�:��Qr2�������D��
���Z����X�e-���M�4���Qw{��uȴ�Z��qI�q$������E�\y:����s~��wٟ������E���>O��P�3tH�	������غ���P7g�p�^�Z�ѝ����sJ�kIy`l�e��s����6{UY������E(�7Q@t�hn8E�v�[l[�W���={YL�5����r��Ѡ/Lf- GT�$8 j�eo+��j��wP�8�,d��cu���$�n0v��x���Q�%�eE����B�}y�G�q�no���̡����g6b�z^L�z-��ݏ���1����`�73;�2q��JE`��'���px��ş�&O��#~/����9!�>SG�웻#\��ʕ�<��ߌ<k2ū�H.5�qGL*�����>�w��g�?�W�i�]W����}%NN��s�(����_o�Sv-���GTa�t��	���=� ���y �<�FA�Ƒp���W�.��2��L��k�k����0\k,Y���ZKo��B\�bh�N�O:���PK2����<�i�j���؛,��\�@��+�8p����եmM�3��B�\)�]O��^�X�]���G��D�Q�d��V
���m����P�_��7�i���xT�Ǧ]�1;J(OGV�p�C�f�8�^K�����k\ /��C���a�3�E}�[�.�\�0�.��Z̋����� �-�)[��&_K�j>~�e��~�-X��E�`�U»�\�̝2���)az�uF6�8�~u�;��LZ-uk��o�<���tˣ{�ɐ�B���ҝ��H�Vqz-,]O�w/}$���+�;����/�=������|�Si7A�mu�H���"i�A�1~*��
���vl��G5'��+@�]���R^��cy���2fn6���ݟ�<amr�O\y����>�>�S�jU�rAs�ݶ���:0����a��	u���۾�48�lׅ��-��)s>��+|�fL��4����bk�8�(�@ZLi:}=��s��~k���tO�e��pu��aA�U��[��fH��i*���F��7�[��hj��ً��Z£ƥ]+�a�,��.�E�4kt�|6/���`#{2�&9����K�1�� 2�.ԋ]�B{[����
Q�1��6��I�r��/��l{4�����9渙jrN�mang˖ܫ����Z���H\��Q�XLk~f+��ke�U�>�327C18�K^M�E��F��1��&g���"^��6|��V�H����p�Lz�_���J�nD��Đ�T�{7u
s1��qh�]�U0Q�[q�U�_�@_{a�dղ���,.)��c,��r*�\��jZ(W��;Y�Yy�Ӗ-��_�j�Y��ۊ���i�t*^��|����G�*�eI��zɗ�6��/CC�8��(���JI2/�_���{��i�{�N8L,9 ,�[�˄w5"Hz���C���[�8�;r�5�6Mb�4&���@=�_~���3�6���L�@ �W�|�`}�����{d�b�DM��V���O>��6k�KPUd-}&�U�g��Ʋ���ܧ3��m��4��\��N�֊��S<Vߜv'��t>��w��n�W���܄�_�~�je����S"֣��sB*���b܇��Z���}�~m���*l+u�MorO ��5Z��:pV0�1�T����\ �?���3e/gȉmQN�2���d!�2�Z?���PY /�G�k%���J7u��w��gX�0��ǭ�)m�y��np�S��jL�gciܯ\�_/�S��r7F)]��Uy3r���@gu-i9�NBi+Q����-��$�>	m!�%A1m�29&g��q��*A��V�)����t�Q0����s�kr��۴��;��)O$'6�F�2�65� S�ŹMɘ���cx��[��ky�\`�O����v����R�߭r1_��9��e��1�/���#�ed���2V�!�k�-c��>��o!r�#��}��� ��u8�HH`_��/�����Eu=U��6k�T�q��R��7��������T��'<H-�˼�J�R��Ky�ӫ�?�';�E�@<�����OF+�a���볩%Q|��t���v�*yoO�����Q�9#�a���&�|�Zok=�O�/]}+����d��t�ma��u���:A���'.�{�ݢ.�SO��)q8��ԃ��������������g���x��Ѵ_vWƩ��V{�L���C=0��5E�9��H@�!���,��� �KiqG����g�{����	*Q��i�ek��C��x{�XO�f�Xs5��U|U��m2�Q��u���e9��@�mV��f�tW��Iݰ֖{H]���.��y�%wJv�����-7�03e��~�A�k�d��>�d��	��ݻ�^wɎ�82H%�Uz�Q�=aӮ ��$�<�C]D��o�w�rd�z����sĊwe^?��PX�0� ��j���@LӶP9�G��F�@�ܜ�V����ʫ?�T"1��P/9�O1��D[�S7��Lm���J�Po����N�Q��a����<>zrw�Qd�W�~�@Ð�e�s��H�o�"��R����Yd�W��a�M�I4��������I���!�-������h������Xv��,�̹�5��[9�G��_�1F���A�Lc9/�T���]���-��-M�UM˓ ��t��Ο^5��p�4j�$����߿1΂�V�i�X�S��<�nK�j���j�	[T��qæ(��A�Q*߅r��f�\���I'��_H-�d���������hB0��}�j��h>�=��~>��C��H���f)W�p+�s���J�u�k�e�$n��ԙ�?�]Oj� �t��P^�]�. 0�`�ti�U�c/:ձ���㷫|�y�ʍ�g��7Gά�MWn�&��/9
�����]a8n?Ɲ���p���c+��K)�J�S\��d���%+c_��3~���m6[/6�S����;�U8c���W*�_�'�f�ךu��3�P�b��$���hTLB,%�n��z밦��xt�ΑR�� )A:� J�f�C������$�$��8�F�D���y�뽮��Ź�s>�'������n�/��CI�T�K6�j��ZjN���ɕP�`���q���%>>��]gZ8E��P���*��|��[�q�ݧ�M0ґ�x�v� �Ɵ��FC���ETnG^��Q����ݑ|��_q:���dR0Iԧ! *�x��{*�|��l29�����f�q
%�2��61�\*�Mg���лlrփ(�r��ί,x�����)�È��?/��s:F�d�A��a��Mcf�Cwo #�['��:�Yx1H�dU�y�U%dũ�jD�
�e����W���.����P-�~pK�V��Ug!L�<.�[�����o��&Ύ:K��5�N�JK��j���DD�]�9�"^���tf��3�NC��HS����y�9/!�m�>���,��I��!�E���.v�x=�"Ҥڇ5�^�:�"eǧ�Ό쬞Ȃ�xk
�Of�3�g�����M<����ٍUx>wӇ���L�K-�ٝ�sv� ���!�G�/�=�t��oB��S ��E��?��`NZ�s��
jFg��R?R� ��*��+�?�㷛�}�r�T�6����l$��\�w�W!���Q"��b��}V	J�d8���-���$���1��9���n)�^�j2	�d2<*|,1��vw=�8�^>����8�č|�@�IRrE?�.����Vtou+���~�P��*�p��\�-���x��xr��Q��D����K�'�n���ʷ�t,�슸 BW3ws�Z�`B�G`Q��\�:�g� giʨ痁9�z��|E6Y
���?�ˌ�R�q-���G4�+������˅��ۑ�,�XE���.�u�.�}���yɚ��s��$:Er�٩��Brض%���	���N�C�n�t}6q*�����Y�S;ة�T��]�|$�EGD09����g�*^���wރ	J�Q	�&Xt=��$�[�7�4�07�E�_HQ�-#M�7���A�-vv���oD���{tc��2�d���`uw�MC�D	�x�R�NZ5���m�6�$�/Ig��W���h=/�o%*|��� /��������X#3��!}��
Oؔ)wÔ49���O�&�=k��qg38>j���HǶ2���I,T~6�p8-h�7=��$k��d!�V��$%9�_�UN�y\�3���v��mqt�g2e9=	�]4����٨�m�J����ǰ�Zo<6��y�!�É���cUi��F����[�+�%����Sr�R�g�c�׃DV�X�qx�XV��s�zUR���2gl�Cˉ��
��;pօ�ު���o�1;U�V>�]�ז��?T��k�5�y;W���ʫ��k���N`ӭ +jt���ƻ<�,Оp\�\'Ul���&�NY\Ui(Ij�%(��^�$夽JS�F��6�ң� �Y��_�aJ�� P�rȸl1�l&�Y:�����ĺ?H����h���K�h�/;��wH����?�h��,��K@ϟ1~N�gOmōͺh戹�ݖ��LI�������v�Y�
b�����Kz@B��x�GP1~���Aē�N4	����d����ާ���U�CQ'��[��BZ�H?"j5��54�C��V�G�ڐ�k������� �~ 5�1��B��1�exȔ��EȊ����A,���V�q' ��]���S����^�`m�ݴ����n,�i�#�뭬�����<kx��Nz���j�/'V�_ 
G����  �w�Y|"C�p�$h�ά�8B_�p9�1HJ�X�V3I��d�ig�[�ԍJ�ޯ]���1r�{e<fm-�c�U�=T(���#d��?�Ң����ct�����#(`m��L�p|Lv��;B�S��d��tG<�9%�c�y|;�aU����U�nw�����\~�3�����z
n]Z'�к��x��P�-j��Z��R��ϔ���dt.�,�h��zǷ����156E��C��@�v��@��h�&Y�r1&��|%LH�+�����I��g8L��ɲ���[����O�!Nk�Mi�,��/ɘ차�!��,����x�`�u�R&HLi2�\�lH������[��N/���7�+��9��F�i$��.FU�R9	M?�9���G˕��vE��2�H!kY_���4�=�r'۟:��\۩�����L�I���hy�ջ���E�O�h�[/����WfY$�C	�g�2]@�E=� �`�М��Є(���z�����!2jWyDj�]bE*��p󅇛q@��2�7�h�|�	K���M'1�*5�G�rxǚU�q,ɟ���8`CCz�㎎cY_L��.� :�z�I��*ǋ�O0�,lU�/�D�{N
�%�K$��'���rsW��xO�g~��F�|�ʗ2~�ړ/fi�G��]��=չ#��	���[����{�yY4?J���lx�)u���j[޸͹�I��O���?�s]x���8�iHs��9�!��=�Hu7�x�D�A
� �W�]����~�8m��>ḱv��S�8�I �����~��X��@2���N��J���ؚ�����[P���wD�⬂�S�����n��m5G(�+(�A����gd�V��eTv
	^SQ3�2�C{�:��霮���,X9���+��Iތ���Z��)�M�8���Q2'�&|4]i�b��[>� ?�â*�7V.��l\��D��^3��E7Q�
��L#�ޢ oK��{��$č��p=nޯ�O��2�5o�J,�4��bge(mRd��_Б�� ��{*'� �!F#e�&<vUe|�iBE�-�o� �H����d�����)hB�����ѾM�JE34���Ȓã_rHМ��	��U�y
��J��<��ɉBH8"�yY��>4.�*�N�J'g?Lkg ��H�'"�r�u�Q���U��3�����(y�e��ė,{2V5;�6s�}Z�ַ%7:��9�-tDU�Y��ql��y��+����Z¢�Z�a`1I�A��h�gșf f�>ņ�I��Tm��{mh�QqO�nOgZP�Gaۇ�H�Ā�(>sbq^B��S �p ���#�4|�]qI�d��N�+���3X"��'��q��8�k'��KO��-謨򘾵��U��DV���S��F�"�����OY�_L�h�u�Q6������z�|�0�"��[�ނ��� �l����±��D��Y�/��ۿM斾Yr���&H�����"���x�?�="���\ؒ�_@�&MU%�=<J>S�y)�LL��6��&��M��u7\B�Q�ݴ��zc��˙�"4��V���B��T4�JZ�`�4�j5ɩұf)��.�d�Бť�R]�e��"ͅu7�l�﮵���I��g�� <ڑs�B4 p�Ѽ��i���5�X�+=�I�ʩ�u�e�p�oc����e��]�咶�d��Ƿ��zض�Xb]b��q�LRo�n=�Ug��2�a��\�.��9��0�}ѦB���Y�!^~�Zp��IN#D���k&ْ���~K��?p�W��*��xw���H"y�)�6Ȝ�����cYF���ԘQ�TU�%�:�mB�k�7܆=Z��
��0�R�;S�S��|x�!�ȫ�Z�_�������vJ�g ��;�*aͣ��O⋭��
����_�̱���t�垄|���&�5�^}	~��P��e�i u!@�mky�D
s�Y��,�/���]�E������h�� -K#����l�{�B��Qk��GV��ʆ�P����gp�`��*�w��+���D��sU�<��$�e��}�!���Ljd���?e�ϛg��q�A�����_n}e����7���]��W!����'fJ!��Û��b0=-��)�c�����B�����!Ov���֪�� ��ɇ?����]gd�+�[�[�_��7D��A��>zi��v5K���(�k3�ɛK�����|���,���Am��w�U�e����ϗ�	$
i�*y)�SS�m�G��h~�gX�l�c�D2ERo}�)��D��fCɅVr��э�����z{��,�C"	���S��?��������s)�X5�$��&1H_-ctwy�� c�B��e�2�Q)�1�K��K=5c��C�gjИS�5��n�Y�&���z�(�s�[�%C�j�����g!���~d�J5t��L �xY�R�����^Qͥ:VM�v��㯷��u�4m��tlh�G|�����"xv���?O6u�sJ�w��s]p����D�]a6����𹻝�L��#;h-dx�x�kݻs��F�����"��:�-7	>N���:Gs�E4~�3hAӡ<9�1(D�(KI���V�i�e�89�~yA�縥��Kf�}|EM�9�K�X��"�EšH���I�I�̆I�d����,n&�n�)���~5�r�@����Z���l �q�2<ݽs~��a�t�r��*���4b��QX�b����zU[���p�����]�1#��F�S���9 ��!�3f��Le!�U�����)�c~Y2l�
XE�DT����Z�T����<�|� ���Ί�=z�}���.�+��S̢����j�迃���@�����SK����OF����5X�p`v�c���J�3/b�BZ�#e���{�fH���Ҟg�ʒ�TO�b����nz0-)6�~˂���#�r��'ܛA8�a���(� ����-�j� -�+4Ͷ6^��ާ��x��y� m�L��ư�x+�����lr�oG��*v�ܶ��!������{�!sxl:�z�ԉK�Pr���F� p�/���2�:��=���Q�kF��&v���_��s�^Zy!z����z�<Z1Q}p� bw�2�n��U��ش�YqLj����.t���n[G7Ѯ/!��Cj��6h�����v���-��+��g@�e��=���z�bn�`����O�x�-`i[
� ���<��_��R�K�]�x�8Fb��8A)�f�
I-Eˢ���.����$�q��>p���/hAR�9b���ȝA���]$�)��QӰӅ�I�C!�Nb$���W�"�}�Tf��rgV��\�<�_���?f�������[Q	�Ϗ����V���]��T�Ԥ{C�P��.�������V��:dNy��	f���B�ؼ}����q���ϱ�6��MŝW��E���pr��`h�<��H־��Tk�!�\��t�p�Ւ�p*�v���]����Σ�X�k+���:t&_xt���������t�{��[�N�S�N��Zy���?��$�{9��Θ�MV�;�	_	yڵ7�_kT��~��s`U�ha��m�}��+`�nj�Һ��x��|������W��C�?����F\� *Xt�ȃ��$�g��e�I>�dz(r$k�G=���j?�ӹSq�ӮJ��$I����ʠf�l]�ɩ0]zO�֖�ޛ �$t�Բs4\�ݲ��T45�4��U��C����{>���Ip��[�5�~6N^Q�wc��C�rO�<�~�h#���~PP_���-f$�/���ʇFD�����d���sF%�*s����r��Nmx�D�kAi�Hl4��~���Lb��1g��=oz���UF�n��S�1}[�:7#*9}�k�C�ܓ�.8���bLCz(�4}��e��T2�#��cfCf��"G�ZIb**����/~$�5Q�ܥ���A�d1���
ِ�F���FD'�1�˰�/ì*j:>�X(�}O�j�hi��Pr�u=��6^ټo�g�wx	�k�����t:c�Y��rj1��A���ư-���D�_�w\O��C����?<�-tQ��VN<�g�<"���0���rQ�g4���Wp�F�A�
�dH�P��TJ��G���OyQ�P��Q0ֹ���m=��Lʏ�:ʎW���\��D���D�=X��b������a�Vs]�Ku�h���+��9�M�B��i�A.�����=�[5L���A���r�p�8�d�\Ž�;�r ��Q)��1�����ݐ��RqA�҄���E�\"�U��ek�v�U�CU��S��,B�L�v]�$�!ǥI{���.h~y��az�����x�'�ٽ��������{�A�����WTj���UK��Ƕd�U����4T+�4v��̴*C��ΐ�ϼß�8�#�o�{ VX]�.�_�oPX~�j�ݽ���{���7WY�y,s^7
�HЇ�[�y��5�|�\)ݢ[�>�STw���?�2(�b|eE���	u� v%_�v�#��UhY%�"��Y��>�D�K��k�Giu�O�i����3��� _�=��z����Y���@��8(�M�	�H,�UT�B ����q=��1��t�k-�+�q�yύ�}�U��MG��6/G;��-R��uV�����Z�~r4%�h8Y!1w��;)��i���������G�?rFL��������03-H���6>��U�c�p4hx���O\��t7*=V��"l���;\��[�_�L�?�C-#�#y)�s�#Oc�>[(I����'�`��~�$����kD���WXQY X�&�H����̵q��.m���B�M���jpx�i�*!	欏���H��36V�~�h\��[��})�<�m����� d��J0�m#��*�+��wZ�Մ��=wgB<�w �q�8���1��z^�T8z�.E��к��g	'>�� �u5�����֦#�1�9x�wխChh_^,žu�o*e��j�"�فrN�>�.�К
�%�;4z/�zA �/�*C�P?�Gg���\�,��^�3-���ŹG��R�O6�"c���Y�}���)h�ĉ�������x��K���F׈�r�z=^�;z����� F��*N@BvT MH
����j�a�ըTi�1�Srgꐘ�_x\�6s�I�Ȟ��ū����ZT��ԝ�=�yz6l��7L^^YM��6�X{���\��T�v~�}��eLuxÃ3��ͧaZR��B#�a��R+O��H��/������5���8�G����(��p�S��Ds[�0�r�@����*N} w]d�U�5�+��0�Eu�R�f|"`����2-mM��1\<�B5�˱]�!&ٶ�@PJQ��b �ٓ���1�}����p�LhFe1������G��
,���K����B�ȸ\��k��SrLu =�c�Z��!�܄s]9<)Op�.���i)^� ��{��v�-��il'��ݰ6�	v�b����*= ��xۦ�(�l�ꢡb`<��һ�^�s�=ز�jb���IF�k���֗Y�y�Yc��G����23��(Y�B�L6u�9&2}X�\ XC��\�ӫI���r�R�߉.W��0�z[����������l�:����DL���x�<.��W&���m?���-��[1�m'B�%ݹ~:�_���Y9?a���Y�q+��Ky�ԁ[7�[���I���%X�M���ɹ��`.ف΢Vxr9	(�;j�<t��%ȓ -2fE�\i���ӌƛ�=�2cfq�Ɇ�$߹Y���x�#�2�C�����E)��9����?5���d��jR��Q�pEG�;1
�1��g��Tf'5��m*� ��B�?ߪ�+=��85��u��8v�_����HS�1C�뛝��ȏB�M��U�uxK��P���/M��ؗ��uÞ2�y�l�T�1;xpKN�N�I�IF]7��}zP����V����w��6;g�c�m�J,�t�0/e�7M(�Ԝ���R F��[.���(m���-���9��g�`(�gG�Yك0"2!���ٌ�X�N�CP"�k���#�i��
����ǠRF�O�,�%���e`e��4���������I�d/Y1����2�}���*Ft�SF!�j���I
���=��V��^n^;a�5>ڬ~W�C��T7z �M.��D��U���d��i�u�},QmD��X������g儘p+�m���q'���5�̫�KcR���b��fZ�U�$��s)�yI�0��&"<���w�q���E�xOV�ɤ[�ݔ/�M>:����b?�Eo,�hRϙ�����9��q�Vy(�S��c�G�@{JV��dE:o����?z��w8.�JM夬s��~�#��}z������<��#/ǂ����-�U*� Q����R��\����s�����%��5L�7�����a�ԦE���n������	�����p�c�5P�/�D꺄&�i�TW��XE邡)���!/ؼ9o�Y��v@��>�ѷ޿{�v����R��R�/�p&t���M7���P0�p�O����3����|����*������ fY2Gз�T4��& D�5Ii7ѭIa�u�	mzz����~�D^�~7��Fn��NptnTc,�Ƹ'l����[ޕ��A�z78���|�U%QD���u_O{ڒ�zF�����0�O��d'��
ri���.�§�W�6�Y��r���A�벮ݷ�+L��ԧݣ��_�=��8�6L��08����v`v5�yi2Z_��#5�'�(N[)\�Yl�B5�q=�65�A\o<��K�W�JH�5��s"#���I&��I�/ ���������O;��؀)B��D���
��s�o�wς�`��-��>��0wCcQѡt����w��\Y�iV0@�����A�t���NJ�.�V�5�jO��d�����g�v��]�*.t���Nf��&'��JY}yU�����2Eؼ#I�4�ʑ�ճ�����/��M#
I�g�D����t2�b�ɡOز�oI��Yz���/FZ�ЏM}��ʛ*uk���G�-�[�d@,��%N�Λ�)ٓo����r�q��93���M��n�>g^Jpv	 Nu�I�@�"^�=u����i�+��]��RLe���f	%TU��~��V�[B�>*+.��ʷ@ԔoC!*�J��j�^_�$�nc�����C��|!��x��ލ{_���W�U��TMͷ�O�[�����n[�sX����sˤ���@��2�XҎ���3\!��Ϗ��V�~
wT3zΈ�Ҏa����7���l��$\���k����	2U�<�rP.H�Ū�ۢ&�r�dxT��Ő|Pk�/����jc�f\��U£���s��]e�Zw�Up/D�q�;��H�q{@�>�ZY���Aw�r��]M��Xx�f"C[>�: �j�P�o��z>��@�՜�V�~��J�1Z�\!R=d�*�!�N5nMD�����}��k|��2�n��(KG�B�~̩�&g�y2�"�&���ze�{M��4��U:{�(���|�<'ٻހ��GO�Ty�2L�J�G'�Sܿ\p!����6�9����q�f~�z+v����Q|��)xH7�[I��(�ꕨ�%Ӧ7$�nO�����/�����D����D�Do�/W����{֖�O�=���(`ħ��e����4���)1��bG9�dd���\���\��gg=+����r�^����S7�V�+�M�fw�7��۳:bGW�,b����b���!/���@i��zXI��QC���;�2�T)����ZPx��.��r�����N&�����-�G�JX�?m
1=���D)��&m���y=�[�;��[��zuڻ����6���-(�����pU���v�����JV�s&�沵�X7t��h��LwO�W�)�P]'��HB'�
߈"�3[�G�U�2�v�?�
@�x�QG�y���E�^����Ǧ��uV�҇x#Nj�}�8�D��#���ÕF�XӢ��� ~<�>��%y�����w9RQὨ�>�� �˸�y��J�SIVZMxۑol�x�@#�����Yx�t�~��H�:k�n�` ����+�hc�ݫ!������	�NC�ݑ[^�\�O&G�'i ��[D���ܴ� R����E��~���:ԇ�MU�U��(xj��?t��TIY3��Vs��сWZ�"�⍌X"GăiP禙$y1�z�%�Kz�\���#LKl7
���f��e�=y�ص��~f�>�`cG��1�z�y��H1��'�D�&�݆<J�_��GA���%o]o1���;���N�Q�����:�bv�\�R��e����·��iO�>��������P����/[���@LvC�xQ��m�>!u?�:���[��8��%�o�c�����գ[�H`ȵD���	be��?�e'CO=��c���/��w�*���i�*�G̫PB��5����i��ŷ�IF�'����H����HǺKDKjco���ܢ#8��/�-���,s�Y�����Y�I7���I{�e2�]}��z��L���U�*{����2���21O�MJ�uJ�X,��z��.��l-f|���Ğ�;+�^�}���ʷ������ϱ�j޻V�k/I�'��_%�t @�0��(L���D|�4����N鿊�Nc�G�U�'!��l�s� �3������3�h�X��?�}�-o!s��( ��'Ӽ��T�e�n��#��z֯���m�մN��lU��iâh�%��C���,AOi���:Cz�˂ E�h9�{�霊]���+���"��5I��6�l�MvKL�:�)�gO9�o�v�aj\�8-���C�ov
��!�8G�7�?��Wi�BS�����J[錘F׷�wg�^��@���YU�d<_����<�	6��Em��'4BS�tCѫb�}Z��$�<�4<��w����~��%U��\m:�]�4oq���d�a�b
��r(���6�mZ^���u}ީ���W@'��23c�ZF��1Gae��d��~�[;y�i�����H�|[�.�Fn��U���z�X�S^��?�Ff���U%)9U�*���Z�w8#�d�?L9�����j�y�=4��`c���Pm|�z�-�N9r�T���L����A�%����Wd���L�
Z��9�3�y5OL��%	0r|���_ϔ� ����p70{����k^o�p���q��CS7�_�3�H$x�iek-XQ�Pe���&���݇O��έ܈mV�T�~��jqǶr��2�y��'�5ǽ���UY�n@�I�X��ʡ�7���B�Q�]�q;��{I;tg��w�&X#ߌz�%��5\���9y���P88���;�4I�OFI��j�?���N���e��`�� ���q��m�b��q��!��d(xӈ���ۆ%vD�b+ߎ�Ȑd����LK���H��,�Lq�e�f��x=-��Y�̔���8S�q�\�a��&��`:��z����n��������g�'η��n�����E�R�b�b�b�bw����*x6pZ�).����i�k�S��$ڡ+j����\�f>}n@d}{�H�OA�'�f��܍��Ť�O�����O� .�򨄈t�����Y�^����|��_���"V��6r�2�B�CA�c�����$Jq�U����z�t�F�bAյGȷ7�Qjhf�H��=e��i1ۤe��UZ,z�b֋g����ƿ�@au}�X~����w� ��\�l��Y3��XrzA\�,嚙K�!ί��-f \R� C�!������ri'a�����^[�V�6����M�'�٦�����IQ�2�^��R��,���|]�y��}�QŦy��a�����+�Ô�x99�]OR3��4�$K�~��w�鞙C�����J�����LcB���3��S|Й�2�;�ع�y�FM����+������8Ui[/Wo��戤&'e��@�z�ZD���iy��TA;@����3I讔�����8e������ɫ��`�^��В�5ȹ�s�D�t���hkd������kISЪ�ɉ�\�Q�&aN�a��A�!�V�WEc�[��#��O�_f�@��9���;X�����/bi�bi[o�>i +�2g_��㉝dĸRȆ�͙�j�7�c��^���²R�Hچ�W����,��q_=7<Y�΍a,Ս�B��[F|5��ЕӀ��HAD��Y�%cչ'�x�-'���m��{�z��Q9	���0���Qy����T+'5J[�t�k�ڗ���\R�����=��\����L��{Y����n�;�c[/�/#C"��*�'���fK(��`N}���!2W�����m��)Ɲ�>�(ؼ~�q�pvv/1�Tӑ@����DY�F9�~hM}��	"���g���	I��p6��OQ$��0Y��/�f?���8Hw��Dg�]�0�N��H�w�p��)���r,�m�/�Ї�_�_��g�JZQK�b��R^���}]���W_1��"��wN�)ND��O�#����F�;�q��� G��N�y" !��}�v��U��1I�B=?�t���mT�4>z��O���VXً@1��à�ܷ���i��\�qaa������;B&0�
�HJ�4�XmI��}��!��c㳈�ژG�R�>�31������}K�9݊�U�	�l�p�|�G��"E��_4C��<��a9��ҕ�n���^ n�c��ʇ���J���_�;Oo��IF2����>R(���`s�;C)�(�C-b��Ӳ�bײ�:�G��^0c��6a9L�������HU�>,��4�f���r�=Ϟ���A���c�����Kw�����Al�k?�a$ΈMP�0x�M�דoJ�s2�D��LvV_��>�[I
� �9?�H��7؆�BB����}b�M��Z��2�?��(��JJJ*���n�u��LEm�5���8���?�Xr4��<��}�.@��ԄC���sB���s�{b��&�z4]T��������/�&EM�[ýX���L8�"=ݶ]*]��IX�׉/լ�2յT^.�l������=M��y��-T[�ۘxs��I�X�/�$��qͿ5�゘��߫wE$S���T�/�?�W,{�<l�t�=̈́Y	���q�q�L��p��䑩�eҟW�69��+��G{m�d�ȁ��~{�J�M���+�e�����"*v�I��� �;�tVɮb�NN��r��*e�:-�3�c�0��?9`$H�Kn��a6����ɣoA³#r3���ӥ]�P����m�7xV�m�{����t1� s��}��
��'�w��(ǿ�6	x� ��8�_~"ʙ�
�<2X�'�ǘJN�rJ^~N#��������R���&_jNT94X��r�eRL�*����^`���.V�{)u��]��Sc�O���ʲ�8�xR�wN�!���η氐�3����q��t����̖88��-�(�YP5qʯeH��F.��2|R����V�ǈ�����l�S�8��N��n%���.̈́޶4MQ~7
�O�5675��r���.�{?���Y-F����r\NKW~�2=12Dwݹ)p�ŀ^��H��#���b���:D�IZ�6U3N�)�<��}}ނ����J�a��75ؕi�q|ax��#^�H�֋�d�@���v�bx�0����g���� �T�j����y\��A-�������t���XN%�_m2_�8����3f#��
<�<>2=l
�d�*��m����6��� ���1SI��_������6Dm�*򍣠C�:��v��{��*g/�TZ5nH�@s�!S{6��~�o0z:�H��������sϯ���"���QWG�t+|���q��vp��g�<+N��>W����m�t�F���5�'�B�*��:�����+������������DR��'�Y���6���ﳾcbq j&
�ˉ�y�hȼn��(��c4�B+_�D��_�.�#6�@�.|�\�4]�f���90�!zy(Q������P�%��/�x���(�T[#+e���!ߑ���/�/�D�)��mV���9>e�>z�*��7q[��	�n�ʡ���ᑧɽ��;���ڒ���"���y�Tu��Ȕ�Jۗ� +�6?�Y�x ��dsj�!O���B�F���[(���
�_�P����|	�R���sOC�����FP��;`\M����yk�ĝ�:�PF�bhU���!-��Ͼ(��p�;mG�Z2�U���p���|L��9�T��;������Ռ�Ѷ������(�@�Q�i
A
�mMS����X�y|�W_�A��)�W������G?���9���?��	E�	�qK�ӑ%�D����_�n���EV������,H)�qP���~F��ן��\�u�ʹ��Qɩ,���&�u��� ).2�q[�:�J"Q�<zE�M[�-G�9�Srɦ]�B�Tf���dwP�}�GjI8�s��?���+�$и	2�b�d�����O?`۱M��K���-�����sߛ��:���;�,��Pt����d$��7/-@r���7e߂�˞C=0��o�e>�5[��#wu�V��?�������C�G?*B=;��H.f�O	B��&��}�T���h-"�`g>�&wCk�&��$��~�p�7�>��|�K�&�Ɛ/Ѓ��r��ҝ�1E�ׯ]�7Wi~���}QC|�Z�Ra%�8G��ƈz���Փ��)���T�L�\#m��~��A�$	���nz?j�o�*�³:������A{���ya�fU���d��4�����R�6Ml¾��6R�[���� ��ڼ�ڧ���U�[KV$��.ῷ��J|X;'�$�{m�|����G"�ɂ�?�,��V5BC�������"�޿�c! �l��N�@H�g�pt>��-l^��� ����l0.)ϱ��L�P:^�5�����|.��}����)��G��G}1T����뭻���-�$��'sw�H�D��#��쫨�Z������:N뭷;�_?�Z���|
L�S,����gB��n��r2xw z'U�4�(j����Y#��H�c�kR"�N����u����%JJC�*z""��=������X�����z��~�~���*4���O��}�JU��(��}�ҿ���/F%i(!�h��jQY�X/TŪO7��ɯz�_6R��0�2�Pw�w"&ܑ����W����q[z�"6����!��Zÿ?%�F�6�O�N�7=@�QƂ�kb����,4��E�R��a��V��'��B�D^=�5��k��/������N6]���T�jA�H_Mw��&@�"y�u��ؤ(�����N|��
�=�C}L'��0���D���.A\�BI�I1IEt�۶�#	oꛐ���x��wܕ������,�N���J ��y
AwNQ$���b��sk�L57���}e� �|�c���%�״�������⁧+�[������Α�f=v,`���g��z��q�e�%c.�oOX��NI������(�/�Zm]Ú<s6�+')���qOk����ۡ��ta��0��Ty,�C{���s��>�w��"��È�#����O���5Ʉ\̚Nlwm�����'�ź�yt ��ͩϦ��eQ��/D�腃7�f|�"OC}֠}(���#���,�c�dŮ�������>�kO@���#[�^/!_�pN��������Y�O��+͘/V�.��qr����m�=�����rmÀ2gK�%kbQ�;������_�À)��)��Q�nٛ���;��ce�^�l/'<}�V���Ɋ��ꊛ�sTz<|�	D�AȬ؝\"�����A�l� ����b_3��
"+��> W����l)��[�T���V�����u����	�&.�|�W$�N{��ӃR�/�/^՘wD
^��͘T��	0:��٧���t���(��[�a�����뗛���Kj������a���&�>�a���6x;�9G����8��)`���/�δ�ʘ��=�_ӑ�a���F���A�1�U��ή�J���g�������5տG��Ȯ	kׅd��۔ � C�H��uC+E�����d��R���4�bvy^����ZHw^�B�Uvҟs�8��{[$je��o�B�u��y$��u�������}Y&�o𖤻�Tʹ�����{�q-D�o�1|,���i_�iI�ZK-8w��œ?6�ԕ�~q�;]l�]�>��n!���Mg�O���|�
b6	Ӈ~g�
��51��t-�$Eۘz� �[�G1�O���4�9:V ;Π8�f��C3B���"(�X`�ta����{q��-yŸWE�O��͋w�ɐI���p�z��ϼ�*پ��tfA��!rpo�'��V���Hyy�1&�t�9��e��+�5�,Ve��۰�`��`��8���E�f?xz>p���G�1P������pf�f��,RG�M�f������;o�/��F�����f�ܢS&�|1\�	FȦI:�u�A�$�:���j*�����5�֒0�:���*��F'�9Zܒ[��w~�a�tF�b��.�Լ��"jv�T���)���!	�ܹ��]-�-��(s^�K���wH �>�?�j=`�����Ú|�x�n����ԀF�t(d"Hw�钔$G��!�-�)!!1)	)I�3��s��c׵w�{�~��y��k�����+�r6��У~á|��.��lK�Bx�1��a�}l��	G��>(�5)��Ǌ��2`#�������_{5�M>֖�zl�L��I���K�_�x�z[gE�E{�B������/L���#�c��<�r��2��]���G�*�-�+�P+�YU	�!Vc��ĝ�w�N��RA���5\��
�m���𵕂Uף$���O���>}
�,+�A��{��Ԁ��bm��g^���&�����D�s�a|�6�RZ5�p���w�.��n��s߹������h(��q�by��ɴ��2q�,���n�~-��"��tK&2o��'�g�S�	��X�G3���9�{�)��S�1aK���8{H�����H�f�� 5��ׯ$A8��xD�Ie�,& �k�(�w����;����fΔˣHLf�pm�f�P�?~�wb��H�y&a��wbR��sk�B˕�̃�ê=��~�*�}��ڮ;�����%���9N!}�$.!F��/��F@5)����b��ܪ|�̦�'i�`�2��.7��M�~^.��h���p�#�;�S=&�G���כ�TL_�M���e�e� ��p���Gb��X)*
-AoU�g�>��Z���.H��I�_9 �U�.!Ϛ�k�*��,{���ó�f�X����O��=�H1_{�䙖*�f���s��2���/�)�=-�A���ݥ7���χQ%|C$}�Dyn�oy*�o��bVOa����~k�E���cPl���ur��/ïI�\�,ȝ�{�C����6eo@o�SL�کH��a+�=e+WMܴ�F���Z���l+����u1����[��Y�%B{�2_f'̞1��e�z����'�ЫM �&��oHT���p�� �{I�C`%6���E�*����	��3����n����B�� ��Am�S���k�;yS�(�P����R�ȋ�>p1C�� ���M�������{gU�����9����N���_Wi�2�4��@ɯ�N|V�"�d ��f��~��j��8��0��3��+Q��u��se�����{����i~1:�^�_2T�jX��9U �b���7���iqZ�6�գ��թ�P��s�Oa�ۆ+�N���*|f���D+�L0SJO���P(�:���!,V�Y�`Q#h����R��B���찂���Q��\OIݨ�"	3!�%!�e�3&l�CЫ�q�g��g �YLڨ���v�f� 6eq�ID�
�W,16O�ܠϋ'GP�sD��AH��Q��-eW��p撮��!7Ce}�YJ�#%��^o�r�BQ��=�'���ݷM.���e�X��!{Y�b��(޹��B�������@���<�D���[�����<�6�ʱ?�y������;""�X��hbw��\���������Fc�D2r�K�kw�H��6��2z�WԒ��#�w�٥Oe�J5{fcA%�8.�/��mj	��p��KIJ��FwT>�Xh񩭒��z$1*me��R��K��������eG��:����|��Vf~N̔�Z���bW���7����6H�;ʡ#�E�T�l��~�{Ͼ��6����aRg1����.��9 ����<�>?��Gt�'�'|ϗ�v\�9�G��2NK���W�c?��a�ʐ�\])�J>$�e��@�h��̈́-���{*F��,y�j��9��Z��>�1큥ך�S�q�cS�|�`e��]�[��� X'�[�S3=*�+�fu�`��뵊������j��vz�<c�i5jU"X׸�h_'����"dj�y��wGh<������\C)��T�i���⡪lc��އ=H��K���S��*'�{�ܟ)	o��5�����H�;�7��1��[��9Z�)2���	�I��p߭�8˪ƞ�e��f�U����D�����5z���P��`����޳К�E��?�OX�Z�6��~�	~��p|�����è�Wg���_l���?ɵG�w�c�	���\��#^�]K��OlN�R��au��}-�M+4���p�I����X��ǉ��1}EI���M�vU:�}L�8��D`Jw��a�ʥ�{xl~jK#��
�� x�)n�oS-�8�	N��Zk.�b�W@9$��|�LCY���=��E(U7n�4������}'2ݼ�F�n��C8�:�u�Ţ���b9�w[��_.�*.�d�2���U��'p�s%qj3��Ls}v��ٷa1��^�G�mԖFk|B�U��Tq�IF�-���fC�&\M-B��M4��\R��l慭��g��r<ٞ��z߃��8�񈣹��ȯ��$�?9��Z ��M%���л��Cc�����^���@�?��aIv���[w���k]j��fԷ㺰��< �3ܬ���M��0����0@��Rn��ߗe��60�?Mg4;��\�+�h E�����O�ȋF_C�8l�lG�^��W��8Y)�kb�dGgL�z6�.%�w��V;�i�j�yG.ڇ����6�~���e�������i����ιCs��EN�4I<���b�G���s� �X�_mZ�R�Kx�w�C Ù�Ms#�'O�+%��W���UT�X�/����0����J�E��}6J�����$\4@k�#��J������V^�o����b����7��,���(���-��DI�>G��4��~���l:��?/����L�-�cD��	����>��	�$�*h� �$��],��ݱ���٦B;�������킦�|�{x�*�i���{g��}���Y�s���ҝd#�f�y!����YM�h�o��;D�[�<�o�ď�[�LΎ`T���F6/�E�f����y}���(�{9lj��4�x��i~s�����NZ.�� ]h9
��X���LRI�!���)Ay�S��8�� ((ԗ����1���c<����>�e�yTf���W��Qlz�T����W0T�����v:��I�o&?b-��zn��i���L���?�dJb��a�2/�%ٚ��OV�8B�\��T*�T�ЄveU��m��,*��}ּ��mL�?߿c��*�A"IT����B\$a�y�>�X��u,К�>���-�=;U�#Z5Nj�CД>���﷝t���KN�CH�~���l��2Y~������$��}�k�	��'��nh�S��Q�b^ZG����r����%p����d��)��"���0�����E�Z(}�r ���k?)���a�K,��8kd������W",r������c��Zq��0�[s&���8HJ�����ȵs����'E�ĕ	0����%��h\.@C2G4�^�ͥ��:)a�^�e�ڳ�/u�]�b;�;}a�QW"I���_�̴z�ӻJ�P��&8��5�o*�9��9꾹����]o4s��c����	0MQ��!;���D��PY�Lt��=[��.���ǳxM�o$� ��Qjʚ� (źN2�����!� �#܄�y�q�qS�7�;B&�Ą|�vp���/uw+���I�i^m��C?����� e���ٯ���p�w��������	|A�u?=?U�n�����t�L��/�m}�L����u-��c����� @[P.J�^'�ss3�y 8�,%�jm��&A���(�����K�߿�U�5��5
w�G��).�F��_�p��?�1��Az�io.hM�J��/-��E�����,��Jؕ�Zf s	`�p���'�þKG:ɔ��)���gS���(Rhe�;L͂,s��y7q��}|B�l��4%f�ы\y���Y�1�����螇`p4�Y����w���n{B�Bk����bƙ�ɒ-�7��e�1�۶0�����ThU8U�'�FZ��9Ŕ��i>^C�ius�n�	��X����݄T��8kE)�4���B�V�Q �-jS�U�-����ĉ
)��&���<,H|�>�Fܽ�[���{��o]�4bt����y��"vnK����Zfgꎘ��u{�Y���`�Yi^+�)b�Y;�������	�h��y�mvr�!f[�Y'C�$ڭ���c6Jyf���x��k�vMj㳒�ڤ�4��U�kĤ��I��X�ܺ$1�����h<�W�^��ʇ0��Ш�4���e�ۑPC�/2Q�&c����?G�ز���Şo�-�xKw|�(��C-�my��70
lAN��q�б�1r��K�喾�+��՗�r`�i����P�G��,�L
z������$��{QC}x���[0:��Ys����"�� |D�#���:���YQDx�}��Z�
��(�ʇZ�� Y\CE��~��dR֓6j<7��_�IHČw*꯾H�d��a��|TX��Mk�>)�@9��=G�C��ڨR��A������P�3�#*�}���b���Hly��^{z�*TuQ�jR1}*�,����f��t/���������B�m�@�dT+bsg��7|
>��{b�G���M<�P��=�Km�[[E0F�q�-��B�D�_�N�$?մ���$���&��A��-'���I�]��,�b���4��}'����V/D�;���!������^D,�l�o����3��ҹw.��n����'�[y�������E߃m�v�ǌY���T8�F�#_�eO_�����l?�~c|͙��vҌk-j=�vb��"��g��K��1f�x���H�ɺ����%9Z�&�21(	Nb/�1��eg:���zS����`ꯊ��ܞ�g��2! VvP>���m��e���g�]�*D���H�=8v?�n���B� �|z���W����,U!�=��F�(�Xtu ��j�~Su �-�OD�_���) |�Zj��-�c\Y����N�H$(�Z-%���D+��Ѿ}����z�6VΛt1J>��{�t�a�Kre�4��s�d{�AOE�,�'��o���������Z^Ts�lCB���VT���:�;�6HO��ױȷ���c(�St>G�������Z~�u��iF[�`��������TŎs�yް>-��Q.�{Os�*�g�S��_�E�ysP���>� �O��i��B]M�wG���������Z�>U�Fymy_ޒcڽJ��me'x�s���͟�B�UKB�+�J�2#[ ӣF���| #�PP�P�3�W��/�N��_'��3�P�Oۨt��`�����\D�h�)��3��.2�ϩ7�0�+P�c�\�,��%J����E�w��%�K�����%�h�e7m�iRs�ݑem��Dg-�$M]P	���B�����&6�������)R�UE�NR*��
���I�;��E��\�8�N��/2��J½�^ёD�������[o�6?�!�&��=�G3��<�,�fx*bG�۷=�ujE�� ק�*ʚlm�\`IlWĺx�G�q� ��>f������_ݒ�ˎm\�&��<���W�:�
�[���\z��}�3��\�)L~�pY��\�)�Bs[�ը��� ���j�k�8���a����J�<Q
ڛ&s������R�ȩݛ}�� ����\���g*v���Y�m{B%��޻���Q���qê�o�Z��(&�]��^�д��y�5/$�*��?�Tŕ囝VF{����a�(���^��`z9��h�|U�����b��SDR��>�3��m2G_����y�����{�1��<mVb��
�=)��8C�^�25�&Y!�!���&)�@Do�!����q4C
�٧��񣨴����h�&ԋOB���s؀2xA� �=u�ILk�`��6D9R��v�����Z'&I�R:�Vc�_��L�x�	� ��E�\쌓��DI^�r���i����D�ِQ2k�Oa�����m���p��"~-L�s.�>qJ�L+��E�	�I���އ�x9�d���c�{}�/��[Y�xur� �^��V-�tk[�K��:��𣣮��F�C�XS@�z�NU^�H�?^�sϙ%7�3�L��u�,ޙ�=w�oa����^�Sb�[��eG�:-W�:�;��jU}ǚ��x�f���<R%�u�edA�z��ot9*za����?������W�?��6�_6dɆ��Ƥ)Ӡ'��-}n������~28�U�%ղ缛�a��%�cg�'�}��W%H�PYpPWW��_���u`�Xz�@�H5����S�D��C�HH�������r�l���ƅ��D�R��n{�
Tu�a��R�J%��g�e��g�1�*4g�suL��:�kJG��y��P��|�aV��qT�EB�u�������Ay�������^7k?�\o������fe�(��>$z��N�٧i�k&�,X'53]�*���
7xؙ,�y!��j0U(��@��%�v��$��c8�/A=�Mv)W��g#�N��N�%�t���; �tp�{��=)���,�W}��"��@�-�&�^�C��ܙGN<��oT�Tݶ��}���o��Q�jS;m�������D V�������o���܆�D0�s�ՠ%"e�����%=�m�2=t��F]5
�f���3JZ(�SҖ7����Zw���`X��O��'��%\��s��D��>���i'�� ��ڦ!��-/��(l���c�ҝ2:�yI� �nY�R�v�{�?hX�p�c�(A9��Λ���5��Ul~�ZiX����@ >v@=�:��}�»Zo�\�Z/^��б�>�nnE�n��?��y��sB�U�p!��3��_O���ň˰:���E��������+#�~'��ǃO�,X7�*X�rY.O|����B4�:���'*0�m��<w��Fk�?�����TP+C�2��!qI���0�V�0*:Qf9�������;p"I��v6����fK�,�)ns��;��B�{vti����MRj�6 ��w�ϔ�*����Z��������!�Q��̆�3~���({��~ ��ח��h��W�sU7�1�W�JM�ch�ǌp�@j���c�,vF�T|��(g� ��3�&�sմ̦ �1��&��VS����:��r%;Z���@{���[&b��!�0Y�R����*X�k��S���/�ʇ�/u����(�tH��н@�}_�d�g�W~<���De�3�ƚ`ls�)��#����L���c�qҍ�<f�U�׎#�׊w�P	ߐ��+�jG�UH��6��:Y%�X�*�E����|#`-Т���-��ϧl}oCy�L���IIk-K�nZ~�������S*���[s�h�ۑe�t�b�5��E�C��Si0#-��]��- ��╫���/���楙L��R�~������F��h���3\hf�]�e�?�܏�}j4�גP+uNЭ�~��v��ܻ�KM�UL�.͐{�J�m�4=�m"�JXwSg���
V1.G)���y���,�*Rw�W�;���ÆF��Dv� %Jף�ŋΙ�X~�GJd$�m��������g^A��n\�n�R�ST�,���
�Y-G�Ʌ�����H�ZS('�XYl���r�SA6BJ���h��Et�����!rt/�7��ށ.�%'�9��D�K^Rp���3|wV� �G��HX�PS8M��;����*����;A�[w.>cݿ��!�tRhO����4�:�s�up�y��g>�yUʙ�.���~��Ҋ��Y��ѩ8�8n���~���~�bkg9��ZD�'b�R@]\{~�׵�؝��L]�#���U��f�~�t���T����֧Ng�d+�$�d����6_&���vy�4�T�z�0� S%��R�~��t�T]��d�Ƈ����F�e�:#2���]�?��qU���V�Շt�<���/��6��m�����Bװ�q�T���lb 0o�5�b�)�ɝ[�֟�J�{��%�h]�CE\�torT��hP`�N��)(�i]����W��ԭ�Nzi�֭b5��|��5��OZÏ*��B �^�fI����!4/�ڄE��뫧���e��B��BJ�l�����ز��,X��>H�#d����w��g���>"�군���c���|R/T=xR�f��pw9�AY4e�i��n �w;x!��ꮦe��W��7؆����`�dV�ރ�N+�{��o�$H~'*�k;$�٬�\o��$��E�O�$x�z�W"cW��F���\ {d8��j���9B�䱥���UII��$<������j		��=d�F/a�@�֚ߴn���Q����D�h�s!h��N�������k9=�M
�N��B.��L{4�l�ڰI2���*�!S3�	��^mb Ś/�}>*[Iݡ�#>z��4��}��lL�QP���LM�W	�6�����������/Ȃ��_�c��SE��ي��W}�"5X5y�2ݐ�%�6@���w�jmY�z�����߭�js������`��׾蓡�T��Vv>x���G�?�򬥋�����hx���G��\�X� � �%���`���k
��=9��7&�B�-u��ka���;u�ߨ��GXg.N�䂕����!@�X@�88��k\h(�Uӝ�	y�s�/&�e��0�spL ���	�����߬�=�
��,}gq���4�D]b�̪�~�9��
��T�eɨ>U�/�¨_S�/��7s�Nʈ��O�=��$�$�������V[XaR�f�Ko��{�)	� p�K�>Ńp AAb���cf�n�Mp1������R�^��ۍ;d���%���!>����/K������J���r��dG��룱$�g\����Z+�����I��4p�C{�}�F�|�'�,=���sW����x�j�A����d`�z+E�@t�{�pi�W S���,�d@�bЪ���M5���mǩ�i�F���ڨ�M�2�I�ISr�5Ce*���v���������e{7bJ�L���'���W�%��턇P���
33S���	�Eg��'���<�����x���.���^O��A�F�x��C ��&'mt2N�lwńh�3i̢h����#�x�I��d#
��#ܕ�آ�$Ky���ѐ�J`Z�ꇇi�6�0�tiD���}�������8�.$5�F¸YFL�s�28�,Y�������fkO���v70Iց�1mZ���e-�u����̒@k�
_�.O��S���2P�G��è���U���W�Ǖ�����]c��F_���o=��>�7��=.x�c/�X~x�9N��D�0Q�� �x7����k%����~A*�+���io�T"���Ղ�y!ccR�-��_���E�x^�E�D���y���S����W:s����6��_�h����½�Ժ��VT?�@O�����	|��zHY\R�6~�.�6�۵-��t���?-\BP	1��v���gëɤ0���4�u?[t�����~+v1��.,�Z5R@�<L��i��W�,N��_nB�ʢ
c��G&��A�Ez|���^��4Ns*{j�/����k �{ˉ�T&�	�6����{����u�R�|�����g
B,��aF��@	�4@ ʜY����4	���
�2'lH�u�n2���઴�F+���S�V����-L<I�ޣ�| �Y4&	g�� s:�S��R $_ʂ�s =���Z6X�Gc���9���Չ�|$#m�t�~�V?�}?��M�'O�w����!b���r:ZW�jV ��:�]���1^�U69	�b�|���v[��=�}[�>F���4�)_&�m	�D�@BM}��zb�6���b�)�7�N	6�	����`���ٻ#J��'�M��Jz�՛�?�N)1 _����|��Xûߦت��B�4���`�Np�|�r ���"������>���8�<s�h�f���3{qMl=	qѨ᷇[~��w��� ?�˿X�n"�����ߧ+-q�� ����@��˝(�-��n���a��~x���'.��}����Z�Ԫ��"�x��4����1v��.�]`^&���b��ޛ;YZ|�-7A�c���qČv�l�:3am��H�ݷã,�$%=�!��}���#|O�/L��
����R�Ɯ����">�q��m6���P���(t�.����4�$_^ �7��N%]��V����.�m�� � k����<���hr	�I�#p5Þ:�Q�7qλcև�|F1����_�߇����.I�A�QT�ʷ���y�V�O������|�\d��[�ߵ��C+�g�|ت���>����;�ˆw���"0�<%�.�yc/��y:�W
G�e�X�63��})��|�qG��M�ml�&Ћ�����(@���Gjk�~��G�0B��]�*��. x}H�?�m�)�}�
e�Ǩ�t��D	bwE&Ak��HY�xM�Z)q2Gr����0�?Dʘ��<MX��#���V��6�����B���u��)1	�����\Z�=�5e�ϚX�Y/d{ M�̄L@���O���Mdd{�8��nMt�z�E�Ӹ(p��WQf�]V�\�+�u.ׄ#sy���:v��eS�L����*X�D�ǀ���u��<��Vu��j���E�S�ץh������-�u6�ml�2���䏩��.?���IO3�n��&�Dy�N���\�7ls����z_�,^��]}
�8�y�3�F:��0r>�X��s3+p�^���?���%�Hc���|�*Weڂ�ly�n���$"�	y×�s�\~�����t�ۋ��f@0'��������N>�D���D����o�#�d�D�^�u+G1_�����9XлW��b#��L;L^�Z+��2����@�,��>��>���d����,���\{��R�u��'�go��TZ�ha~��xU�,�U��"|��Y����d�nߣ�V���h�:��o�b��P�W�N�}ȥL������jTdF��峧Z���f�S���"���cb{���W�mB���[n���7�`���|z��E������VC���A���e�d�E+R�!����L*�{����YJ�Ć�p�����=���	�I�7�P[?{i��di����VVq�0����5�NN "$5]g콸������-��|�jd����Rl����Թ����O�=!E?�-#�4��)+mzec)'Cr`�0� �g�'����Ѕo�&�~�������	7a�s2�'����J���h��W��\΁���R���ݴ#����qs��5%����k�\��([:Q*�H��у=��o�WS�% y�W��V~j��ߙ��)&�Oš2[��w#����4����3��V�"�@�=�F��u.���GNc���SRs2�x�Q'5��D�Ե����63�4������LB�kR�����]�d��5����}I�H�RM3���_W���e��[�as����D�E��C��s�=t�Z�*�w���3Y�D�bђGHH����q\�XIm�qI�g����t��q��js
� P,���G؍��뱤�f�ʄ(�h4Qatvr�d ��/(��U�l���
��������x�������;��_�Ԅ I&F�6D��{��}gi&���[����>�Yׂ�B���gH����P��s-i-�n{�L����ṽ��:KiJo�x����`kdl��f�u7_�7Is�1k��5��1�Z�]��5��R�i��$ى�i0�َ�T��7�$0d�6ZE	��e��ZG6f����E)���QS>�<!��NM�r���B����d'uqO#`nB$���80ć.�L��/.��q����ᦉ����ā�q8Qƈr��Ě��`���h!Hn�ߓ���S�:2�^�la��
=a� �n��l��� ��f���%��:��@�#���b����u�3�|�EeE>w�5��"/Q}T�L�SU�{b� �q߃�����Y}��Kp��/>�^�=	��I4��:9��<H���$Y����-�Çs��=��"Q�vx`�v�A۱������V���iN�zp8�#!�n.����`4�[�4'!���/��E�>J� ������UD���޶*��H�\�M��)<�է-�VU�A��
!q{h�[U9
#f�i�����P��5����7Ip�`aJo1&���͙�(���"�G���N�N��J�/��0�wXU>";��uyb|]�	`D����l�����EIx�����D��6��3=�����%��np�=N��X�u>���X�13U���H��w-��gv��}����/Ѹ��u�D� �??�PG-w����(�q�O"4�d�ʮ*�z����
�u4:�u�����]&՗&[�9� 1�Q�������,j2��3*v�|�e�^Q6`���� �5�Ɨ<x�ը;��2�����mql�m��2k|�͕kσ�P�&zSO����#����K׆A��^΍�14_r�>��JUE�{���_D�!��j]�N=�R�^�1�VwO��q`�p׀nI�N��'���o�[��IJ�Z�x:���J�Cl.��T���p��:Xܚ;���� 0ɱaTDj��#H���7��<ŕ� �W�tTZ��|����ؖgJӺ�J�������A����������N��f+웘=�������,��e
ɛ7l��j!oP�CC|�����傌5o�3�$c�$�@W�|z�h��o�d��)��	�%�	�P��蕊����󻀏2:�^�~��2�O�|��~����x�qc����@��܎�`qLre�Dʪv�=N��Vg�\z^�A��ćK�6���o ��ȼ�c�����ؾyD�h��I
���h�B�=���˰�xɢ�KTc�5��`�Ԯk_��w��&��ID�[d1{�bnv��>7������~� +$�0�@�6Q��d�FL�>~�<��@��IW��$��%K�d%�ϡV���#�05~Іh|�;�|nFj�c�O�;s���A�E&�|CPמfr g2�v!V#�b�!e;CI�.-
X�3�D˲i�KE�	���Yy%���!#oR�=�UX�i�[�q���o���~f�/�-�����Ŏ������?֖���[���FY6�t��5����5ս����XC�Np����tn�l,��"5��v�Y�/��0���������m�]|w�c'��������c��-��Ŀ~\l��v}����8�,0�� _{n�H*�V|/y��T`��E��Ex���o���;�yN���>jur���4�>�ލ��I}�E���K1Y22��&�J
��^�n�|��ud]�)y�{�{��>�YB�H���ZC� !��p�B�$�v���;���3�sF����X.R�Y�%�!�O�Q]��px��4����=���p�|�6�V]6\�R5��D�O&]�#cS}}�S�$�z}M>�;��UV��
೩TH�tIj5�{��FwD�ǋVA>t�&�u��p��
������d*k��b �������;k&,��u�e����K��*�uz�%�_uI���˚GՒ�	��i�g`Ͽ�����U��MI�a�~KJ�`��x�5��,����N������x��ֽ���{/�M&S�Ȱ�J��r-*�GY�ڲeA�"�I�-O(�8�_��ZCa�k�Ǖ������R��s��bdV�Ͽ���<aZ��w�������NN�	j6;����#�a_z�W:_L��ʒ�\���N�8�-����Z��B�my�<�A/A��d[�:�A��׺yۚ+�X=X�ڇ��7���E���	/�Eߡ.#:�K�,mߊ^{4�n��W�m��~��ɨ�|�����!���8�!��֗y�ُ 2�B�D�ˏ.B&3Z�eíw���7��O��ߔ��Ą�<������%__�6�C3 VYJo���Z���@�$j���4?���~%\���ڟ�+����j�K�}���\�̲��^2ZJ_��]��X�&�M�$'F��8���o���Z.�ca.�M�|��C�����aX��h����jY3@M��:����R�I��������}S��΁NbK�)�m�pO��l��Ǹ*>�Tk��v領{Y�"��ʩ_����*�0y(+�56(��ūK�#�ցp<��O! �yA:��Q=�'ٺ�ߚ��M�l1(��I����ǃHI+y���jBN�]Ӊj��O��v�f܈6�l��V.~:�\ \ޢm6�p�fiX����|r�`�͹E
Mg��n{M�_�ǒ`۾�G����+����
՛�X��tˇ݋�?��!A %7U�s�NjZ.B=QS��窰�u{�P����?��l�lh��1\�� c���A1�Dď����W4j_s�~�\�0͏�)������s$�����% ��-����P���p�d��jBݫ������#�EW����0�;����k�5`��n��j�	�����㙛��zr�S��2���̼Ͽ�����$8�/l������f���=���I���dT���;�1fG��E'C@�b�C����UJ�N�@�Ωϸ�f��4�`թ����;�Ǹ�\�D��.�{��|pH���eM5�#�������͖qTY�����]6 4��Y������S��{
���� :Xf��FwX��Kl��4�i�I�Ɣ����w�/�$u��Թ�%ĩf�k,J�%�~��24��Wl�t��OyJ����`W;�d�Ŋ~Lgk���L�D��Ꮡ�Bb�̣h��w
~)0��J�h�� ��w��f_eD����{����H~�
��r��V�gJ�4�+휧����s�%"5k?��3��C�Z"A@6�ւ�æ4d�	�
GJ	�����}ڮWۙbi������	��?"�?����3��3p�=�
�Q]��;V�R�1�}�/6Ԝ�T%��4_�����%���t��:�[���ọ4����=2�$K�4�:jR.V���Z%�b��9��~�?ֶ`=�dS�;�D3g���:N4�6�j����S3�|j���T�7����^���^20-M�iM0�q��Q��²J�P�1�E=Ȯ`�����B�f�`_�puz���	��3[s����O�!�|S-m�tm0���'��R@¹�Ɩ4���k���_��Ww?��WFx�M�0tl�z�JBD>��ն��@��0�xP�9v���򆊾C��u�w-�i��2�0����ç9�b\�u��PCI�Q��W<����&���w�x���st^t�GL�H	��!BvI0x~�r�`Қ�J��7��	I�2�6���yF<"��"?�.��E|E3Bs�Ĭͨ���MQ��O閸XЫ^O"���xi�ĬrI�3f��\w���Adp�@�Cyz��	��W�GޗI.�__��GZK9��a��e�.�9E=� �j^MV\\S9Y��8�7�����Q�DI�_~ԡ�<4���`�.�LB=�2b'�e��\&���	�����l)&������%g}��|`S����s����a�#^'��E� o: Fq@S���2���ҏ�C�Q��è���v�k{.�9���U-��.�yV�J)ts�4���K'�? �����J���Yn�R�}���5�L��0\+� ���%_t���Wڮ�@+�	"���%�L2��v�_�
j�0�(���{
w*v��r����I#��=:M���t`�g�v��:h�� !ʩ�:4�5#1�f87`>|`��6�쀤�%E=��>����Pϙ�:.��ܺ��hT���ޓ6F;Q�o"sT�d�u�z�{M.�5;�[���˵�`��ۏ�zʫz޷�������3a�My��ǹ�e;_�_���Kb�i4[��.M0�?�QYz���~�`�-�v6�3hT�M�gN�h;Y��)�:k���^|�4�����b� y����=�S)���B��Ŧڎ�m��K�WRuu�u����
������?�SJMͩ! ,����&�[���͙��OC�Q%X`q�n\7ֹh��e��.$thO͟Y��O�'	�.��P䶂��=��EƦU*�~���L@ØSݾ��X� �6,�d��"F�>�x�P�7���]�Yj�;4���2 �!�`cG���f����,�����#Ql�Y����
H�'�t����z��A��w-���3$%��~�z�k�HZ��ə��?�&ǧ�%���R��4�������2`o��6w�p�Q;�ͨ��V�D��?�,p�F�+�.:�$�rW{Z?P+�	T���@�8Ev _��5TΕ�'��oؽX;>چ�4�^;Y�h���83�i���p2�<�:�H�NC\X�M�߷� $Z�b�c�c������g��cojԈYU[R��������5j�ޛ���ҐR%�޻�������_|����<���ܹ�s�s]��}��^ίd���8���9:w>�W��>�y���P��n=q^D �0��2�^��W�0>�g�8���h�g�vm袒3ٚk{��AS?Ҥ�QX?�3��Y\v*r&��(�)a���R��A��}�
(�؈?֔��E�� �U�>eT��w��'6ۏ�7m��p�DL��L-KH�oĦ%�(��ȥ�G��#�L@����	���F����G���6N���]Pbc$��9�J��yA[��;��h��|��֖��x?f���Z�+�cߣ�?\��}K���#"UWM�ۏ���R-��h��U�f�����~U6=�_]�w�����$#�iA=m�381��ޘ������jM���M�_�,��f�"%
��N��I@`l�M�iY#b�;��NI� ,̕Tq�������Ͽ���ۍ��Mv ���՝#��Z�߰m'��x8Wr(2 kg�g%�ݼ�2��/��񋬋�D�(ics����vs�R�b�%���6�����q����'\���ȋ�"���^�� ����z�rվ��p˛�"���Ҽ倐U�*���*%L#)v ���AՂs\�U�lۗYn�^�������Ś�a�h�K��t3}V&���RA���%w�����C����l-g?�L�]��(�]�����u�b1��S��#d~=)�O��IǇ�AH����v+C�H�[��{�vo�~��5&�3_d�3�f�ʏ�g�F.9!�Үx}4�ʯ.��*�N�PQ�M�zXb��O�GR��?�sYՉ:����@i�Й��k��d�c�)]T_��7Z�>��a 9#$1�I�%C>+WO�Y`�� �Ql@��.Ay�F�;��(
P���$ P�Mh�azw�$\�e���]ŋ���ק�J?����0�/��$%WKX�>���Ɲ�h���C���2l�O�q�0�ԛ�Q����إ�@��g���[�{\I]�ZjfҸ�0}�#�g �z�Ra*�~L��{��|�]��[�q�����[Fi�ymж�S�Ё�����o�v�p�.z_�g��Ĺ�E���@G
9�Pa�g��M較\w��G��E��)e)2��"=��K�e8�$@����u�ǥ@�%��˵
Pl���<M�dӮ5{Q��p�Nu����kPV���"�ߜ��ְ��;�a7�!<)�A��1���ښ�v�/�L�;g=�ݓ?�.���W��
؎&p�x>��:,R�u�yv�FAZ$�F8��c-�!����	U��O���-3��d�@�Y�I}�ߒU{&��Ƨ�!$Kۥ�Ko�h�(�Ņs��J��v��㴊s˛^�<��N�g��%1��o�)���.510d��	|�c��k�^�
{���J���r�))�������:Cl)�6�-��:��׬/ǖ4��)(����I^h�o�'y�"��qy#��l#J>3J�%N���������5�N�=nG�/p�C(͠�3�r7��¦9�������ӿ@3��
[��a]�!����(�<�0;��Д,9 �'��Z��Χ�����\�<fN����⶿���+�qH��� ��ѝ���!3D_	�Z�bu;@���(�)��2�ɪE�7��}����i�R�����P�D�/��˼T F��C��E��� >��Z,��L�%I�H����</ݱos+����`��.�	E��9*�c��J�'�Jb�R���-�Q�| V��Jo�O��OZ:���P����5Jo����_>�+n��S�[#��Ms4�v��y�l~> r�F��!�8o�s΁��ml���QR�xF�%	RP�r���E;!�t
T��8����e� 	�(��G��,�r9Ki�$��{pG[4�@b�Ǩ�)����A���L�iNB��$���seȈe ���q��
i9u�ST��wE�Nԩ�f��Kf�*LeyY
8A��t@u!l�&�nH%K�{V��l��`D��=O^_�T&�	�;�#W^��5	"X��P�o��J4�m�̭_��.E4���BBU�Äo�&�Q�f�[����;�u���v�XkHI�fĭN�\������cgDt��K�ͪ�uɨW�ҖcBw��<؅3z�.u��gd�#��Il����.�/�"��G<���)#�V���@�u�#���+�0j�/থ^��c7��5X{�d���wnB�=Ӭ�i.�md}����<aS+o����rZ��r�1���/�'����g߬�W�/��桌�!�}���k/$���Q�$]�����d���%�#�I��%h%$�`YY�b�"fv�q��2�"�`8 ���9HPf%YA
r��Q��xSI����i��ݛW/Q$�aaw�br���Q	AI��ܼ��%0�tEV$���;P]H�Fە��	��n�ӫ�Ze97n����Պ�V&G����hX���T����F8����&L�-�ưr��s�c���͔�Ix464��R�Y,�5H��	�E~l�J>�{�؂+e���j�5UW^�?=ɑ�^���#��d�]�E���z��)��|�>���_��,��h���X�j��Gt���y�x���c������f������8W��@\�6���Y�� _
,r��- !j�8�7=d�^+ �\+�=��D�gr�2e ;������mTP��ʿH�>���K%GŸ�qVs88�4�)�JO�S̻����W#.�Eĳ_p���(���['��HE��΍���\�P��]
��"nJ��`�ۣVx:�v;.����-B�f3��RF�����q��D��չTn������Ec�=�A�B��Q���=E<ݷ�88�%P��^�����L����RϾ�f,�������`�_����#��]�'��Ϯ�`|	��!�*�c�)�E�x$�uC������%#�X��Q�3��m�+(������A��q�&�a���0��J�C��
]Cwf~<�(<	��)��+r�6
�8h����{������d�5�4�ūA��.���@$�x����+!�v��N�@d/,����DrD($�is�	&��"-y�FA�{�-��S�r�Ŭ^xFpё�ԅ���n�}�J�Im#�R�څ״LV�_Y��5�BW�]y�z��A�_O%%S��0:�;+}�w�l�N� 2�M۾���`�D��)�B8N3����v����g�4Sl��1ĕ�~&�t���מ������Tc�H�7q�:Wp=8�#X��W�
����n��%�Z��y��������#-Fs��5ї;�t�lm�����	aA���ON]»7g���v�\
�~��X���N���~������x���	���&~�9����\'��4`�b�=*�d1���!vz���C��=HUS���W��_�&�GT�&����՛�%�qI'N�2P�&6���ov2�/�z[��h\T�-ٯ𤳉u�kU<nK�#���^z��$��@��w{i�)�j|X��N��@�=(������4:��b�u"��=����}.�Ԑ{�B��f�������c

����Ո�ͥ��/%����DZj8��� �;�6D��T���ѭ-�ֈz:ƣ���n;�?����.�Љ��S4V����'�Z�� JT�6"��n�����<sK��Mu)�9f2��h)f�~�ѹx���{
2�H2���� $��4�b�Fl﹒�\�C��T2��6�?���TC�߮���C6��*�M.��f*2T/�(R���y�IMR�k�͙�Ћ�z��Qx�l��H=2��Vͯ��	ƾ�z�˔4`,k�:���q��kb���ۓE#�k�^����Һ���PZ�����y�B��i�޳�`�����$���Lz�|������ggޯ䀧������h�=�H8u��/�-�{��w�#K�� %��q��1�|��1КcPy�nû��'s-\A����@�=��9�Y߯����eS�}�C;��}��x�%�fy6r��f.����Ǽ��N��v'ڡRy�����~�<���N.M��$�G����v��:��_�!)S
�L��N�R$�%vx���&�N�xv��-��>f��禮7ۊ����G�˰Jp��|"[��XZ�(a�j��"�[$s�g�jН�Lr���w��"�b)M�p�N�t�(V���3Ғ�..!Y�X�,�m�ĕ�N^Kb)|Z�H�ʢ��Y�d)c:v5Lς��a��$�̃��29��&U�ƗO�ð�Ճ������;��*�3�x�3��L["�/m6�f��5.,�h�ض�<a�9Q;y
�N
\�r8:�c%?��111j�������6o[u�Ϯ�v�Y�>�Zy֝%-v�&��D�{ ��T��':�}e�����Jh��Bu�W����{�����t�ڹ�O\Ol�#"�Vu�mTHod�z�J���>���n$��rZ����xnȷ7~��TH� |�NF
Î�=������m��[��7��vDj��ط&��@�,�����k}@�q��a��(j�v1��E���'�zVw���!|n�YA��>4�ڳ�ܺ#1a{O���J\f�0�$��뇴G #�F���Q@����َ���˟s��@P(ұ�f���ό}H�I(�:��Q�1�o�A&
��=����h?��Mx�c�%��#kg��ۏ�@&���_�SR�@�����$p�@�����z�j�����$5�-�P��9t��! �C�"� X{�&|^����`�9�h�FFt[�A`?���_~�֮G�Wo�B�"
�-�(�����.l�;=K$��S�W��yg�k��$e�FPl���q�2؈8g�e�S�?kY�cr�T��}�^�k�:��bF(�u���}@摶n��<�W��\�^>|t�~P�$@h��Uci1��V��.DA��II����"��X�E��NqJ�a~(z�5�t�aQ�I����p�i�=eG>M\[�c�0�ȇ`,#z���S�5<�ݚ=⇥�bC ��Lv �m����|��Mv�{,��@�I�OɅVZ�s��*�zk�������tl�����|��E��S	���u��Oh��{��j�_�!S����?������w_󺬫�����J+YȆ
���?��w^�EE9�*��ڛM�iC���&o�2"�����T4�N�f/_.*'��س�����=�H���?��3'j1�ʷlŜߍo.}��l8w	�M�<V�^�A�6�^B�Q�֩�7M�}@�y<�o/�����J��3�7x��h�A@���Ŏ��MA��
54Hu-�,�P�a(
�@��6�9;����Jb)H��2o�$��}*��V��{�|;$��Ks�\_�ɺ*o���mX����$��{�^%h0���ɱ��m�0Q�����ק	#�{�D�@\r���
�����UFW	Wf�}���������&��Vo����K�V�BY#�zڣ6W�㦇�I%�VKv�	&���]���f H�?��l��+�u֨ ���Kh�bL�{�6��nqw�6�C��˳��٧�V{~|���N���(�>�ؑ���xĎ��p~�,�W�n���+��]�R�؜A������}ѡW�Or��X�Z'�x�xa�&<3��o��P��������}�Q�XL�-û��4y�H��[��+�4���h$��	PP�p_0I@�ဥÖ�Y��%��C��xqۊ� �D/��;$|�m��ܝ��3w�̶�ʋ{�rY�I���L�[��)Q�U����w`�
� �R$:6<�3:0#��2��"����ά�J,Y�^�X<s�-Y�(��t_@)�ݶ�	_Z=���%�fĳ��QK�"QA+tA��ˡ66�����i�;0/�܇ѱ��Y@�3�-.�p|P�>�����l"�^�1G0�u)dv}�{j�CS|o$G��
�F&�Ң���q���?�E����v�+���be��k�=� Nse|�M� ΂v��W�d��(�����N�`�� ɷ��X�'ln��T�z���KX����b}U�s�:q����AR�0'�Ew`G.�}iNg��oe��ts�N��P�>?��.=aʥ
"+r�z2���/��W����޾� GZ4}�~��N>�Nf�`]�E1	]�.��4+�\�i�� ��$�I�5�
x؟���3S��zt�C��ꋼ�}��������W¢�߱����(��Dw���l�� 6�z�/�	�V��X|� ���n_vϸ^ %
I��V;��0YȚ��g��t�|��(=��L1	T���vtd �z�f���l�(⓳h����L�A�*Z� �X?Ӝ�dY�G1���(;2���LѠA�5�B�ϐ���'qZ��b�8УHc|F�b�M�t��*ү�yפ!��h}ޱ�`�s"N����4a��hB�������=��h5��>��7�Fl�n�Z�Z��JJtE/�	U�q�(��O���8�� Z$B(���S �*s�� .�x�����&w%�ǒǬ�IH�l6�ݘ��%�.��67�)2n'��v��������e��8�LB['�q&;�1}��G�0jL����|>�	����쀍�Ӭ�y����d��)����[���K�P�L�Bph��"v!ԇ_�}G���Nlne I��[��m�"(�x����2�_\I1`�����oآ�(zj����'�-�&�e,B4uq���-�0�S�t��B ��>5�NxE������-�i^h��&�R��Ǥk1�7�+�/G�v
�>�)�JRא�s�,2���b�G�?=$�p��:��+�����A�/��j�����+S&Oj��o!�͍5��\�S��~�1ӿ]�y9��������j�m����0
��Cr�M�H/ѣV�,צJk·�������:?u^�B"&� �������U���^�|������1a��3: �cJ��<��?IB�Q���keZ���E�{���������ޡ��D����%��=ry�XlO���#/LmJ�!!\?�u���<7v�;�xz�K�*H����$���Eֵ`��샠U�#г��YH�l�����x,�{4�>8���DF{Ծ�t�OW�-��e��A�-��-����܍�l��P)�>�U���dj-�H����hE�ά�4;[.��~<yԋ)<bqF��'=�Va1���#�H�n�y�^~�u�)�h#�H焵�/��
��?d��K�>(6>x��E:Z����}eι}<_�ԇ�7���H^�	�.���-�!�a$ψy�B�-/%�0{�
�p{@�",5�k�{����xd���HQR���UN��VQ|6�TlRW�g��b]I�����ÞQt� &�����P*�G�i�*�p2k�(w���1��֘���[L{2y��8s阗P���6#�VB^�������Ǣ���[��U�=8	J�|� |��$z�4 ы�x �:ߜt�Fɡ�=���"S����:�x����I�����߿�ݗ��s
����[�pDX4e���9��C;��F4��+RFM]U���ּİ�k`�����̝�@�uh؏E��ȵ���׈�"kap"��"�F'��#%�%�o'J�!_Rn,��)K��Դ�~�dCeމ�ѱO#�����#!x.�G('�����gV.�Mu�Q)����Q�r/K+�RQ��S�V��.��yW�<���*Lڮy�ox�P?��~n�4����ӯ�X���Lo��b`{����3�$:N���7>����INo��9܉���� J���[8�
$�u��
��^�q⪑+͖<z�H�zO����q��X����'�	Q��3O�5{ ~�x�H	���a-n��d��"�	�Ԟ?M��oX��,����A�4������6��Q`E=�i���ϫɣr?[J�i6�i�����iaW)k�W�;3�>U��)��`(����-�C��N�_z}/��/���V�V:49x����Jj����4���-����O�[<�¶��T�]=n��s����M#C�">��i�n��t�=ތ��w�R�{���x~'���N���d��|�K��@�4�sC.�.�����Y�ٴBN�v/�x��9i�=���i�f��2��1�=�H��H�j��Փ�-!B��pn�ফރ��%�~\U��Bm�sP�Ō�(v�fM��f��_Ns��BZKW�`�e�M�RW������Q�E��P;��'H�)Іk�ʴB�$
��5���l:��*�η(��7���3��*�@j���/�{))��`��8N��/��6�����ĳ�	-�X�د��&���"%'�ͥ���O`�90��{�x#�����
G����/���Tk6Ք˸3���92l�xْ�$zd6����H��^���,-~<������A�[�p�����R�q��a5��k��/d��{�w*>��ք��1?k������<���'�����D�C'�{�P׬�� ��	������p�������U�jY��y�Y����=�c���94�Ű_�`#K85Ӕ���݋ís��ĸ�/�ݧy�t�sP�%�W�j��ѥ�O5�@o'YF(]��o���m��)ﭰ�;�K`�Ȩ�¾��B��r�ѭL[B05���ٛ"X�N�KD���������	��{ѱj��2#/72�L�K'��n7�&K�M�Kߕ�q�:��̰�9�1���rj�j���`؀ ����	��x�P�`l�0I��-�o�n =˭��Y�7{>����Hg%KG���oō(���Y�B��u����`8�D��giD�t���<�o�zj��oݨ��sY�#b�-6���ۢ^�Wl��F��5����|����Τ����ݬ�W���E/�3)mɃ�Y��mԜ���n�;��B��� ���r���ȧ�Z�({p"'h���'���x����(cޣŌ\�
@��f����8�YPw2=��@�a�7�����a}!�ܣ૝�|A<�I���H�)tD�"o���4w�����m��6{.�;@���_�R���y�(�ݨ����_Bs�Ut���@�sG$�5�֗��5t:͍2�I������°|f��Bƹ�BZJr5�/}6i�����K��_o('"���\S���W� o��p��u���1��`���FR�����ىΝ�<��|�z<uL��p��4[���5�Fc2�C�f�8�����^n;M�\L���5�4�O�2��>Vq�i$�VGp��|'0�
�������=ߔ�9�aة	]5!���|}n�C)���R�E}�{E"1�|�m�u'�O�X/��J��ZE&�p�)F]�8>�K�+p�	P��M�cXuj�o]�]��ϕnw��R�О��f�;O�߸o��.18�J˷~O+!ԗ^�wg�@�%���rćIw����|��P`BM�Z�S�����k$(�[UYRp��Q?3\�-U� %�����3�O��J0/�V��Ȝ0�uks֯�Ӈ�,�J��pE�F����k��}��Rk��0�}�@rO82M3�J2�<�Z�*C�Wۻc�L�cA������l��fl@����Гo[�CӒ���Ejǋ�R���0�vE��Xi���?��2�ȅ���̀���b[=s��3$��r<䘦�|��4�k�<]��j!����3��#<����	�j�?'��J��D
��������� *>I-@+N�;Lpn��$��9���r0S]��j�w���"Ҿ�!SP�x�y��� m�ˬ��Ϥ����yU��QEu�S �H��Qm��2a�G��L�U�� Z�A��:ę=i�e �4�D�K;��((6?��L0��,>�:�TВ�5�c�i�(����-'����Q��N6����i%:�5Z1�Pn�F%K�����@x���L!����#**e��1b7�����8�ƭx��>���ў�VO�$1��+n��ʗHY�-�A�%�B�_������&��8���.�Ǣ��=�XB�Q�?ܾ\͙��{��A��=|o<��߇Y���>A,&����z{����m��}�/ lC��T7ɭ9X�}���o>���>�{{��5�O{�ɊV�h̮�͆��<����yXѓ@���0������jq���aS�3l7s�+T��[*ū�&Nd�[F�*��t��b%ꇯ��FTi�i��j�,���ٷ@�"�_<�5;Ko�*<=1�����؞�N��Z&�4��]��N`�GC/U��z�?��F��p�F�;��O	a�.EK��I��SM�.�ZV�k��&�pFJ	;<��+�2��Y�ɟ���3��D��a6P�D�����F�ܘ�H�5�tR�&��F�n>�>��,���&#�g�F%�z!ĥ��m�W���5�CiTD�H%FI�/M_��֬���rO�ft���M7�M��y�3���V}����>��!����@Y�y�����cm
X��Y�"4w�Am�&1����y�'��f;"����l���T/�VE�^��?뒝� ��UY�?�n��� fy������2Ο<���&����:�sk֖D��v��p@�����>]Ug_w:����ʹ�o������p��S�͚ �ߑ�c����K�
�Gr�����y$�>o�S�$�^�¶oL�Mh��a����ǰ�oN���Ꝟ�]}�P�8��%�v\��3������[��ȇ���ww�L�F��j*�"!�J0[Ā���@�B���qx0����0?�pC��5��駿�G�w�X^�k2���9�D<�뛫F`��%�%#��3�^��1�4�]��Ʋ2-~�ʡ+8�^�K��$�m,�MT�aݜ-`��!�?q��ѵ�����ɒ`�܄���������+��k�wk�=�%h�v�6�G��ғ��Gῗ��H�`2J���&�g��%�����X�1��uq�d&�ӑ���=�śm9(O�l܏��3�sx��xᓅ�W��T������B�{�h�5t�;0�xIS�)uT�0#��E�a��,nf��̉D"��xݷ�Τ��I��������<��̕-��L�'�nV��a�q�&\����_�Xʾ[�!`K_9z�U3���(S�B��aq��j��ݕ�������d��.�#v������]��?���p�]ݞԯ'5����2�'A�+3VK���P���a���x���}F��t�zr$�|$҄NA���4����Mk�e}�r.'ǈt˶t_!�I`�>F�z�-�<S��%���;c���Rg ���U\;����r�q�+�Ya�@D���}K�Xw�{�����7S�_E=	�h1&uI�U�AZ 7����P#7
+�7k��W��i�Al>����� y�s�%mэӆÄ��-��'�B<�r}�nvжq_��Gr�+�t�y
o^$�T��	��^��N���_C��Be7
ܴ�9��W�1�x>Y�4�>#
M��S�i3�cw����y���P�T_��|N!��9���uJ	�������ع�cW�BT���`<��wN7H"p��"M�~�^�@ܵYn�ߌI�I�'��p�w�V'�ٸ���g}!�����B�&`������	���yi��3�gY@�֍c �z�����j�*�'�K��1#����c��E�eE���UW!J�F!�
>d9��F����p�G����vJ��/�L�?I���T��c��S���|mo��KN�t
`���Z�΋+�A=�)�m���kx��o�L�pJ3$��}Ep%Ļ��q�s���:!�R���e�t��0-BK��&&�p��Q��dH<�gb?-#�ȃG��p�.0thR�a���a����t(���CNY�Y"v.�Qk��k��݌���g��F���j��ڃ���W��c�,�La�ʭ�[v�@%��.��S96`�`Pd��m���bcE�l���N&��c�~Uu���ù +���w{|u�{{&���^�1f���ѽ�޽q����ec8�e�%���4cwcy�y5�T?(~a2G]�ȉ��*mVFSp����N�2�.�]���?p������z[�����h;���n'KGv�*�z���9�)k����=��&�Ǻg]3`��J�����OV�%���y��2�:�C�%�9W,��opɎ+E��ZKC��xk��3$sISx�R|0�a�h��:�������t��T�ha8��'-8ě��)������B7��wp���$�{y �]p��Hw]�����z�m�&�Ч����� ���r�m��uY5��M�p#"(�]�m�	s��L�#������?ō��v�+�$X�*��Ǉ0�+@Ǜ-��w��"t:��#`���&���/y1����pA����oD�����{�@��y`�4�1�A�?�f��V�	��欫�mf�k`ɥ�e��$asJ�{4tPW�о����Fɍß;o�'�����r�}t�&���5�¿�,�����ƽ̂ٞ��9�������H���K*"�7�|����jƽ@g�K�o�F�ʜ�5� &_�ZWm/Q��5���J�E���r��2���u�%�-���R�Xj�3�� �Iق�H7���`&BE�]�u!������&e��j�\h��]����M[}�.����[����e�m�e�+��\w���W�+�f8C7}�[�\,��9�㳴�q���@;l�(R�>kV�37�t�Bd�E�&�����,��籯�8,����(R�mS NFκ	�q�G�SPe4_��f߯�#W�Ŧq��?���Ἴ�Z0�������G�^֌�{S˪ӫ�G�w�e�sI'��R}YH<%P;��ܩ{ӹ�v@Kr��b�"|Ї�_�|��@k�lE��}Dm����(bz��N�,���CJ��4�t�~�@�{�j���mtO�D o�V"���F�ã�x5_\�Ow�<���%́v!�����V�σ�dMә�M�
�>�:�6���z�ps �[�Ǔ��<�<AͰk��j�7KC�!�6�H ��Db���B`��eڞ��Z'	�%"xg�z�eL���A�ni��3��4�=~�gv/a�8qĹ��~��)`�R�2�������	���I]��Z��R�"�^2Mi%�[�a�@&�x'�e� �T�����0m����^poʷ\I�_{ނvث#(��#����v��!5���?q&^��1Bs�^��X����:���u�Q� ��$ҋ�p�U��yl�mFIʍ�M+$n�6h�<Y��
QK���if�cW���m� ��i����q7T�l\K�s�������M�獻A�>̥ڪO[���"V�u�\����qf�����ۈ�@��m�n��N�yUٗ&gp�!�`P�L��&��κ�f�uW��T�թ�K
�n{��+ ��YE̡)i������#����O2.�� 求x�Lҟ��#���2�d�"g<]4�7G*lm�A%(�^�4$J֯�:����}�I*�n�؛��q���P�b�z�e��Y�H�����Ó3X��Ol��w�V�?y6����7�S��H���~�����?{��w����#�>�S!hE�CY��Nze��eAÅg�B#���D�f�o�5�a���W=���i6n$��	�[�"l6`5�H�H�^1�����xS�䅽��o!�g&�W��nYmg�.�_���k�����d�����dE��G�D\B+����Co�mu3�����k!*}3����m�}=���
g��ES$eYd?+o�a�����)/�S��Ґ���l#�j��G���.�F���X��Ϥ0���b;��<k�$�#Є��#��v��(�~2F"��q��-h����	���p�
��N�&,0w����+�ު������@󵊁Əa��_B����$g�Bu=�"^�ex�����}aO5�;�	�ڧ�d� u��=�<�?�Z�$����{C�ӯ�Fh�$	�d�����k±87�3ū��^D��=�k�[9Lb
l_�c�%�L�4��j�����n2r�m��{ޝE
�X�@�{Յ����k�,���էk��Ғ��V?%�**�^$�,n�I�����@�A�&I Ri���Yd��E/��R6�=�����<?����﮾�Z	�� ���� ��8ްyk�|���.>���|�ʼlw<I�H��R�	s/p�Z}��"G�����\'�%������N�Y��g)g2h�q��ߋic�����77A`
h�x��wb/����=X�E��w*]f\3��^B퐥$�H\!Ѓ����UA-�ލ=\;I�>�Tv�����v����٠v��؀�E��#W�E��&������8	��֪�Y~p鵞B�$�bK��E��,�O�pt�k�� &��#�U����j�s uG
,X�Ї��q��������R��s�勼��9�����[���c{�	d����!��{�F�Hn|bo=�<|�`Y�\Z, �]
8w'��9�2�j~�ƅ��Wo�mG<���
���޵��]��V
r�<���O��Q��I8zĶ�0�D�*9KOj�OU4o�u[�I�����	�7���P�9K���r��{��P�\4�.��-�.�^`�	dۿD����5�����j�>��5 �T���P<&�l �u#�*��$D��y��$4�u��\V �PM�`����ᎈu�Y��-�����e� May���b^����"����)W��*7+ݙn�oi�jI5��<��5WQ�CM�rٜ��b#�u�ů�-Á��%JU �6�����������E,³N�2ܶ��<�[�ʇ�^�,'�Α�:����.&)ʀ��IF�W�4Q!���:�	1!Ī�.܆/���v�Rn�
��nC�8s�X��=��o��-���w���yi�װ7�˷?�C�l�:�����y�Ecy;�p����Z?��G/>V�&�G܌�Si_�[<��xA�l�ڍ�<���2�f��+s�@�Ī�.��ړ�-qC���9�г�m
DWw2sl)ٵ݇��l/��L��]'e�g{^��ـ�bn��;��!����%*������������S]�5�rn鵶<?űK��,�����p���/�����*'l���F�q�m��&��,\tc@���e��XR4w��� �������e^����7a�mX���H�&nVbM��uv��*fj I;��|ޢSJ��Vq�����t�w�Eաt����䧍܀݄�K{��|�	��B��֞cUH��=�Z�ӱO~��WLz�^g�K�-s��4��S�����3��-�=�u�$)zXqu�`7���8�FR��<�
G9��9u��fP�Yu���i� z���gߋ�d��nN�wF#���L��/l���wG�������u���Q`O�Z*�r�i�r��/���}s}Q��h�¥\���hz��0���������`�xw�tw�p���v�[����U�� ��6��Ȗ���!ҋ���/��o'P�H�׹��z3c�X�;�m���Ի'�)���X���ݓiZ-~�:�E_����F���������F���G�,#���G��Ռ��6u�(���z?�3�v�5�q���Z�TDp�����Q�{��p]E�� -1w
��3�{=J@�15�'hU�H_�T'�0z�N(�ѧ�P�`��B����f��狈�M��7t	hѩ���2���7D�����@��c��2��;}|~`�"|�~>����Un'*}D���z��[{�� �\˂�B����X'u[�HO���wi�RQ9V:�����b�L��Q�W��W����5��R� Wvlt�(p}��*U�A�	�����B�X���ؼu�(�=�5�k>�k�2����jևR��@�$$;!��35`�-"|�L������,��?/���{D�N�UZ+����-q�:5�Y���֬q�+ZU�[}k:�d� �	��8�d�#HƇ>�ƕ���d�U@IC$�w��}�:��É4��?��>�`n��^A�lA+$�#�ғg�=8�w��j0F�����ᄃF����J@���&��u�#��SRq��s#�'�3iEҾ�P	�^#`�kt�kG�5߻ĭ���]>����}�v��+��ϑ�������UȮTchdk>� \�Ҭ�yu����z`h�"�X�,�_�̵8��6���Ú��,J4�䟄���%E����s����� s9�,�Į��,����'��p���EuM��Fn�K�򫩼�ݨ'��"]r���]/� cԁ4���Y�j��{ qRʮ�o�M��U�"g�I��by�41���ogacן�9ЍҎ������B�w�ީ�/��ߣ�߭�CK����j�y�} A)��P�ׄ.�(�Z�i!�һH��.]z��;��A��p���sun�ެd��bf��g���ȓ�^7O�=��Y�_Qzh��Si�~d�K8M8���=B�G_��e� ����jv������8����1��Dsi�U1���C��g^�k1������n�u/� ��x�o��&�}�\~<�r�[�Ƌ�<��<�d��{�fbU�e�S�m6!0�vl�����=�s:(� r�7T�o�3�\�MX$e8��c�); p�Ҡ�&��t?�/&v�J�Wm����Fc>1wp�Ƕ�R�v���zM8NO�[�(��kçy�Q�P)X&�{�i�����}ze���wj��-"61��o���d�O�������յ����<�ڬ)�����G���HwZ��U��	�=;v�f-d��Þ�e�1�5$���j�3oK��V�F����ʎxO2D,�a������~(���,�R�mK��=�j�53C���K��N	C�	@�[��,�ɏ?���%o�n=J����y�����=bo��0Q��w�3j�}f��S�;'V���,���47:����dC�mA��wFIl�z��T���x��qh0�ì��ٓ��rB̓�&?��r4�'�+�7H�c�G�n:��¯Z�J@���E����i� �������������m��.��������	h�Հ��k͙�=���˒W)��� �4,��1*|c�LҠv�OK?�d�dq�u�ţ䃐b�~PX��7e���G������9}��$Q����$��-6+��3��戀�H֭�s]���t=k����A1HȖ���S�NTO�7#?��З:�㌇(�:Q}���~k�q�&��P��R����ղ���,E�w�ѭ��邙���Vd"8ȹ���i���'��Hv�������D�J�gm\��_���,�A&bl+]C���^v�|���b�f��)&��#�?�%��aMC�<~�98U.�ܙ� T�d�Z��M����&O��6�]4`�ݏ���J��[(����Xa�l홁;�'��έ��Q����R�H�ٯ���1d���-�>�$�/݊��M��<1�y�2#�+�>.��n���X"��h��-bK^��p߮��B����D�\�{dӿ�]R@�V���$��]	�Xn��`�u.�Ά��R�W��h��H�7�4`㻧I���,�\z��|�夁�$mȞ��o#��2��W���d�߭+��;����>��R��m����Ӳ��v��xG�����˪��d���[��z�[�+{��y����1��/iPg��8�U�Q��B+�e1�4�L� �.�Hz��"mvӖ�BP�q�B�Bd����5���Kzؘh�8D���Z�pΘ����U���E���Tj�%����Ɖ�������d�"ȇ�r>�ߗ�?]w�t�]�Ɠ�vF���Җ�E�,/R�>e���;8��~9H���������G�n�~Ǟ���z�2�[���E;��������
T{өd��ou}�8gh����0oH�`ÙJ;��=H`%�&��?F��J�U2��w�G�qo��ӣ���b�	�}@;�bn�d��n�j�������id&��)�v*Ix���� $|�naYS�|��	X �v<�����yg�ۜ܃�y��h_���q�0$����U��c��P��K'V�T�9����K�k�_��=&.x�`I�=�]�ޒ� ��|����wc����娳������c!�o��x��?�=ױ�ٌ����;߯x�=@�Z�H�����^��J�*��+�W)Ej$ՠ�Z���$�%j�>�O�n��B�{�ʓS� ����ĠP8R�GW�k|"��b} �d���{0�췇�f����?�]��w�F)�A�QV��Q�F���j-n{"�f&��񜳿rV���&H��_T!�;��A�Kd����{�	��h&{�.D!�ο�!C$��R�Ga� ���j��k�_��%̣θ4���f��%+���>ݞ�"�\����XAi�8�a���s�}B�����j|�����/�G�V�V8�����'���+�'� ����Lʕ8�o��c���.��o�Q�~�_KU��^]y�z��.�7d��\�3�iV0�m��g�p"qH ��s�	�����O���J�X����r� C�ڇ��p�2��R!����d-S;�1���g��;[�UCq�����rȽjf{D��WfK�e�ƌ��(���؊C�������RD�����+,H��$���F�1�f���)Nw���1뒟�W�9�6L`��mk����>�kn��NβjaPB����N_�X��-���-�.X)ȱ</�d��Ԗ4K�8�K�}���~����P��0�iM����
�YA������jf�����``V�{�K9'��p��|79����Wƈh�2�ܛ����"�e�P0��n]���!_a(յE5 K-Reai����^m�|'���=j \�*;��Q&O,������ZQ�],غm+�z�L'�xg�SO���2|o\is�k^tG��,�g���Ʊ�c�Ά͌��(�wYM�״���W�W�)(��r/%i��mFUy���{�\����p��,T|��*�[��#�t�i���</-��%j�|��^/+�^*��_@^�tB���$$}�e��:'w��ѭ��Lsg��{�n�i��?~�d=c�T����>RO�,!?l�\���J�g��o��&���.F���kvV/8�h���3qy��衾���z��g��E�3%\al�d�rQ,Ė$���>jڵ���>����c=H�jR5_o����ki���]`v����6s5SE`z��_Q�Z��䡻;��x@�/�u$���h����@�N��,f��._����[m��N����M�\ṽ�o+��8D��"H�(��9Ϻph�5�At}mF�c���(�A���"c�yY~�u�iH/�f��p�����체��۹PU�Jeqy�Tf@e��K���~/���@E`Х�u-��	ő�� 0����;e�d<�����a�7�`��4㈇K5�Z��(ԇ���
�عw�x����dPS&.��?�2����� ����5濕v����P�PQ�t�E��<�Wز���|$ɮ��x�}�^$/�{�_�fp#�(zh�֭��d�d�iT��K0/��{o?��
�b0wP��Ɔ�%*�[v����x��94EF�[�!ڏÈ�Q������>Έv���%��	���%�֌�d��0�̳�gU��jO\�!������OW�ƂI#��~�I�ֈ'цɎ�\��9ٸ�J�����Ȑ�+�$;[Yvza�1b��}n�ީVOX�z]������y����e)�z:sD$�}��>�4���R�� ۴�+��ʵ��i�5����tg���:S����]�/�l���í��#����\�"�E��_�H�7��+�]�tU�]WJ��xx�����ot�<�������
��������T��S��|��?�Ҟ���.⟌������0.�8|T�]��.�)z�����O\-�~����d؆ߏ�������i�i�NL)Z���l��dce���x�sը1�r��3�=h+��@�i���M�v/�s -����"g��Qh �Fi�x1q�dt"�� Ǻ�XW6�
@���D�[/IZvx�1��,�Ҹ�ڠ9H�ζu� }�F���"�%l!��
�, ����Y�T�Fb$\�
xK�ܥ~��&�x@-��!�1�5r�?jQ�9���f٭���UQ(�s�uL�.y}���p�|0R:N�P��C::�:�g��������Уr0�b�=��	�/S0ŧg�5y��TQ)�Q&&�l��~VR�£�*�8��G����wv���qhZ�R6z���Ъ�j&�M�|������d�4��Бe������D�I���'�M���`"W�LŔ�K�I�4!��a㍞N���W/�@-e�!m��2�zh�w,��[,�B��ӼP:���c�A4�	����Ll-�Ft��i�,��?��挸�R�[�̩Sm�þ���iM��g+��{��86��W�WYu='�T�r9"GT��;N�;p���"�;V�O7غ`a�K�[>-:{mj�h�y���Ϭ�[���pe�~�b�%�?{�!'��l_{��,%�t+�����%�k2�
'!8�:ȺY��~��`�tB������e?��)�&Z@I�Gk��!��iUΕ�����73v|+��8G��|w�.�Y�S�q朙Ol���M�>���Sۤ�g�%��j�jn#c��9��b��'A�䊇&/k�e��&E�3�#C�q

�\���[՝�nE�:	-Χ��E2z��-O�O�����u�.Q���/*l�Q�i)� �z�9e^{���L���=��r5� �6B��F&N�j^�C�Jg���8Ρ}=��ɫ۪�,}Oc��Es�r�3�>��r�sؔ:����S�,}g�W��7���:o�ū��S���8�9�i�p�XǔȞ��O���o%e�Z������x���8f��e3�},��
��P�k#�:��f�K�>���>���Y,�仕��vOe^��8,�>�>�nK�'J�
��ج�
��o8���� +����d�C�������?���9�Z?�)�c�퐬���w�l� ��%������A3�͌�ӆ�d�̄E���Ű6�|q����[���:���"�A�,Z�Oa0S�`S�aҫ�$��}= �U�ee�iyh1��4��&;��uۚ�]Pu���Wj�v��:�<uWF�uP��n�H��ˡ�H��т��P�t�(˂"�g�����W��I�Յ5���_j[��@eg�X�l?�8ZU��E8M�T�u��My�>���� ��>�j�N ��i��߰��!h^1B��:��TB���e�8��"�m������O������K���<y]��Oo�GFUFj�7v��t���A��5kd)����`/�w�
)�A�^|��H���5�j#��Q��O����)�nhg��x���"�借�Tm>z,�+�W}�OyF�y����ΈvW��d���	@v�(����$I����K#�cՕ�!./Jx�Zs�@`�猌������s3�0��[V�T��b>�ߢ�ю8��흻{ �X�r,ߵ7���b�_;	,>��Osv������[��yY��9Ǹ��M�ѭ+2NX 79��L�d�+_I̽�)x	s����&�
�EF'���-�7�-�7�F�>X{����/:wUNg�m<���+�y�:����[���B�KM&����Ƥ"��:mя�jx��5�Q��wu�{�|_8��A�������m�������:N�g��KfS$���E����R~f���P��1����Ӻ�5���Hd��&9W^zv)z�Eqb6�PZQ�����v'�C"�E!��RCh+�^4���-�:��q���T��.G�����	�	��9���JI!ї�"�5A����Wne�#���v��/mͭ=���*�d�J��Hk�s�-����EbI%:�q�HŨ���5˫�+S+�A/4�> 
�?*F�N�i�˺�����
6�D8_:<����a�(�G>&"9	��a��Y��� �K��0B+��%3�
?�z�PQ!~���۽Mb@`�H��e$��l<�mc2>JH��9����֪�������5��a�_�8�#�4l��"�X.kiC����`�����ys]l��kw�}:��h�����|%��
�FZ�A��pa-ѝ�]��{�Hڛ��<(�Wc�����5P@ߡ��^����̃�c��|�HO�qp|��W�����ʬ*r�T�q�W�9�Xa��o�l� ��E�%!ak��h�}�2��i�1� |�D!�OYC[�Ӑ���ǥ)�`��RG��i�Sv^��%3$�ݬ+��sΩX�G�~�"�oR�i�L�:���G�r��e×r�l�6�'���H��.����&"̀�P�!ū��9�o�Y�ܲb�G�U�k7:�v��3��r GEu]�F��ŀ)e���Q�3���6@�A>�~�IC�(��#������I���lL ���US/��\��:y�F�
����.S6F� Iыߓ����E�SP�u���7��S?�f� �28g�@S|�z�%69�X��*�����_͖�7�J��B��qz?�k�owq��D��[R�
�Q��H��Alwz��0�b����,̓Z�6Z�q,�ǿy�oq�ֶy'yNq'p܂5���N��9���멏>ظ=4��=d�l���l���.MrTY�ia2T�)>�;S�{�����w�_ea�yb�`\j�a<wD5���V�K��ƾ������!�J;�O()i5�dJ�\N�F �x"�ސX���Ŋ�%���m�X��Ml�D�f�x��nF�yM��RS�ǿq������)��ESz�P\�R��y�r�v�|7�K:��8�㸚�i^�)�vD�w/���u9u[�$����qkktkԍ���H�)�����;.�2�x���B.����84��j�8�#�ڏ�`���Hd}s��F���PE6`��գzJ����཭�}�/��:��鈧U3B*�]�b�_�d����{v��	��Y������]�&��	Bg݃ڪZ������*��n�����,1���:�����=�j��������P��T���S��c�e�����!#J,��Z�n4�=h�%����0��-�M�����0���!�����
�u���Ag��V�>SpW3�x�{fz.<J�����io��"_P9(K_���/7v���'V�rQYW	x:�^��5)1#3�Ģ�R��y��hp����0#C�\�3�D�B�_Om���%FS���Y�l��"���g�SVJk�u���ߧ����T-��<�7��'
9<I���>��X��j�@��Xh!�̽P�tؖ�!������;�f@Ǌm+�&��C�M$6f�1]��e��y��DIIh�A^���SV����,���m(�ݨ�U��h>�^�����\�=��a�X�F-+��[���KFv�cU2ם��xt:y|B�2�x�|��s���6��� C�pQ��abQ�����_�%Q�6*Jć
���d%G���U�qR���_�K����L%<�#j�m*KYj�W���t�x���@���?vI 	Wؘ��G��ݸy�Nq�������Q�x�;,�Y-Y�hE$�i;�OL�B�<=a���_ ��t$�Ƹ��حh�×����;�%bi�z��`ѽ۾W�d����5zx�"�V��X�}���e�ta��%��#��c��lnOrvPL:Rk#�u^Z�C����7E��{t�^y�V�EH�ף�����u�;.�{��٢'~-�q�ҏ@g���t�N_pg
�#��29xk09?�4|��[$ŕ���4��X�lɸ���\�˒������;��yu��r7�t��t;%u��w�|�Yzwx`�;˼㻎���1ɬ9��X��U�Np�+��nf>���ư
��|17ų�����cg��ᙟ.�����H��u����%�k�Ҫ=�h���$&
q�W����9�a1�X�4�=%���s���u�&=Y���8K��)T��wFL�6L%�4Zvn�+(�j{ ���g"�8%%��������0�"]j�{�H��DYh������{�N�"{ �׼OQ%�T}9P������A&xȽ���g_�!�K'�9;�h$����I�mh�����-�	�I�$T�E!�Ehrb������k���NR�c�/Q�=���)������FG�ڨHi�^��u�մ�f`����t⛈oP��]r�^��d��I�/�3c!"yª�m�_Q5�Ȅ� n������ܛ~����?07���щ:(��}�뎉f"�����r�1����2�9%ќ�r�#�����9��f�	�mF|��vn5�l�����((4��t���s���r𒛸���Ǯ[+A��hڷ�{'���/l$ް��ǭ5lW��|����D�pN�۞]{,�&keZ"�����z���x��E���@�eϮ�3^Tn#g��%���]�F�	�<�ᶦ�N�F]�r`�O[���^����d�-y�T\h�Cw��몳��HRF�w������ˉ�Cs	�Q>
}�y��p�`����G��7��@d�۠L��OE��u����3�b�.4D(ָ�����</�N�m����Wֳؿ�Ďe|��-i�l�*<r�^,�uir"��sr;]?�H��I(n��I���7"2�9�������ӈ��;˕����Y{'G��~�2���|r�B���'I���M]��AZ�L���6�(�M�e�xXG�m��4���2Ј'Buj������K�Bg?o�����c��~�C��)�]�7woh���ǶW	Qtlޗk�ˢ�\N�������^�{��Т��#��`�;�q��İ�|W������3O��ʧ�uU�8�t��*�?s=
���U���$)���3B�t�����z��;~W�IH��9�����cҮ����pISڊ���Q�N�^N҈����y#/dE���(�6���s:Dmzb���.���n�U,	��?����~�LLqh>֑��1����O3eGM����i�������Y�^�y�26o��7i�!(��XѬ��]�0�Q��϶����6!o����
�,3�1&���8Y>���IR����t��|�h^���h����g[����c���P���m%�K���
؜�T�-�J��l��6<<�_r�	�l�/2΁��������'��-��z�:w����DǕ־�;ZL)�g�d�L'ܛ��R\�|���ȇ�Ÿ��Wɘ�������v3���t:K�ܝ�m1��D��Dg��6qOWZ�*,�h�Qˉ���c k�(;`�t�.�}%Ry$]tu�r�P��(��	�d28m�-�ǅ_��O]8zv��m�fe�� 4*�<�T�}��s��Z�nk�-���ERf�X�4^����Oؓ�q_�D�ù���ƥ��ݥ�������;,�8v�/I���0�{�s�W|���iwӂ���w��l	����b��mB�������a��e�����Ew˵����-�݉v����n��/u���;���'�V�4x�Ja�����6t2�1�����[��U;܎��I�Ү�/:�o4U��\v��gP'!���Xok�o����ɨ��n��߰7h�Ԕ��7!������������l2��<rp��.椰�q��.��0����Zno0Ԑ��d�1HmA������s�9�Y|����$�V�g��[��^���)0��{cX�d�LCW&���O���],��3�	gֻ��ҷ��܇��������Ƶ�s��bd��Q�{
���x�v�ӛ�BZ@�KO;;X�H�0��~���B7d�#����ĢBC����ОT����hO���o���U�W� �_�����r�fQ��G�e�|0�o�[�/.'Lq5�����4�D^R�D�ǖ��k�I�Jk)���$�`qL�e��4.������#�O�$��9���\��n��k�uBMк��=F S'R�,���/6gg����x�J�m�>Le�V���!�1Ù.B�e��1�|�J�iFޗux 1���Z�ᛪ��^l���\�F����Br��iaf�}#w�G���D��SN��C���u:�zr�����mO&�.:�8>�|��F�{�4���_}g�t~�����!�)Wf�w<�:��٧��M�w���]�ë0i�;w��ʐ��R�M��*����k��e-�xڎ��2��BߌSs砷[�{���a�zJ\�<��L-k�C��~�ih+�H�HǮΨo	�&�J�E&u�0
��f�Xp��1'��ƋGl�_�@��b8ڄ��m?5�cx~���<SD�@<��%��Up��p�IER��W
$�x�E����{z���H�d���J�{��~�������D��hb5��C�Gw<���X���ؽ7��d`9-��ШH2�gU^�f���^�6��++��x����K�?�����֌~N��9�]��"3!联�b�JD��j��0�9[!ʊg�P(���{*�� ���T�{��X��;Mf�~�����_�fz_�4N�q���S�=�1~��+$}^��D�i�pʼ����:S1h�u�+� �s�S��M��&�F`th�,��׺++6���ۗNo1>�;����| Z4d�2sQ�4mV�*m^�`�J ��0����;zF���f��-o���8�#/Nw�؋ڱ ��-F�Y_��(�J�:�ԓ�{\匭�xnѻ����N�b2��3-o��PwF�7S~W��wXኻ�Q���y)l��e�_�ϕ=��IR�9��f���Y&v�{�<*����{K7;���L�;��6���1���"n�Zn;��~ث̻�һ�w���3�������񥻫%��y�ḛߝѸ��m���^��<��z����o�䅳w��eg��N��&o�������b���q����u���h�ݣ	��fm�1�����f�Ȅc���&D[��f��~o�g��qϖ{�3�:��B����m%��16z�6�������N�N_NB����b"J5b�4EV=FQ�w�Mw�8��T�mdr''`��"���u� ���Uq��E��8�nޡ�9ٹ|	}�Io��HLM��ӠRQm�2}o�(~��G����xu�$��C��Ⱦȋ?�KI�e �Ə9b��FG���tס��߈:�рF1E�O�l��1.g˻�<أ�%�����s���峉�����k+��+oV�A$����0�:��g�v%�����M���?��
M����	���:�ihR��!C�hٌ��Q;D���r�z`K�!� ��
�B9K� 3~���?��jA?�	0O�Ap��+�am|���ͣ���n#z;X�E�h��.���`qBu��^�g�Tt���ɛ��հ0���aG��ܟ�66H��5w�'��2��2Ӕ(-([�z8�z�s!��t���O14�<��*�G��j5D�Y����|�>�D����otü�sn}������x��6����Z:�Z9 ��N��9.�1?R�U�M�����;���ႏ�,=o�e,lO̼f"g�O��赆 Yʹzj�y4�vr�_w@���˫�VH@}��=���4���==Wq�A���5���ckn�t��VH�(�8�ٹMaW�N�/<�l)y���`5x����^#����u��#I:�h�B"sX��c.=J	9L8��e,r�[��dJ��jQDm+Z́PC���;* i���� �i}�>T�Նt�i�@_��yY���ɍ)�}�˂ژ���( FZ�V
���z�@�޹UH22*)�"�޺������ָ��#�Cvc�?o4��:*�Y-���6����whb���ч�����,�S �?BOvw��~�tT�.�OF�dڭ�����JI#�H��U�y�((��#�-�5�Z�*0�$ECԽ��b��X�H�V3�Ty�.;ơ(h%�e#Yy�8�]�c��h���G���l$���Ι�t�I�3ڄ��.�"0Af���uZF�0G�)��z���`��q}'�H�1�:ͺ��˱�8exE�GF��`����X�1����&)�إ��?м3�c�=�4���y��Ws~�#��{�� ;�/W2� �}I���V����ZX!� ��h*�`XSmR0�e��?(����a2��&��IV���0�b�K�?|�@2V�P��U�,ɉ `���^B����'��v�T�؋�)I?��B��'*�%���ج $�6.u:9Nt.v��/.�<U�)A�\�үۿ�dY^  D��c��$����J鳹S�#QÊd��=*����S%���B���ϯ>�k7�
fZ�`�P���~�q��p��rsxZ&1��ׁ�|t�}�G>�Y�ʣ%$�qN9���c�ra�v��d
��5;��;�<�)q�_�m����d�8̽䕏��6� ��#��X/l�kn�:���Cܵ�����GhÎw7��Q�o/�DK����d[:���Q�A�_ ��=C;D����<M ��i;�'�˾[Oj}j�}�u#�۹�`�J*��MA^���gQf��@�BU�����=Q��W���l�b�|=j],������^Z���4:����Rq�!)B���TLK�����'K���V)g������{��Ǚ���h��Y�'���ߓ�f�$�]�c�(������t�Rt��C��ü$�>5��HH��_�3��;�f�+�Sf��ʉ�dG[�Ǝ���\��.@J�]��e�%����5)�d,z$�}_g[���E Ԭ�
L���GIn�$�pg�Fm�]�'&m�$m��
�e��!@�%�Ή�,Ad��Ǌ��V��[��'^S~����?�_W���ֻ��v0�����_}R��O������ �t��Dmh�ע�"P�=Pkr�`��5��m��Γ<��ee(�����t`�ɠ>MT�&[m�a�oh7���VEc~ݭ�v�@mTublW�=�(��d��!���9�%�AL$=,f�?�Q,~)6�@�*B3Ub��N�����7ن�j��4�Y�x�"/L�ǹ�<V��7�L�6F>��۲.���+}����ա1��
�w|���f�s$���������^b�7�ͱw��ۀ�p�!�"rJ�H&e��`>��ү���Z�#d�ڿXqP�,V�W�	�b�j�V44�~��ܛH�
 �̍�o���F���>�5�I��7��f�vⱚ+ф��F���	[��N�;J�~DZ,ch�4��;a�X���.��A/���� ��	��`��Hm�@�_���J/�C�pV�v��g�a�U�����J�#x�Ñ@H��� �?�ڥ��[P�-�S���BE����>٪Y�� �8��""7at�E7B�V���	-��wx�GxP_W�W���4	��D8�c�%Py�J���b�I"�R�F��2���SۇJ~X��/1����Mz�l?Mc0�Q�L� sR�!/-�^�����N�/c*��t��Ȥ�Y���Ϧ�Ŗ��o^�*5/F��ostaG�y���aq1؊����pt]���ⶥ�����--�����ya2��>����#Ds=�`r��~���!�綢�
X*B�i�������;��A��5�\L@e����t�{;�!��SA (��`�vWZx�c��JC�lW��zr�p/�eQw��礫OUm��㩇�Q�
���^v1����vJJH�O�-�\���U�����#(�:,_��2�gGƐ,e�?*G'$lϩ�~���&� d�Tr�Dj��-�;EM*�+��r�s���J��.q?���>�D��Z����Y]@�Mw�^�S^���`F�}]�����f�3�/d��w�V�Ȕ�&(���VʜK�^��HJ�&U�e|���}.s�B�*��:�ل�7�E�^,�n�=��g��ms�ؒ�#-MOQ��`�p���`[�8-����R1��ۼ�[�o�ĴV�KQ�Y�%z�˶1���n":m'�1�3�"��$2x�A �˚���G�uN��j���*��o�� YWd�A�E�oY�]:.����j��;�1�0c���#�O؁�?�=E[B�A.`}h��3��'��g=�y4���
jR	���"���wh@�3@�'�i���<օ�^⩫dS[L��G=��'��*�@dy���/KY�����3WĹ�?׍�l��,�v�S���5���^>ULl�$�A�A�P�"�`�f��L%��!S�j�7��kC����xX�4t<���)u�����6�S�T��<*�F��VƦ�g&c�E�
��,hn�m������2G����#7���(ū�F8ܨ������cL�3FYu^!A�8#� �4g#Q�L���Pw������?�8��F��i�u����[=�lϪ�*�w�9����CD� � a��7�Q��ٽo�e�VoO9b�Y
���<��6T�b)D�xg���W֫�<+)����y�ꯨ��H=��M�/`�xR������[�	5&�O���&ШXU2�(�g>�G9�dڳ�e�`<����/��5��б�B���"��=�bh:_�*�4�&�����]e�nT���Q.�D��*�BߩeS�hGG����hxhA�^��9�J���&�K<��cC\9l�Z��W༶k���մܞ�
gJ^ެ�������s�6�'�J�f^^����g^�w��l�`2�A��4JV� �^fT�Fua�%T2mC'���EcȤT��p�p�%��A(���B�ј
q�~L|��f�T�����l��'�{W�PO�O����"�f��ٱ��*	Uh��<�x2�9��vJ�S)�ߺOE�������-��Ź��!7!u��3u)'uۘ�ޓ���ۣ��ح�ў��[3�=�Y�f�))t����s�6��$W�8�'-�~��8�y�䇓_��ύTL?r3��� V�~�
\[fa����U�y����^�(9fb�_������!P�_#]Z-�H�o2�A���+|�!�$��) �8���*�6�b��T"<�y��Zi�	e�#�3��!T,6H��5d��2��HK�I�����Y����98���p��ߘ-�3���Ez*�7L-��,�&H� ���d��m�SX6:�YK�b��HT(�����τm
\��ݷ=��}���#��X���e���qn�0փdƓ<v������j�{e�\���f��4�1?$���[1��ɠƸ�Nk>�^7fْ��_T�`^�`͒���RT�2�ب�ҹ�w�W-�44(zc:�~���3���^(䪶���� r��
�c�@�oH�B�_Gڱ�2�U�;��$�N���=�{I!��+3������	IpZ�qE|��,�{;�p�Ý��}*j�,a���?�5Ze����T:��s�ʂ˒qО�$f!RH* ��%���Hi+9�4q��V���XX�R��ސ@��w8����}�i��r�B+"��/�x���p/q����Tv�X�(��;β"��Y>i�%j��j���κ��&�jw>�tM�SO���D��)�҂B������~˺%�����~��F+e_���{^n_������*�eY��s^C	�*�����i�����j�g9q��##g�?UY�\��7��T��M��_�E��T��� �SMDj䬶˿�`P5NP����ay�6��^���Z�����3����Ty�_��
�Xܠ��:Չ�����Y��-��Vy��*�i��uS�R���&�%	σ���0�^�=H9a)�_�<�Y�H����������`o8���lU��&c!����h"
m)����Â�_�Ma�P���!h� ���a2�@��ˏ���C	K�坜��@��I�>�9ߩ�#�z���̼���؆
�XH��@xJgR׾��jR,�z�@X��@���\�b�Ks�v������ز7�<�7�+��Λ�1��6��6��� �g2F?˓3����?mk��rw�'3��vg�����8N?4ݗ�j@7P�mS_l�[�o��p:�kĔ�0yc>.Αhs��j��I�ɞx��i�ú]�)�t�����&��R֌��.�x69)��Mϊ[�&#�̒��}.��?�Չ�d���j�f���c���t�-�a�3*�~lHX�Z�br*�o�3��A��&?�ehG��%ɿE>���	NZs�A��N�!a}]��]�?p�\������c5����x�>At�Q%���I����%�X�� ��X�H#s��?ի�:r���D�ab�sY0��ox��D>�᳖��p���@ik�#A	��'w9Q�g-jÝ"�S-@r�@'��_Z2r����ws�!L��2�@�����Rv�o�iʁ�#$������x�6'SW�_�:���ʕ��ɮ&�."�r��g�ҧq�1`ܟ`�3����'��ݻQTX�A�muCZ��l��F#���J�b�_��*!�_g�I�}���VluXI3���؍��0��oĮ��
���N��|�!O?���1~�l#�kܯ�Е����pю���%蓤����JGvٜ��$����V����nDيP��1�Ah۶�A����+���ߢD��\TQ�9����@���S�b���=�h�" m	�s���:�{5g☊m��ѧ�P�+��DTk܅蹴�����U׹��:Zj.�n&}�􄏚ZK�8�WX۔���^��s�t��_}��	�UA��Y��h �Nd@9�ixt��U
�Ka$�e������j���	$F}醍�����)��H���r0���!�[�S%Do���s����Z����}]����z�޻��M�`�j+���;b3C�8��<�%��?�1��&:�L���ǳq7�r��)XY�<X��7�xR�2���;CX@Jj��SD.?WEf&�C���9C��[�ߡ�I���i�����Ԝ����;>I���|��<�h���֠�!2�1=�$~KUXeoE ��z_����6�-_�nN��u��*��~�{j�r�Z��ok!��v~:ޤP#��FXw�@y�ꇰ���5Y�D=j[��߼9 �e^�R̻b��@��ߪ[
j�����֟	1���k���s�l���P@�Au�;�w�U�⁡��qϿ��<�������$�����#�k_^
b,�^�D���.-�mO��p��P�5}?\��_���	R`(9�S�u�8&�QF�<ѽXt��Z0c��}����h.`�����̟ݢ���/6ܶN�)/���/��p~0��ME�|5w�S��#��O�VEQ^\��^h��J�<��=���X�޹��M��7/,��U���%gc�}ڤ�X�s�$��T��\4&�u�}�r︿QD���{��3OE��b��,��&O'(͘����^?�����lc������[�G؏Mb�\�7�4�~�el�!HO4���E򞁒�iH�I5�g�f"��y`Kf���Hϙ3�00[�KMR+^�2*.Y�U
S�i��Qk��3�[иꬸ�"�Fjd���N��)���X���o	Qzs�Rk������@����i�S�&�5	���G��D�lqk�kІ =�����~x��?3m��F��Ͻ?��[�� �է�n$�0�)�����\�Y���VtOn���sSH���������)�7��g��V�凉�7zq������uB�ǌ�S�Q��8CNi�ȍ�%T�\���j�?T�k�q{��.���<���� ��W1�dDr8s:��$�p��ڍF8��QJ��K��LF���������#@;7x�T'���w�_��5*]^ha �s|�O_�3�/z���j?��P�U������d��~R~~}�8pr���g��n�����`@��
�kxT	������8@߈�_G 靴8��ɷ�>�U�w�Y���\�.�z�o����v
�䢅�H�j��<������sN k��M�噉���U��3��1Pf���y_&�\����ZN<�4��x��`__8�3M3�C�w�rP�b����A#�2����U�#C�\�<.�Q����)p�3\P{'0g��.��M��K�
��B�V�z������@"r�-A}�}�O�����궀�������C�����X�������r�g�a�f��l��tF5$��k���F��v�O��}�E�?-��8 OGN�X����������/���=�^Jq�Pw��o���^�ү���Lt��?��Xړ��'�<�^��k䧍7=M�h�,/�������T4 [���gH��/gX�:?�&���Z� ��')�k���H��Gʩ~A�Sxw�Q��#����<�m�Ͽ!��F�<�4����f�KiΥ��Ŵ�K-�n|O��e&gy���{�m!MG�����h+2 �J7�MqQ��S�/�s��r{*�Q:K�Ƙ~���S|�VJ���,��*�c`�`�@����Mt�w�	�%�U�]1Vrھ��۲H�Ĥ��/��ң�����.���r�JV�J�F��ަֲ5�<���+v��y[3��c-���>����������cosۛ.w~[wA���y�@^Ѽ�X��P��\��FcG�*^G�M��p����Q&^���M�+e�m�	�?A�Q9RL��3щWЅ�o�J系�T����9�]�8��x���[�����D�|ҟ��pz8�m��|E9+�R�:*�:��n�f�<ʦ�egqB��nOg�z�*1�}%?��@� Ұ�q���w.2� KI�Gڃ����@�)`L� �� �=	6�6����.��C;��:��B��$���&[Syծ(4�k�F��.�;޷�W�RI~c�#���w�"q���ǁ�����	�\�+�v�F4������J3�8����OVj���	�G�k=[z��Х-Qq��~;/ύ	AT��(���V��[q���'��_��npe���?���)�j��#�^���;����R�t�$��BE�5懻���~2w�vO�ܒ������x�K����$����:��<��5�GwN	
����9j�C�xz����/>��g�HO(#�!��F���'��RَS��0	B7�t�KBdJ�R{D��1����ur�}!�D��V��������u��$h���cy��q�ߍTS�Ҍ�{E��fRp�	�/�W��e�ͽ-edp���.N�D��"G�w�h<78��P���>z�ϝ�N�����x�y.��Ą
�chK��u�n kX�{��Vl��=XJ�d�qiϦ����Пz�?��Ӥb8^ypf��(P�قS6�XN'aON% N):2��F��2`�c���4�X橣0n,��Y}i2Z����Z%�L���}@v��є	w<I�F�Ӧ��̬0�H~F �@� 3���E���C�(z�՛e	X��=����0��ΪNg�\?���R_��\,j)�h|�+���4x���;�@���:��Z�X�q�F�#�� �zZ�B$<$n�t��	��|�! �<�T�iq�1u���}8����~Ebň��ÀGQ����{���g߅�CA�*llu���چ���󾦾`(�Y
w�J!&X�ڑ��4B��*��+�*�B
?����ц�zd�FM{��_��:�
 E����4��^TO�1�'%mDvH� Q�Ң�&�)U��p�ww�䅧��ڰ�pc6��?(?Dv��("��I����I��{�u�@𯉱G����e��zz|I}��*aޑ\[ �.%�Fl����6}���^Xi:9��{�L���Xې���/���΀���N�C4�]��*��X�z_K+�z��p�2C oD-V�1>�R��Eh�k�.�z4Y���ly0��;Je��]���wH�R�!��%�.1�dm�!t���,�l���(:Hw�f��٤��j\���]��N/�����,L��Ư�U�QU?�NV�O,i@#^R�<?���e��ښ	s����-��_���BK��n�0�Ů�M��[��QBB��-��ij�����|q7���(��$���^�����x�n�Ēm�K�D��/���ƺx�����!1�7X�Nl�w��⇯����	�� �}ZRT[�K�s��=L�w�C/M*s��\v�>CY����Ф�<'���<ׄO��4������u��Q�^�|���sv����(����� � K�{�BJ�9���ed(��ۘ�7�z����C��R��N���M'�z<�x\'V`\Y`b`m)/�I�$�lھ��om� $�G<�3��@�-�Ɲ7�%]�%4��s._��I�
ywڄ��EݝH�e���x#��2��swf��/F�*]�"�h=4�?���^�?B�d`vs��ƴ��}�d�/�g8{x"��� �c<���LB�Cg���E�����m�[W�͚�Z��
�
Z�q��$�A���E���0O��8!�K�s4J�(#tcs���x�\J@*���P�|��_��D��d��_q���J��ݸ��w՗'
�٤�U�g�;������[������ �͵��]�.w	�A+�VB#tL/ql�id��'yk#]� ��T�Cp(L�1��u4����p�+�H|���� ��M���h�{BEDf��*IG޾}VyO�Q��ϫ�S��X>�?��Jq�i��^�G�MC�<��JN*�/0���b�fǷ��v��:I�����5u�C�ݷ�z�i�e��&��:�DS��P�HQ���,���_{mH�n"e����G�~"���,�%�0���NGd��>��D��jY3� ��֏�����-N�L��+u@QN2��!?jj�����cᱺ�xm��@^��_dk\�R�sx���A5f�|d�`İ�~�U@�D]#,�ͽRO�\�I���������O�}^�P�#� o�CW̃!����(�"��k��ٹ�<Rs�� � �f��H�TmT���ۄ6��x������E+�9]���7Y����Ɗ%32`v8�"@�)iY������&�r���h�:��J������!��jkx��?I�枋����ιQ۟4��jb�t���L��ޞ�̦<��9[�y5�z}6=�Y��N+��'�,M�SS�*h��yR���NEbv�!k��a�m�b�6m�����S8i�ʫ7�o��W����J��ce�C�b,�����΋X���,V�ˠ ����>.�H�� D�TJ�ۆ���Y�n�N�L�������}4`c��^w ݇���%��OM"歬����;�6sӳ��};��9�V*���k�k:G�2p���-������^������m��ѳ^��=��i�,�+���؟ަ��M&�����	Y����Ȕ�������]am	۟�g�L�4���E٥tO��2Nwj����R�2�6���8%���j^�*�f�7/�{Ejm���MW�^\L]6��%i�O���"�L4��V&8�mXpn��/ʚE �>#�CҨ~z��o���}�fb���>|���H׊���.�����J"���4{��K���ϝSC�lq��/ ��L�SQލ�9Ά:-��h��ZN��������٧C�� <J�c����~�Ͽ�y�k������/�UMKDJ~!)�$p ��e@v=F�5S�J��'��k���[s�sd�
e��% y&��,,���	,̉̌�YSwIX���,R�8/7�6a�%�(4W��o�RH�RXmzI�*�\��!7N�ۥ{��eE����هO�}�Q`�.g���ڏ�h��� A M!ċ��T����E�� �kA�g{Z0�Q����=��\+:�q�9P�?�%�����ҷ�!�(�o�x�9���2����
���fz�k�
�ň8Q�]�:`&�wG���.���ݻ�M��-�� ��ڀ�",/��n��z��M��t�x�bEq������"��vϺ�|�q5���hϮ�i���e_�Z���A���C�	E��gƀ	D�I���Acb�d����Bdb��l�9���6�Y��W	������47���~0�f����\�<�� pyq�-h�HIb�ZF$g����<_�5 �d��L���c��Vi��<B��þ{�����L�=J�"�"¸�`�QcJ`-[�'4�:O`mbk��FD������� ��,������	2#�d�H��ݚ�:O0�%դvw�̚�N�'0Ś��Y�y��!�(��&J��/�SSdF�uc��x$�]y�h�S�N���~�s�)a?��a+��.��C��WI{jG;��Z|�d��_Cq�;�ҋ;�2s45c?�R(}EW��S��06��U�~�S�W�Y��Y��h�����FFVV��� ���iff��P��)�OR��좉;7��c�^�V��7��
"/��k�h�rO	�;��"!�*U*�Y��d�)a�&��(�Q�����r{k2.}�sݙ�JxE��?:��5����j�-�E.D��1�|��~�^�O�P��R��?/C��of6C�d�O�7���J�Xd^O�>�tPWX{���APF���jU��b%�jń���Pe��y���b-N;d���[E�N��ޕ�	��S�*7��˻�Y:���#�_sA�5��or��sA8p�nQ����a�W�͐����P��2G��~΄4
�*i�v�X�����xb������~}�5@TU�c�gP����M��U��Y�!��a+�e_��������UI\�p�؃½��M�(IE�=*���T�W��3����,��C�­P�.}'������7�ʴ���m�x����Z:A�*ݐ��)PC�2v���hdu���S������s|����6��%ɩh��;x!M�U�=*����C���vJ�L-�ل{q;i���a���_����� O��{&��Ÿ���*�����Nz�@N�����.�㒒�{/��rz f�yXjX[X��|��������* ���cPS�U��5���"�ę`m�U���*��jA�&̡�
GA? x��t��
��z3�	�Ϋq��d���~���r�]ޭ�ߋ�≽O�K1����w�U_8`������=��x�͖��-��3����_A�h�VIV�-��M�bR��+�����=���N�h��|q�7E�����jX�b{�ɪ�����۝s�s� ��ɶ�u�~�&&�"��ɂ�H@RճX�C���&��5@�Fq~9R���*�*���<�U�?�8�s��W�L{Z&��-�'�p�}s���SēSL�>
���C���QaHϝL�Yu�����̀������k����;�r:n�Bs�a�H��Յ?�q�&����5���^�����}����K���]<���#�<_Q�}c�zQO4��r5H���֒�ji)=u�'ac癟sD�u����cwM�?�/ϫr{g�"�b)z�)SF"=�K��AR:���1|@��tM�������%Ͻ���vˊ��#*���f�B6&K?b�>�o�Ql]��Ŀ��2*�����S�-+��%z�k���(�/�h��]d��AFoeG���P�(��'yM�Aaѩqe.���o������"!B��r��)�シ��v�S�����>�N��$d�j�m.��O�9M����T�X�=W����o�4S�v+Z3:�i����C[8�o�3!�6*�>o���PV�`������o�_�:���2�'ijR��?ςC���!�+!����������S��A�  ������dը��)V6�m�Vߐ	�48'�k���V�)Tԙ�/R_�����Ex��j�S���ڰx�>��9�8���7fU�I\�g��{��_�?����Б�X'x��&v��)�J5��{<��7?�z���?-:,�ߦ�t��^��K���_"������Q��:wb�ꪰ�7��8�����3V��u����Ա����'�Nw���c���p�a��a�n1/��M�%��o*Bm�"�3}{���@8��Z$�"�xZ��r�JI2y˵����u���z�|U�e ����e�l�dFL� �4�/�.!����nM-T�Dw�B���;*�s�L�]�%W��|sF����zI_���y�
>��]&��O4�g�>��:�|��/��l��v�so7�~�2�II��8c6{�/��Y�K���C��[����͚,��Ά�n9JTp23Y��XͶ7u��8ݹ��Ɨ�}����;���J{�
ʘ��Ct���Yy*��z����__}��v��1v:��o����v��)O�;bn�Ⱦs��:��N�j�GTgtH�ru�XY��R�Ʈ���}����U���D[��xuIUC���Z߲��ef����Jf�L��aB!Vc�,-@�11h,�K$n�v�ċ�4R�z��N b19�M�x�g��U��j�:35R�D�鐽�q2,8y�K��7Y�C	�~� S���U�^T!����:9P�Q�w��r\$���Af�nzi���B	�:
yJ�d�H���hߟ�M4ް#,�DNV#�������v֞���o�1��h5���ג�۴�I�(b��-�gA�5�ք����^v�)ѥ�9�--f;��=n�A������aU���<x����"ۀ+�Rj�[��`V��\<�E�#8\�:��d�� nrJ��>nձ�6}Z`hݠ���Ԓ��=�w�ok��^��I?<�>m�<�������z�T��p�k���!X��'�箯�W1��y�w����`=��j9�O�ݾ����W��P��)ϴ�t���5�������񋅁�\/]��������?��ݷ`�!o�z=]�O���5m�,R�!����3����+����$�nl�o�ܨ���Nؽ��*>�X7 �o����BH�*�{�ɨ��N��w�a�{34�>�|�l˛Xd�,8�y�
a����!�p���!�@DiZ�G��I;c�j���E�H�� R��5�\���n-����3;�Mr�Nߢ��&����!��C!����Y���x�c�gdE�.�M��.��d�F��ښ�aw�]󏜩���$��K_���T��BH8^�G�*"���ӌ3��7�����{��2[x�M��k���Xv&�ٟ�d�e�S�u;ұ�Mr�7��I/�P��I�I���y���sX̬KfV\U�xb�����`/g��jޠ�IG�j�����-���}ja�� ��A������#�����y�A\μD�9{��GJ�yB��z�M��k "j�DL�T)����B_e�����U-����#W��%wK�_�V�erG�����TfD��HKlF������`�V�:�Z���=E9����	��6y�
�dZZ����U[{u}���v;�YS ������[��j˩s�|/0Og�B�i �X�Z>Am�^
A���߯%��^vt����(蔻D|�E8�~���*�Q�:� �Nn�X*Q%,2��I��m;$�d���{	Y&�́��z�3l�k7�>�da��ң��
�I���m���7f%~�|RN>V�\�C9�V�\�?���ߜ&�!u'��-���7�G�L-���_+���ޡ�U�2�ȶ:U+�/�4-���)S��S��t��4�P�����]�#��[���d�W���m_���Y-N-PT������C/R��`e�hռÛ�����~X7d�S�\�"��_1�feݢb��P�y?���4Og����>���Z�9��e���S�pnY���`P����	㄄j�h���:��SM��.$���J��#�����͏Y�G����4���lhI�Mx5�����Gn�&�0��F�ql�'�����?�O�t��3�Y@��C��Uu���� FJ`��É���q��Z"k���)0�+�����s�|�=㓠X��Ӆ��ؽ�[m��Z� >VB[K�ON�U�� �x/�@h�յ��쒻��}8�e__���h[��s����>��/�����n��O��r">��c���Ƨٷ^~l22.VV����������B��N%�Q�Ĝ����;�p[�,&>x�5��Ϋ.�;�&�� g�ꊭ��)}7r��3)�3��z�Pi'�C��C��+#],��Z��澍I�ϑ�[g%n-w1qF�9�ÁwX����W���w�� n]�H��]lE zk������T�����u�@��R�V���e{�EV�x��'�8��X�7|`�sґ;i�f�g��Pz,gGr���e��C�'�ncY�۷�W~�a��An=u�#�N�
v�s�Vp���O��{B{�Ƕ�z��Es��J���d��M�@��|�����:�r��܈�DǴz���'��1�IQ͆iu�l�׭�|v���@��Cp%+���7��>��H_:�PN�����{D�o��c�<�f��uQ�^@*����*"��[�.��~�g6W��t�<f�m(v,j���0P!w�fU���}��jҚ���'s�gp\�.$e�:�Pp��&`l���j�qd����4	L*���[���Z�_i������,��0Q��g��}s=���nGbXW:�}
�\���U�+�<��������Ǚ��$Ou6��|�%�b�5FAK�	��V��5��BW����8� K�>���o�fxd�O�ޭl^,��a'DX�����ǽ�ԫ~�^�W�\
��F.���.z�՟�#Y����#�ʪ�>p��h���!`�5V����r�u���á�����	��v2r<�]mv)]��q�_/wZd�l�Q~��㻘N�74�O��8��	�9p-*�p���_����~l���u�Y�Y��ڽ2���c���H�\���������
����gf�l�OZ�l�П'��i��r�k������îiIi�E�gݜ�)ͮ����l�ߖd��V1��>l� �a	�Y�\?��့H�F1yն����_ɤ���ć�����W��軀��]:a��h[�|>z���K�|YF���'$>x�TfF��g���=ˀM3�������H�gɣ��zu�e�����G�е��25�q��\����L�}��;*oys믊�N�s�)ʼ�+��Ug��s7�>Z�5�=�����v^c��6����Ҵ�Z*�����^\z�A�|<�߰�*!�)zC�X�M�[�r�v�T(G������u5[w�I|I��Q�Z�hC����F�l��YB�4|�S,�G�z8έ�6�A�}��T�%��:�?��2��j	Y�^����A8q����I�g�a��G�~���斲K<8�R�zg7��P�v�j)e�A��C��"��^|���I@j�N��+3q�t��v�A��BfW���%�8��Ҳz��t�	��	Avh�`	��m�s�ȰFg��9���(����*j����'��d{T�~�,ӹ���f�e)����XP|��v{ꠎG�� B�`��<�>�xk��Ţ}�7�g[�\PS���)�3H����-U���4��n�m�$������z?#��˕������I��u�T�/%}N]�Nў|1-��Ѫ �Λx&@OX���NN�fNZ���)����*o������܋Z�҆�ҁ`W. n?�/��_���g��@�z�y�O�����}��]��9�[*\�EދM��x�����};�K!��C:: �8��ޛŋ$��XG�9ޭ$2�=sӕH7�qJ����
�S��
�Z�i�>�d-�u�[ʜ-�9��"�pY���+��m@���F�e��Lo�U[����hܗQI���E*T�����?@��ќ�T�G3�8RʺS{���K���xO�]��[��ׇ���$���<L� :"��yd5Fv#���ǩ���gFW��F�ֹ�k�PMwK��iG�D9���Mj0RЋt\��#�>EÆhޔг(������Eܛ��t���h�w͎kE.�;���z]_�������~���)�D�PְU�����=+*	OL$}���^	v��n��*5i̳Hs8E����j�o�������{+�46�ø�a]Nbж��رq}]�uS�yy�L��`�i�Gm���4�%:\������Xt��v�8R�
�������ޟm8�Y�H��S����+��f˓����r{�XMtF%^���ǣ���E��T��u�3}�L.�ʋ�?^d�y/E�L�y=�w&U�}xٵv��gw40Л�Տm���SS�R�P�Y��؜�?������;��\~'u�	A
e��cY�Z���i�zG*��Ǵ>�w:Rw���������WNhh����1Y3gR��i1R�g��1ps[ع���>�e���-+�vq'O�ܻD�ǅ��_+kqE�Z�<�[D��<Y����;w�6��gX�,蹝�o$#�{i���un�7���|��K��*�	`$��`(Y����]~1�}5މ��}���݁���`�0u�1^�Ϯ���i��H����!��|i�������&�a4D��I6�wmuOi���%���F(����V�mʫ�FF���(�d�e��,H�m��p�O��'��4�Q��g��2��0բ��
:c,�|Gꙃ�8<I9�F�cl��ϴ�\�΃�Ylvm��ͫ1U�p8Ů���S2��Ɋ�&M��-�;�-�B��5��M���dw�ޣ^/=�0޴�XvH�H~>�"��Bþ���^SI�l�Z�|C�Z�$�Oȕ�DKioE
�=>J��:���{!�R2%�I�%I�ߝ���,2-�4�qȼ�'��E{�8�@x!�O�t4�B��S}M�;��n}���H�eC��	>���^�L�!7o�=� uM�ޏ���J�5�7k�<����q��<�)�o�]���p��Ob~��:�Ƽ#��2f	hT�`<��i�A*���Á�&9�R�D�ӗY�H�rJ�s���S�"���K�X�ol�(�qz��y���,\\}������d�ㅝD ��ǾW0�OTXC�H	2q���P1�e�:ά�@�s$拥�Ŀ�+��c���}��<��ٜ=���_5I$89NɬqrzV<w�:� ���T�=���^���fa{.���U�����o[^��A�ޮ���j PK�K\ćaP�� OM�Ѕ���4}�|���3��|�AK�#@���m�
���i���Bylt���[>��w1�K�x�4��A���:�d�M�,�L�(��E�V�<��}؉���ꧫ��mm��r�N�_�������4Jy���&��&M#Ly�-��ǐ�$}�LN>���˚��:�-��27J�P�W��/�O%m�9�G��Q��`-<ja��rR�o���UY�z�I���X�>q�"8#]k����4j��`�4���]T-���9���]��D
s����R������C<� -Gl��;�(��G�	� m&�d%"2��U9;>���PՇ�\�ȊcN���|�i�=���__�H�P�d�#�!!\�'�-Y��k �a�Ɗ� %�j�>�s�w�4�k��;b?C���=�Ȗ�k���T*C�R��������Q�44�<�6�o�8v�⥊�O�(5��g7�	�dI"bEkZgX��3bD*!������0�O�?y9���TmJ���h��!�aU��2t�����
U��0�ߢL_�$�PQ#�	IA\�N�}��~`- ������Dȧ0ٷ�`��:�PQ����[^ i�
���E��B�k|��k��#�j�EC�u�����De?�|sn؈�4nj�u��y�W�Z2z���f�Ǝ��Ϥ��ȤYB֤���0��b~���HM-o?�&�L�l�HOB��ɬc���NS���.��5���3�(�P��q�ښt��M�B��T~rݯ��V����A��A�t{��V~�����Qt��)�?��,U��NM���z��sK e��NOK�/��6o|����Γ�ͅ����d�F�N���W�;ݺQ�
$���w�s�R�%Ma�<�X6�����j�œB������6����巣㉵��wX��R�FAg{��oqX������k�ϘQ��{;c��{)$������g�x�9䶶����G��C�����ۭ�!�V�a��ā��7���$P@ѣf�|�_2�W��ĝ���|�ׄ"=�Z�da��6m�׊�t�/��#��_K3����;jC������g���eȺbg˥<����:����n�L��F�>ګV"��G���������`�C�el5a�t5r��ti��$�tD�N���+��٨�*��܄֏�T3�����C�g9|�U�E���.s���k��A�/���W)��	�%B����;�EL��!�Ϫz����YD�����FK�\d�KH�b�Y-y���Q����|��\�J�p-X�d�*���=m�4�����;��gv�!G����&�I�Qds���l��:T��F�:����1~.l�*U&�C�K���*|}�j��f��0+U�h{f:=�7�F����]�}5���$��בk�wa���E�EX���D�tc��͝4J�;���N�~)��)�RB�x+�,�go���4aj���u�3_o^�������W��^�\�.������.���c��f�J*V:�KY^4QY�x�U�tEeB������`jN ��w�}n����'�/�ۍ-��#CLm9L����.f���?�&���G��hw}�ӭ��0��K?۫��X� _�T)@��{���R�=�N���U��I^2�+EI��d*$�V��w�F�^�qђ
��2��x`�a9�-�g���.��>e =^2�������S;-��u���G�f��E��p����r��2�r��� ���@_�����%�/,b!�R4r���RK=�'�ZR�Zc����W���=��t�sٛ�F���X|�'�����>Wն������fb���2'��Qf�rdE�a������a�;��z,���靖/�W�6�m�Zbb"=�=G.3�Q�dp��#n��5��8��s��F���JK8��&�v,��ڂ����5��ֱ��nX?�%�&�h(���4Pwh�
R�:h�V�6ܟ���Pd��M����Ҝ�5���[�O��D����7zq7�z'̚[�O�onL��nn�7����T���:���3�z}=ͧ�`3�.vV#�y�?�]�⭝X�(�A׾Ή媦�D`��R��\Z�J#脥�i�7xO�ymu�e�c�L �I�nzqɉE
�"�fN�Ζ���)&�l��< O�b~��sٱm��9��&]І�ݼ}M�T�)�H�v֒���R}z4�N������Je�����ιQ��@i�s�_?�\�,���w��,P~�yc����%�����N�ݷ-����E���9��ʇ�+(�KR�%�y<�it���Գ�
_�(�=��3�3�z�d�i���\��7���d��]H�U��>�9�A�a�B]#`d1����0�D�ոě  �r4����}�2�.���� �a�
1�Q����K|�4~Cܰ����-�1q�Hs�6������?����������>���b���F(k�bϐ�1���L4P�^i5�5� k����Lm�X��!>�P��+��E�^�*t}.ň&�I5]���H3k_�aN������km�oda3Q�ĎW�Hq�v��Py�b�m/�TL���&�W�:@��(��g$�E�x���쏫3��@��!�hC;�F��Z:&�h��Y�ǪL���6�'�\�"�Ms5�,7�2�&%�ΐ5)�?�\�V5'���N��>J��⎧^���	�\�&��	<��?�n2�|�ui{r-��%����O��K�c�1��R6}�86��q>(�Cm}���8�~;��1�S�)G ��x�!F0N碈��z�Ķ-��ӹ�|hی2YL˷�����������g�����g���Բa/�=���yYV�SG ��X�Ò���Sa�rA��g��;��O�Z�5\���}����i�6w(P`y�[��O��}�a�ț���a}�������:C���5�Aî��a0��+z奜q�c�ҍ�V����0���.�3�y�D�� ]c�{O��E��'�U����$?��evɣp�ӧ����q�\�����q]d@Z�����W�{y���'���z&��ڞN��|v3¦m_���6�;��>��6�;;����(-&���л�ݿV�^���+:hm("����VD/ֲ:��Z^eڥ����R���xǽ�h|TjY�2�D;u���a~�g�R���m��6)u�@�D]����N��1ʐ��=�p�M��Z����1��}1��h=^>.;�0!W�>�5��X�;M����o<�0�x�y�9���m9��ZG�t\;�pq)���u�9~�B��^��u�,[�[EE�]�ƴ��l<u_r���.^̨g��5��g}"
35
A0E\�E����
J�܊���;�Q���.�c$OJ�/��G@����&Q�6}�߾�~r{�(�HB$a��yh��+qV��V`����S��F�����R4+vcռ�u�=9����� �F��($Lac�|���i��L��{��W�ٜT�w��}�	A_t�x^
`�~׊|��z�`�O�z�����;�l��W���N+X���YEGU���Q��=E�ń���0����:�ShЇ�Ҕ`���3��!@�n�ZR^j��Ek��0��?�+������T�˄B㞽�q��	��q� 6�F�)�"t=�G��V�E'��I���<Ŋ�ëY�,��@�F���pX�=�!��� C�C!���W�F4���4�z�yD���7@K�D�EnF�ӷcY��,3�Ӱ�>�W��*��||�/�
��8��p�ld�v绋w�Y�P�ԃ��:�H���1u�6��:��
ˊ2����G�O�|��	�]^B�Gzd�d@X��v�<_-^^">����3���ʑ}��'�.��S�Q�rz@'�N��*�U�3�w�Cw3c�V{����ܼ�E�#!D-�'���|=q����z&/�ݟ��֢�
�	�:Lb��ft;h��ԗ[W�=��wa�aY��i���]����X:�@6߯�E��ڢhk�"A�RJ�X��A��U{�H�+�������UjS�6O�����ʝ�|���u�'v��r�f�%(�B�pAԺѤ�~ƙ����s�!T�yKJA���8�&���ɆҤ
��m���Ҡ�P�<D����
���<���$~���9wvsw�_A[4��D:�Eri1�BF��?��U�U�F�"��	$-P��_���Y������Q R��.!�5�U�l�6
pC�H��-$V��p���lPw��Q��a�k�+xE����C��_W$��9����s�t6?� ��ª��KR��	�D�1Ц��Q�u�Yy��/W�_d:�+Q��Z:Q����&��C��ҳ�ٝ�bx
⻶��XJv�(�@ ����ŹK"w�"{9���S
B��O��"���`��m�8��������G���=����D��~�����/4��N��j
���S @\f�-x�IQЕy}J
P�\l��CԬo�~�O�FN�U�Ҕ,��`���BȨ��������w�k�O��;�j
k*_k�'�5S��~�D+��1g��e�3]Vyœ��;�ZXt}���9ǃ9�0p?�|?�g�e�ؙ��"ғz��?p�`�].��J**6]���!G����������}!����m��������	����mk%N��nk���U������%=��� yd��,�t9��� u�s�'�53�~���O���u*�vB1=�h�����R�jzjǱ��U�;:��G�9��s��q6�cȰ�.�T;	Xkb�����O��?���?����H���+�����I�c�5>��Ew�꽹�_wΆO���oNV��n�3l5;����q-f�x(�#���_Q���7e�].�ں9����|��IU���ŵLYΊk���c&�M<�C�@��A,������0�l�~V-W���dQ��|z��>^��1 _��}^E��]��:DVߍc�i;�<������=�Ǿ�]_\R;��Q�<�	�m�_>p��	�[�J �!'���6`~�����Nb��x ���ׇk�Akz�#��3��bBq���a�A%��o[�Ҡ�.�����T�`G��`���U)�܍�T �,9���3tԾ��8��tu�7~jr���>o��������y'�`���Y���/Ʒ���,�y)D���"+��S���ぱO��*��̸o��UƓ(�4�&�����I�/��~.�f	�Wz��@r+��Y	{dY�h�(W�=�KSmL�L��������xF���K���v�Z'�\ޤ苎�5�/y����i�M1U�U�}�)��-��.֏�__=/��e&��$����c�_�<+��-������X�A4(��	���ht�V��]!]�fbV񠞓�=�>Q5�%�G�+@��K�Jh�3{��P�In�~ʌ����aB_s(������0�r�xҫ����� ̓�X��) �q^
rx����CI�{���X�v�u�x�$�\vU�<�>��zW�( &qb!ܐ�$!���W���n=����N2����j��v��v�y���M*���3��߁W�-ǟ�z����b��N{�����Y),�w��6
�Ƙz��w?��NЌ6@ǽ#'*�Ei��h�L�a���HX�S�.ؖ�,;�^S�"���
�V�斤��O�t��'Ho
	V�[��������A�q	2��{+���� ���Y5��8��LjQ��_Kڄ�Y�ԩ��,�g���ax�����"�:�6`��
�Z�K<�B��C��x^d#�C2�j��q�d������8o}�Y��Z���)� �9�,���}� ȗ%��67tT�%���):��/|�tC�,�����y��ʪ��Iò���x��ⷧ��03��>�d5�%�^-)`��h��#g�I� �B >ڭ緱]>:�����I���\3�^҅�⭌�؝ ڍR��%�(����9��'2/��h�3H�X�Y�z��ըg_�ڍg�79z�*�B�Dͨ�H���(K��Ũ?��ĸ��բ>{!��*k��j�-�ň��$�a��u�)�˷/�M}?�\��<�"��q�'�uPe�����n$\�Z0��V�������x i>eT�s:E�b�N�4���@w(��V~S�-~��_�5� ����'�&�;@KBu����G�w��^�y�����ȭ��j�L�����L� uq�.	g.�b�]�� �}�Q��|,j �1���6��f�d�}���G��<���)L6\k!�<	A�!��\PŜ���qx(׵�l�����l�BK��d�fx�^�,����@%�!��=	�\���ܸ�U���t"�?���:۲����4������ ʞ85�O��-/3��4���5��+��HnI�?�1H�Y��m�}�"�+����ͦhѱ�6F�L*�Y��05������]|Ϫ��SD��:B���nZg��Vwp?D���djV�c�|H:t|?Q�̖�S���B������R��8�̺���m�8Uum��a�6R�]*�;'A`�'V���� T+_+'Wc�
J.���ȥ���J� ΅l�ްIu(.��0@<~v�z���Z�����f�w�}�C.�2F�_t������,��<��^�Z/SFcت����9�`o���ѕl�=��/�>Fm����R��#��^����Z���� ������^�t�-�("׿�X�=�w�r�m*��s��%z���'bf�O�R�s���
��Bb�kF���i����H�v���ٓ���m+y�JW�3��{���97����f�Um������fL���˼�_̺��M��,��?x�}���x���41޺�F���0D����>5�PW���j���P��>vPLW�p�꺮��C�ct��)%:{�`ò����^�<��Pf���k��-fn���=��X��]|�l?V؋�a�:$�!\�ZfD���/L��p���C_�a�v��T�M&�@?��/�

��b������x�P+?%C�����3����Z����"3V�ݻXrR��ZV.�}��ާ��g�ڎt>�8[��K��G�&�{M���{W0Sܦ5���Qf�ŏ'!��O���f~��u��p������iO�zk�Ji�N}�H;��6/�s9��G��q࣯�o���`\Dnw.�V��ߏ{����P��"e|�2�M��&8Na��֛K�O'�@>�x������D^4�����r��#B�xK(��˂߱[�5ߵU�����!��I#\DtR?�E��>n�32�*a�k����!\B�`R"i�">��^5��k�s�<�&�����e��k��9I���������^���5��D�@q6�Y�3re^d�3 Fep`� &������Y�������"� ��,�[���%�:��%�������"���+����m�,Aq��砂���ޭc�WBF5S_��R=�,nB,6z&��X�\���i)�<-�L������<��C�?�l҇����u���}�&5p�Lf\r�;���<S�����lј���/���Z�|򻽢��ٖ��G�S�U���CZ{�����1��6������|V�K�ΔI�^G��LP7I����)��1�I�����ޑ�z=V�)�51�՗���~͉���Ή���Э��>Y!�����tt�����+S�����y+,t�N�RcdF^1*;9�D����]�2�;�ɝh�r>J�WmҀʞg�� 哛�
����<�<D�`~�F�F�٥��h90	����>�ڏ'	O��䏏�q_͡W�����	�Y�~Gu=5�1�E� �S��V$h$��w������^;;�~�V��zB��y7>gCU�L�^;o�R��U�N����Oze3:��:��\��;ϐe��uU}�֏D��-�W�Q����W-=:�꼕�(���(���G�<�S�Q�
�����Z����^�&�U.t��EQ�wc�Z���t�|!8� ��*VD�oOFG�7���W^��n��Ǿ��ݸh�K��w���>�*�	BJ�J����!d���r��K+�6�__L���E:��Sۿ�Ӣ�^���fT͸�UyW�X�V��D��i!�j�)�Bὓ�?���w���(��)H�v���7+��ˊ���*V�#VTB�t�i����oES<��SO}�N�������YZS�p ���Da�H*���	q��(�~�P(���>*x��@��G�V{�R���J|�I�<걧�W���!�QC0,Z�i�C1CnT��u����-��9vG��Y���/�ǧd��Y?6b���QdkP�Z��*7�����]ϯ�������9��Q��ᭌ�R>'8��7��j��,)}�m��2�ڊ
쳶V�v0�s*��)0z���)uQ�5�T�푙�	a�d��Q�؀����f��k�JH�e�ɘ$���M8N�������ƛ��j�w����jbAn<.z�Q���s�MP!5c����i�됪6b�����0�ڻN$`bv��wR�R��ǐN"�kw@��Ѿ�ڥ��s)yܣ�}�?���@�3K�6�x^<ێ:;�Q�>���s�����Z5��8�ZU�'��b�ބ�7��L
pX|3 �������ɲ��Z=��ƢU_������=�T
�@��I�2��u�����[�ʲ(�4��<DH��P�s�ɐw��h�w��7��}�e3��汴�ni�Ũ+7qM� �ᠡ�x�r��TX#$Oʜ�'G�V��FL�#+���$�P�-���I�,���Ԃ�,��}���F\<Ϣ�,&������K�����j��;�d���Cf��zËC�Kh+D� ����?����7�aY�D��2�K�G|T�j��l*�9���dk��T�&�PH]�x����LDd�U
=�,/���_�������&����Gd�T^�.�;j��_X�ΜE��*7��f�9���%��+�t�)Vd����x�@�����q *�R�C ��������o�tz�`6˩#�s�YiQ����7���1�Ģ;\|��3��[�yp��[�y:H���-m���VP��j�������L�ۿ!�j͞>w��+�fk^��6�幏�DW�fo�_]�f^�	lq=+���G��S�VS#�\��V��1q���ǨL}pξ�]��K������m��㟚��4��DWq� &�0�������{s���;>d�1d��[tP;0Z�B�[�?m���U���.�z�k`-�`�%�~p���bل.����+���'��eh�BE+I����In"	YZ�6m�P� ^�O5�G��R´��?��А��ǵW��������{�p���Q9#����ў�Ջ��&���ҏ�C6+U�a-^��Ǟ�L�Lu�K��N�a�C��=�R���c�������i<��vs�h�z��M~-���(!Z!1[z� � 2�Ы)���kP�j���z�lfV§�������F���k �E��<]R�#2��v+��nǱT,���n'A_�Z�A�j�O�w:z��Z�*Q�UɅޒSk;ٝ�C�O#�M��oX'"�v}R���2s���j�̲��Ϛ���M��#��Cro��>+J���i~����f�=%�"��r_�h)*��y�Qr��3C�b�j�D��W	�x��Y��\�;h�UĘK8�n�	"�b`b�)ý�B�fl�}og9��u:���D��d�.~�mYz?p�G�c��ީ�'6�Sָӂ�X�������_���V��Q��w�J�f{OېF�U���#��b��E���K����D�x}J"5r#�����c��a�n�!��@b*����zxf�&y�V�5�����ȕX�c�������>�p��Ha��C̥h��$���W.�=���Y�}�	*�8Y�����8=GbC����P�b�0����O�hX��,H|�>�9�;F;C �,����U�gE=���S�=^��V�W�A i����s�`&[z�����G�c *t�F��LʷO:����h�&�u�����脣�PuE�vh��`[��n@d��w�Ш3\����>����&�C�ս��>�\_�^�LO�I��c�"&��M��#�����Қ�s2=����5?�=elSe���X4��,���$ϔW
֎����k��3!,J�B�ݥ����&�@ 3!kՅ��TI���_l��nl�kw�2���@�'^w�e��|�u���l�yI�mL�����#h9������ӻT�}�di�T��V�Z �ʦc��}7����e�\y)[�V��������8mho��h�7 �tj6��>�M����rV��b��	�Ϫ�����Ze�9�yU�
CK_���Ν4>�!�'�tc�ݨ��sK ������A~���?�*	K��x���V� �-L����2qRV�D��2�E�W
>ӊDb�#l�L'+�@n�0�S�Reě��i:J�B�s�g�JQKϊ�XKf�Q�̅%>Ukc1��)�����z	����U����\���p_A�z�碀%ꬉ;h��qꐥ�r�t����ʴ&��eK�:���؄g]�y~�� .ڋ�a붝���ƈ����2������H^]ݭ�^�H������4��Y��~�jZ���̆c��nr|.���U���W睙7'jx�%�;���5;ɇJ�8�\\�����&GVq���)2=�g`�~Bi�pB�86��1O��hM匋s���tz�Ɇ����2����v�R��ϟ�����*Gk��X�_���-�E��Ύ��ぞ?����2|&���G��Y���bp�MӮ���@'%$�&�tV�@`��1i��FL������U��w��m(7�4!�.�]*����D�]��x���c��.ӱٵ0v�A}J����C5�3��+4�~K��+�˓�C�q�����n��\��dv����曊�K�K�-�_#��
�Q��3���R�LREZ���}��c���BM��|̊�T.$;k��{��SVO�`�b��G�OQ�[#��d#h��%p��&Ӭo���S5��:bB;�H=QM��֝w':O����'L.j�9�d<B�����Xt�İ�	0O��n�Oc��\�s��ʠ�	�Ƅ�#���k��������\�3�Aa_Gu������Z�n�~'�1�%vf1��i҆j��pE�.�(2�n�ٴ�
Й��P,�ބ����	�5_%�F?�x]��	�C �B�ڃ	rS���@DI��S��+��o\�{nvrߑ�4�sݰˇA��(ŦL��wH�s�x}1��ȼ
��M[k�@g��VՁ�ԁ��y�fv��tX�dY7ΚM9 �T�Z�)���'���7��6�<l:?|����0�p��S����C'�[��ЇET���j=�U��K���?6\~�������U����FqT�Ñ+?��׆>o�q����{:+��d*���"����f8�x��r^(�t�>t�q�;6�*7j'�+/�9�ņ�j��� ,�[�{J�Ys.N9��F ���Xjz�� �/{��;	�;�J��v��1n�(eO�5�(�����l�g��R̭������M�1�y:U_\��q�08LT|�i�� �-�)/xہlF��;KR�%g4� �T�&z�c��A��{�X����0B	�F:�.?AV�a9 T�Κ��#�	��(i:I��&� ����O&�+�(,�cgz*�\�͗�o���>�jo&��	r��|( FϜ�_�)��f��I�2	�1c�á[&�[~	Tp�/�%Y�C8��:��`U��n�'+� ���(�jV3o���C�:2�s�������k�[3�]R��f`�uZ��4H��J.Șw	��-)���^`��əM:����(����#��\��,��w�����섰��	#D�ޢ���`8a�z���E�f��F��jCэu�5�|9\�"b�8��a{_s����3���n^��	�����N��/���/`�L�=�C5~�r�����Dd*;x��y�U��+ !T���E)@.��]�6
Po)��Ƅ�o�+����]2�*,ܭc�T��`��a�Q�t�́��9��ލ�wi��ӿQ�wN�7p҉6����x�#cB���&<�t����n��n5�����T������{�ۑ�������۲��e�U���Ү��6y�柧��������B��:����3r�>�J��_b^b)j2�ۛk��tM���n	�6V���oW���_��чO ���ɼ�������k���5���+SUW�->o�Q�.W�k�L�H��W��g��g5N0��E���T�֘�}f�>d��T�?Љ�H���h�ac�D#۽�9���r�A����><0VA!��  �5���m��7�׈i�j���u��z� ���+���P϶�|}G{���n�L�����}�ڮ�"�%`�`h�\��a�|Zf@8��V?����G� ��SK����������#��z+	j����i�9D{B�(e���B]Hr�Ș<D�6�����'�_}$[-�Y��#��}��*��F��Ď�q���pL�s���̉���u�b|�(����ι�u��/�s��O
���H&*�*�O(͙ ��e�Ak�����qq�}g��Q���'��Ltl{��^G7�G�>{�v
\3Z	�4Oޅ|$�e�*�R{r8����-�/*.��?�^e+|��/�#i3�5���g��� d��?���/���%htRS�UbH`(E0�B����SP%r��{�
!�I ���G��_J3�>�!�b�[�)��yU�ٕ�E��9?��(1n��U�n��Z�%J����M��9�$ԍ}?D�tر��gIۨp�#5F��c4��jC5�A{�\R�=����kq��>��=+��M��6�(���gxcAiV�HmDQ�?�آ�i&o�Q�ə-<��ew���4�  %��!�'n����r!���8<u\�0]������N*Xx4�&%E��#����:!æӏ�wHo%n�]-߯���mt=J�J^�� ����&�~��;���&�r��G��2Їr�|s��>�b2.�,�W�����Y�4d�*!���*��/�U�01��K�!����C���ap��$��X��>�Hh'�?_�.6Ӽ�dm,�A _�j����W�\�C���N�;�w�r]Mv��8���-[�`@[��S�D��5�7syCާxLm ���G��"W��{3�B��ߥ��k�!��uX�#^���*��Mj��kI[w��~��>��	�،,���0�jJ��l�����~O�u�w��
е�)��٠4�+�S���E��5���#�g��^R�nO�z�o����s�4��t�:�ㅚ_�q�Brqv�C��Nb��ӽ ���#�'�*�E/��82Ċt[�6]Z��29Dز�**KtB��Jp�祻�\A�Қ�ɣ�L'`'�o_ӌh_Ѫ'֠��l�$/p���-������to����͆FU�zPl��NN�	���I��ҥ*WL����޽���Dk�3�Ҋ0�ٝ���3��Ag��-qF��F ���-�7�F���Vڰ-���e����5/J�����v������^eޮ-ߐ��J��u�tp�W��� ������mc����ͫ��L7խgӭ~g'�n�_�A��q���w��/�Q�9:�h!`�I� �v��&��lu�B}F�$�V�����m��׭�ً��!�ҿ������߅Ai�����K�d����lP(o�c�(x�
�1e[NWs'p�3]�����'�.�5��Qvb���P:�����PI^�{� _߿i�����=�/w&��Rn��v�j���H����K G�V���!��Y�M����C���Xn ��]���� �ƃ����W�i�@������,D{7����W�`�����7��/ϖP�҄��3�y;#����{��_pX�7J+�����JFy`=B�3i��'��R�Dhb�8���'nD��v��ow��6z��]�p���g�66/��V�7�w޴ԫ��;�����Q�%=�ݗݗQ�o�"��0��
���bT����&����*��G]U�'��
b���y��AN�� ��7�{��\D�=��'m��Jl������Y�o�,>���eM��R2�TUȰ�+�a@���G{�F����Wݣx6�����uׇ��/Ea�'�vU�"F���b���A��y�5UU��s�]e1��Cx������ۧ���~3�I��&]����]
՟t�q�|^e�P��|׃�赏�W�XD��89��gL~5�����ؗGjy]����>��N@��2Lb�Fl��|Ûn�9�t*��Km�򡢶��8>�?X�i%h��s�D�K?ji_XK�mD��9�?�AR��,�@��T��;�Zi��I ���E�5�|t�x#�<�s��vq�����p��v��7���v"�Sj��pG� �5�E������=�"�%�fyԗ�O����J��f��|���
O;�Z��Q�ݢ�C�Z�\^�Ѫ�)TU�5}����U���<%����ѱ�yl wP[���s���$�֫�ۺ�c1����g�#(����I�k&V�F����F�};��s��ׯ,��R]���yGV����c���׽2��kv8�vA�sZ�F�A�Mi"Ĩ�BC��~�{���5)�����2R��%�C���NH1���C-���(�uR�?4zj��J8�L���J&S�;H�d�����
'=�gf�����InE[,өIT&��U��v�u#י^B"���Pe�T [Z?9�$��2Å���&N��A;v������ꅡI	gK��~�<�~������鰩xROLӰ��I]Œϱ��)tqG�/F�xy��8����?_?����3,&��� ���JΟ�u�o�����n/xB���]�m�a;�/w�i�m��y�NX~�;����K�܀ڑ�k��
�HV��������dȷ�MYæ6�dT�z���JUZ�)���(N�/�L7}�^��P�՚߯��HA�ֱ|��nJ&8�y�c겜��s�\Y�Yݓ����3ěaAÏ����{�d��v�ٽ�Y��mo�[�B�{�
]PE酰F�����6�M�ZQ�AMK�.�j�x��"!��&?=���0�"�����g#0V���Q|	�X9e�Lx�o�6;c���L�k��F��ٌT�����{�C�J�6�J�W�q��N,t�)�����O�.�OD#H��HY;��:є���+�~+B�;�:��Y��zw�N{jTځ<E���#59�+
�G��SZ�)�K��Im�:%���e��6���g�^_�EEEmoÂ��R���888d�7��fF-�s�J�^P�k6��9(��e�e��뻫�����Ѧ@7���ʰ/�;��6��֟�J�!{�S�/���n��Z�l����g[o�3��]���^�	��z=qw��:�n���:�PD��x����!�u����-�{������ͭZ N~��X ,�.?���J�95�v!���8S���;	�`�Jyv�C
##}@zruvvaFh�C�0�YQ� N��|�6�I|e����촫eÒ�'����`�Կ��?�U�-��+;=d��]�I|<�j�cP�x@��I�Q"�������������%�wf{4d���h?W�Fd�[�`_g�~��XF��a�e3��|��c����T�J�y?8� %�'*�Bh�R�ʐ!e+����� ����Ꜫ)= ��Oz�������[E����*[�<��md�*e:�à��-D����r�)��f!�.�TP�C6G�
����Q�_|u�T�N1fų��XXN0��+��z����A޿%�+|�ш�X6��Q%��=�7u�#ԦC#~�GV5k�B�ԧ諀�[�k�������ǣB�C5f�b�a��ס^<��8-�G8�§U��l^��I2e0��tl	R���:N0�+�9�|���Y��1��/�Jݡx��m�G��ΛY=t�!���v��}%i��"��#S�R��QY�%e�Ha����|�գ��8'�4�|Va�ðq)�C8w!U�d�SS_vo��6�"��It	i�W��NoO��i`���wh�?}z˖)�b�LX2*Պ΢�6��(6��"�$��(Z]��ѻ�{�����˜$iZZ?�QIg��4�Ke���1y+�$,�g�MoP^�D���f������q`V�:��G�u��br�2�j*��Zdy��/g��e����N������e8�~�3#F�'��/[����^�h�d�!�YُB�q�^�rY��Jd1*�~Wdͪ����t�ch,%@�"�5����'��=+�vf#����//k��@� ��C�����ևdi2�W+�����H$�y	l����]���c���V5 AÊ��zD2L~
K�+T7Y��{ҷ�5�6G��O��X�9�0f�%�m,}G2w�u2�W�18�����Y����ю`��Y�8w�C�U!����lLV�h��~ ��3�/a4n|��i�e2�P�B{�pƪo��V�*Ý�o}t��y	"�����{�'���X�o�J9c���MYD:9˦��O)�c�ٝl�����-����6��v�КpNk��B��0����<.�s:0�(V���[jO�%Uc���i�5�o��s6ԃU�mV򐏃�Q&�X�Z�*\��qc��:�?�O�/8��E�+>��oѻp�8\xc��>q��A,���BH��5à
)�X�R��Tb�Ql�Ij�2�O�~�R@�@ ��\wr&B}��]@5�U�'�/�%AH|}\���:i��;�Z8^@��!ƍN�4��h�ƀt�.~8|���M�_m�c�A�
'�Kz���}���w�y������l�ղ���S�����w��W�i���]^��]�ޤa������)�钯o�8�;�,����n��f=����'U�y(��f+�?�������7t���)�$qa��yI	ʗ Z��}:��`$�+���6/��װFl��z��{e�*���Y\���n����q�y;�5�B2d[�*��y�����R{�w���vvm�TJ*�r��*�����Q�*h,Ef#ú�Ia�ft��zC�'���'�x(<dd&[�zq���Ez��X����:+\�����5�ݎC���M�c��?n�E��W�P��Mpm�>����s��8c�������ğ���,5th&��s�?���mn�/ug�w���f|��T��m�D�7FaȆ�e$�h�}V���OV�3A�$H�>������C��C�#z���W��d�<�iN�Y�	�ɽ��4٦#Xa�o��Չ�bT,�8��y���-/����mLG޸���[��N�Ex��N�t3��H�'`�'b,6��>Or���'�k�Kt�3^|c){BZ;�w|����Y&F��Y�{��ՙ-���a���i։�9�,�%��|s�ǣK�-<��f�Q��t����|�%%,��P2CS�%����pv��+�*�b����kЪ��|��|��������>��AX�v�6�dF,U�adhYʙ��Gp֍m��J0�J��]��e�s�7�m��q����?=ş�5.ڇ8�[����,�����j�w�:͏ؾk��	�p<8�h���,������Fg%�'*�iD+d�I6w�<�o2�%s6ߩ�~�b~���h=h�� ��S3�w�Y�@��4�`����NYeH\���$�T��fY�kc��f�>ḙ�v���������U�����b�?�8!�'ϋ7��qQ��X l$~���-F C(�#	���Ԑ�S��<�-DF�GlY�Y���VC�����Qr��Y�"ZC�+���N�4&BDet��+�ϐ���.b�T��F��U�ag���%x�[Ap:�w*�V�n�Z��&U?�����t}ϟ�P�c���0��T`��nO ��j��M���@��ɧٰ��R���	� ٞ��9MG1���؁�:^�|E���b1V�lr��� �6v��1y/�|ɼr�$��$Q�Q��g_�X)������ƒ��G8E�d��F�R���'�ʿ�G��<10q�'"���� �&IG����Dc}Un���ƶ;�1����;��
��Rr�%z����Ӄ�7*8L�5u�F�#IRk8�MyaR U��1�IU��S���a��<��	Q�ٴ&/y]�ѫ<�E����#V�T����G줎���O�EZ���`��I릚���}Ad��}�=T���j�2���|04\XȬ$A�I�?8�n���.R�A*�Ef��5��E5D����Y�F�"�
'8 0~{&vKk	���Ӹ��$�
�1��-uI΂�f5��@C�?�.�
���$� ��X���V��,=�c0�`3�p����r�z6Y�Q'J�%�?x���idx�~7�xs��"�n{���b��6�������������@2������n���`�.yyqI|)�0u�%�ןW7�[dG��I1��r��	�L����W�c�[#P �a��XA�Y����wr���X�{�XL`N��L�vTBw?�q{�8���v7����|0�+�1p��JD��w����[�SM�����"����,��� �?�&Phi<�9#������wy!�;2l��$B�M�I���j�I��x��p��e���!6v�n:�X���Ge�"���	A�'��*Q�SIyZ�}��t��V�2��u� P�A#hH�$���f�ˇ�c����Ց���;gq����c�c�����O��a6f��;�"��G;�wE�����2U{�
����LuE #�s4�y���}��ׁn ]�9�!bc��^K�z
�k�縒e �#�^�=��i}�`�`�cJ�X=d17,�r�%]��sdm�\��Æf���,� %�J�X+ot�ik��
vuu"�|-�-愁+�_Q�?�A�4�p�<a�#b��7XZ�I�O��^��噳�8h��s�x1r��֡}��'1c�G_<O-T�^�J�������$�x*��lk���~�������83�J5�ݑ���� ���^7����We�&�N'����Q`Z�o�1�*C�c��^�:}���IY������VC�HsyS'X��&���(E�@��Аx�ʐu���%0O�W}��ۯE��2�=���$�<�}�_�"T��/��ۤ���@��D)گ�Ŭ
 /��x+�%j�XSY���ʎA�[a��K߂��B�o��ܖ���������=^j���AF�*<1����8B�W 1d��J� p� �'B��_[�	��9��_�m"�������_)�5�y�ZEe��^ݎ`91����_O���E�#�LvR�[ ���_D�4:{��?�vN����) ����M�G��30�ӳ
��5ݯ�B{��`m�3
0X7Ϊ�ѡ�a�h���1����6�Mr\/�LdmW�G�Wp�]���P�a�#�
@� �(�Pu�E��[�Y����
fݦ��i����_A���A,ǮU��gA��b�Lw!�d��?�QM�5�^g��ƪ���a�f��`�ڀ�73��3m*�������P�����7���/��|gh�x����4VƇ�ckmî��3��:�TT�[|E�����:T�����Bqa�@o@�[ڊ���ʫ��������z��V%&U���L�#�M��&�j\MR�[����:Dhc��-�����Ҍ1H�Af�+�v���m�8�F�kMd�f�?�G=�92��ew|�Fz
���fM�|�B�c�+��ۉ�@Ê�R]��w�1�c�<1��rq9�`�;;ovՌ������E��_�G�>@j�{^Hz�O���u�)�a��9�VմM���tvI̧@�f����	ݝ�����K��X��ߝ����
�L��z��z�v�x�t�xIv7xM��|�fz;���4�@l��X,ͼ�=��ׁIm��tU�k������%�y/sK����1�N�E�c$�D9�I�IY.)�(�mB�*Y��B7ՠ#�+V���{���t��I�Ev�I�Ë�y�B�N�{�u:��2L��O��%�@`4���p���c̓��""l�T_�`Rwv^E��YXf*C�L$����E�y����ͺj�gA�9�)t.��~���I�]�"À�^�&`:"L���邈l���=���`AI1F���/%0ƪ�0��@d|Ӗ{������55���#Bh}0��#%��õ�`���
������C��i�h���o\ws�욤q��!��1c�F���[�A�x�h}�Gn ��k��M�O���r9�2�ל-�c=��t�"k������pʕ~D,��n���U� ���?���-������t���3H
H�PC��0t�H7�5t�����
���9?��`_�\k���yf��1{8A2:�K8��=��Kb6M!��|	B�������1B0,[ᘪd�*l��C��t�@ƃ�g��uQ����<��8�#���S=S�ʙ�O��T�¶���K
>��$ڠ�S�����PvZ����B�ߝ*����U"g�R^��A\� \�AOs��v}=��O����w���㳨�)/>���O-N�f�=��{���67�8������E3'��H3��2���y�j��'`��)�:-�h�O� �i��T���]�nF��d�=�W�[�`n�k�c�!�U$�{���(t2����rB'�Fѐ�����{Xz<#�ҪY���LqkU�������\����pŰ[���7:����	��<�Mb.�^���an�RqwZ�m��Nٗz��s	�0�U��:��h�z�ڇpǹ��l��}yQ������L|����s���v8���-������>�}Ah������O���d{������󳾊��,����c��Z���S�\�*'��X�7��������v;�����Yv��H~c%�':��8R�X%�J=m|=�@�x�$���r]�k<߭7$9׆"��߆3&&�'0~���q6y�8�=�N��|֮�K��� 	yڤ*!������퀨Q���4��&��q��`ِd7��J%x�jWb��:��̗���E�����(�R���I�U��z+��P���Ӯ�z;)��Eg�W�O��B].�
�Bԍ��`�oX�����ν�Y�PxO$�3�`���VsD&.��d��P$�j�5���˴�%����gىX����@���a�6�9i���ˊC��Y�(�=�M�E����!�� ���eRi�TFK��� �{
�C�/�V�o��R���_ ��]$�|�}Q�;��1ނ�+�WQ{����x�׿F��ų�:0�x�y�	sFj����{)R-��F�p�/ �\�]��4�?��	X㇌$dh,���f� V�m!����-k�^����g��/G����/�𳜵ՔQ���)�n7�<�g��P�0�O��9��6���%J��3�Gu-\��s���-ѧ�	�	)H�U�&u>��oP�!��j��z���������_��)�����x�^r��=�������)ǿ?�ߞ.�^m��,PGX�E�cf�"�Z����yك��=�/δ8������ݿ��9���_թ7��n�L� �!'�@P��}��8)04��Nga��[WY�zu6�y\�m���r1�#����-�tꍄ�����E���D�s���([��ʤ5/�Ȇ��-.�%ϪW�� �p�HS�LX���n�hb��T n�?�]��R�poN�پO<�2�<D|{|�u�`|�p5�\�<��RJax8���aL���|4�c��qA5��	TG��_+!�<�'���?S���S�n��?�ז��M웠��*�����g}�4�L�S������m6��˦T���X��x�O��k���^b3ة��̅+��Λ���4L�b|J_����bm�֨Z�h��4�Ѐ��(�%����M� r�/p|h��՗���͓������/�1�b}�c����y�D�W���b߬Ǚ��:h��:�K��̩��?��[���� ��k����Z�PB�
��4a�]�OW�F@&�Ob�?�������i�����]�����ca�Vern�dq@ME��7�*����:��l��L������M+�\�ᢂߺ�F��36��lQKWm77Kc}YS1�^QQ	XN^jNVf��<�(^>bt,|:�hc���2�#���U@�Ԍ�knt�
�4�x�KY�V����Y��_�y��Dg�j�[��$&�شJ�4�:�C2�`��H}TtHt�=�d$���,���d��&� J�_��9�Wp�
]�tjn��#��jj������9ߛ�FA���;PrJ��{�G��G�7�DaD~b&��IŶ}�o���ML4�:b5Ҫ��z05H�A;��b���ΛT)�T��l�4�4Z6�:.�L˧�%`!\�.�"�4{q�n6jh��Ψ��Q�"Q�b!K�UJ��Ⱦ����?��� (�[���P֚�V�};]�;o�`���ܟ��e�����,m?���\=k>YN��3�N@)}O<m��jDԩﺨׇ��������>q��2�����@n�����9�y_`k�U%�kځ��0���2 ��V?�O} 6��?u�S���K��;WϿ�W�� ������pSI67�y��	f�d3*10�>��
&Ƕ��#���ۖ�ξ.Ӧ�}iT�A?I��.��PѦz#	6�ԤL��A�"ԗV�3.m<N��IڷI谀��+Q�sʇ�ۏ25.t�H�dU&�u+v�	�"f�_���.�y}�9����a��+[�.Pm�	��nDARf~+,b��g8��&��f��l�%+��{�BC���ySv��P,��T�'`ͨ��x_�OՋ\wQ�|gMQ*�P 	��v�`��2�>�8��J&�;� v��D3�	5���ϖ��gB�j���:�l'�}��X���,�����_�n���g}�u2��i��?'���������Ø��*����~ծѿ�)�/��0'd �m�>�U#��c�`CwkM�{/�W��؂qj�H��Ę���M�s�S��FH���3A�Xу=�P3h����$�4��~�(]����rb��'��^�� �o���v˂����Q��;���JMQ��*f��Q^|�pq鴹���0��Mz�c��;`�*�2��������� �����w��[N���ť�>�W�5���*T�D�r�����K��mm�2�"	��ʩ��(� =L*6x��q�dl��.(m��4{Sd��b�#�V���+���}�GA�x.�l:�xQo�1�8x!S���(��Z\\�+(�,d��� 'ݳ�E����$u��%��_���?���azf@�6)���Գ��s��,2��~��1��xa`�*^C.�,2^�X+���!������k����ɧ��U���
 �L����N�N�f��cm����cJ�.*�Ç;�B0�}�'20�����J��K&��a)��EQ
�]�w�/(����.u�U��`�ԥ�+���ӧ�B�����Y`���[F�"M��T��l�T7#v�� �mAu
8�6B��[�����I�;�-� ��zW�y�$��^UX���H!󗏟��WPq�Dٜ^�����N��S[��K���ja�������K�.�^)Ay�K|��_`�I��I���{��:�>�N�"}k^�;�8�����J��q3��?��M�'b;$������?Я�p	ɢ��y�{��͋����̏[�:2�q�Eb�6�6D�K�^��1#����!ry��5~V�'Cn��[�L�(��>�)6�G��Ɵ��=WGY��F�ɪ�kp���{{�{q�1qkW.]���B3R^�(���;�NP��C�U�Df�N?�;�?Cyƅ4
�%�+g�B����0�s��v�O���#Q��e�B����Ҙ͵*���>��!�*�����p��QO讙�/xR:&��H�����>���`EG���W��E	D~ݢ����y���s����|�i�x�I�[l�	Ԉ��G�]*>�I)A^2N�/M�� ��XJ^ ��dvi ~�L	����G"�n�b:�� $�@�Ǆ"/��X?�+�My,i�5����M,31R�S$��.#��/�;>o%���.��Jy�c5�� �7�^��� ,���-��ANLe1B�^C�Ze.�o�?ԭ����0�Ѻ�6A������Fp�+�6?�y����	������
��tHY������Qn䒇,��p�.ݭ���6-�%1O�~� #B ;(彎�F
�! �9�n�WYӔ�T���iߓ�4SX��_w.<�rB�ŭƗj�ZG��πQhN.�yE���#0�,�M*5�ٽ{�e�BǙ�Q|�qy������+�@cE1�*A��f �$ߒ��
� -C9~P�#���oi!ۙIײf
�Z �>�[�is�!�TS��H�����|�q��>F��Y������N��Q���/������}�S�����ڷ?���m:Ų<L���uZ����-]��ӈU�3u�Z��@nq��TXf�,����I���>:H��B4F���'Kqr!�� Ό�ϗ�㺁�L՘� �z�O��� o�9�!n=j��}���N���_^�[��
y�]	�����4Xw��ީKN"���|�F���1������z�d�|�^"��2��&���d�I���_}�v�ײ ��Q��~_I1OF�tt�x"WX��\�Á���
wv������LX����<loR�����N�Z�v���B�+���qҗ֚���~yu�,�������)RT�+g� -f1҂�&�L�G�Z�S��)GW�����S۝�NN��P;��O�.R��:B;~g:���*����g8��A8��|���N9�0Q��_5��ߊ�^�pr>T��ч���qyB��z		��I�!nab��k�]�V���W�6���k\W�YN���+g��a�f�8 $
���'��A�W��:�Hj{���[����z�*�Y;��X�6�z̶�Jͬ�%h�$.���]���K�ൺ��l3��N�&��ZT��94�ћ��[�]EJ�Uچ[L\tN?dY:M�3X+*ۘt�tn�Zb5d!+��(�dW.���� ��M5���V*@��SU(��|D���+N�7�x�| �YuFJ<�'���C��3�lO#t�"��F�.�*mP�Ġ@}�4#�x�*�1(�ä��.���E}���s�"P-�/
���-��<��	�)X �܈G_�xH�Z��"2��4s�ۗ���$�u��N)/����������~�y'�bL<U�L���Jز	��6�l"��"t��2����̯����\��%Ë�:����f�hQ�d./e�����A�JA ��YB��C��^��� k|nq�-��Ԩ�M5)ԇ�,��Yu���c�tq�'��ۼ�`a�gĔ����9�~J�����i�$iX�\����{���Q���ݿ`�_�%���y
2�zBV�h���L&c��b�e:���dM6��P�f�c���C��)�I&7V�/k��2`�t̅�q|9O���mĠ��W2m1?r�W�U_8m�*��r�ۭm��j�@��;�^�[����n�;g�sC�wdbQ#�)�Ѡ�ek�7z����ߺ~Db��|+p���+	x����ǶL�\��d���T��D������Ij~�)�)�O�"�<�8�EIigW�k�f�� �^�Ai]	���n�m�a�ު�#�3�|�+��UX�L2���x�:5��4 ��/����j��-r��*d5/��d(eUE.n�C%��u�R9�ot�	3��3~eae�ڹ�+~��˺V��IW�~n��BI��+N/�ܚ$�%�;��G{s��%<��&u���g �?�ޱ�9I2&���qF�x3�ri�#5�cB�f+5��>=c�쐞퐞"��|�Q<�rT૭���^e���i�Od��'s��*�ņY v8s�2%\nʤc�d�؉(�x�te�+ݿ��O�e.bƅ�Mwk$��0���J|�����~����D����K?%>�Kl~���������oW�-���w}���@�\�+�]B�'�R�.��e��e��_o���\UZ>��#2 Bq�m���%������
���.��ࡅ��
�2�kh�T�8�y�&ğ��P���`�y^~��!�R�xZ�cM v}�5J}��'���4�_��\�m��m���l!u��2	a|����L�m�fu<Ԗx:L��Kp����E�6_x??_q�]<�����s+�O�A~g������F*���`:mAx�O0-����#��zLI0z�7)�Ц�.m�gTnY����|�C���	$p��+N��xu�p�-*?�]�)���Z���W�8�	f2�ٛx*��9W�S����E��R�V�5TVg(D����fL*�	��h��qw�h{�2��ڰ{R����z�~��;���VZ3WLE �)� ��G��2���ҧ�����R'���Eh'�Z�<���˲y�������U���I}�c�u8l���z���lbB�-��gŤ/�Q�ĀA�"Z�T�N�Ԇ�1�W�z�iЄ9�+ RLz6: ;;q�M�e �D�F�)fĐʺ}HpA���*۶����Z�w��/�����D����tkPY�.��/��hGuy{}#'�;�ˇ��zŪ�����K��؈�K�$fo�K��w�U�l����<�"�R]�>�s��Vhc�͕i H�sd,����!S�H܂��$(O��0���1�)��Q��p¬Ff�m�@T�"?|!�/�;�AN�0�3���p_�˾��#��Z����j55����Խh��ݽ�p�w�7�2��v�Ϣ�����+��%�uz::&@@LxC��D�CCƝ�\'������X�Yff�����ڙjÆ���'[�>����j���ך'���ʀ!{o{{�)s��มj��-��Q3S�����D{ۓ�g����z�4��4��J�0	'�l��Y���|X�E�=V �������MN{^� �g�Y�m��"�O�"��[!�f�d!�����kj4X{��ׄ4��� ~�	fZ����q�{�1��v�p���O������oGDT	����'�{9��;Έ���S!�7~��thA�2AFo��^T���E6=N�e�%Te��O��b��L�"��nBDkr�[����%���Y"":0���3��hж`ߴe�Ff�3�e'��¼^�v,8��G
|Y��/k��x�F�����jV�ˬ�~b��✸�s��!_���*@���Y���X\֫�uqf��8��_=^�T(�j��	�oe�0^�Mg����fY�+4��w�Տ빈��F��[��X�&�n&�_�DHO9��;�l|{�2K��tn�ܹ$<8K��Jڂv8�r��-�6f��|i���
8zz�Z�e���8Mk�s%���>5��/bQ��ݖ�z:��
�2��ѕ=ل_x�|<��F$H�_BQ���J��~�Lo⇴��r[g~�d���`"4�w�@�;�)@:��#�3v�!!�Y���G%�����F�YFb��$�,�#�v�6��{�=�~n�N�����$"Vw� ���e�� H����A}�e�;���̓�cK���4I���E{�T�.1c�����(ǨL7O�N��QB^�^�kb�P����6�V��Γ�(��V��{?�4�(�ѩ�,)EJ���zQ�=��	^�`
�pC���
/��	|�t��i��ٻu{���H���(�r�J��U1���yٴ �jW��[_���VW�� ��f���/bs�2�y�r��kF�8w"�g��ثe�
��u-bS��]X�|���W�[n[/�R���1ufgy1�Y@L��c�JhA����G/��������l�#��Ҙ�8�k9�=Z<��lD�ۀ��q�~c�s�G�̞ ��m.�0�r����iA��'5�&p!\���u,�O翝��m������������F�w��M���<�/��c��m�V籜�?7V�վ���x8޽���#�yKڦ�&�^�c�#����}���[��9���!�a#���c�c�b�l�T���(�c��q8Y���-/Bћ����ڃ�V��=��>�C�!��{����鞺<���]�~J�?��qʇ�˿��JsE>�\#H�Ui���x�����
͠�Y��i���4R�h��6~F̟�r�#��2�z+FH�s
�zY@3�_x�r�b��FZ<���}�-�S�ڢ���qX�::@kQ`��,�C������^rVi����ӽ��E��\��c��ދ�����3g��������9=e�2��%R\�\�D���V/Wc7���U����=$�0t�g�ae�)�,��*XO_#����2�6�μ��H5}�t�SE,��a6kb8��}�.��AYEqD�T�Z��Oh�rj�{�W�b	�P�2KI�Z%È���4i�����Qó����G��v�rqÕ700j�❷���'ֵ7#�/*v�ʽ�;kY���o��ݿ�����B��6�S��a��q�ټEY��/�0�rhF2�?+4P}��8���s�l�^��KI2p���8���5�(��t>'�5��)�ol�WA���TǕ���Xi����K4t�ٸ��W��1�ٴwǏ�? �{��B��*yS�)RM��v`s�ϝ���Z�`Yo��e����Y�\u�k=5O������Z�J��|�����/��>f����@$�J/��j�e��y�8���i�-���I	���Nb��1*�8��l#76ԮU�Ni]�l�; 8��E�y���OUl5��*
�˖��D�NPg��"�����ҙ�f���f��ʳ*�J�N8�=?@h��'�}��0JB-��p̷�aS��
�2e2#�,�ZPp$G{�#�q���<���G�XqOP�XK�I�W�r�IB�����o����������	���z��O �I�� �������-�̗�0�Z���8��NN�	��?��^�ݗ���z�n�"�X��㊺`Bn��6�w^q����C='G�/|l5W�j�L
��!`�4x��8)�6�g?&)xh׿�"�%�|�f�\�}'z$���h�ӦS8���20����A�xo�^�(o�`_�b�$~y�qG����/H��8E�v�x��}�$���0Ҩ�:�� K8@��X����r	�i���nac�X{��Ho/�\\��IL3I�����D.8(��@A�w�(#�e$�����d���~�Kq�KW�BS�\��+f���_cp���0���lN{��T�v(���)�G���J�Q���,̺��(S���u88L�P<�s���d�/�M�F�p�#E�ܭ���I�e���Y��8�q6:�>�=�K"��N�e#L��y����?i�q��#@^l�<ҷ��3Hx��ϣ�
1ʇ�!���\^=����@���n�M��FfBTe[6�&�M\ڸLg��. � ���qI��)>�&*�����c]�]4U�C��w���#�w/��ާ�l9��f�$�E��D&x- �y��"m%��eT9�J�7-����f�- ��2��Q]�k����U $�4u$��	,��~[�\$�К�-T��c�E�� S�Ο����i��3�7��^&ݗ}a~�Mw_����O{�~"ʃ��zwY� 
�w��ٕ�,bE
����m{�J�B�p��NPJfm�4��X2x��5�����ۙ�}�{�G�����N��}����ݨX�yXEGR,��G
��<�1Y1�h��=kk8�0��-�7���)�-�w>��:�#����ol�l��K	xa��0�^����%�z�S��!g|���� ��x��)�^���T�+Վ<q/�:��~��O��Z�_/�riШ3�C�#��� �<�m+
K�ΚA�,/{��/�×_��?##��Y`�d�_�D�����˛3�N���S��L�p�}M����C�����6����cB�K��S�8gQ�	^,�C:��b�{[�cZ�a�븰��mIG���/:/��]֌U+&�o-Ĉ��E9�"�J�R^!���E >����p���bY�k�V1)v1q�QŌ��}�p���M�o�Nܰ�uJ��ٳE�qW9���Oe�>���H�bZ����M}}P���P�"��'�0�$��2����ְ��)�W}�����L�BA�(Ҭ@�Q���|�P/�+�5�:�Jݮ�pY�B�)"���  O?�)q8�������v�� ��$���m~YеV9r/
c�)��h��^e�?93�#��@�V7�j}ˡ�@�=Gz ��ʏ��}����_��r}��U�z@�b����"�OT*��1r�1Y�Xi�R��5!v��d-^�c�٨&>��`Ȁ��ϓ����Ń��.B�	!ҏ�RVk;5!"�i��3>�%�hB'Y�kYė̂���񳱪��<��`�O�מ� �LF�U��Z��ne�0��Zw���3�c�'s��l���� uie�U�8�0��%Ю�4>��S���YZ�g ��3��Ħ+sjvb�d��9���aVJ%���,����� ߛ2�#�)�^Paai��Du�!0�ÅkY,��@�l!�<SW| S/��,@Ĵ�OD�p�m������[S�� ��[�JA�`�VO��>Y� 0Ρ�opu&�-������裆*eZ&�s��?��c��m��%�,}�Z�(��d���Ӗ�͵<Y����t����ZH��Bx��j�b��Ɩ�nCI�LE�e�r�i��r1]�@Mb�6}G�u�3JL�]ꍊ�W�!�w�To��:�$ZH��WTb����lm;s��:�`.ԕޗ��ɴA��A ��w�L�ܹ�	��΀n��<�O����otȝ��어em�R�DWB��H��;\���Z�edk�[�"����$�E\�pt�Ԅ~�?��?�]�����*�R\f�?UefT�94.d>xlθ��|�8>�	W�O�@�#�A/�%-�1��Bٷ��g0[�nB�����	�	:٭f��&�J"�[�Ln���X� ������~ܕ�|ygΟŘ�o���y�}�6xr��%�	8�n1C�l��[�~�oh��+t��~A����fS�f�
e((/*Z��#��ӡ/Y��uZY*[z��uڹVv��M�z˻��_?��{��0�^�/q�M�hח�),Vv�C*;mu�އ�-|�����r�.=�-���,�"�4��D������i��6�G�Es��n0 ��s��^j���/ݮT��R����"k��H�pԙB����ډ݁�p)����!Lnڈ{�G!yr+�ŌP���А4u��໳�񟂦��J}����sj����a�5�M|=��bTzz^6���K�N�@���f�S
#�����7%KS4���5F~��A�����	��{is��wkUZ^6������gB .���JJ�H��r����'���I��-��(k�VJ"�m�3B�0�Gi�dpk#��~�\�n�%*p�L�?4|�me��}�����|j�i�}�5=�7�f>X��*Ds�-NP��'4'��glM�
6\�9�zϛL���Ċ�	��&�N��6C}w�|�|\�8Jsd��U�E�~�XE'�"��o,G�d��[��ju�(��np'����r�u���J
i�f�I�*m��{�N]S���m���.1߯�h|۴Ӗ2�-��V^��mb��Q=;՘�0,X8��s�koO��c��:v]xR��Nj�lel��*Dy��F�!�T˚"�*�Dn�"�s�fė���SqdS"$�Pޓ�E�� �y��4P� ��`��	��i��ͪ�%� �0����^)���[�Ad�� My�8�o�{��Is�������2�����/u�Jd��w����g�{b-�¡�o0�v��nmH��B�{����sLW���0n�!�H ^� ���潴
��4�����v ����%l8|X(�w�$�YیbMB��~lwS]�W�`a�J�k��"�+�vnR�i\2�߸���"yX��}rP[�]�H��;�Ga@>���!J*��o��}0[��tT� �WBѡ��,_�_�&Cg��+,h;ڞ����_f=M��m��E�1�z�yw��>��B��2�=c:?���۱]A�(�A�0<֚v��ld��eߥ%��~��t)��s����6�K|NsUۯ���Mf5JgZ/�5�a���$��b���X۳~/����6��T8��^<���cxu3� _R���m��8�h��뱈����T��KZnR>�c~�ޙ�O���G������W �aP��a�E���k_`������\NC���O	e�] k��ݗX�Դ.����KK�l`����і�f�D�H�A`�ϣ�ˉ�␌�\yB2�:ì�@�w|�!���� B�
$9111-M�]�
�q �����'s�*����Z����=��~úL6�I���I�`�ӧi�sG��Q�]�}W�ާn�Q[Tw�W�^#�q���;W��r���簍�I���$���ǉ��<�Z���ǝ���n�j�^���r�l�cP����<^s�KrًΨ��8���k��Ts��¯}ڟ-9Dpu����!��v�)��k]ϴ�qF��{m�r���n�T���v5�ע+o9|_����9�:�$h^�X��a�'&�㤠�ki���i�4������U~L�/Z��i~�U�߂=��>a�9��Q���^V�7n�#���%��G�w5�X` /���Uu��y���������Z\|m4�Bc,�-����l��ߡ��}o��)1���S��<Of�)h�x�O9�w;�p2������F���Q���+�����}�K�Ry�d�V��m��s%@�Ǫ�Ȝ�'�e���"h��v�f������rS�u�g�&{V(��c��Q��z��M:�q��9ȵ*�'�V�f�Gx�I�J�3` ����7�p�3A`�.��j��Zj�c�N����kõ@?�C�>���+��I�f�2�X�����`9�T���Y��$;�6��^�Sr'T��6u$��*�r�*V���|o��$GU!`����{L�����S;�K&lG\�aF�y�IǋX�0���w�	Kz���y!Z��	�4�=��I$/���saޞ���b5���f3MiESFRώ�]D�~���k���a�}b�1pϊ8)��9��b"<9>�P(�Ox	�Pa�]A�Wg�J�+m�����^��7�~� �wnyF:�y�2տ�P���Oy������>�/���.�m�T��k)�Vz�xA�<"�p�/�6��e|�K�3���3S�]�`k������Zs�ɟ	�L�.��Z�+jά�t��kN�測�Ǭ]�B-[qB��ak���~z��N��o���s����LH���2��N��_���$Ar#�&-*�\�s�c*N�g�G_a�2?%�0oWp�Ճ&���C=��R';�xOt�K&���z��Gp�A��DѦ=HB�9�����u�3���oS��(	d�k�OR��"nM����:��4�	g3Mp���.L�,+�e����1Am!�g(�HVI|��6٫�O�=w	�*�)J���[�!���f�$��Fu:"2`i��r��jP�?���i�/q� 5Ϟ�}��_4>~#���++}��	ҕ�rNɏ�8�@Y�m��泺�����m)�4j��g$��1��)����K���Cbd_�M��E��Qï�A�vJ*��i)�R≒o	gw���bV���pD&����@�t�7n�X������� ��+�Dl �*YgM?)Fkb��c=�:�â��^&m�d�c��e*�V��GY:}f��:L���iT���in?d	��7�#�;3še��_��ĕ��g*�l���4��|��fs6��uI��.'-�mƂ�����x�(���b=���u&���l\'݋��,�"�[s@�����:��r?F�W�x��������Gq�����tU�泥0��_�ˣT���ɰ���xD_�u�@E ui����Ղ�ϛ�o�����6�6$�#W@�����Dt�hB��a�\�kY��P�J��S�i�t�H\�Wj@�P�
���4����d���l�$8���$��g���E�:蔚��J���V���r}�z;���s�ys[���q��>���V�����-�_=]��J<n*y<�����jR��ο��!O��?�e}���p�&�j5Z9F_��M�a��%E���	6H�/�+2ԏ���R#}7f��T !\ַ2�=���D�m>��AڭM
%�����G*J�W�أ�ܖ��ժ+�c�R�҇`�׆�0����djXO,|,�ҾR\��#cN���1F���,��Հ�
5"k
���}B#N&.Wl������9�[�E�D�;��>��A�1<z���j�����%���x鐪��3f�Jlu���f��k��%�I0m�?�V���{U�U�]_�ip"8l��C�2f��*��`��$����Z�EO-M��%�ES����͘���'�ͣ��!v��0��)���y�.�X�ܙ��k����� N�"|�]�]��p��fZF�?j[i_���DkޕPw�Ј��h�?]G��p凯
�ԟ��������+��ݓjo���@	�P@�@�ڳ�P�C_��Әh+%d�o�}�P"�v|������&x�U���cD��<�w�\1���ό�ܚ���oo�Q��?i�0���/,|v�J��P�� 쩂�d��H�)���_���ЊtW9���'J��S.\�M�~rVT��=��=�2��؂���͇�kal��mP�!�ئ���T��؜B�J�+h���RcD��K�@�����!���,X����_���������<�y{����S�׏e�y�H˵�������<1>�'�1Y�~'j#_y��J��=����*$�A*� ���.����z��N0J8E_P_�P����������2�'ۃjX�ᚥXL,n�-�H��(z��d��j���ߊD����2��a4��%	/��P�(��_��گD�ֆ�Rh�n�q�Q�`�b_�U;����قw�\�
*���q�_�O�4yӇܗ������'��kk��� �vs0R/��ǎ]��w�E?��Yz��#t�S�WÖ�q��� E���s	K��v-m�e���Id�قc�����݄h1���*TTTb���g��<�ZQ�ԙA�c)\�o�0�7�%g�/����%��;쭖	��JR��(��ۤF���Y��k����S� �f79�I���JH|����<ߣ�cy�Uᖪ�j� ۡe�g������6>�����S7/e.�;��1#�I��s�X���)Q�h�j�9�Tb�4�����|�>Ƹ�)k_-�*8Uc)̀��)�d=��2g;}���4���D�s�Q5#cmP2�z��~5�~N@�%�t�H��`{A�z�c�TB��
�p[��zTg�m���١�Ϛ�ꄰ~�M��{����\��2�:�58f�����)�+E��x>mk�C�-To(3���K�/��� �H���r����Q�E`�����(�/;jh��M?�D,m~9���w��M��ķ��I�?�_�}��)���������}xJ��4�������XV��k�������Qr����:U������rv�,E�&ʲ��rUA�_6�J,�A��٢�ZrjAS;>s��d&Ie��z�(#6�QY~l5F��J���Vn�ūs���~�`�D������CCs�����5�V�it̴�s�,$_I����"� ���$yא��2f�h��*�P��{[���X�R�2)6 dn;��Q�|�x��xQ虡պ؃Fա��\l�f�`ٞ@CŚ��DC�����Ƕ{Us�����yb���.�X;E�G�?�L�Q��?cU�7� i�A��l���*
߸�|ٜsA�=9��ݪTK���#����z��`vI���T��ڻߕN�i����f�y�玥+m��%]����톘O�+�ʖ�A�� �@=�@�:���i��61��W�)��>����ϫh�:Q��\a`blJsr#�?g��W�:��SG�t,�� x���#�����2HȌ��:<�`_*�� �����rm�|`� !�c&ڱ$V�B��!7�0��N;#�?�`�����B�����ѳ-c�c��G(����#��ڃ��R�Æi_�v�d�pkyd�X~��[)���Ϯiq��o�z�؝t�!Gj"��A��Z4��.�yiqI-����"�A�-f� xV)�8�����������2�l������s�J�6��;*1*l�1S��:a��q�D%�ӵT�ᯓ3]��܈��l?~~R�M���o[H��R�DBG,��i���J�ug���>�x�
�eM�Q)qd����s�_���/H�|0He��2��\�MB�B���R̙R�1�{� m�ڑf�﬇T{bZh=�{�dbM�EI.� =.r����C�Y�م�+w��Z$@q+���)R܊��@p���`��P�w9�;{���#2�y'k�z��^�5�I��cqx�Z�5����G���Kbb&�0�\���t��o�l�6��>������#�v�m޷�����edZ�}e�J��eQ�$_�HVS�A[����!��*+ǂM��f?�����SZK3r��us0�(3��q�"_SV�7��PX��x~D�0��Ѹ!�M���[���0*�v6�=��:���T�C"���o܄����Ж�S ~Z
%'A�uQ�����S?Z��_�3��br�r��)O�^�2A��kp��������i*�k'�}x�n�(|��Đ��=�Ds����\Y��h}ʘ7�ٌb��}�G�<��"�+�)����˩S�6<'�BT��u0�U���e�+#��ޗ���t[� ]:��@�Ę*�WC�u%��"1�4�(F�.x͆�@RU*�Dz(*h��Fy2��^;��3�r�������Z���1geMV��^K�5�Z��_���)�z����dǛC���$XL�ʴI����%�EPL�o��|�MN�X�R�F��i9TNU!��T���U_�v������@��Z��j��ՠ���qy���剓�Ո��ӝ�Ө���Z��9�Z׭?�����ӥ��ӯ/�7_���U��vL�n���pڱ��L�ٿ(M��8����\yw�X�v �`�r�x �W@�D���n'�xZ\����b���Dh����������'�&{�����8<m�
��*�\N���Eoc�L}oa��4BgC�Į?����m�أ��9�%1�g��ͱUU��U�m	�?�H8�;�	�Dɽ
B "B ��!�а�zX�SK�N$���3y�M\��Cv��,�m[.�/$�2�i�|P�["�<�ڔ)�/���:<�ny; �H?��N����S��|��hV�{Aa���[ P�݀o��Պ�������WY���c�8G}?�k���<'����"���d�����
��ꯞ�Ywl�O�h���Z�8��Tσp%���o�h�u�UQ���X�������)��{}��	��#���-�Ӄ�(L�q ��*��@ Y�E�L�~�?mϖ�;���m9,�9��%��s0p&��.Cէ��\����B9�c|�ErX����Y[�K<�}=��c��˱�:�c�b4�#�pj���gZ�Zx��82TS4�i�eN[��mn(�Ç x�  o�y�d�ы�7��֨��K�TyEa�K�z��eW��	�(���1lHT���jS�Sv{brL+�߾�Q��#��S��Q�`��h�jjh
.c��(l���bl�@d6�8W	h�7��y5Y���?��Q���+R*ݿ��k/����VP�l���(�B���Px6�+��HAׅ4��r+u�~9?Vo[�@��,�A��|����M�̬_Hd@���
���P�|�-\/�4�8�ҲD@QR�{�j��'�n��-�b�\h~9Xp�M�g�5���j&|�\�86�^�[F�c�{ڃ�;*NSG17_����`��D�D+�a�Z-k�B�r���N\���2F��iF�I�/�!="����2��(��K���W�,۰�4��w.3��v���҄C��ܠ�e�S�
��T�rt$�����<灬��d�,�k����@uo��7�� wǆ�;K�^����l��/�7}����Iq.U*a\���m,O��#Cm���B�;vʀ���#V :ӄ��s6��_ŢI�w�i�&K��E����y֧��g��-��_��P�Xl����i�{��aޒ�������\[�Lo�9������"�Ø�p��;N3f)rEy���d��K/�!yws5cH>�P�u��ۣ!���۱�Ԟ�dK�	�Ȩj�"�{�l>6"-]G�Ak���V'�X�>>������b /	���ުTWa�䌦��x:D&�$�NA)4��Y��+�H���h��+Ɋ�ǆ�^T�.�B��Q�_����ܷ���G_&�)����c&#������;7g�{�(Vܪܳ�9*q������_����N�ͷ4+qa^��\4���=�����w{��9<>��&"8���-F�;��FIR�<�+օ}y�}��1y���������レ�����(E*�JJf\�-	�Z;�A.���`U�\�XQS��(�g�+޸���uu��ɴ��X��a[���y"���~�o���d�h����R��i�OON�q��;�J�O��u�<�/���Ϯ�g;d���b�q�ǔ�y\!t��&S�h�I�h�V���;b��2 ��&��y�b�}�����G$�Z!�Ǯ�f��-�v@�YI	6�:�f쭍����U�8�~�o`����'�O>� ���������ՙ�l�Q���#�cw�k��f��4K�e �xN秹��,�������أ!���m��ȿp���ooZ����X�G�PQ�P�j�(�R�3���<n�.�9�L�=���Z�l8�L	KH(��3�9~��]�*�J2:`�����קe8�����Z-��\�ŏ��Vd��B@��W�a��F��|���G�W>o�:ͯܥ�]�_�ް����s��Ê��ۂ��쒼3��EX�Q>?�Aw1C/��~�hȲ��ca���w���56^�p|AR��#�]#��r_��<m)��F��%�5��û�l�r�@��n�HTxD�}��+���Wu�L1�߂1�v�e�$���hu��?h�"v�u;)j�s��u2����I��|�9�,8�<k�`_��1[
2>?o��5�T����ީz܋m�@�:���iW�o�b���:����3�%�a��Հ��y�`-��_t{|���6�՟��@�Tٓӕ��RA4�YwYYYo����G��Dz����,8:�kƯ<$Jن傺}"��3��+��<m:ژـZM67����B$��ׯ��;�{�IB���\���$=�(Sk��(��]L��������|76�ה��U��=�
N`���=�6����1N�ӒS����G��Y't��`���K�,%QrG��A9'#��qSdU9�Sd��D)�{��\�Q����M�)J�y����Z^CU%Ќý�\�Q���R����c4Sj�LK1$=�_9��.����D�ej+�3+�D�q-tN�r� �#�͌)<�66RY�Þٴ�x��Q6vW3�HK�*.�Vh��H��Cac �F�5�D:�
�?��Ⱦ��>��ugy+�=�oy�rIbܯ��y4����׳���&����KT�D~Oq+̄\��e�S�f`���zHM�p�4�n/[�hF���i�� ���U�GQt����(�r�::�e0��k�
R�i�
F]�gߍ+bQ9���wCa�L�-�����1�E3)�$q{'3[e��ח�� ~*z$�`��!�rnR�|����t��;�g��=���ĥ7��\��n8��_V8�i��Yb�i������ ���WT�ㇺ�:R��`UT�W	T�Y�n%.�+�p�:g��q4�{�w���|���N5'�̙#">G�켹~��:�%�A&�z���>�"�M��˾����N����v��d�� �a=�����Ȫ���r��]K�<�z�i@�>��_�J�����Xt� �g9��%�FV���4�����'b�(U`�ѿ�P)%��a�g��b����r�y0��\>`\�Êh��^w� ��}��`���S��TIg@2�������>�ǥq�������8}1��1hz�O�\5_�$FZ��y�b�%��Y5<��q&3<,�d�t�h��;�Ks�ᦌϣ	�ʦ�Ӧ��M+m@��C�Y��X#��D�p���*�\����������:��%�Ǜ�����U�����3�U�
��O�s�[�Z���Y�ţ�.d�Z��g���Zd"/����������oPD3bd�;����X��-5�߮�E�'�k�n*�r�9]XG	\[C��O�=!h|�T ���|�zf#�9ޠ��|cU��B��ǥ��M�P%`g��㕱��ωCl�W��Ȣ;�B���8ї�D���ߕ��D��!����V]�^���t}��u���ͦQ��o�7ͣ��r�4���G�/��_�n�q+�|�D�f⊷��j~0V01�۫K_/��d ò w67�12�� 6�=CD���NA����	�A���mR��Ű�St�u�u��6i���c������~8���쾝ct�����|u_J?�:��bQ��ޞ �>0���/FR�5��:�+�Q3�W��|¶��nF��&'�]�M�u,�~X0h�_�ۍ��&2�B
��n�k�d<��-Ms�����|U��x�p^�,����m����Xud���g|Nf�F�K��:�;���5��l_�|K6?�ӫ�HG�VW���@��q�ǵ�}�������VX5Xڴ��j5���\�f�~*)�0:�ux(&��׀ڠQ�^X��G�8��ܶQ���b���u.$<�C��G,� t�۠�Z�o6��-���)H�h��^)�*���d��s���v%�V��]?g�Ty~�8B\l"�I����^��9���޶I6~�Ɏ@i`�:2
�g�>)Oa�4R����G��Ʋ<5�WR�B�%B�-1Q���9��d_��`o�+��c}fF����@a�C,�Ip���EJ2 �مt��r��j#�?��b�'�a�|`�?vFB*Q�@�O�^��4�@�7�6}sb�wE� ��4��ݺ���]:%?�8ʯ�o�ė��;&�R����P1H2A �k���ɰ�z-����T������f���l25�S󡒚�H�t*4֯����jG��vل׾X��	�R�X!(L��d�i����v�"��������=�A1�E���)BY��v3ts����b�����htrB9��.q�_�c*��w�$ŋ�)}��R�]N?a3�6�]n|�^�\���r���J�I�2�{�IKb"BuRz�t� ��?�tȈx:�
���+n�[�@�0k�l�zg٧�� ���(k����f��g;Þp)$%Z2T`�2�������t�gK�= �c��'s��O}�V:N�gC�H�BI���0�`
�٥�$��ݓN�/�7�%�����4/���d���_pPU��
�E[~��~y��j���>Fȕ��T�^��Y�XԞ��O�<�d��'�Z2�vs�b)-�Pb�J���N�^����p����1[���n���EK��_�<�_�1S���q�.U��sUǧk����r%
�m[���Ox|"9*��m�Lx�J=�Y4�7�{�]D�Rr�k�|���B���2��f��S�{{��t�d����8�}�I)j0�aC{��в���h��T!���Y����cS��E�o�˾������=M�룮��N�_��>�����_�B�6^�n�>Km*�|��ޕ�%�Z�-R)�?���s���I!Vzf|h�@�΀cmp�H�z����:����D��uX1*�&3�mBV?K�ê{�Q�ъ7��n�����6�\��F�I��b%
'�Ij`=�jm,��B�֥�ȿB_�A�Y�E��eǉc�CY:)90�Od��b�|����1K�T��U9���"��{����y��d�0Rw�yz��d"rѻ�6I��xS����"�2h]������0�w�G�(u��818��(�R�uB�N���t�8E�]UeM�f&���������o���i�fG���W�@��ta
��)�'5gk��S�FVD(T�짦��S9��#
%���U��vac��I[W�r�J���͏a�X���\��F�^QQ�{"�;q���"�Ѱ+�&�$?�S0��W�M@�;��z?s��-�t؋FO<��N� ϋ%Gg!�M��� ��~y%���K,�I��*X�/	.2]F�(LJ|l��KYbm�z�#2� q�S�(��wޮ0j������}�Cσ�y�K�Af:C�gB��uy{�pf8F��E���l�#&�b�Tg�a(GM6��$A�q8� P�P����{�V��G(W���� '�H���b� XU�����h�n�E5��:���YB��g��$w���)��l���9�o�I��Ėfo�N�ĢF�u��u]^�WN���)����
�@>�{���uVw��p,�Q��IZ߰�
u"/Y��4��e�9�x���2zA�=���2��¹xn��2Zs��
X��J���9�kQ���ϭ�D���^,�:0��lP�7�UHka�YS�5�ĩސ�:m��GB:�=�w�>�����K�A}���&Ե����ͪ
��[C���ŁbvS����"�2�x�I��m��	�ǋ75���L~���М_G�m\�����ד{�Ó��ȄA�E�L��1��!A��$�$g5������;���*P��N�����E�
���h��	��beǸGP���Y�Ӵ�sF�E6#���{�l%�4��Nޚ9k����v��E4z��?�H�R�j,T'�L��q��u��`:Ӟ�)L/��Z�O�8�#����cAVG^J6;�9n��������<��H��>����8��V^/�b�o��*��#;ru.8��Lg���:�&�w\'hV��V�/�l�pr�7�]���*������/����O`Nj@���Q��}����v������-8�����$v����8)�7�*�1r���ksZؑm�p��ao��@�>�%	��5^�B��<�J��I��("���P�ٹ�^�������F����X���1����:� R%�5�|L�68T�3��CA;/n&��7p������������K���>^��wފ��-Y�z��61Y�/�u�|��pC
L�P*�Ξp�Wf,1����b	E� ZP�� q��k0̜�zO��5$�!Ij�U�)�Z
��p��F�G|s���D$u�����O��8�7?cz�v�?>:��G�{������j������T-~w6�����d�u���:��e;��Β�[m�X��^��P#���b���o�t��鍑E9p�k	������� ��ul5��M���2CV�W��c=��nWն�i�{��B�Mb^�J:��+�i��Y~�_�ӎ�x�J�ey��@nḣ������=��VbD?� �MQ���3� �E�N�ce��V�KȀ�|��V�j�Ն���h�o��|%����-n��2ڂi�������#�UG-_�<�Ǌ�?$�0���j	UB�X� ���Q
��S��@앾<� ���Ā酈W�j7�5�!����0�}�[c�*b�_9�'Ӗ�.����?�JؾV�Nd�G����v����� öBf�0*�ncN�Qǒ�=���[���'�c*4�j��|��RSѷ�,��b��d��-��l��a��� �m��=9�Y!D;: ������֝0��yD��RڐK7��P�o��zX(:.�^c�Ab�c66���/F�%�5	-dw��u��ʨ>�tKk�w^��ҥ�V�٫�iZK3 I��H�<��:q���qE�p���J��������i��e� i}��s��~���d	��UlG��򾒤n5ovoN1F�*Q��Lj&��u���n(F_&]kܱ�+�`X ��9y���v��"�Ŀ6�y���Cjh���`�b� ���T���.z��36�=sK^�*�G%=K�E.�g���!���k���L9b��Q ��-�4rL�����(��^�KYq,I���B���&�b)�L��B /�R���"��ņ�&���N_Z�>A9F�s~8��3
���L��@�\"qN/�����VU�'��G5����
��k�{*H�f<hڏb�*��.�{T�:{�+�R\v��n�|r���v����0n��qm:iw	��/�bG��~��<s; ;(�~)*;�[:D&
���BL&����`���$PTjJ
+��7�����y\@�h��� ���SAb�r1l�%�����
��n�*�Ou:��P�g��v7�}����M�)U���m��t�s�Q��l\y���i!o�d���1iM�˸F�1��@�$g��#[�hݺ�e�N��;Q��*�C�l�9]����R��l�X^�XL�Zb�e�Y�l�]�d؂u<t�Ӫ�Y���入X��U�����\!i�|�ǶY��v&���;�\�bΏ�%h���}�f">bi�Z(c���#����)�<OOZ�p�;���j <f�5�c������w��n?H"�b>���M���B9h��þ#r����y���z�k^�+��Ϙ����g<�'2��q?��7���������a�^KZ�������P��������l�+��������k}�n��`H�Z���(����I��I��\����U���#�J��i��7���|�C{�
a.��I�V1��4�c��X�����4J#��&�F��Pf:<���3�a� >3����� ���}�x�T�j�E^O��Y��PW���9���s���?����]���7{��ϛm���GM[\s���ssi!opbFiyG� t����ʱ�T�5&���3��od5����Bd���5"��5^{���r�|ȊW�����
{�������h��b)�����M�C�����VlWs�Y ]�� ;����_�Ih+��9?d��eCrH�~?�":���Rm�����8q��l4�Ċe�ON� ��۬��Ж/��n����aR������Pܵ����Os��O�9�ӆ�]�s�k����\4_oώs�{��L"R�2X�����\�����#A��I�����L�2g��ka�ǀþ⑩I+�$O�b�
^k�U�F�U�j�u�Z�.^�'�=3H�z�z�)B�8����\?J�l�*:�7��tZR�5 '$�px��m�.��LA�4)��<.�P��8o��{�!�7�.aO�9�	L~)�CH�i>�ɉ=y��t�׃�^�Z�9�'rN>��i=A WaR~�]R�.�͸�H����Jf����Č���rd����\�, O���S��G������M��/�����fp ��d��_2U\0�sL�g����>���G&=˅ӷ�cJƴʣ��<���D��GS��~"�L*E��)�<22� IB�0�)~"�LA�=1�LI2@;���-wy�u
�[�w�(�����Ϣj�tJ��:3PuD�ʟU�3uF�j�I��S�2���i��@Ǥ�VZ���yn{��Z���+�)�ډEz�pO>�8,1��Z��0!�|��'�n1�Χ
a���"xq��D�vn�������Q���rr� ���rL.�E�4c�J���D���(���ټ������b��:�'��~���q�B�N�w孟ae� ��G6LC�sL5��Za m:M+5ӝ���(�">l|��`�0��bG�)�&���It�m�H5�4p�c*MUZ?/����?��u��4/V.�°�ɑO�$�F���������}��Cge��I4IJ��p�(�][�6Xx_�8�>q>x�u�9[�#�"ZLG���
�J���x����h�,����6��Br�S��nA�n�=b�~d=�#E1�i�XDY'�;q(�Gm���eJ���C�	�+P����%�K��/�Yw��~R�N���FBIcE�.ևKTr-�������x�Y&D)\@��9VӕJ�!�
��c���ÿV�����Y��@�p��DvI���t@ �N0Ub�w��{����;^&)��t��>hu�
��J��Bm�[v3�k%���F�5<�SҤ��@D�7��,�<�V�R2[{��b9��>v=�^fv��v������ņ��u�m��	<_̮=��<��W	ϑ�"Rg/�!֧�(���*��*=� ��U��aMԊ��&U��U��[��Z\�R5@�|Ѭ!�,��������Z=e�5]�2J�+����8b9��Vxɼ��I�Ï�BS�?3�/6�-��t0n��ڴ�)m�wk���Ĵ�鸜�﬒I��S��oKu���Z�+^���,}�J9���Y+r�VYzͷ�>[e���Q����O<>"�M�V�F� ΄R���Rg��h��,��r����b�=�d��%��]�)/1^����k����X�� �����y�-�Xj�8�)3[5	M�����8��Q��7]
\�UeR�
q�7�ojygKRܦ�;��h�ts�P������<�iʽ]��^��81}>���{����h��������j���h������J��Gz��TQ����WVr���8��wp�?	�����)x�mxR4)Yˉ& Èǌ"����=c���?�6�,��TO������`��D?��>}�蟒:�'��N�埾�������04;����[J�.m��d �&����Ejݿ9�i
(#_�7���"�ph"ǌ��m�Y��Ox�_�۷��=&�"����pM�<(�b��k�S�sQ*D���gr�`�]<P��ca?<3fw���6��C�%���ʥ���yty��I�����P�?�`>`�����rOg�_�J��[��5���kQVpE�;��x�eݳ�+���	�%�����ڿ?���~�lt`:�|��܂��&Α��j�0$�(c(<��,�	5����<."��E�3�!YZ���)�|�*�|�bp�7C,E� k�,GmهFs9i��i��mM�Є��6̓�����F ���$`���W����� �V��~�%h�P@ؖ�`���uh��M��mr��t�u~���NJ�3wnd*Ni���M��:9F��S���=��Нn������YNm`H'*��$\�5�~�(�1ed\9`y��˯Dx���*�j�����T�q���lKS�
l����䥯5�Pc����_����Z�Yz0 ��[
e�����+������]��ʽ�I�%D*<Y��}b�=�a,'?�
6��_ ���r���$`���'� %p��c��kҝͼ�G��QM%��6o�8c�~9Q�7��TsK?����6D��o.Z
��l�9GqnA�J��t�-j+P1W򠉜àEq���8j�@��>��1I�5Kf8��ZP�`x\`G�
��7��_����agk	ԺhU��<?a����^�anb���4�Q��y�$��	�g�a&�.��>8�A�����@�8�vo��Y&c�ӻa�����;��l9�mw����%�e-.�1��߹�d:��������̆���������s(x���:�V��L��@5Tł
���ת�W���'<��L�]��U�nT���@P�?(���*����53>�$�||�4}��9�|'$�u�����?�v��c�t�K�p\���M�����%S��Q��'v�%>���|5$Δ���$,f�j���J���p�<:��K0�$�U3���0�r�U�,I�pغ��mg�,����G���P�RIW��eE�����NUI�E`��M�S�������k�g����י_�~W?�.�>�:u=\��?e���4`�?� ��<�SLR��-���gwĭ,\�_<̣�,��\$[O� -�7�}@o7�^�(�Cڢ�9�*fe�B��\��Э�n�Ȣ,/r�!���E�f�4f��c�f����=X���K���n|�˽��v�_~#-�`x���q.N'5u�.�L�v8��	Oj�U�d͌��̻se@f��qG񬰺L�]l{9�1ꪊ�T�r>�s=-p�v�޿��5���\ǧk
���J�.�ͣ4���q&4+�NF\�*�j�x��%GV\�%B�*�3��3�hJwr_1�����㞾�|v΀�i��F����Ag�ApQ6���'���o],*0���+��@-.*���L����^j���[d�"D�L�>���j}��fzs�Ԣk�0m�4��+�@Sel�(T݈�ChX=�����A��?�q��v�ɼ���qn��H�F(��Jz_Y+J�v+Y��?�*��{��M�2�����`1���&1ۀ�Uλ@/��jԯ'�!kE�F���^��Ӵ>i�Nfb��ʲ<��4��F�}%��Zj?=��xj7~��d^������j�̬�/l�k�eVӥ������#1�<��������+��j	
�	ZXإ	�+�T�R�q4�*S���<��$7s��9�6칣����-X\����18)O�Y�J�J�?s��+&�D��]1AmT�`@M���BLפ��&�AJ9��_KQ�%0'���J������`�0S���S��L۫»ߞ��P���;��@��_��[�J�ޕm�o&���� b�Tl��)X��	��a��ת�X�� 2�b�@u4!?*4��m���AM�(�l:3���r��W�V����3^W�5#��ㇲpK��GE��!(IY��e���)�)?��prGɝ�߽��c\k�{j�1{��ȇ�č���)x��%���!�A�R�4��_�ηt]�C��$h8^7<s��xL��9(��ل謸���6��+��!BJ�g,R��L����W�V�+�a������a�%�d�F.���t��ć��7�݅���4�[ �����4�]�����h������+��;J\��&` %oa�C����9~���lt�e{u�$�Ic}%��c']`��It��1��b�Vpϱ��e�8�}���^0���o�@��!P����g�^`��a�Y�ţ$����Q./���N-~[�,@�S_w��6I�R�@���G3��m�m�۵L�T]މ�-�XL~w�� hE���n��G���+����L��%�-xwC�}�Xm�ݿ����0×��F����Xf `vSp�U^� ���3����D���i0����0���4A#	�����敱�&ۭ'W�]@ݲAt�&�GG������-�E�DEa��zR���W�ڟ�!�l���Kr��٣���l�78��_��>���t�%��W�������H��t��ڈF�����ԢF񤛗;8N�@f���L���I���.V�������*e��B��M*Sy�K%�u��10�I�cp
\�#�,�j�创=�s" �{�2B�*OP��i#�/��}ϱ�{���v$|������e������A�_�����L\��l��E���x��#~6���"�O �4[�?f䇠��d �a�iU�g	��-ӃҰ�v^�������
�a�;��@j3���5��X���S"���7D�e�V�O�R�4Mr�_�7����\6فK :��t��/��� ��<�������Ͽ\`ϙN���V3!�Q%�|�@����8d�bovkIB��2�M�o������Ԥ������W���yu�ϟ]����p���`q���L�N��P�r��q0<x㺃�R��ѹLۚ!K�����^m්U:�SA#p= �u5[���+p�j�N�F�g�R��o�)��p��������+�2r+��H�
��K����Cb����ۂ�iͱJ�f$�},� �O/�z��nP�@�v�LM����vi��+,��_����"�J�vt�
���k7���V���q����`
�;��#�U�W�+�/Ξ������y�Og�}C�фޥ�Vb No��$#�u9��0 ���)W�Q�/|#���z}�q�ֱ�Z�Gɾ�AJ?˭�v���u���x,���=��s���i�y��T�8��`�������S{���|�y^�M[L�d~+��3��g�H���EҒB��@+)Y���~u�t�-� k2�2+|�=�y�0$L� �Rch�^����@�J$���b�p�����M19��,�Bb\B���He��"�r8Ij��<��=�e�큷��NM5���|R�����Od��{H��Pt�qJ��]�����S��`5�)sY�{�bȎ�k���!,x��b��+�ECgv$�P���T���u@�/H�(�[/& �\�OHb6�/r��E�0��[z��
o6���)�d珂U5�����͞��k;�#/F�6��7u|���J���1k�6��PY�::�H�6����L��������%�LR��L��ד{3Bx�~c�97��O������¶������g3,�2?[��|c�ۏ(Y�2E*���t���L~Ȩ����qn�!�|C����o��*�	� ��#��]u��z"����7{�����n�����d�H�Z�eʩ�n�����Yz��v��fP����ׯ�����$/ȁ%�qa�i��o�=�ؔW��Mv"�%J�l��i$�#��d2�;ۚ"��2s�vb�@�\���->�gQr8&�^�#�y���o�R=��!=o�"^�Sjw�7l?>��T�4{x�g�`Obit�V嚜�ehk�1��T}��k̏�
��-� �r�U4G.�X��`�y#?���_�þG��1 i2S�A�	=T 0@���y�l���H1���|��{t+lgo���yT]sagG4+��,*�k))el!�!B5�6��4��:t`�+��Q�
}QIǫ��������r|:0��� �����ƫŻ�-
Hl��`{��d��h+Z�x��b�����M�i���n���.M>�#b�����L��������_,<����}�^7���ջ�3������:#�A�s3n]����0��
Rf�0Y��S�v�
�Ou�p�
Զ>��uhQ*�#��i��dfm��6J����o�!�����h(���ִdW������d��x���D��i�X��
u حfݺY����^3�}o:�V��˟�6��/�3�o�v��NT�<��Nήך/������Do��)8r���x�:�>������:��&�j����	����h��|z!��!\)�ݬ��JC6�C$��j���=m���+n)��#�D7��ҟЏ���l��t��q��i�ٷPc�j�4:?�Tw�W���$5���}�Þ�X�V�[�AB���l5�=��K-���R��X:��b�!а�����|@CoC��������U�6�/��85����]�Wz/�[��ǫ�~�O�᥯Lŕ����i.��z}W���_��������O'��O�]~;���wk����]�/�t��0���t�&�u�k*z��ve*ܹ;�����ʔ�j=�L���zh�4a��(O9я�,v�E�8�,�	��������͆:Uͤ
��]�P����A�����qo�,׊2_��UC����d��Φ� �_�*��S���p��-@o3���.E�8��?,��e����jN��1��KU%G�w����^{�������3,�~�;�qC��e���X��x>��bg'�"�`D���c��a��ZW��� ץͽ��'R��T�d�G���h�rj�\��%,uR��[2��}<�?�(�jA��9�Ü�#��@����3�a�����q�w�\���.�콨���� �'!�����ւB{̸
� +�����nr��I,1@;��P�/އޠv����꬗��_w֚������\wƑv�:��X�Y�Z!)�{�C��!o{����Y�H=�$nZK�7�C��h��Ȝ�b�|5�E8���q�c�]G� �W.Z�~�rC���;�T��H.���=�O��#��oD�CV��=:���*��(>'!����	ŝ]p���k������z���������D6�S�d�u����d��$�hL�Ld�9�t��;�m�f#����Gw	zP�Zp��A]|^&�G(̚Y����1����A�A�uP��@�8��R2"�2��tH�>��?�e��|�1cv3�'xi
�)����*�רD�+�*N�,E����-���������&��h@�����{��?KR~�n�)/�+dm��4�p	j�^�����|�[�K@��\�*K� KVs	b��
+����,T,�cy�O��0�: ������|�F04#]�d��]��@��ӎX�RG&�Рu����ޚ�U�t$�F W�ĤKq�j*�bbU�����x®b���@�a��D���Wk�����ź���<+:����������zeq�HE(.����'��,����`$D�N$�ƌ#=/!%��CI,,*M�f0���+\IR=K�,��������K\�u
��Z#8v3���/-�r��Cu�-3�R8�ZI�d3YCSl�Eۋ�Z5D~f��]f��̸����9���3���}�|�Ǭ2w���~���c�-r�0�P;�^8�9��؎�'���xX�6�-�E.��H�&���f�����* ��{� �� �: �KI��-0t#�Cww����50twHw�" �����]�Ź���^�Y��k��v,-g^������x%8��6�@�}��d��*���f<���y��옼W!mBM{RM��������ǵ�n�u���������pӃ(�z��8�X�WV��Y,�d<j�����Z[g��w{��_&���8�o�˕�YV�	^�3�f�m62�_:�����L��I�a�6c�53��]�����ح�V��QK���c�S��/��y�F3���5Ɛ�~nW���_1:���!������/I�K3�[��~��W`�;�å���Sي,��j�4o,��d/2]P��M���;Q���U
����D�:������r��^n��A�����O������D��4m��|���{�(�m�$K�U<3n�3q�J��6L�c��~{�"܎j�A�{�3��w]����L#�}��}z�[y�pkD
sY�Xj�?��`�5�o�9]i?�?��κ��h�8�t\{x��}:���}����=���J�j}����woX{�h��'@���chIՈ���ŖW�x	x�e�X �q�1fR��Q�һ����5�k���/�5^ĉ�L�a.NyD.l���d�̓}�ɫqr�K ���~�V�)���� ]��
S�0Ԑu�곴PS��DML��;�K�Zf\�Z���?��=x\rl��?����������tx�ǻ��WW!��{�==���&Y��`�m���;ւK�I�/�BUK�Wu��l`10J�7�VC���F���x�I���k��m:1�h��:��4�w�ϥ�E��\P�"�]b�y��;[��N#0W7�5�WL<λ�!�wx�Ȕ�!Ŷ����f�]�1Z�b�%�w�֐�1�Fr�eE���P�M��ѕ&k���A֟U���]<��{+���J����lm����2C0�5��m߮+�^�o����_�~k�Z���x�2
8O��{5���85�v�p<��0�#��xJ�zv#8~�7���t�	l�̯c*,��f�}�T��'{��D�J�K�O�0�U��I���%H����O��"I��0���c�?m��_F9E�&p5�v�b)���0��I1����\���đ7��0&	�_x�����erWN��S�B���L �����JCjrV��,]�	��k�؉ ���N�@=t�#��ٳBK$�64����DY=4���a�
 ��_��F���w(�i��d�eK�.�VB b�}��Z����w~�� Z.�F	�<*�E��H�g���5���I�D��)'̽zXQ$u����".]�~��'��ʭ����\���%�� �S�g�M��`�H2�v'��_�r�[���;����`�z[kIq �Y�_IAZKA�Ŀ��K��PC+(�㰀��?ϟ(�k:	�h����ֺ)&���?���t���mdI�\�D��Z�)�6��[�\X������aƙK��Ɔʛ�`�[x�ny7%bx�HcTF�[yk�;�O���K���i��C�Q_م�m7��L�]i�8U3�ȓ��F��2�{����n��lm	5��j/���#B2�^p�煷Y
��C.�)����K(�G5(�QK�ɓ�@)����)uz�#1R���4Q{-���L\$�{�����)'Q��RڷI��T���e߰�B�i�iU�~��Z�E:1Dg�(�TU�s\���?3eR�x��sS�>^h��.��Z��42��f��*� a���_թmJ���?����1�/	������6p���#Ysm(.ĺ���#x�j�sL�U���j>�Y�Pͣ��Y�1������w!&�yo��4,�II��@.�����$�����y>s�OF��Ƕ��
Ō�~.t�#9��?�@�z��eF�G�B��by+��w�1O��KinO�Q��e���/L�������!ϳL$}w��)�k�fO�"e��Qz�,�q1����K�������tȤ����3jvq��լ�Y���<�V��W�Z��Y������]E���H�xj���qݓ�ܓ繦Ր�o���1�t��"$l���{�zK����捦�(��h�Cw�G�{������a)T�<�V�F�L����{|�b��'i,��i�<6J�����Be�F�G���̷�\�g� �vW�4��T��!虜�j�&.s�H�N$��O� \d&���-�����,�1��.e&�<F5 4�=���Q�}���X}�L�H-p���HRj2�A���ݱH���Z��cQ�ӆgWo8�>�^�},�a3�9I�H�P:X�*���8�HRu�CNR�$���=�W+ͭ�����^�Q28��b����W^E7@v��I�&�'�����Z ^����$� ���\�^o��:�d��ɿ{�M�{���B�,>zCt-�u�5m<��ЄϷ�Q-�]��_Gq��^,��ER>�����d���xrd�0s���4����O���m>����� ����%R��6�#�B�V�B"FN6��K����P�
N�+�4,WC��P� �� ���{����U�)�L!<Fy<%�����ǲ	�Z*�Z��0�:Z���"U�j����/5��mg�re��I%tB�Խ�r�i�3Iz�ǰ�eߒ�s�$��Z4dA��@�i�O���f�d&%��ȜU�  n��vB\�yut'�#
p�n��q<]�i8�L]���"�)�F߁���B�x�,5�Vc�KV<I��/��<��7
8��%�t�x7���7q��ikmU�C4��l���Y�;<l��И_R�6��+Ȫ��YK�Q �o�UU?cH��2����c%���"ݏ�p�O%��%�S[�;X��T�o�Uѿq����2��t��1��ě�5���R-䢜��zc��sg����ąix>����4�D����׈�vS��XˁF���^@'�qA�H�j����4՘���rp̼;t��̠�Q&&�e��H�e�xb�L�qW��)���>����X޹6��?x��sdTy��1�Ÿq4`��N��M��@��O���1*�IZ�����B:���K<`�B5�/1=���>��DF3ڞh��^�I��1�O�"�1N_m�쬦.�~������x.����s]起@���Db��k]�"b�
�9'����Δ�to�ʡ�'\�=���GoG�gqZ�X��`�������I=k�>w�R�Tsf�;�2˪����\-��g;l�����<����/�$8s,�5�kS�+8-V�6��YB��Zڥ�=w�B �A �Mj$���9M���*6o�y�ʜ[��T��1��y)������[��PR���\�ؑ5���ʑ�4�OJ�g��\��ئ�Gxv��D �St����l��ŇOas���$TLrr1�YD��Gc����K}3?��Y���o-�_;v��J�R�����;߾o-T� ���<��㿾�+��E�2k��]�Q6vk��C��"��*�b�c1��"�/4��`���>��'��R3*�Rn�C�`&6�Ë'Z�����{��J�k���_l�[����/�񪎥2˽.,P���i&��v乼����o�_�~w�#����W�����q�w�'��������]���7��8��`��r����;�a����ˇ�}R���'[jQ�J}��	/ܐ))�����4��Ѷ��w$�K�;�ّ�ƀ��s��֋���sKŒh�߂�\1�R�qfv*G=��c���=4e�%Ŵ!�"�l���#��դJ��\,�I-N�!ZP���;O��+�p�6 ߵ�x��V��oC�����c CAn/�bp����H����M,A�P��WyEQYJ�q)0��H����O+�_�AF vM[���NN��	���J��DW���mh �����DJ|Z�F�j@lF��%>M8�٫8��h?�[_�2f'�L���OL@$�i�%��HzT(�+-�ʹ�����_*?N�^�H<
����p�oH�D��;�̞��>9��8���2����	�Zdb�.�[�_�$ٸ��C ?�#0��v��~GtsvP�!�-�ʆw���ú�*i�>�Bf��F����ޚ
 9��5��=��0��8��9�=��i �@F�5g,
N%�ݙIc$��u}(��F9ͯ���z�����8�^���wl�YMړ5zZ�ߠ
<���/�u��ħ\m;�M��r������A���
����%�0HJ��w.M�e!s���_{�PZ
�c�yz5�ʔl8���m����(^�Zi�&��&�xj���i��HS��.�"�i�� Ւ`��[�*�`4f���;v�`���H�)/o>�-�n�"��}%?��{N�Rt�g:<��M�`��۩pK_���US�{c+�α�b4�J{��z~���c���7��
�m%��$KAP�[��o����$2�^ׇ��!���-[�����7G5OMO7���1Ow��Y�=�k7�
W��r�#�2�'�"���lӗ�����t	lc���gK�HQ?t��q{��V��h���=c�3 ��f������Q��.K"��X��*
?�+�L"'<ٙ�}Ťe_~��́jzV���!1�Kݒ��gT.���!���2D(��K���/Z�P/��A"I���<���F�_MႫ�{�3��&60����W%4Ro>�1�%�
��_�E=k��l6"�-��Y4=���h��J=܏��#�	���O3.�Q9#4"��<?�[+E�v��6��켜@6��6	B3��[.��,���𪊬�S`�������#ci�H���2+yw6�`藳!3�S��}"N�
$F<O�Cv�'���p�O�����[�t���6�c7c�PʤŬUm��=[#�����N�{����Z��k,-�b�U}u;��"������~z6m�}v�P���r7��|������FӅ���x��&()��+8{z����m�Z������q��Ϋ�1��r�G��8h�z�c�> M�O5z�%��ao��#jR��c,�S1U���J��ns緬Q՘<復��e��+N|��(|b�%!BH�w��i�y�����C˿XT�����!+�L��-MCB�EB5�2)I���2��y2"Б��`�=�_����GRT�dָ=F�6�V񝸦��"�q u�N\
�Ͼ�f%�r\�9�)c��P����@re��*�jm
)�~-��j��:~��H-���ҦY5���������n� W�	Q��`��sw�$�����|�6>�s�/�fm<����xu�Z����q���ٽ��b��J�,��r%m��y
��0�U�����8U�s��ɮ-�{����k�����<�N�����5�VcT�Gd����k*�ܠ�EU?Qg6�_,!	�F\���++>X9��)�9�{8hIΦ�ӽ�]HcG��t��H
�M��j{����ʋ#�������frұ�c�2 ��z�ϓ2�������*����j�A��H�~�L�����`�¹5�����#�g�K�yC_�\�e��KRco��ڎ��9)��<�Q�8���2�0����R�)���u�D���QK��Y�y��;--5$�3yR6M�9t�.��Z�qc��SK��{{�%���\��7�k�.��.�Z��k�Kp>��?Z���#i�-�4!RSNPLߤ���Mk7�j)�9�!�'�|�jWS���n?j&�����qp֪��V#��	f��%���jG���p�Ƭ����%I<�-~��؃o7o���I�� ����B�C�I��x��/g����>?�6�vkߠQ�+R�n]�w���ݷ��hw\-rW�<�����_Z�����oU�n���S�x{�$i
�i���;f��@%U�i8�Ŵ-|�q$#Q�\h�r?�H�z\�N� 21�h��¸�^qU�RE)�-y;���[c�=����q��@Y����c$�hF�v [שU��(�|2E����� ��dK����3��,��H�	�����r<���Q3�Q^oY;�,,�5�txy��ZyG��Fl��[;����B�1�|�6�V,WUz̔v�&�m�6�O��M>[���L�ot��B$E�ףv��y�q�ɣ�'�������ݬv�;��^:R<m5��?>�������-�)U�i>�<��1h�(!*�%�Ccn���En]{�<,&35�9
&��*����I��D���u�|����a~'X?_�.�?tbo�j�oW뙔o$M�6&%�ӈ��ֵ�:�l�@�͡w�u??��tYCI��]$1��X�����x�&Ai-!=H��a)T0>�H��_�r���K�55!����<����R���(�~~�������-#b�Ra����\��_IfX���)�x�C�Ⱥo���A�p�ָ��c���x
0��8�WasF���W�!��Ћ�Wk. �%(ښm�L){��4�/�clz�ZVPq+W;�����Mi3�V9� 6�����r��a�>��7 �:��|z�|�=x���z(s�x~�7��F�V��������-��9��F�T*��^8R{�0�����������w���Lỡ�U��݊6�C�
Q��9�ƻ��r#�ˋp�J���A%*���y��,YӜy�{��o��pL{�U�^ܦ�,ǉ���.�:"w�Zމ��Wv�M$��C>b	D&��pD}`K�i�T�K��W���v��]P�i��G)F6���ns�t˒aS�e���s�d���I[U�q#����F�7t�$'��u���,;���zPjݜ�i�?��|cx*CQ�l,Na�R~�N��C����ɃA혒L��� �)��NS2�o|�S�ecڏͦb�8x�n�����n��(�@ �\B#؟~J��I��tj�R��{�x`�b�g�$�@}:�}9;��;�'ǈ�����n��g�)>����Ng^I���ˀG�Vr�"ۍ5�ݍՐ=%����x���:����8�WfE�D�έ��m�n���^�	�ޔ��\Bx
?��L���������� R�lć���k��&՝f�^������ߟI�@�f,����P�+ۓ����yJ�+)�-o��mMgVO"Q�����t��|Ok��]ɔ�Q�aԮ�	n����vIr)��q�b�e�e�{IMs������Ԅ�WN�v�����3��Z�\�Y�p:<]@Q� ��f�E�::��1Bc; 09�^uO=
�lNi�T5���/�uR�$����Ϗ<�z�KwS(��>���U�Le�7���f���-KaU&���1��<!z����2���G�}t
V�u`��N��f��~qЇ�Ĳ����J9cJ�_�hi�;㝫ࢯ՘u�2WYN����������/:���&�Ԧ*k� ��Fڎ�Ң���\.�|K�h�2�]��Uf1���� �/)g�x�E��L3(gp!��[�'l�H7��e�0��R�����೸5��yGr�#�Q��y����A�a��՚����Z_�}��J������e��a�4��U���,��mQ���K�N��4=�Vr��ۯ_Ϫ]�O�G&uh��
�����S�K8F�Q��R�ZK�OU!�J;���1��u����A��v�v����ɹvc�)�
��hY�}aa��*��[jG�ACWH�z#2�;�GJx�1�,6.?]lj\{��cq�5��l_��0�q�p��Wnk�9��)�޳x{}܍����!u�c]�Po�P�\���+�|/hVtB��)�r�����R���3(�Z���μY_�	���9n�>Z�ȼ����8���(�޷>��r�`	�⩾��?���0�o�P'o�+說r5���ki�b��~r�%���	�0! �t�C��t������M\����%&�K���I��ƃ��-S�Fԍ�۵b�;�_Y�j9my�+&��3��蹐�e��s���[D)�F��n�E�0v/�}�2�VZb����H�Z�l��Q܇kv �y�<���UY�	���;)-���M��O �G������+i�{6>GC�Ӣ�����0 |���f#��o-����lu����I�1>�����j@ؠ<̄�2�-��r��ncxQ�.?�2�k�W��ļ�4�S=����C>s�yl��_
0O�P�[	,P���}T��� �-YK%B"�ڽ~�������e�kDN�AP��Ι^1s�خ!g����Ž�������,��K�L��Ṏ����T���,��^���)u#��;�9���>���C��t�Zϕ)�6{��Z�b�]y�u1�cc���8.꩎��@ֻ�[�TC�Mܖw���&�����C��w��3��o�(Z��EW���`�s��?�*JaZ<I��PB@�ⴊNL�k$�44i���t��
d*��Gf��݄�E�q�(�,�i��J �L���Z _[���A��Q/��n'4�sR���ߤer	��B��`ƭ�_ ��0��J�/����uC�8�cW�$�  #iT���p�z�r�
4���p�#�	�ɶ��I0�`ʥ��D+�����[ıV:v���FLN���ݩZ��^3c��*�z�C\�H��䒚�%߆�{!>
�B�����'�똾Jؽ����lt��˯�z����H%J����6�k���\��ܐ�����:Z2*2`Ɣ��^Ą D�ʪL�F������]������;��`1M��]�C�����9�wN��nG�?M��Jm���c�?�e/���E�z�� ��8���܅v�Qn%9����7]��i1��PI��Dѭ�<N%��cB��}P����3�d�ӴC&�e
����6ݛ��/�K�br����L���&X��L,:��?	A�a� f79����8%>�"�@���h���uJ�&�c�ԏ4�|u��`��H(����v�y[�����\}:E�@�w_N����,�1tϖՑ5��D�0�L�����H�m�ꒊ����
�.�{� X�;�\�v�P��&m������Un=E��.h$ztd��=�72�8e���|��2)�~�V�z��&���S��������3��g��r�{�~�Uy�P�Y��t7��I�G��no�}�,����[����B�"H�o¬QR�+������KQ���jB �։�a��jh��L�.�טSY��P�P!��Q0�h����3���X|���3�BH(5���|��l�v�&��5�8}]���~�~=k�ti�;N�\�-�$���[W�@�1a8�����?���ِ��ؔQ�����KM��y��ھ����۴�{�<���N9��|�REW�{6����7�����(�b�?��?r�mˡ�i:�#�EG�a����B6�P�6�$P�����%������{�1@�!r�d��z���Ϭ�Cf��9b-��p��`2�雓vG����Z�%�����.���Ue���i���}����%��R/���)0�n�rq�x�j����`V`��Y.�O��L�=\l�znŌ�?>0(��y�י�+ E=��{w"�߶y��o'���h�G_����ky=����������X٨��O�����(���l�A}�\�L	H�1N�7�����6�M�.���Y�����d�%���4�V�$W:��~�#	�e9���5����a��H����Yp�I��5�:nY��9^ӓ|�����9J��#(���/ʨK����,����Rr���Xk8��45������S*�����'�$���g�O\�Z����C�����/��D�֡�k�߾}�OYпF� ,�	��YPY?�=���'�X���U�Z@��ݴ �HE1�����"���J�A{�cW�\`L7�ŝKڬ=�� �R��L�z�q*�N�W28&7���������
'3��Ld^]]�}�C����W���d��*9�4��!<��p;�n�?F��{��j��`v��Q�o仹�vs��q���~�5�q����'��<�a;Y�|A�����J���m��;q��,{/���z�u~V�3�&����eM���v���[���?h$X��;2#��|2ݡo�_;�2�%*�ƽ���u7��B����E��-Ń-�"b�U��<�p�:_�ב�'���Z�r���1	B?0����\������H<��O&#ԓ#WV�O����7a�|���9ztSg���oݔ�X����)�Zq���XF�9�1$DJ>3�l��n`u������_@ >:W�d���K�N�hI��{�9���
r�D�٩R݌e��=Cac	���(�P�e1*n�㸪y�DK������yH|��}��l>i5v�iT��Zx�egcY�!q�5�ɉ/�i,�{�-|�exr�,��H	��R��0W9�<���Tt��W�5�@�C�����5ӿL'���}d��&�Hb��vD�nv�� �����U�IMߧ��o��l�yb�x�}JX��R[W
��C��*eU��X�@ 6pjWQ<#9SI����p�%�z(� [8~�C*����G;��/�9�����0��;bc����e�,�������|�k?�.�F)��*��$zu޼�����+�����T|Ax�D
Ef ai=у���[������]�+p�iQ��d��n٪� ]Nn&$��N���"��&�&<z�P���;�v^����19+9�M�Mϳ'7f�-��JR����R�6{j���v�W�`B�c���fd�w��n�&�x��1������9m�o@~R77wU������R��k����B��Y��8Tּ��ȺJ�IjkCi����%t7ϓ�1e��0q���~R�T�b#g���3u���̳����eꨋ�-MV֪-����X���-�X�w��K͋���
���<����Z�[��p��hk��4��/�W �+1+��M�w�������g�ƀ�$��Cb�jm[l*ޣnm#lx�t�:1,�-iQw5��7���w4b��߰T�秣sך�1���WF�Հ]���ᣴ����'v�-W��[�_��Jj���l<|��ĳJ�Gk�<�\�?y�4��c@�ިp0�2oىA�M9x��)_�W��b���ab�tإ���6����g�\��̬o?����=%�Jg`�qL�q���<=F2�ȡ���x��K��z_j�A�K�J�j�_�&�ʏG��;H�5��l[��������0���,)��qw�.�(iko�}/%�w�f�W(��9��}����UK�&y�0�s��0�w:
v�<��/S _u�L~���#O�~��^�c숲��~��������4��k��F`)V�����"�A�����[j�Y�ؙE��K #+�\�)���3H�4����U�o�^pK�\�[��Xˤ'2�P)ߕ��?p��L+9�G���
�dHXg�Е�3�@3:0�9%W��H��R�gZ�Eҋ=t<kV� �]#A(�u�шC�S�GC��j,���D�� =��>��f��=��3�%�����價�5DzkK��[���-���	L�&��0,==��f>a*�`�����UՔ�קE�5�t\󝾐{��NW���]稜XᷝM�Vt��f=ܧ=]�(�_�?]�9��f�L|������.[��.�ջ�o�{3�+M�sOӲ����k���s�o���Ŏ��`mm��^�|9�S��w%��a:s�)*����h��������&�M�m��KF�J�:��K���<���HW�i
@H��ӛ��c,/�3j�u�׺�L٩@�1���;����85;6'�|D'A��uH:�Wד`"��zx!��j;q;�S!o]��0-g�����,b�D��k�NIUU\K��e�KS2bF��AWr�se=�^����S�j�f����\��M��ƈP9"JD�SC]�_�.9 ��1��߂�ռ�UO'�J&H{G���4��5(��՜$�����D#����j*FCA�D���IGS�+����i�ޤe~E-�UdF��8Y>�7�-��׮��L:��=��(��\D��H����[e��A8��ޮ�mo�@2������7�7��x�A�f��b����)����>f�A)���g�<:ՙ���?��18gϓ~�o�)t���9��[�����Ox���ⷹm_�N����L���g�z�t�����^��.���Y��`	��<��)@�t��ֲ�����YK!�q&E��i�%ԁj�2��ie-���m����*���W)F �~|��^o2C�8�驊<����F`>�j"��������$)L�h���Z+�ل��S�Y�\��� ��`��W���U����!t(��'$��l�|Ek��8�1������F6S�lg#��|�-6v�t(3NQ�f�P�xy�֐^~�3 @rC}����F	�������SV��,<
�����j|%�,-�f�π�Կ+*��sn��+���+�����:����/���f� W1׵<��9U��/*��oa����Ev�114<�#���4w��~���#oOXe��|Ki��]�Ԫ��9JH�v�O���<ē���J��A�U��+i��ez~N�m�����IuZ��>��+�$�1��wb�V+����N�I6C�7ш����B ��3���{��WA�*���T�M�%-e5%uy5Iq���]w{�0Nl�FG2 �cSr�maĂ/y�v��E=~��L���Vw7��St�2HF+��z�����'�s�`���nH�>f�� �����8�*�#(�
p��ch��x��@��F�Qdsi��C3p����X
"Iҿ�>s���yc+��ZaW,����k�4ބ<��Tb�JM���K��m0,���}:l���ԗ�5��� $�T��g�����6���V.K�|xƢ�R(uy��=z�7��U���G��cG����x|�'��Y*��[��*{R�_R��3����}hNgc�����uئ�$�吰C���'_�׽��?�
\��|��	.*m;������,ֹ���/@9^�%��P�]g���K��n+\��ݠ���Qu�v����!�4N	jv�k�m̘�����yt��?���FM�Qr�h#�}a��J�1�Y���t�a��1���9	�EbReDR�l�笧���Q�c�ͳ�k���6 ͇�����y3l�v�}����j��e�~ӊA׿I��X�
�7�\[uO+I}>W�����8|�×�ꞑ�f�\ݠ�C-��dc:�$<���}�q�,W|I��H�)G_�?3��@����R��օY�e �[���@�W�yrc��Hi	"�M�|��Kr���F�K����ۤG,���=���J¤���s�)��p��y,�~9����t9�������ݚ�gK��T����_^����h��7��N4^@#�������~`��������8*8xP�6R�Z@GԬQ��\E�wȈ��II%2;���LYï]Z�l3�U��#*V�N��r����~�]���J���T��kw+��_���D��NΩ�o����=���T6�wI�iw��t�4?�`��Q�9,w8_uE����_�v�B�<�)�[�YL����1���)25T�d�� ���Hё�E)�$��9̯J�:��ˇ�)�	��F_�3��"���oن����B`�J�ݟ_|�LG�?�*�Lٰi
��l%q4-"4qv)R_>�ɪ�K����G��=I��8�r嘐����"���0����|���]���/���X+#�'��b��i�������1J�R�N�{�4W>�u�&?2�|qan
T�=^�:G�+?O�_<���S�_k��X0�����s�d����������J]<��o���Y
�?R3cʛ��\���)�1-�f&�ź\�������urA���,�A�-�jn�T�(�Q��N����R��v�zpU>����G�eT��[=O��̢��2�K�nmO��n#l�����k������O�jjj����p�����w���3��2> e3��2d�L\������)��^k�:���$���٪*�E6>��lXO����@�WG$�t ��s|���"��[��YZ���y"?�����T|��d�u�Z���7/�,-�oXD� /��/m��f�ڇ�t ��j�*9G8L�q� �i��=��6�VqA�
q��=����1�\��jL-�Z������(K��-���k_`&_�a�/�D��6��NkǾk�y��"B7?fx_�M��}�'I������-�c�%3�w_CF����I����P���M�ɯ�n�f�#tsS_���2|2V��zj�2���uN��&�.�����wP����`�w�U���bmB`�z�f�T/=R+�M�x�𛩡S�����(��67!����Bc,f�۳��7/�|�}�h��߆��ܓğXU�A�@�Ȯ�8��q�8�ڢ*+��T ]%�s��>�3�jvHes=���ژN�+�Lڄ��75��4M���� SSr@pyfqZgE�u�	�<�2O�&�l�1���F���.�~A^UuI�OQ�����o�5��S��ڼ����������&Ľ���6nF��_L���K��ݮ���1���+a*	��ˢ��5,:R��aq.�0�*1W�'<�z����J����!���C����5TVh�����q�
I�mI��`�@��а��E�e���.��B�s@�ŗe� 7�@7dt�R��Z����t��x��mGu^~䄫Ř&�̞�H�=�u����5>��T�=d\{���Y~�-�0��{�\,i�1^ �Q�4�7��Q;<�)���s.���eh�X���Y�[~�;;�T~�÷t�%�"�xM�n~#�2�+�R��XC��>z�R�40�<7zwF��SJ���.��m�cI׻S��z�j��-B�l���&���х��"3� ��́G�,����������Y�u3(q��$޴6Ʋ;T?~���������~�9��3�<�H���:H��}�^��CM3f�n7�O�'J���=����d��3g�5���"=9ԍd�1ܵ����4�'���&R���)�����#l2B��2��'��l�.���0b
�ς2��j�����u�����<�R��C	V�ڕ���4�l� 02�߃����G�������8��L�F���<�Y�>'��:/��$-CP������� ��]�i��������Տ0`z�!=������Q�	3��������@W`K��y��&[ٳ랢P�?��!�s�v���>.9�8��!�>�,�=m�m�w<�-�>LU^%��>β<d=����w��ޮ����?�g=^�_P�=��[���c��X�B�h(�r5��������), Z]���>t]����ʴ@
=R/�ʰ)�VwQH(��	a��	j]�#Q:�A��U��?K��k�j�*�a���H)B����y0�W��g�	)7%���-TeVhiD������ƙ]��x��
R�6:��*��ULWr�$�3��� F:C�?�^� t�jwAxh��2�Me%M.E-΍�E-�������O[OW�@_������	���;��G��Yg�&�5�lx�ނV�!�oä?[�A��̶�)�E>0��{:P��6�O�FR�~�z]-�*����S�(�4��8��y<�������B�b��?���J����\';�s���u�g���E%YYZv���H�EH���P�eӛ_c���ߗ������Xj��ۢ ���Ɣi��M��(2��Vtt?�]_�\B�&��l�o���,�%��}��lT^��m�>�W�2imྱ��ya�<och��la$�>������߱�����Vj�Pv�\qt��\"�'( ����̙n�0D���ީ�s����Y�Y?�3�$�O�{�;����e�W�����::��m������a�B�2�!��M�M �����3c*�<�M��	�G���s�����A�X���ʂ��!�*S��KJ�u]]�Q:��m���������gC��L_f�y�Q�.՚��k��8_)�0�O0��l-P/a�ԑ��ȣUᲅJ�N�ͩo��,i_26���uE޷6/��L����������� $Q�����1��oG�W5M�_�J��s#�;I�I+=M��6�Y	Lt1TwpQS"4����H�r֥6!KM ��A\5��e�fM��&h��6gr�2n���l�Y�/�`�-����vo G�_�����P���""[|}���Ɂ9�T!0xy{q��YE��^)���c��#�V_Sd�.$�4�!(>�^9qfqR�^2�'�~&�'��G�?��2��.j�@[Z(��iq�	Nq'@q����P��	n��Nq+��H[����M������Lf��$?N�Y�Y��k�� 1��t<���,+���H"C��(�py�s��V�b��Mͣ�O����`�@�O]O�QipWW�l�;]�uܣ=ߢ8nvc�� Й@�/��<Xxp�����Xl��'W�H��Z(A������ZI���톬�)��Vd9������ݚ�B�Z���\��yչ?3��'����]\@���z�j�1K�·�/���m{b��3|�v�r��W���=���
��3,�C$$��AKJg�s;\*M��5�C�b����]�*e2
3��O6��ɻk���2��3�a��Fg��)��ie�pn㎻]���x�ڲ*�Y����M�c]:{��x���1�F��fc��_z��k���4֕ڥa��ܩK���Z����^S���j��y7�٨�#� �U
�%Ok�H-�V�WJ+�>�R���mM��G?{�F�z��V�'�@'ӛ՘�	C\��J�zZ�#5ɠfvyl�ܯ��uj*�0��w�>R����3�r0��L!y��2`�q�p&T���~�0���Υp�2�1�Yc����>�]��^�%�����RRR5	�2�C�w0������pϜa������ݓ�q$8���I򅔍�[N�~]8��"K��C�b�ΙC+�������"�'�\�~�;�����{c;�����y���;n�����������s����=�k$�Gbw��4�e}!7�ǘ�tM�xT�Y=���R�|���T��
�Kb�WN�GM�5L�Z}$D�>�@�}�<ݥʖ����?S��x��������%�6���c���w���l(���IsP��jn���T���?Mg��;�RSN�|�+1h�(� u����)}�)S��k�4f�"_�T���b��e�eJ�6�9�0-��]�5�����;)����v�G33h��F]�a<�c�0�,�~��D�-�ӟ@��1�����̊zCeZCC��Ui>�2/�>"$s���
�R%��s�b3)�Ve��LrG�k��Ȭ��<L~֬y'����cL�NG\DKD����΂�ւ���Ca/�A6~�k��~(.���%�8��5C���l�L�K,6\�~���B&��J�Ɩ��v�1��U��C�1�9Ӧ�^^�������SS�$x�O���QTS��dژ���Q�<��&P���q��mT��Ru�7h�<�.�����=�+f�0���,�)y��m��:O��$��C����\R�b
��Ɯ�̏IU� ,$��j�zjJ��X�~ܺ?sT���P���7CAnŸ[��@p�墳��X�H��)x�pM�=��I�쳑駬n�Lo�B�Ŧ_��}O�)��ǎ����I����bOA�1P$�u������֒�$�D��osM)eN8���pံ�:@���>�	��M�vp����v��O1Z-!3���������蔆����˛���ҝF%�!��gd�u���\����cgH&ĝ����y v4Ni�0��HD�n���ۙW�WW4��W�t���mYYK�q� �,N�G[֑H�J�{u?�.	F�sHD��N��y	���-n:AS��13��W76�L!O1Z`W�����,��{��q��K�P���J�'�|&ԼB��ڷs��[�i��J�����E`��C��ܨb��	�e�X�5V�`;��p�h�������������Q�,������[˞~��+⁄�uDݑ�����[ػ!q��	M����0�Ux�X��3o��=���c54�~V�7���b�8�P�P����5�}�����QQ�c�]l���G�c+W�V�J4_���s���u"��2fWP��1w|�Əx�6��b!��C��ę�I�@Bh�2fd��̜��Z.g�H.,������)���V�^چ(�}�S��3��M@]��%��ϳK�ţhQL�w~�*�/<}9�������x{(L��T�!�j��~�5���K���C��W�^��P|'�4�N��T`(��ĘO2 SP8�K}���nw�/�}��xG?G� � C�Sw_�EB�D׊���V���7�y�5�
��n���3H��p��������5��K6�9���jo%B���٧�
 b�*3X�4Bo��㾵|TQ������.]�E33&�vꗵb��C��p��E���h����X�׆����PžK����?'U@ `�i�����+1�'�_��<x���@�W�p��+-4��c*������n{���������t/�RA;���\i=�����#�Bsz�� ������0D q�����g�(�� `3���ٻ�y[�آI���o��:	"ǭO����e=�g���G6Y��M
{Td}Y/����߈}��~|�}�1����������={��nv�qz㟻{��,������|�o��+��'��>�ӕ��M)YMN����~6��.���N����(dH4���з��ͅ|#���~}����=,�J�t�"�UCQ]�&?�B��)����<�;G>_ڿY�o�j�U�Se�&o]Hz]�P5 Z�2�����S�cm�`~
����)���}�Ö~�S���oW>n�ֺjѧC���V�h�m�z��H�����z�����|�f&���]�uk�p۫�oOɊR������d�$�ǿ~��q�e|�!� <y��ς�Y�.�'D� ����Rk]���ݯ,��؂�IU}�����+7��.�=� ��1��Y8��x�/78/�`�Q]�O0Yù]ZB��\�U�Ne؃�fp���aq���JMMM*_����ao���Y�d�w��^N���+c1.�������\yA�t�㈈�-8�Z����{N��SE�j�g���Z��}7�]���}�'��ҋ�Xz������wt��
IJ4E"����pz��2� t�Qj��P9�y�n�A��C8�Tt�yj�������<��S"��*�����c�I��.�1�wqV����0`Pm���]�8X?�A��IWq���I義ocL(ht%+�C��r07�YpP[���������tU� ��ir�K��z���TF�zL!l������6hg��:��"��Bp+����ļ�KK�\�d6Ӛ)��ׄ�v8�������?M'�Y�-��k�<�|a;�_�	vr��.��)�/ÿrssۛKk�r:Z*k�s��k�$L�>�W4\��"��^��P:�Omu�����VS@ ���/����-���J嫆?]�k�C&}Mzco_o�HP, 8%ԇG�\L�==��o?� ~���E������`Bk���8�W#D�ҬK&��m�%�a�z^�9}y�[����ݠ>�D�bC��>D�阜*aLaܿ�ut_h����D=�n.C�;�b���'�?�'�Kv�"وa����.=3elHnu��)R���5'kro��Kp�ߤ��w����6��/G��Y��
T}p�<��4�Vἷ�4��P�}V�t�����=�dE�$��vg�YIWsuz�d��_3���O��NP�p�Rn�z����d�
�t<;7�n���t�p�iM/!'T������ӓ��S�&�&&���Q�d��j���ώ!oL0���+<b./�Ajb�4hz�P�]?[Y	^)�t�^�I�#-8�i��}?�`F;�p����� ��܇O��� '�i</�9&�?�~���+�5面�"���EP��=P��
b�*�_�*�o��m.d$���c�7BP%>�M�q2�W�:ftۣH:��|���WU�LF�;��谆d��pS�%83n�!f3?�������� �S;D|�a����s
W�d�@U��Ϭ�$�+��8-R�T���x���� r}���.���޲><��K�Ԟ�M�wټ��X�r����ٗ���ōu�n�MsL穖�h	2J%���L�!,(\I׵�C�6㒂�]�$1b�	�C0�r�K���k>j]�C�,�<o��{?��N�Ȉ�~�8��f�ߟ�m;��;�|���[��^�}8[l��������}�ڭ|8 v�_�7�]t�?a�1 ��{��1����z�ˆ�2K������B����;�N�Ͷ�I��J5ly�q˩�UZ[�WB��ſ�c��5��M��j�0Z�L鳁��8��98`�:�k�1e����%Gu�|������*��b��D�UP�^��F��b��m���⨉���k�/	G|��a]	R���H1�$�Y���VeZ�/�R,�H��x�)�V�I���^�^˗q��hqR�Źns&���j��gݥ��������挙W��������lc]0e,s��r��$�ϫr4/Qn����^X�+��G��$�� �qԥ�`��� �>g��b���q�~���ki,
�ih�� �UD"u��YG��%Bȃ�zDG>��9�5:����7r�0F^pj�и�yA����{��5�u�����W��� �:�ԉɜ̮��wb�d�M90�	)�d�d7�%<�f�k���mj�B��k������҈��\����%1�M)� ӓ��b���j���p_,~��}:��r�Q��?�'v�Z�[�:ep������ʵ?�C!�	��
�Ō���1��	4���Z�ޤJW@���j�=*����/˲���
�
fx��U����ކ��b>����,��!V��&p�k�-��N��kN����+�R*7(E����f Z�o���F��4�3o�_G_����w�h��E�����T��u���ݖ՞&�ƀ�S�`P��m��]���l&�#�:�2H�F믡�1������P�صM��>��i�M���
(�a�`I��=��q5�{8��H�t,J���f&�{���r���4������E����gz��=64Y�v���++�z>�Ͻa��m��@���/�zhi=Ӄ�赴,���tɨ�L�^Z����xRn�v���S&�����s�>Q��>�/GKG�e^Ť1I�ξ�׎#mF�^����ql�QIyss��P�"���?Pz �B����US߹��)*��r�,?(.�ƟP�@�~�\��gO��Oʞd�P�������
"���|A�9]WpGo�l�P)n���pwo���:�N�\��J�rt���*�B��$��k���l��j4Ԗ����5�C��*��&f��77h_���f�4�O��g~}��B��UBg����2�N\L�K��q�a�!�X��=�*V�y���13�
���ϧ�����M�eװި��5Nff3T^~S������#�(.�M�~�ęϖ��r���z����Ðq������R�]��Uq��=d��ng߶�2E9�n�p>S�޸,�s}�|(n�q �V\%1��45Sha�R����BVt�jS�t2�p8��NH�����F�	!`@,��m�ڌ�q	,H8��eZ1�Q#��-�D���7�'�i��I��W�۷	�P$72 ֆG�|����n�r϶`��tQ8��J��\�.�<-ZK�e���3f���c-"s6<X3:���ů�gT�� ]P��}�<\/R��H.���Q� ���I���Ms �A��lK9�	�_}�V�S��E����c���?-~�.�~�9��{KS���W�A���=(��=J��Z؃�HF"�%=��C�R�.S�3nߗY�鵜�5�Y��u���X��c�wۘh�c���N�&��P����N3d!��V{R�n�$�l|��}"pC�ӧ׉�f��?�XxHp4���͡*:��,.�Z�|��j��x%�������E�릖������~�Ce�#��C�����/-��a��-������oF��)"�k�w0ءϾ���Hy�o~�ݡ\���L��v�����j�k��}�׺�%�-t[N]j����$z�Rq�vg�Pw�PRUDM�4��U���n8�㯲6��{�(0�~�T�\��$�zN�C��!�{/ENN�[���g#^_N�,��6��� E'?�!�|��'��/fOO��	��5�_������}o��N�b�{�ہ�ȗ��M#K{Q�|��ϭMvT=L͋k��Ks�g��c������\��/�}�{�˃-��kg ����\�˗����v�Ryt�e|��c�wkkk�솊�a:"���t�2���H�e{,���^��i:	Aؖ5kȧ��?�w3`@�Zq8s�~(r���baZpn[q'��Wȹ��:��!M�Q|tR*y5�DlV�T;ů�v��nz�]����|h���Q3��������$81%%%;�H[;l���)@��ɏ?:c\�`���^p��Ĵ>r~���%?7����^~��4�	��� ��X����(���6每#��:w��d�MYo���͏^�Ǭ)��|���i�{ѶB�b���@����$x�͊\W}X�>q48SL��0�q�h�ǥ.��6�8n������fQj����fxW���z��]�[�O���@���^^��V�U�\�J\�;׭D������hk��S V�Bkz��-!ї=�����^d�k]67(Ώ�=U�\�k��AX۷�t����@��2��;
�Q(�S+�@ �6���q�q�u�3v���!�)&I�q�ܿټ�.��O��Ih���M@>3�XY�Hb{b�9�4�B�t��՞f��$��М��A��y+�m�h�H��7��ixj��U7eh��>M�n�����������yA^��T�=�SSZK�9zQ{�U6�t�"�2���;�MI0�М2�5Z��NC/������j��s����jj&WU�����b�^D�&�W��͘ӕk�sEC���LO=�-hh���J�����jv_BS��wl�`�n����e���^&>&Ǝť-������1']��/�\�p.\���x�Þ�$����J0����L���_s�?���̏�����o�&W���Wm�L�SO�0Wd>�wmP��|\lĽ��|�S�ㆼ��y��kИ^���7��Q���(:�������'u�%���x�Ƚ��k%���lfQ��������&���7��>�|*���l�,� ���Z�Y$׼���� ����E� �}�|�������t��R�ζ�e��E�E������C�P�K��~4]���c>�_�D�P��*�4�� ʷ�A�����w>o�x���%g�m��enOZ_�y���k>>�#I�sQ�in`�|;��f�Gy��#��AT��	�o,c�fL�u�Nr[Ab�%7)NO��e��P���U���έ��X�/������B����Nd0�z]��f��Ƨ�r��I�(<��/�������n˫L� r�w/��7��E�}���w�*�9#>4"��x�D�R�w���{M�U�j�u�,k������Qf]�.X�������T[ION�SΦ�_�	�@�>������8 �ٙ�U�X~��z�$u�v�������ؠ��5��-�A�Q�a�0�L��d<����n��|p���Ͼ�㙍��a��y�����݁��6���hz�}/�#J�6���T���׀�)={w��x���{3��q�Ж�XA��{�5oz����|���m+S��ߢ���ae��Qɣ8��"�	L�TO��8�Vq���]<���]���*�Z'����*l�BU~���5�'#��I <��yߞ�O۟�?��'� ��ŧ���~T����1(?Sw`�X�
JH�����o�*Z� +S�t�����$�?���]�|�T.��	ͳ�N�6v�*��W�m�]�Q�v�G,rݫ��qK�ذ����{���M��Q����¦2���������߻M�2�A��[h��]H��pnP-��g���yi���H8\���&���$*A�>�Jf��Uf��2̧2�j2�"��������%9����pE�]T��k���*` ���T�O:S"vO8��JkaaaVp0��
U�} �̠0�y�Nf�Pz��8Zc��gWj��Sצ-h��2<wPN'��'� -~�"��1N����F���}Ms)t�Y_�c��ƚ}���,�-�VkQ��1��(�>�@���ܿ^��Wb������X`�4+�`P��T�}I�++�	d���"���g����m*���8t/H���d����T �s��������?��q�Z�d�wP����>�s�7f��=5�~+��߸�f7Z:����#��N��)�J���so�S��Qs�u��e-�7��a���oȳح��!�ٔ��W%����%Ksa���a�� q@)���J�P�]������N�C��սЛ|��8wY�6������!?l��Z���I�S���\���ڇ���'$����n4��&�:NR�Ƴ'nЙ\cS;����������Ħdy���29%���N)q0G�yԂƸ:���$��h�F3�d�W�����F�о��Bi��yݴ�J.�)7�$,@��B�Z���Q��lc��-����J&�JvD;�տ���ީ���H�JȹM��M���Ƀ��1��q�%��ll��`����`�(ڿ���(����m)���7�@]7R��#���T�a �����ⴸD��V�5y饐ID���tZ�T5��KwB��<��2S�G�7{ߓ�הS��u>��2�,6�����EG�}u����AI��UWV�.,��*�gAeV(1��/��VMF�NFn�O0X�M�� �ͣ�ͱ�F���ȷ�L�(vv$T/'��^�|�"���] -r޶^ǀ��h�s��z�~4b|UVZ.�6=#w�ckck]f]V\+/<%�[Һ*-�zD��UG��t�����*,�k'�@�Z)SFmU����?~�P[K��֛���6C1XR�=�z.b0ʼN#�b���f�"�K/(���|�0�6G� ��9��<�G n��� ~�w5�'ǐ�Y��8��K��"�8������.��O���V_>Z� l�B�}�f;JAJ!�@YI�_^;@�i���sq� 턊��������z����'�v�j�_&nL��a)qa �,�P te��bi���E�W��#���p�%o����N�{��C�}rZ{�E/��=�x�m�wf�z�}�Z6�ծ�!ݎj���k��j�*���t��O1^�~ �D /��r8������$��v���L|0���T&W�-�=dv�(-fj�5�T����h6]���q��:��e7�xw���1��s���pSt�x���>��q������W��T2lE��?>k(�-���e�<��܍���G���4���.�8�.M�3�����|�	��{�$�N���Nh A�JvS%I�"�Q��!Z��y�i` ��?�U'dX>#��fUR�*��_��C��&�$��9�����GEw��	��,�X�O}%ZI�&E�W�UpF!Bu*���������}�+��>����S��&���n�KN|X�����ꒊy�z'a)5�L��8O�0����7fp�>���N��?z��ߞ�l��aOZx�ڜW_f7_6���:ߘ��Rn��?c�󽁒�Q�y�L��Z�Q��]�٘�Q�3s�̧鬬Xe����3l�Ff��=��|��pD���3�K!�3D��[� � ȉ���%�9	5�3oZ���z),3r��Z�����H~����	�ƴp�iu�n�u1HR���Ur��4��ǟ<��n@�9귳���B�����U�Ϛ@~HS���$�)A�Q`>��H�P��z��ݖ}7��>͢���2��@>����G���Y��a���nT�rN��j�R����yJ�����K�c 8{7�Ů/ԌU�Uh�.��T�,�
�b�-d���*Vi�n���h~+����"99пK�]��Z��3���P�8:�8��9t0��b1vk�s�(y8q�Ѱ�x��P����:&>4�?=C03`���@ cRљ��-,mq�n{���b+��*��S�%"r?ԛ��^���u2^����->
�+1z2���ޭ�p�ĩH�����.Gq��ƺb�/a�߻�)���탸���	����ܝdfz���v��K�RL��ܨ��Jc*,�{�{=��8��eZ-ߦE� �I�q�k��s�OR%�=���3{Y�E����V�@:�TW:��Q͕���Ve��U"*���zA�h՗�i�}&-�F��]���v<���k�	q�/E�����������ʙ�#�X�BB�U��Sm5�XF韔�"� ���=�;o��?�[��%9��rf}��K��f����T�1v��t[�	�i�2e�%���L�wB��m�2����'}�5v��2���S�\���|� ��<�u�0X�>8��;����]��,.�����pk�~w��޾���ڗ�Ǧۓ�'���+S��t	 �@�0
��٫�i>5��b___�E������[Z���b2*3�զ�6�3Ūf ��E��IK|��9`HiƆ�i��́wU[;��3���{��ߵ�CG_~��Y�9�5�pDRE���x����s��4�ـd��ĕO��i��KG|�SHw��@�jθ�؆��~ED�}�3RFͯW�i;Ӡ�v{�;I��$RB�̓�S:�]e��9��	 �g=�E1*��M0�����. of��Y�|q��M���> �����'�n�י�Ѧ��}�E�j��n�7GwK�Ϭ�_#�F\��yD�%�F���c��e���ȕD�#��K�O�<7���������K��piZ�LԶ��h���&W���^�����N�A������9`��0������pQ�r0-�	u������ruDofJF��]Cc�����v�z��mN
�T��axŻ�wU�ζF=%ˋ�(A=�\O��a���u��X�/h'q^T�һmYU�◽�*ץUyN���g��*VH��cK��Yc#��A�Ú3�xʻ��&]��2�
vM�UM�k�r#9V�e���R�g��Tg�(��%	�y�xW�?y���0�����V��*8���>O�{�{��E�.��/a�� ��Y���f�K��s�w�FWҬC��A��V�h�<=l���J�9b��4����QJ(P�N�Rlfݿ^E"������Wz�9������)l�������,ɲ��!���Z�%Y;q�Zl�^��V���!���%�E�c��h:�]��x�ѱt[it�h�x$�J�x�����e�Ы��>�����g�2����û��?w��>+�o_s����1����W�p�>8����r���v�q0��~��8Wi[��yJ�Cۣ�QM���L�+�e2��W�Y#��+T��
�KT�њ�q��?1���Moвxl�*�(��!�@�����\E�MݑM_ǈ���=A���P8.-^7�1_�Ÿ�����	�Pt�f�Yʸ�����4(]a@��6ԃ�Ջ`q*L�O���G�&yx���_��T'%:=��5	T�!6?Bu�L]�s�f�!-%==->3+/��J.��攦�0�ׂ�V�I�������q������/�w���_�/�Zx�{�u�G4��m��?�6��X9�1�AH�(��a�c�l=�rJ,t�@,t~�2�m2�@wtJ�:�)�T=��R3��ԣ�]��N�D#>����;0��I:G��F�X��9�c�9�W�r�ۧ��\�(�WT�+� �$=4-*�ɴ�/ T�Y��ECIt�e�f^���3�;�O�@^f(4K=)A;�MvzR45)9)#!.�q�+�E�3�J7L�JOe�jHϹ��Qsumm��m���>��̃=U�2/���=����U�g���xx�q?�#���ϑ��9i�_Ńt�'2�=3FA]��8$��X1����h�u'���-��J�\���s��1n����(�
=�[���Q��(ti9�X�#]+�'�VA�=)>r�C}ʔ��sI�T>��Dtɓ~�-"��zj���4y+S!��V�J����g[&���E��,�r�Y�3g�����?L��*���k��~O��t�N�5'��?ƀ���6���O��S�nL������a8n͸�W�#�(����r���>Cx�v��T�k?���y(Lr��1e�Ї��2*��º'��w��-L��V������qNP�jW¥%�2�M?�yj@�tvx"�i�H]�Ŗ�
�\p=�� ���q�[��df�d.��z!�I��f(�=�˺!���;GX�l����n�8�c�j�l^+6Tʲ�l7��lf
�nfi��?pյ�M�i&�V*��&��'�o��&^;iƑf)mh3���+��"5�5墱s?�O��� /Y&�0t��}�����,!�@MϢ������Qg�s��"h�Ŀo��E[T��2t	�t�>t�r�!�C1n=R��y�Q�p�:��;wo/jkj)ǲr@8�,��FV�YGm�Z�ל-gi�х���7��2h?G��$���(gQ�d�n��b�]bk�TI��GHH���'�\�m�T�=z6�^C>R��_6��j
�:)��]�I�����x�2Y�����:+�4������\�y�U@���k���!�;��T�R�6��5݋[�9N�
£���gk��Ь�])�5~P��v\���ߍ7
!����P2:H����`$^c��m�VE/
X*�[\Rz�!ʗ�^���׮�<�Љ�/��.F�UV��h~�����	J+.�b\/��J��K���QH�y�	d�W�a�p��5-������ѱ��u3���S�k�����b�z?	��E��j�����h��#ʬ_U ֔�j�6󥰫�E:2A�J�m�x(�=�̘J X]��(�S %��<^�#%̝�m"��� `��;�J���1�Jp2P@�M|�X�p��@4�|��� ����� �ex0�����"��y:���1 g�uA	�9�.��yT>,�&GB#��e& ��Xt4��t�._з6�W���l#�� NH�두)�I��	�~<�����GJ�J�C�ļ�E����(��|�+!��D�=o;��պ���2�н����+�ݿ���a�L[/�@�F/l�:U�4�ʝK�j���@+~+����"""�"�����j0��*_س�[*蠙�{�ν�FE�r	"k����P��`�!�ذ���2����ݦ���-��.��E��A��+������s���*����v<�T��l���%��o�:��/?^d�P�q�w�6�p��{z����B]s9���B&=@�54��<����%$������̘6��D	u&�bs�b�2^c��8�W{bI���KF�I���9`�O��̂e�c�9y��3�.'�.�B��R���#V9>�ө�$�, �&�v/�M�(�}��	�z�T6rv��i����QJ3��N�Wy&��˞��H�������ս������o���e��u��Ջ�|��L!����߸� ��8�����Q�YW�����.5ev?����W��z8`�����=���#-��y>�`7�1��7ե���.g�l�.���)
�l��u죂�	%;jO��$�]o����)	0p��'�f$e��%��e���R�^�I�N�ss�\��GV�u�����ud�[�떐��D	�J�
M���=|�&.��PS@�A"ȼ��{�h�ic��Vh
�N?��\l�j��'|���*������f�]`�]����;z��Y�}�޽;hټ�X�5��Ȏ�ojq7]g��'qJh8����%|��#�5S,]
�Ѩ��\kG��)U�~�U���mD(��]e�8��#�m�f;4���jk���=�����ހ���l�T/����;�
���TZ��zۊh���C.	7^��ڠ��<�Q���J@���O�X���*���!�� �d����V<5	/��|�?3 � ƚнKI(�Ǔ���W���t���E�6?	��,�O ��gͮ$�P�.G༒-�hҦ%�à¸>ڗ�'��`�$3G�f�so�	@r�%��]����
4�U�!U3$J��^�R��z�>{ʖ�x�zN�q4g��P��w�{��� �i9iO��h��V�/2�ո��U(���ث"Y��:^�+hЌ8z�k�6V���'��Z���[�k(�X
��ͬ��ǀ0����֬���2��j���,�S��R��tL�R|%_/��z�\5]G̈́+�_�-h,/��Z�?���m�ü ��8�&'~]�v)K�H��ڪ�Sڠ��A�QY����h��4����{����"�d$����"��tI�ۇ�[���;Nz#.I��.U��R;
d6ț� ;�����[;N:�������+����I�
��TE�O��+�z�K~8��E�j �H�ƴ�eXD^�f��YGv��`����MV����J�3�K���:��	�/�����)�Lc�e�{\���ƕHb�~��x�R����V}C�Fv%�����S���.�e�@�a�r���y�U%�ߛ?}o�j,�ii�� G�b�O�.�Vv	�r0�p�iV�0��tE�B����"jAO�%��g�v�q
xB�d%�#��/�|Ge����}f�|P`���G&2���*���F�g�l��m����i�ql������
���{���t�	B�*�3��z�z!w ?׳K9ح�pb,���4V��d���7T��U��|U'0�:�Ү�"�L��n-:�5K��CHDZ�5���.��@��4�q�G�ǁ�r �(r��}��� Xw�Ո���=�襨�<��]FֲW�^����= N�ޥݍ��ey�g�Ǔ�����S�L��S*U���'�Y��%d�5�|�yA�yi$�t{��ft�5�?���M�x��{�^�|\�sx� vX����{8Kw�;�3z���~���^��qգ����{�\�m�I�R��m��K=�2�j���EW^�H܏�0�s���;���.�?<�H�3�W�ҪJ�4b�?=�V�vz�����C��K���J��]"ب�I8�ͻ�<�7�q�eb�҄s���r�19A��q �oBk�_g�����f !���n�+kȻ�+��l����-�u!&�Bg<3��M�n�'�]�cе����KS�M�[�7f��?�Tvx]�k����ڕ94q��=�5˙^�4I>�Z��ڊ�����I��CJ��U b5��C�m &��k/O\����Y�u#��M0ʚ�庸��V���څ8� i���D�h�����/�e	����W�H�stP�'����5�{���c��j'�dG�N��z�!;��##�:���\�N���ː�������	�YuQ�r}�)����/G�������߽�W�����F#^WG�&�PeA�������`�O���z��4y�?�~��Q-$��<e|��js��åR9%�WGP�鋐�eDر��I.ӵ,`!�_qԪ�3����<˜�[��k�q/�����ѡ����kz������=�e��ŏS�	�����,2�q�b���pp�y��������gV��X8�׵��2X:.��C�n�~�J���r��mŊk�������(ڠ�o�d5�_ˤ�R����������5�j�Ix��H1�U<(�Xe��ֻ�y\�|#p�UAG����}�I����|\����M,�q̯{2�-k�lcz�=�)�C%�<p���R0$�;�`��Z�\��T�"JiϤR<i�2���&u#�Ve (}*�,����դBN�իf�X֌>W�[�k�E��s{�!-�f�\>��e3�ׄ�6���4�C��3d�^� H���m��GU�J��na�l;)p[�!�`�|��i�\&����xD�j��m-?5ޫ�e�����lS�fG���8�T�������a��&"�a�A��6x7������R�L�<1aM���d�J"���f��Ao�g���3D�3� �S����ʔNz�ʭ&�s�d�g�HZ�I�#�-L���
̯m�܂� ��\��	Ԭ&'Τy�1Q���Z�;�ؤ�T���]�Y⌑e�E;ʟf@R�u5wN�[&ú��(�7��FM@�˯U��U�'��ѱ�U��k'��R�L�`�e��	�.(z����h��I��(앚�5L*_/ }:��<��������0�Q)/N��̲~�=
��\�F�<�H%kˍj�d�����-� uv�Y*�I��T���`��a�p�s��B�MvH��3��uW4	R�N��.eֱ�u�"d�Ž�}ƿfL�L
)�r�I��J�pb��meص �Q�;~eu��~�c�m��ZD��Z�篠�ԿDf�J~��wE�@>ڷ8#���=ҋyژ���ݯ%u?�#�({ˋ�ub�ׇ�k�`O��}�
7I.P�t��7��}�綂��V���_��0X�����������[G5�����PI%R���n�2J3��K$� =-�tI�蒖������<������p�����^�}���nh�:�@�!�~AD���yR��j1���ay%�.���;o���n��^:��)���ތ:�.K�u�=Y������vj��A�\�>}�P���nW�Z�u��\N���.��=���8�qd�A����x������~5�נ���.:M�aeU�(���(���@�vѐxP�p���6:i�9�yW��t�D��ԯg�y�����t����Ԅ�h��XKy�!q"��L��|�	�܃)�����Dc%,�6��Ւ�仾?#������`��G�zE�i���'D'�����)
$�lfWo6�|˳������MN�p�]_����˼U�2����)C��^M�k>�����e��S�S� ˺���̥e
��C�D���_��@�$v����om66#5�����]o�׼�Qo;o,8A��x`�����7q�cx@��|HK{��n.P��8��y,\6>�y�|�4ԓ���z{C�$a�Y��WVh�PO�� �n���.�T������i4��m�Ml�?��d�Im�A��������6�)�t!����$Z�����)�p�%��
j�::
G��	+y\����S����^��Yѥ��b|v�&���j��霣��h
���TT	A,�n)\�W"��dFy�q��4p_S�JEҿ�.f�^��}.�0[���-6��cɶgG`��]�n�ʏY�w�X9�1��~܏q�j#^���:���-��||�~*�asrQ���>��t�N~8��ݲ��zE�p��:�~���g}l?M2��$�`�-���ֈ0y~=�g�^��H��!����~*�Ho-������=�co���ߵV�&7�r�B��X?D�s�tU�^=(6ǄS�iZ���GѰ��������k?#g��B\�C��c-�J��Y��ި��3������S��\�޺�X�9�����H���7�s� ���e�N+�����Z�`׼V���yB�%�3�u��ƾ�R�B�_�M�o֑u]�f���>�пÛ�o�2�d��c�ʓ��d_���a3'�k�b��v[��%�����ou�th��?����s0�,��޺�lZW�<�����N)�enu��.�I�!k�S��B�7�숚�n��)n�dEs�����X�`�z���>�7�l u�9y����W���(��hus�?�Q��:<)-;���ed�JI�ϙ��0�/��� Tn5��f����sFe�ȓ �1��e}�����JH�| �L��eOJ� ��g�7>�g~�5�8"��|rd_�9���c�� p��nh$jQ�yܱ����AKjC��n��UE�]���G-z�#.^��=s����*��N�	.��+
B��﬏?xJ:��Ӂ���}	�G�\F�����B�CyGg��W������$�ר*e�\ﶂZ* /wfZf���J��Qj���j��:�(u.��?	�oEb��j�r���Y�W%u�G^� +o�F��;*DY�p�����u�
��E���� �-Tu����{�����n�D���8�s)�c)9w��VL�:
��������m�^�#�/Ȭ��������A���{�%[��o�t���85!$h���R^[JO��a���nF����!0�M�A^ٽ�Kr/.�y@�������(d��BbǷ��Q�ռXE���4�6��h�+:�M%H�cL��kr��=�;o�Ri��K�;9.�_w�/�w����~w춄{l���ޱ�?P�/�wRﵜ7��jt�iK��+��w,��z��~�C��������⾼��h������'����tVa����!j̴��p/G|�N<Ў^mR|E�C�}-?�z(��u�`$�(��p�b�^�Em��,j�v�fՕK�R̘N��ȡ��8�!��I��ϳEHPy*�'��n!�ޝ�&��7��T7��c�S69��E�ݬ�gx��[���܌�_�)g�Vy��켿N'���[��U��6��>�1'��;��{�NLu�3;�<������O{��$'�;N�[���	���lI:����џ�ODX^�Z�v�p�����:Q_	1gp�Dj�c�3�^e�Ф�S�RS�QRD�iC�3�\{�Ү�-búQl��c &��������P)<)I�g-��U�� bɐ�:�i20�n��]�a���t�1q��T�3^���N���[���RLX높�I�;.���8b����&�t�o�8��cd0V�z�t\?��w��J2���F�c���N�]���z�7�%AJ�MA�*��  ��0T����x�8A0��>,��9hT��U�D�ր��r��(��H��Q52 ��d��X4x�:ҝR��hs����ԼP���jQe�_8V�5(��<��0'_�M�τ�X �X�J�J2�ϡTe��笞���P�#�����hU��MF�;s0���-��%�aA�GH���g���_WDY �� c���|2�C�Κa���k�n��Xq�����X��t��iHq��	�Q�d�$n�7N���?h|bG���/�2���(҈.X� �Y����>�ds��q��S��'�\ᰴ���z�����HM�!S�F�;��RuV��,�?#���������^wz������b��xh=k�뭷�rGdm�`�6��v`&b�H@�!�c	5}���i��z�����LĎ�輆�+�f��Ê�8�{�z�Re|&~��&.���ͱwzM���ű�g��K��0���h�EP�q��]�yr��2x�86�	��`ǀ#��F�/��z�zy��d`pd��v��|�����Ǧ��4թ�7�8�j�~`�]��Ǘ������n����?�2����1���/����lbD��e�/�>���vO����� �H+U�I}����V�����=��3-���S�_����	�hx�^ی�V����ąa,�냜�$���-VQ��K'��4��%�ч�����"�ݷ�KT8�=8���r�|s����@��K��wi
��4�F'��s�MN�f���&��W����L�t���-]Ht�z�]]**��y;�t�%G��a�� � w629���q�*d��^�f�gJ��A茉�4{���ض���se�ܑ{�%������!5�t�Bā4�|T�;+�še%�������_�m~��z���;9ɻ'�2�O�� ��M_�� :T,���4A�<Hj�����^��߇��mQ�s)���^߃������HB�	�âO2��l���"��U�E;��E+`>O�F_�l+[�v��1�b<x��`�&f�:p��ix�+W�}>�rw�mx�o������,����O�������������6�[n������&j�.����T��,O�����4��뜍�#��E,�^5� (y�Q���vՕ�������s- d���%��NG���%m�t_2�<-|�o9V^���W��8<\�_��?&��Y.��8�uM�κ,���E�1�ċXwP�f<W��E��WK|")��KC*$���ܽ1(�ip�:\;;ʣl��K�U`*�#�r[[t�i�(�����q�d�L�����(r�4��`AI���������>�|�⣈#5�U�UR}����]��0��DT�_2�V'"?���w(����O	C�ES���{�vԋ
Y�`�����O�bgV�n��(��kwo����ZW��J��a`1���0�Ϸ��̼b��|���q6�DR"Łsb� �nU��_�(>�#e׫�}�/6�������u�������3�?��͹HZ5b�f�K�~����}��G	���F2�&P��aL�ޚ;S�c��\h��I�Q4<�Z�i�������NX�ݫ���87�&��A�a��``n:��$�4L=��o8h�\"�o�G}�Ԋ2�V����n?*�G�[q�����5`O���A���~���!�Ȕ�7�b����"�PunYF�qi����|��P��ǵE戜.�4��W���8��m��A�����.�C�c���O1��µ<M�{Z������b������#^$�f�'Ŋ�J�+�-��Pږ5�à�C���-9{�~m���Neӗ�	�ۚ��Wh��9��5�I��2�=�.S��T E��-��� �5�-�+�c��|�0敟˿��^���%t�&�0#��z�wT��ĕ�N�Ĝ�
�U�6=Ȟ?�W>�P$�KTA�+�L�2ԣ���M�ӸrJ.��4H�
vT�`~i� ���{W\sd������c�>�����Q6M/��c}We��&Q w��S��N�{� S_eW(��4[�k��l-��{��^z#�����L���
^M�]�#$21t���VI��d�$8�:��g(br֝x����&�3�/�S��'zJ�`�R0���˵�� �!k>(]��z��z1,����~�4|�O��G��M%�{3DP�9����r��Az��ؒV Ǣ��5���� )5ݧ��,�l�<�vݑN��39���Q7p��`�KO�N�����:#�:�Ƿ�����ԄԌ8�dM-�'���R��B�NG�R��f�$��+��z�aa�Jz?�=Әyr���}��m�tC��oYb�^�T�?e��)Itw��Q�,=gP�����\�����w��Di�%��b����V���{�@HU�y��2=��8����{6�
�;�fyU��%���|���� ��!>���_Ϛ%g�y���cRM�u�pOG��*�{l���ŷO>O4����å�k�,������ c!r�тW����&���{�O?aiĩ_5�~����X ��kRBT"�(���!D����a�j�&�]f<�C�@	��}h��BRnY��	�۫��a�ݝ�,u[V/�7��SG�S�AM9cz�|�@�d�`"8Т\�oU��R�@ J��k�� �n-��٭�����1w�����Q�T��f��������qY�a�a���ԯ���31��}��c����7��K�1-�77rvw�2Dφ3���/2�&Ta�4Y�;�D=S��;�������F�\�ݘ�&������JW.CA	C�
Z^z�ȸ�`��ێ�����K'�92�l�v�MB�P���۬�Y� bWпHv|�m9EU�k��*@n#v:$��L&�L� �<���8��� ���~"���g�p�2d�Y�(�RX9L{I�J�sVll����M��C�x}��$z;��@�h�Ɲ��A���c�Ò����-�[�sm�p�`�J�=�W'��xŘ����2"I+�{ǒ�$�R���EDH�K�˂�K7��iӭ�P|����%-����Z+���-��Ǔy�w�T#��g���Dh�������H~�,�;����������iSK�~��w`mҸ�H�G?�`�`���4c���$v}�M,�����o�^�Ы����P�h�{ܲw������?qnv�ܨ��s��n1��+7���yT�'�Y:p�v���8�c�*��yl0�{RE�{�*�/
_�l`�g��v�^�z=�d��%�(.��V-�FN(�v�4��>V%?�}�{��Q�^�����Vl7^:�-�b�����RU�k�����~;�s.iX_��=<'؆>I���T�������2;]��5�e�Q��૾�>��/�y8��
���������g��A�M�ȗ�����m`��ڿ�����Xp���� 	-�3f�}<�SJ��'��xt���QI3�潵��x'�P�R.P?30_�=?pS\5�vb��a�hg�|���dc�{��)���\Y����o؋^$R�I8��t@f"�ђ�bq#���u�X��)u����i����䘬h*���aGB*`����I49��/��I��=�-�ƹ`VD��>����V���ڗG���Gjߓg���m?�~�%�������?��G��\3]2¤���/�zha �'?��)Ic����y+�^��<�mӨ��PbFk�y���؛�)�k�w�K�m�/�^Η�Mm����_�ջHd���������E�O���z�(��0չ�
�\r�F8�����ZL�:��o
��^��-�D�2��UܹH	�	��a���'@4�����1�`�����{g6r4.��k�r��貞yw>��87���ƀ�̹Eޛ���?� �����'�Ą�� �\����9޳�NpU��<!A���[LL���T�������c�#��G(�M�B�X�6�tjR�$��X���Ro����s����=��l�b�]��^��|�A�b.�b�~�M��t�����FV��h��ڟ�]&�>�Đ*m*�5?���	�&��26�_}R{.�.̓���]-RJ�5���/X(�����:/z�o�w�n�?���-&��ڮmt�$����8���D��^��kU�۞���C02���F� ��#���I^���@k�H�x���f!���H��6���@
]fQH�K�-v�	7��W:!�l��<`���A��T�����K������W(q�ފ
%,,-r���H�����*/(��ћU�w;\;j���6�s�)9�g(p�A�p��'v�p�mxtF�{xjx�U�wR��q]�r���w{sw���f�ɮ鶃���6�bw�|ͧ	*>�qYH�����ڒt���ɠ^>�j.��q����}
,7���i�P ���'�UZ���ǀ�0��徉tNݿ0�4��S@�J7^��"n��A�2���<��̱�C2:*�rbL��@�C����\䜈��=�8�f~�820M�"+��Z~us������h��������m*��%єA�:xp�"̠���Pt>^k��o�sj�.�SIs�J�;�*��J���Wd��ڹȀ����	�N|V�E�wŶ����rW��0G��A�#��U�w�$��|t�q�@Y��m�XZ��+0�$��ј)�"���ß�+\
�uĭ Z�4�v �:o9<9����Kp�2CY	�Q׿#��e�?m=���f��N��o�; ����$&�$f�P����(�������POW��e�9-����-6�������2��[��NV]����Z鿦8�,�n)�Xg~k��Ŀd��D�{r�ږ�
��ϊ�ƶl�����-M��z,��\�s9�%��G
��&)Pw6s�6\���:x�Td(ڲ�XOҺP�o���Ǒ<Xb,��D�"k_E=y�/�Y�W?Q��(b)�����k�g,���T՛�z�r$����� �v"a����C|D�ݵ�|�Q����4*�<Ej�w�Puc���d������?>�-���Dy�؛u����<�ױ��&R��W�c��[O�����1�B���=��+ed��Xj�dJ�����觙�[^rjɗ�)l���6u��.�$B�o���\���n ��C͗t��(�h�� ��Zښifl�W)�y�H&�|��lI��D|�`���i�`I���5�O�c(��
�^�7rٷ�k�԰I�Iؾb��qa� �Z�~W$� )	g��!z���䃴���xI>����Y�v��fIn)����L�Lq���G��o*0:���|LbL�=Ƹu�<
��$iF�Imd嘒�I�|�7F���=���F�E����o�q�z�H6p�(%hSS��l�����['~�t�d��I6'1Oꩼ�m��}8�i��_��$���a[�%�M�2AF�9F.@��l�I��m n��- ږo���ʦaɽ�`4PCeC�9�������H' �{F�V����:�ߟx;�2���i"T���eVh+���:�#�I��f>#S�`b���a�Ff����QR�G���n���Y'{)#��gJiРz9�bV,G�������tC�o�w�>�
�1����� y�hT�� ��%��3�䥟���ѐ�-���S+�},�/��������f�Mod�.�sT"�h/�/03YF+W�>t��g$-��f铅�'n�]�g��0�^����$z�Ρ��ɶ8� f���@ @k��' d �PD�����|iyi�$�W�|��I�
c�qݩ�pv�����PUK�:l�D�᦭��'��K��!n���@�$��Vg�szt�E��{Z��pL��{��|��pOO<��#u�ϣ���";r��=7��փ1�����Ƙd��y���wyd5�m�P�0���W5wL�j?�"�=��ٺ�mY%�*���)P��������,˳'yz��+�KG��y�鿂�N��vB͏3���ю�?N�~#ܽ���7����ty�g��B�S��&f-��9����%s�n�&HK���akF	�O����Y�G�\��c�Y �(N���נ� [nW�*��Y!ô�4"��`�1�Y�|�N���'��qڙ%�j�/컎�K5�{39��{t��|���H���0���Z�z�MP��|�m�w��2��9ľ��w�ox�{�|q���&���:I�nV��4���{=!i��y�/C���>�u�����G2/�5����Qt��%�?jJ��l� �F�N���c3�u_ޫw�e�2�� �����2�]�N�/�����)o����qp̯�P�����aZc��YzB?���Q�')L�����B�{�+�A�M���}	�[Ñ�Q�&P����4I����:0�=�]ӞWm�����%Q������wټ���X����h���!�2Zh��Q�2��̂��ֲSj$A��23&�(���N�?����H��i��O3�+
�3��(|�,z�"����b����k��c(����i@�Y�*@WF�ڻ6~�86��h���A1V���Cv��x,�pߗw
��S�߲�~����q��A�-�%�����������5�@���50�lYRr�M������M��MsC�>�_О�3ٴ[[����9�`0�S=�$:nߢS�:�;�l߸�����x�����J@:D�rt��$�o2�kW:�30d�iߜ��\b�����>C���G}�T���v��4�(�OjR&��R�ːz\�(�Sϧ
~�CU�7�N�M1�.?�r���i����L��E<~hn΄c$�����BvSL�t>�,�aQ*���~l�9�u�*�$"]�*w+��n��T�����P:wO<��S��/���.�.��{֣��b �15LD�B�`���"Ǟ&�5?ڿ�8 ��Tי9HO�#���"9�~>*d>�<�r>Tzs�4� x�f�ǧ�XtFw����^l+�{@^��]�T5�z�"'h]]Hj�<�E�ø�Q-a0aP{�6�B����Of���u�6H&�K/]��]�69�y"���7�؝�_3��9�}���7��;�p��M��
W�<�SU�x���dov��՟��O�3;��S�b�^e�T�V�R�Z>�B�p��ĝ��&�R�`݄��8���q��6E+|��]+P��e@)��ׂЌ������F-��;����΁/}_8�#?D�*�˳�)�n���U����gS�0V�wի���<19⊋8���xx�8�ö��s��O��n�52҃#\~��]�Ͼс)���3��aU=���̓��
#C�]k5y^>��"�b�����3��m��a���	k�qk�7:	;��;:�&o�eD&A��X{�?^�|F�S~�}mOَRJ�����/���w2�����%�x�6Cc;�"8tt≺��/���V3�R[���(>	Nȝ/^ko<i�%����8���{�8��ɝ9jw*��Χ|�`Y����H[aZ��)�����@k�Ϥ�L�z�8n>a�8b��u39۸��٤@5߀��%���5�����Ѳ�?���"Fx>C��(&yDp��M�2<��ID�b"+���5>�`�<^�@��^0�<����jp˗5iwO:k۬��:
��p�0�$Z��د)P9$�JE�*��p &t3X���4pY��GV�����&��lz�#����kz1~kS�8u,֩EL��o��H@�uU�]���:mT�#���n�%�0�,$�K����#Me<�mO��[ M��̞Y�4�=��Q��Mb�#_�S�r��Tg}S�����O����J'��-B%>KH��\g� ��q�����҃Ka�$C*�T������.{_o���.���"G�sd�7�bW�[n���v��]�e��u/]'e��1��/�;�+�ߚ�?�6���=����!vݖ��s�+v}�kws�J��u�x
����w]�znk��:DEa��N���%hѪ������2���m�����1T���NG�e�y��:�E-`϶?�å%;�wKhK1�p|V���Y��;<�	.9>VX-VްB�8�| 4����;C�-n�
pj��9Af#J�F~���� ƨBa���=����Vv�4g�^��r�Ϟ)拺�۽M�~����U��-���t�/��;2<Og�!�a:�,�hI�5��#w��1�,��p���@0�.N��#��.Ij	;y�����{�3N"s-8A�#�r%��q~�7�~���Ъìd 'jy���Y.��sJ@,�TA�H�*��� C�#��ېWE#D�`nG���x��b���T�y:�T�4��u��ѴX|V⇙m���fV���Ѳ;�f��E���~���mDN)D	��Q��q�.��(����mG%������S��iq�+G��z��i��������cð�����9��BYLx ���^N��X��n�:%���u��-�M�iT�����,	�LV�o�_���Pw��%�7����|쪔cO��N�طx�yyݍ�]E�"BY�ހ�@�j=�skIC'�	Tl ��������X�?����z��F��F����
�#㝚��:�Z���օ��o=N���3~�aUck1][����b����Q���MWeWzʨ왘OXX�gf5���|ʩ-�q�
�I�M�WϘ��`������Ƣ��kX̭�r��	��%�)���V���w�`�[�~��4Hnq�cU"�`ca�X+ݥ�W`\��㬯�u�_X0-�I/�ӳ�o�/N,�M4�,�H��V���*ސp(��{A�g���9��o�L�6���q}���Y���/�Y��7�x4�6��B���jb0Rڋ��P�ڽ���U�ٻҶC��ȵ�n�V"�e=�t��D~đp0�C+����l�T4_�i���)J���U��1P�*�G0Zuv� �&�)ݰ\��A�nR�<B���|��˯0:���T��I��6ƌ������sq�u��hL��a��d�.������?J�0�n����u��>�g<7���eN��:MIk#�����9ӹi?	�̌MIjgb�Sf� ��~��H�[�zx�`�����L�ցw}J}�Q�ҘM�`O�IX?�B��ߙ-�����Xh/Z���,��(�d��^�ZA�̗̍�,���4[�8�[�E�'E�,Cq�@�?bF	^��W����bZ������Q<ꐠ����� �a�FM��������W%JVSg�������~@M�j���٬�T��n�=w���kyZ-}��5L�?�� T�t@�:��)u�2��G� ����H{M����\ވF��9(��C�b�Jt�b���c�&c?w��3�R�NS�Ǖ�#����QYn�7uؠ�x�(��Pj�3+CB�),�T���S߰����
+�m���I	����w��@U_�~���v���J��ܾ���Uz��妦ߕ��ոJ��f��fL�����
������J���D����������4-��4�����.��'h|�#2�n����~y�maȝ��4Y��׸�?���Ӽ �|�9��*����cP����2P�B0#��_�L�k�b�!	�ȶr ����������8Mi��i=�ʯ~t�1�H@08��p�|嵉@2��@T9<,"�p�}C`��˄\
̤� ?`E�����PEM,/_CU M�6����9A�ⷿJǯ�צ�-v;���D��3_���t%��J�A�����-m���88����~ܭH~���``�����S�˶n~��&{�ݐ�̱\I"����Xe��$�H����>�Yg�o0`�3�23�������|B����5<b��n��8��ؼ�M��ތ�lU�������y9��0��X�����w�]�� cl����Nh�������ٙ�f]FO���<�$->����i�#=��B�"��Sq��]���������xhBF��/���u�}=����*b.��}Ѹ6�qs/բxS�S��Oy@$c���A�<�\5�^%��L�������NT�_L�q}i��(�"υ'��=�|�̕��� �M���8흌Z������F0Ťy\� 邑n'�?��i_S���S���#�OZ rU���;����>�H#,ÐY��,U���k�.Ԉ��������.:z�F��4t+�7��P�@.W�G"�
φQ����J;�"�S�4Z|uN�S���Qt�E�V�n�Pg��ٞ�-�N�ធʩ�&�5�O��*_P�(]�{o鈺��'�ߠ�>A��s�����2{���(`���CwJ0@��#<:�U�S�D03���1��`���]�I7�)�IW~�_
���%46�pK��xY� �۰����g��}��4��Mt��۪{���P�4kq*⤗��/�$�A���d��޳��8����{����T�H8]�H�������̼��R_���=�dÔ<��ײYW���䴀�Y\ĄA���V`�7ب4�3iܹ��4S.#?��=�S Ecޜ��Efxc?�D��x&h�h���`AlY�n�ɯ�Ҽ��e��y��W��&r���bq.��oR�,����U�i8ˁ��O9��?=.	��H���UEc|���ôFbY�����\�d�r;/���YyA���
�z�����tz*E���2��?�z`l	�$M$���G��J�.�66��I������u1���z=�Q,·5��-0��D~j0��[���A���%�vA�� �+�^�,%�ʒ���<���^��Wm@�U�
�����8*��o��$z��D!�� (�4�Li�3��%�m���$��?��(ƺ�} 3���{�$���#%���7�(!�k��"t3�sG۱����c����"��X�Y���8g�F	L1o28���ZY>o
�+�0����F|8I�ɍ�FN�Q'���\P�w��9S��ǗI�!��enI��?�7��7f7~�Z(����k��8��v[��V�v��^�����P������V��7����L2��'%�8J��Jh9�@�w�/vy��r<�wy"g�X���J�9)_ה���$���0�a��J8p�4P�����ּ�'� �`�3kn|
Q1�*3��u$��#F^k\���c�.�x���+ TH��iH��F�4,���84%���s)�S�-ZN0��UXcR�V	�@H��&�)V���8�[���خB�n�`d=�vp���E�R��Ze��Mg��������ϘE���p��[��ǲ�ة�\����lOv�J+���y]���`-����8D�󋟇���R�$��q0�q��� �g���E�Tf�ZEY�N<ux�+���r�ӱ�h:�!�j:�^,˟�h���W`i����Nw�i{��ImR<�dVņe#=�f��M�뺒0Q;��*G㟸��Lh֠B��'4Z;�;��ߟ<��c9�72�),D�+r�Ik�Z�o�QF�'X7���/����BQםs1����^� Ʋ�J�Tj1(
&� �)��-�VV�?��{i�X$����>�����;�(�4Xh�+���+����4tR���mN�Nb�BN��[qIo�)dÔ^�!����R�-~J�M��P��#,4$T�`�]�J	 o�c�(<f�s	�%��I��?F��xý�ѐ�$�s�.��3`0��$�`�p�%��U!����d?��_R���VO�ٸn���j����,�7%^�WZ㫆Sd��Z�>ٟ��E�]�	��t"�)K�y����p�)��쟖�d��N�	?I�nl~U�r3�H��i�ш���0�1�E�o�Of��t�����'�oĠ{�7|���=��M�r��:�/�cM�:Tr��=���NWn����#t���߫h���*H�pOUc&��R�t�����Ɛ8o��,��W�#H�:`���a��[<0Ĕ�eqhZ_�K����	4�������翥�gS�a� *Q�Z�iB���n�el������j�.����2��p=�P~�b˂׍������U���)�d8�c�tC����4�n}/&��!���������,�A� ��.��m�m�94uVꪔ�\7c�_����~]��J�C@hF	�����gŅ�,���JO�����J4�\^/��  Y�{�y�+�x�>�aM_��m��k�ɮz�T+�4���yHE-��wX���B�ḍޜ�����]%��Ij��LZ��34�rc�j���<L��6��аT &���W�%A[�vƋ�S0 ifч���1N�����u�>�FX[d�zj <��@��D(���: ���<��y/<�Hw�b�"���~�,�W��)�����S�nA�����z�Q}س��Al`,߯$�{,�9��Vl���r:h0b5����# �c}�c�^y���X΂�m�����'ݴ�gwW�5�@'�-�Ғ��4S�`���< �xP�7>6����<���+k�8{��P�`�����]�#��ZS�{��Nn�>����%��^Ŵ�����0o9\���a͸�����?�����\Lj����;I縹��_�Z���j�@�,58����`2n��^,:������O��\{�o��a��6��mQeݖ�@͘��Y�:�k�ȿb��k���l:ژ���%�N�'"{փsŵ;���t�*V1�Y�������0q@�f���3��y􉭄T�F����Y�g�};�\�#r�k�#�o�"�㔣��&�۾�	]��gMI�/��?�-w�כ��"'G�݆nG�rb��!>����^��n��C�მ�����xP�3�x��Q[TDx����V1��Yg�����C��0	���/�A����bK�
%y���z<�ފ��Ͽp,q���y�����T��*LG�xo��Y��ă$�$U���W�X�}ed�s�y�|��y@ɉl�\^�o��򀂋��ccA*b�kA''��-���+%���>.�����O�F	mW�7�8<]g�˓�B':����Z��O��o������R.�^��������e/c~��g�&cXmV�̧�OU���=�DJ@����:%�H����АQ�D�BM�������Q��to,
xPh��JR9e��U���or� ���e�܎fS I*DT�C��J=��0�4�?��, L(O���D�_�`O�/�ũq9��0`�%�0��K����'Q#<��_Bh'��_mp�5��<'�Et�ٷE�`Mj-����֣�,� :�'Kˠu���=ݭ��1/{��eP��$_�¤���ڞT���ub���}�Q� F @d�«�ᷕ��
j?�p�6��+a{�
Z��;Se�q}���#k#5,���gǳ�I�8N�瑖��J����ߜ���������B�{C�;�v�v�v�F�{��Lbn�w���/��m��m��B��B�9g��J�Z/�2s��#��vzΌs>D��ٱ;M��Q�e�b���T5ũY"A�r��"�ѱ%]�3 ����Qt�����~�[;����tׂ�M����P�%�M�O�M�c�0�0�\(ȠLg17��c��D1L�-��^j��.��jmYʚ˛�-Y�4$�X{豂���n��+�:���!��:���K�J��������;�a����>�p4��d�N�3|�QX=��p"E�,ɉ:����p(�)�'-�I�ڙ�+44�"��-���c��o%����y�A�EdI�!Ԡ��������c�BW���_�"lVi�
al��:5��Z�l��b��W�S��%��M��[J�Z�TZ�Uj��*K��8�tA�M*��<f��*�䛜��p����L[�60��	HĂ'a�SX>��V���(�!�O��$���՜ ��ћ��e_�D8�Z�h�j8%m�6�"P����}<l	/�8P�Vк��J�ZJ�ѵC�HS*�\(K5
P�����y������,:k�j ��@6Z*���W,������=M �������W�Ĭ�yd�t<r�<�����W"�G���?��U�+j/��fc��u�Ƴl�&�����z��
����߿''?S,6��ҷy�JA/:�ֹ<�ب�&1NJd${�ѳk������n�So��e{�T�{��*�?$�pV�|K��_#c�;�t��/u��a�#u�1u�@�W_��\{�ή�A�H=��t4�/�NCSS��cڭ�z�mE$DB�J�H�F�C��H�T�a�0:G�`t�%��Q#����������<�y���s�s�������]���m�_����^�D
K�4���ܯ��߷Jݵ�߮z�����V4�������n����6�x�S�w���l����k��Ք��-��a*��o�7���}��*���{DI�v̛�EN�C���xbVzVrp:@+���/S���+��ydB*��KN^�U��l��׽�%/�M�Q# p�+F�/��2�a���z}i�����7Q�E�G*�����Pm���k6o};6|�该�c6�`�h01[���t����+�|Ns�{#�q�q?�4Pr�x�#!'�! �R���j������T�1�hKި�-�l�H��C�1:��6k5s-l<3c����	�J��Ã�+xD.`��ŦJz�f��e��K� u݉%8KŁ�[@އ����	��{}�V�4&{�*����4J� ��1��3ߖ�~���u�0e�ET9�m*�9X���L����b���
-�Rڲ`h<0�ڰi��w���)��#�)G5+[ۓ�7=�rT/�aw��;?��v2(�;\0r��O��LWo�qz��ڵ����w� �����a��w5�ё���6�e���*S"�?C�>��np��_~�>4C��Q�1�̞�]�*�!w�S�v{��O����A��)��Y�s[����@X��Ǥ����;P���Fɸ��9�3bk��g`94眰��M�	?�㇀��f;���_#x�ݫ������/�:q*�K��御��_K-������]�(X��=�
�]h�¯￩�l��l�S��ѿ�͡���;-�L��$��ΗZс�J�ţ�v�ha�l��n����AE�����l�E)>M�es~?���CS���'̧����chw�9���޷HHc��R��Vi�JI� �cߩ�����p!���.8v�$�>����D���G7ۛ[
�۬��ڣ��Q
�#��k�^:��q�?M3&�3�g��t3����?�n*)�)��)ԁ���=���qbm��pz����?o������>&{gz��e�p8vT�yX9�"x8� �d+��ɩ@��XA7�!�1iQ�.��h�/jHciH��JU�LU�f~����4�n�K~��,I�v��W��ZoH)X��đ�[Fa�>ˊ=Q3�N5�<z|/�y
.�J�C�(,0�챙B�k��y	�SY~e,wV�	��Q�ːW|8�;�Ĩ�d��,�u���Y5Y�S����6u�X������f�x)mz�f�~$lI?���:�?]���?�]�yV�a	�#�����9������w����+����&;0:gd�r�`�������&�@�lʜh@�Y���^n��k�tBIy�g���^��b��g�i��*]Q�=K(�,P�U�EFd �������������va[�'G���h�
?�������P��b�/�k�C1'��/k,)��*8���=?�차tM�w}�{���!C��� �7�E~��Uc�H��������)+>����×��Y2��o5���`.����m!
�G)�T��U �ڈ���1�=�A@�Wh<��6�Kmd��:p���$`��[��'W<q�2���yr¤�������6[�	�B޶�I�����AWף���?�c�b�'�{僎�*{\´쎕H�9����M{���f�1ב�����ӝl��{�������c��w�����o�r?�R��K��w��:�t%n��Fzx3�qq�$~�4.���,op��ҜF�4�5b���2��O�������M"����/\�1�d�W!�Ԃ`�ddT۴e,J��-��� ����@���<�MA�c�>�����$J�~�"�t?�D'VL�:��=��Y��Q�1n!3��#�C@�$�OY#D���XBr�$�.����;�q2iM���t�sFj|Z��b�{8�8R~���!��9�鷓��¶c�p� ϵ�Bc��Xb�ßZ�4�� 
���#{K�6-���D���9�$���,������~�
�B�l$���ٸ �=dθ��{66}����, ���M�pKH�N�����v������s�ܮ�&9j�>���ĠPOQ(b�'1��ܣ��|l���~���^!A3����\�q���L���/FH|�IL|���v�M��I���$����]EE��ȹg��˸��[VJ[�w���Θ|Zu{�T�R=���H�8��_܌^���$�X�r�b2Vu���E��K��}�nd/��i��=Eפ
<�FK��c�o����æˢھ���y��4�Y�o u���T.5��/T�[Ź/u
�{^�,R�B^T�>�Ķ@�SS�_b�̧�!:u[�������MZѥW� �[�&�sK�Y�2�70(�����6��d��c��5?,����3�?�i�v��Z���(2�V���c�Tlq����r�`���}6�NG4�����Z�0�u�+�s��DeԔ���n�D^3�Ս���qN6�Q��FJsHIbeC�t=(�@�.7��W,�ӱ%�䜼J"�.�� �5}�d��Vǲgb���ZauF�e��*^<���� ?a�<\n:JN7*l:*�������D�׳G0߀s�;���^t,��Uټ�������&T��8\��h�D(?�nD;���fs@�c9��*�<?�Z��8�J���>�p��	�Aވ����V��'fژ@��{S�Ie��*b�L2�
��N
uk�6-#U���I%�^�1�Xۜ!w�PQv{���s��E���!��9�ź2�vϻ��G�eA����U��u��bȱ�(�bO^g_-t��3Jq/IU��<&2�X'�Gxݓ�4(1��Y�w��H�`V18-EK6�7�F^%����?QR�2�;��'^)���7'+f�A�`/�Yg���T7w-��ԯ���M�ޞ7[SrqS��Ёj�O���q��ŝB����b����Z��8��`_n�1�\Vu\��K�Z�{mU�-Bڲ'�Zv��b{8��Z��3KI�b��K����R5��i8��P��}���jSP#��z�o�MY{��s5Q����RF&R�,�q�*����.����Ųj�U"kk��
�e�㿗�҄1����ZL��t���s��ܝw��t�[�N��n������ƚ�RļE�.4[Ƴ"*����8>�� �W� ��g��ś�%g�Y@S���+0�<s-w���
�Lv�ۉ���xޮ�����)�5y��E�����T�ՈYR�W�a� 55ZZ�O����)	��_݇��$J��{,4;}o��2�r}�Oꍒ4h;��"���|q�w�i縩��o!�y�����`�Q���e��טK�ٟ���W�-W�w�X��>J/.:�4e2e�kdZ�8��zV4\���^���U����k�Y26c�7�z}B��*�=�Ě������ס��WQ5d��
�
�\}r���N��>߾|nÄ�d%G�h��񭉟�89��mG$�4¡�)�<D 5yfkb�r���4�e�����xar~b~�Ap����;[��e:c��Ý#�l�;Q�˨(�WcA��W+ؼK:��Q���#�fY�7K�\F�/P��%��U*:��UW�%���4�l;�	�}�X��"� ���>�;H�Z7,��P�_�̩\w~�Y�L�C=��\T���8$	[مGԎ��8�f��dL��>�!���qP�׸�FM�'���4��;���/i� qFct��ҧ>��������i,��j��o9o9��6n����~�d��R��wO������v���se�~�����թ���ߥ������4�k��F���K�]��Fa��RN� �S�6�4��Y�*���"*�F
3�:G;�?[�h��7�5#��/�x.82h�o� P0��~Ic�&��<����bs:�����@;�����K�_G��|`� _~�>����}&�k٢#���T�9<R�G~����Rf��e~V8'-�;��]ʬ`f?uC\ɜ�}[#� ��}��k�U�b���@X4��n]�vh�S�UL���,y�
��p�䙾~WE�3���&��M Ů�ͣ?�r���2��ǻ�G0��3��A|@�� O�O�/d�L���Ĵ���۩�ƪ�~�����ƨ�먒������XS�X:Cr&SjI�Ʌ�׫���K6�Wf���C�tW�����TU�̨�صڪJ\1!��9y'��q=�,�6�;r�]��Y�w��������oH����$�(��{e�/c~�ۉ�����$�6HR�n'��ua[�y��,�qE���)>��.�R:�r�Q�,�j�Md�GC�m�n����Gu��l�a)�\��G�H�K�����wn�[�2iU��W�;{S��v����2;�nR�,]���^�[���Ҵ�W�q"z�|�8�u�3�q������֐C�=ih��J�q6�W}9�Q)U�dk���;tzr�-�	�Z��MTb��`�Rb��)�-S�N���W]����ǜun���ML��p�/$��c���[���s�¦�[ȟ��?ؼg���p�Q{���� 2gUı�����R�����Zɜ��u������_�d�r�/E������_�G(<C�>yv��8�0&�q?���/F�dX�T��n��$15�'_��W��<�s���C�2�Ǉ��o��yNNT������G�c�U�t�y[5��~���ߞF?��|B0��I��^E��4u��B�Q����à�d�m�Rݏl�|+��5C�U�!ո�����PM�[��|@X��?]�=4�	u�T��$�d��g8t��#�;~wG\�^>�h�]�uB�:x:��bKw�k\2L7-���%f��!D�w[��5$�B;B�[��a��4���/Q+����Os�R�e��IΦ+��0��Ն��pF����\�H�,�'��>�AL9e2
S��	��)��Y�GJ5�|k����vhCi�F�Yx)6kzK��߮ɫy���;<� ���fQq��17g``�il���"   ���Bn��?288����i�E�g�kY�����K�%>C��m�E���/�P�74\$g��,��N�۹�����z��1�V����R���ɩ�W�:�ΖQ�M[.<j?�2��E�2��Sr���(д���vzZZFjN�Kz��_���%̽v�uq1�������������o��.��n���{��/��7,�N�Jw���6�m?Bo\�f�|F���36��ǧOm���*�O��ϓ��앁!�Z[`u�}-=97����do��>?*`��1�\�D��,���:00:<64_�hc8p,���$��bVq����d�B�+����.ԍ�۟f�Z�Gi���^��~E���~k����ƹ�5���Q
�dK�,)�d�����&���uv|���%K�m[O�#�f��8_o!/��,0nO:��ͮO�<"���N(N�К./�.�.FM���E��ch���9�`�1�r��5��֞��٥6;*��Q��R3�q�'ɷy�������n���"�|��pk�N���~$�ׇ��>�+�$"K굌��d=���
��3n9Ft~�Ed�UL�,ٻ������@j���i��i�u'����G�.ڽ^w�x/#�g*�.�����3��LEO�w^���G޵�y�k�*[j�����ޤ[Q���������֓Z ��:�[0���KӌW��e��&S��?p��/\2��@�Kt�u\�6�j{�s��|m�;o��M�	���?ij�Aw�u tىq��r�����P��Mo)�j���r䧽?�|E�*�6���г�þ�������$"��[<q�i�w����U/�[UsrY����?�rؿt���ms�8�%{yg@��mu�t�h,�����Q�<
[�:n�S_���֌�0ޔ�}��b�؂�1��x���&�sU�k5����8�Ⱦ�NP����O��}��b3H�w����5�e����*@����c��X�>R���;�ә΅�e�%��'��񜤉�2�V�#{�����dw�k �@D��>_�	��n�p~@��0�^�@! �S��v �1!�l��w?���������"�D�X�4��5�5)��k�Fz�ٲM�u?�)|W�G��l*!�`µ���������=��-{]�E���!?�R��ʰ�ny! $|�����Y����t|Z6[���i��a�z�����Hjw�.8e�Y���qH�۽�������R6��h�.����`�t�|��	�w\Ә�L�0�Ҙ��)�iH�xj�����5����$���ރx~\=�M>�<V�p��Ci/�F�?��?�`	pt9DMg B)�x��pxTUC�( "����e^q8�s�h!B3C�؜0V�B'D8���� ��M�Q,��R�KQz
�����<r�Ir�
VM�Ι?��C�F]Z-_z�R���$hG0���	6Ş"�p����
���7�cK��$��<��0�5�p�/�����H���&����*��z�Uk=�ᔠ�5��$�����T��BF�f�:.;#�����v��Â(tx��h�	Al$�N�Ж+3l�
����ci�y@ۘ��.d�����F{&yr@)F=�8E���Axqy|~|�jW��{țJ����7��l�4*��	����aa��K�����^Ѥ%$'��������5"lRR��B|�bl�����z.󣒠�)�;��4G���ڀ��/��V^��k)Di�������3�Û�D�7�e�Gˆ�M����fz^*��3�p>}rP��P�����;u>3�7���Pf��Ͱ`g��MĀ���n���|����ug�EXc��^ShT*�Mi�bFJ�jx�q������j��Ȓ�l�������ŵ��v�i�d�\ы�3�a�������ǀL$@��?��KH.��i΃�0b"��4�Ս�]���@�2�_(�t��a������͠ӡbd��]$
��G�	j��n��n+<	�����T)�K���z`/�i�΅^�U$�F����;;��
�P�ʄ�i�~NIa;C$
~�%�,��VM�����\r:�k�P͏��b��*j���-�Tͥ�^�	���( ���
FbX����m!�6�̸�4a��|��rk��M��AӅ�1�zhE�����i�ސƋ#��ex��~������7�)1Q4+����;D���oѐ�?W�8w���nq�NT�Ɲ��IA��wA'e��t[��B�\�@�����QG<�7�ڌ%�$����\#Ft�n�A:T�	}��w�)C����3��d\@�e���������]��X��s�ЛV�
��A� YЄ܏�L��
dq���0��0V�Qc�4�*m#�"������XX'���8��幕��sl+�" �G���,j|�����;HU�����O����DWf�
S��a��\l@�J�j�׎�vdj3��@�_^��9���y���3�WC��+��U{A#Ib��5�3t�*�[�Y����Ŗ�`���u��?R{Y�����Z��Q������xऻ�If~B���$�&�$�ֈh�K���J�WO*���������?�V�||+d7yd{����a@>��W`f�c+�aHb*�qz�(&>f3�yCC�d�� �9��l!|"v�v�M��r��������t���R�$M��XP�����a����x�8���B��ul�,� ��o� @��p_}>t����Y��{v7�:�sR@���V9,�-!+���P�"�ޔ���@kՉ�O磑�U��de�B�ߨ�h���ʇ[mYҕ=֋���� u �H�?�:S�ֈ�-OΟ��?��'#$�ǃl��>�{��Qj�ߚ�QJ��@��q$x=�O��ry+X~��X�1�ߤ)�?�9ê,/���l�'e �&j�Eٹ5�rᬎI� �?��.�*O���q�\�\)��}|�[�sB#U'������f>���~ps˫�U9����O �L"�K{���������%���!���Ps���Z���ś�]�8~�Q�w��ɠ�����`
�v9Ig�qJ1���_E��l[v�6so�Bx8��Ս�_^���R ��|*�=]T�2��B�5���4+�Ӄh��*��,\�0Y�qZ����
�U�R���o�%��I�u`
{g���{yy���7nll���"�<T�f��[�<�&��)z�bM���B���'gN$���O��<%�r�Dd��ͽ�`���K.Y����JO�	]__7\#�����]5X	�����Nּ�<��I#	iM�Ӊmoj`�[@�g�'�%a���I3S9;��/-���v��u����w,s�u�����<�89ӻ�x�B���Ӹ���a9@���(�s�3����ߜ���e_U���
;�2�S%�kv?�&כ�O�\Gr\�̳�W)�!���{G�����ϔ:G�|�څ��aMl��*�s���R%�5J	W D�,����A�܏�&�c���
5�*�l�<���U(Q��U�?��C�#�z�e�-�DH��E>߭����ޘ���~ �2�-�5��0�d���i_W\i��D3D: �#O���8g*MB�ч�2���0�L�,t�M|ɠꪱ����!}�f���햋ܾ�d$ �M	���#�d C�C��'��_`��O�Z����a�:ʪl�l��������;Y�wuC6�T����>���8�+1�9��G��Ð�2��g��r�!��/�z�#b�wj2\�9K��6��1��(��G"���
p��{yO�����krmZF��vt�S2�5���!d�NFM���ƶ�~�E�@�q�"�O�Vc�F،'5�:���>� gb���S�F,̆S�FO�4�]T_��Y�0	�jf3Y�����v>�	��٫�=V�;m!���]�˄�G3��)L�%W+�n?��ՕF4�=Mg���o� ��'��� �R �pyctB�X���������P~�����8������L�SX�ϵ�wh�lG�YoE �A��I���:��d�6�fZ�Z�� ��d�+z��/n~s�p���:��v�Cy,o�d���i�6�\�u�.�)�cGyR�v�}f˷c�U�5�3q�JJ����8��<�}���<7\�����h{�Oi�����������@
�����eBK����Ά���/:aOM"��fP���e�d~j���Mbjr�ؓ�2���j
����!.*~2~3�ኬ�޶����ų�̏^�����֊3�o89~���T�Ď(� zFU@O��<=;?==a�$!Ѿ$z{[���� 00X��F��m�
���#@x�_�ǎ"J&�mN�:R�P1�${.�ޜ鸤'`4��ДUYY��I����eu5�g�%��e�i=�yә	�������.�E�Xh�:�ud���)�|&ij��W���Vy, ����V�l>�Y^`'4�cL!Lc�-}� �%O�#q��5��m�k�Mv���LE����n���
A�66���*Q{gB�L �0�x��P���_�ĚEE�f�+���'o�Hb_̐li[��G�����G[x?�-�:��T�̈��b\G��	��ÕƢN冷���v
��\�� �	�/����I�9^gv_νO�U��ƞ\��|Σ��H[�ĭC@�M�f���t�,E��t4d�
��\�q�u�y(���=z=�pL������t+b�.���n�W9�0�²�^LP�V������j�������#?H�S���~`�ƹ!I����ʓ���ER?ԑ����)|�51"��7��-�c����^fu��E�<�� 0��lD'�!}�l�m����hDa�ll7�i�A�vB��[e��0�ۆ�&,�l!�uPф�O� ��Է�en��7|G���S���E���U��\z7�s�'���+R�-�yh��6Jv���#esS��m˜ǝo2L��m��!$ ����e=�/����RT�#�ŊV�ִ��R=��>!�)�C�qd�CUF���N	�_U�����ԉn�_�_ĸ�e40�z�N��r~h�D&�?�{����M6�:��e�]��U����_ը��+������\R�0��R;����3�Ο>fK�H��Q�x�.9>�x�� 2��u<)|���) <c�є���i�R��=4�M��B����3�l�"��� z+H�"�a��r��7���Z����¬|�V�:��?F4��e#�wlc��n���e���0<sEH�����8��#��LV�G�����<����\�� o`�U�˥��-�䫭���&'�ߔCwA[�Kbӯ�����.4����o���%�'��Y���!<O�>xz���}�v���Ĥ��BX;S'=fdjjj��v	M�7�?���s�_�:��r!Q�ݼ�l��^�����[g���b�_��H�O�i+�m���䵸$����;�7�̯{~H��4s9�_~�Ԋ�le���;�^���ܳ�@z�pz�~,��[�L*/(yY>!	t����"��K�Rȁ��M�P__�����PT�h`�&�Ƽĝ�Q@���3'�Bk}��ϐII�F�Y�T���&+� P�#�E����1�[,����55���m�n�G�u�����q#�@ J�XYV=��R��`.eB}R:N�l����ãrx���){?�a1�t�d.�\B�����E�H�hL�.`�h�r��g/z��:�w�mu@l�y����@����Q�3*�"�旨�S�<��Ƿ��@�qa��F랎N�3����b�S)d[�u�4�m8�a�A�(�����r����]�#���I����f+�e��zfz�D՝��BAW�2��]*����e�bN����Q��Ҥ�gm�r��}
K�f/C�*���J�	�����8��G."9�^M��J{��*����t�or\OMj��kM�����`�.�����q��	���q{	�V
/Sax�6!���w�\�%�u�Ѕg-�B��pHiz�Z|��ow����x�4�V{����$��vco7q��Vm�u�)_ne���2�!+��CA��G__��D��&�L������Ab��M^C&���t��GùN�`�mb���7s��%�2�?{H�3��]q����$Ϻ>cD��6���d�᤮�>�4��l=v���R��Z���:h���:ш���(�_Q+�W�W�[�m��dl�ZF��۔�����/P�kĨ141�0����J��G��`����>`9 _Z��|�(Zz�ۄ�|e����c�o�3���v�AVY����,���A�j����e�Ǌ�8���8	H�Yt"�ߪuU�5!�W�}h�8�o�+S��&��6b �E�KTȡ*ѿݧj��y�^X*r�M�"r̣���ʇ�b����H��!9���'�G�T�K�����!��a�F�Z{:�&��\�3��'�@��p�o�P&|r�6��v^��X5���<�y@�Ӛ������&�M�pONN�!���I2���w�����#��BUU�>��6�)
ӳlsR�{y^��J���3� �m(���WC�g]m}}M/-?_a[dRtI��A��AO�C75�O:��p錵��mJ����t�伍%��R�DtvN����óG�h*"�ɪ��'��z�o�+�eS ��#� �hvL}F>(unգ�J���Lh�B�O9k��CV׏EϏ?0�T�ŴEn[o@My.+U��m�v[!��#�XH�"�t�h�E�D(իqK<==�x�8�HN���$=���c�٪>E���x3w����/ٰ]aު��G�H��X��G���O��*��˫�5��x���s�u�2�q��a�կ���ʩ��
k)��[���T�.�1�އ��\v9K�6� ����Qr\� ^�1f��v2`L���k	U�o�����z*���Ĳ���N��Շ@�İ���t]b1��(�vws�_ɣ�E���~�I\��n�w	��ŭ�`5��R�x陳���W(���`�����d\�mk�G�mP'�3���4\��ҷq���1�F,�O, $b�R�"��V3��^y�H�:����p��X$!��� �E�mXK����l��Y����/5~̳J��J�@X��#�q���$9j�ߦ�3k� ��K�X���������������R���}�&�4�m��`�Ȱ'��[�֢�S��:X��f!��d��x��}�TJ�qN��p#���)�q�P���[�V�R��dSH�P�Ab��;��~n���J�K�E��:�"��X_|����H�Wl�fs��L/�wG��پ��8)Pg�1����|�ǃ?�蕎���B��斵\��ގ��/{�䡝ev��pU�X��܃`<B���"	
���l�t���?5��Ý�l�p,�,}s�|�n�(��ۄ��&�L�$:ƻ�iS����7��_]�74��|p�������y\��4�;��t3Q�f.�?.�O��}�\	�sۏ&��ߪ\�\�\؟�O��J��{9B�B)m��OG�gYs��;�G��}�N��r������L���+��S��SJj^��v�}�澛������p�L@�2g� l�����U6տ��B�HQ��:
Y&�g%F?�e&�a�<�ؙ��4��G �����!X�Xe+�2�[���_�k�,;��Z���z5bYS����ao����+�	$�u���F�L�.N�NO����>vK)�h[���%��Lq}o�?&I6q�����E1��o���WRP*%�k"�Qm��������o)!iZ�&�LtMܗ��ʗ�K�C�<3���`naާE�ʷ9��B�c�~�b��b�^�^y�"f�b�_��M���"���\�e.S`�b����e�}�+ ��������C�!�#�7�3ӑ�}��I����L������¸I�ر0"�#��8 ���`�FDCTټ������<+�N��ΚC�D�a��1S|"S;�G�S0Dˑ�v_^;dh�O�B��d��ǫ�o��b^J�����*'�a�F�*�C#����H��T�^��`���On��������:;�Pg���L��h��$�_���{=�4��5q@r��A�6�/Hˇ�6��A�wM~�t�HG�n{s;�؝�$w9�5��#�- �0�F��i/�٦0��0~���[�
��������������<����L�N9�)ǜ|��L��Ϋr�?pb8�3:ǁB>��c��Loy�0�%j�o�V�B�-7]T����>s͕l��O^1���4��-˩��Q��KMj�,�	U������ �}qI�FC��$���;9)�����}�,3��B���xp���x"Oxr����|���_yd���6��ݴ�+�x�/qS��~��4�U,�5Ou��)C_r��\�[7��}�d��#ܿr}ö>#��OƘ��d�I	��C4�BU�e�t�"�k0��Z�d�?H.a	:l�:��I	�}�}����u��A{�փV��O������x�7Q�Z���1�%>���F
�\�_7Y���Y�ϣ��KK���D	
�耸���Ԧj�D۲W��q䋵E�.�|�c������N�?�H��_�l�^���V�`+�8M:&X�4���ic4e(8/3܅Ǜ��4�!�.d�_|���t���?
�ly�лn���%<;"�8���i�g!9T_<�ID"�����BR���Y�J2<A��㌁~E��so찌<b��Z+>��h~�����{�~}k����T���0]��ݴ�;��R]�|��y�s�����Ǜl>�X��s�i|vhvjdi�ka�e�g���Iք w�d{i�.>&����� pM�Z� ��Ɏ%[�0�Sz<�Vg}�%d��d��!y�����Q��ᦫ)L�_^^�q��������ڡ<!�htQ����%Ê��ܪ��G�=��zA��O�jO�=�b��߼��,����Z����H¡����ef���V��^4nA��6�LD�@��3�'RQ�|(���/��\,i��������ZO���@����T�x�a���e@6��%�@��S��_Uj���-�ϟuhSp2 h1���������=�ʨ�O�E�,����j�=�irk������VȽN�@u���R�j��Ŏ�K��	l�4��������§K���Tf�A^�G�L�S�e3�<2��	8!� Kւ��@7��$�%���+�;��aO7D9��:���>��7�y��}il�5�!�,��+8�ǭe5�WHѰ-�1��V�J�^�խu�_-Mh����ie�d�S���_���O(*FF�-���W���P�7=v�d�fw/�7���ry�ac�'��.�F��WY*�>'��rBh��~�M������ts�.�5��	գ�s1��,�9��;z/"`�'�b�ت��AS	rޒ:#*���TT�%<m-���5��W��T==H�ls<�qط~�w�����h^�+2i(�Mu�k�������s�Oq~�tJD�V�M�*�����He���6�С�S�rU��J���� I���G�ƚ���m�v't��D���l�:j�
��F��iJ���,X�N��^+�!��6�y�_R����]��xVE�i%ҵS#��T�j��Q��8�����#`x �xb�����T�9�o>���5i��5�-qf�3Ƴ�1p[�1���q�T��k��-5y�OP@���8P�bM �1��
nXNT�[UR��!�R��BP�lޒ�Tȁ�R��1\�,Dq��^���r����)�F�*���X<'�	K�"ie�Q6�q����C٭���y���Mf�ɇ�G��:�	��[�[@���|\�@��!�'p�lJ֖֕���Փ�U-�����EJQ��6io)����h�'V�gkq�C~G!�����'�rN��J� �q�nE��#��M�x�W�w�4��*}�f�3.��e����:�eXb"޳�ݝhp���-rpop-�|�5�aטb=s08������$���bD��n8[cs��&WZ[yM���tt�땒xV3P��7��A%3�Iwpxd������֚�W�G� ���	���Qh^LR�$�d��#&��Y�{l�	���U!������\p���FPX�cxdhlt@}LIC]YYI�K�F,:.:*:�,�9|���,��Y"n�K0"�\�P_!c�AB�Y�V�nr�;TP�t�/�UMp�x�����*�|�4K:��B�N�na�ö�;��BL�5���ݤX����7�r��~�$������L�f��g�_fd ��3���	�dޗ�+����>��YU�?Plzo���� ���p,J���z-��4�78 �Z\�����'�D���ex�̈́{�xz'�{'^Ʋ�X�.���d���9��Y9�=Ӑ��$�vB��q�����_�<�w���lF����` 55{�ּw(��2��b�cZ⨂��*���5A�&�������>Z�
�7��11j�� OL�j���q�ձ�p�i}�uX}sj��B	�������c�%��w��$o�\��<�K����>wp �Ȝw* �-<�������*���4â�b��\Ҟ�r8s��t>��e^��XL���ڐVtF���g���)0����Yl�ܿ�?�u��r0���v5O0ҡ�h�B��[c���z)3���s��ٜ��4�EH�3���ק��?�rN"���(6���k��B��f^I��kGz):��?��SW�%��Gc�@ i����	b��c��Ay�b�����V ���m풵��O��GFb�{�`�B�x�H(���N�a����Þss�ǯ/x�mZ����*�xh<=T������V�Asj�%�Q����i������Î�����,�3��.Ab5���y���8���
��U��#���*�#2�^��ljE~�&�G9*���Oԏ���fb���;~�2�O��~��v����C��I&�2 ��#���5~��(���qY�a	Q���	Uq����]qR��&ەv�p3د8�S�()rZc��5��M�`Y�O��q���ױ�` �PR�ED�Ǒo���SV����8I�y�?5)J�v���~�H&�4��{}l�fkH_������!���Qr�O~���l˿<su��r����2e1	�N�D��m̕�s��Bd�0�/�����ux��Gۤ����,�B>4��cLmD��֭|��X����,�����/5�Ed��� ��Ғ�Đ��tH�R�!%0��4�-�9�E��g�~����8�qζ�������~�ܣ��&�}>h!�.�w�"$��U�0�jT��n�.�@#-���Z }���'�cB�A��H�x � j�;?"��;�mX�)�:�=�OC��g��.�N����}t�5���K���/�S���ho���$��kLx^x$�;�*H`��I�8sYu���2Z�����ta�B^5����7�Å�V:;��$��A��x��LTϳz\0�����`�AO=��fh<�g���\�>j����\\�&��U��NAFr�������ӊ� ����b¦7�%�05)[K�\��1I �;���T�,����8ws4��t�(������W[8Q
V%m�VV�UU��DEE0"��(���������N�ez�"������M��٤s_��D)8��k:O�JЫ�D�ۢ��K�_/�93>�.�`���`�����Α���_��;l"�0E?R6}F��F�T�;ca�ӿ��;�;�����s�RU9��zirM���}�A�����B�����1þ���	z�����5Qfn'�lH
p
���f5&��p��c��p�IS���J_mO/�G�>��8�F�`t����ן{򩄣n���`�d����o�"���	��-�3�����M���N��1oE�n?�?Cϣ
�s2���CF�,�%	��)���TD�c��a*zJx�LzL_I� �~ބ�X�����_���F3�~�̰|�����旕RR;�]Xx�!y:���)�(ne{Qr�݉G��n�.+O�vҴ�R�	c��U���)q0Y�X�Oym����v�5s��4���F���칟�.䷙��=�OU�Ԅ�>�b�1�<w}���ƴ/�A��j��9��Ѷ�D_�:�cJ�q��Z7�(3/1��n���0N
zb+?�;���g>L��4]p6ԋ��}`�{�ر̐]K�t�0�{����*CtϢ����a�����"�Q�[
�z1�$����B�A�t+)}%G����~҃u����ʳDr ����G�{��Dc'I&	(!��2*(�)��J�-E).����s��'54����Ocr����!1�������Cm�&|~��^���N�1��q=j16(N�'J�"1�'O���� 5#¨�����$8m�8Q��eNV�Oi@�і�o�Q'����gL���<6�4>���]���KJN!�o�������C��#/|/�`_�ڣ�3�[�
������˯8�Ҁ3���ܯ}���D�#Q����Q7;X�p@����!��R�}���dܚ�0�6�knm�j�Tv�A*;�������@H���df��Y���11��^���mE�c�1 `#]����-2Z*aâgn��Q��/��H�;-�>}nI��˛e>ٖu�Au<�b�Q-`�/=�=���m;�8I�wS��?����W����e�_�r3D��f��KP���O_��m6Jz��f��]��2�;$7����1�j$�A!:�7��<´�|�%�*���W������HΩ���d��i�D�l}��;ʽ��ᆝCCr�]��y�r<~���b��4��R������٠�wn�}��C��큫��1:Xh�PX+R�#��=U�6��)�I�̿I���%b؞���%R��>u�Kz?�O4^zb���� ]���� �����|ܸ��P���L��J�1��%<�}d4�#v��'�Ǥ�kT2�|��4d��dB)<�z��㺕���c�s���N�O]��xu�zA���?��7ȵ��N	��s�1x�,��~�n��1�l}�����M3�T�5�2�
$��f}�Ӈ�fb�L�M�V�����֪8*S�cm&��5l�`ϝ�I�ӳ��G���5t뮹-�>qA�Ŧ�,����@���p��EM�5X(�+�"�j��h�g�q�;����soM�CS,�H�F����w% i$�\/�\� a1h/��m���w�+�N�"�	��`%bbHl��ah���m&����|s���@9`Sz�3X`ɫL���?��ތQ�m�p��zU/a����b��6Q?���9���R��H;`~��A���J*�����z�iSޥ���%��O.φ��o�T�x��~w��(�]�vi���%��7�/V{I�yhbJ�VAcp�}KߝG$��|�/�	>$Fm�F>/[o�LL�? ��e�]^aZ�Z[[����c6�I�H��ș�T��4��V��M��B·]9��Q�|��ʮA�J����#E*�����ОQ{Q�$Z8����E����jc�6g&rN�cp�_��c�9�������
�+s_��N�p1JX�r���_�T
L����z@B��0�OC�Ӎ\Ѕ���G��&�]�Wx��46���z�}$ �
�9V�Y�菉��֜+�ǇU�4Vu^ b�=��mP����Y����L�(�A��ōU������U��7 �b��� ��O����;�5\V��]��bA�u�~|��7�ix{�H����|g��WF���p��8���E�U՗ф�)}�Ȥ h� �8��ԯ��Cd��!_?�)���-|.c����=;r;��k�/�h9��f}P<�W�wp�_��{ JZKx�����a�b�Q�օ�8�����ǥ�@br2L}�&o���arH�\$�W'/Q�l�6�]�[ ���%#{���W���vi��C���g��yt}ԇ��+{0%�B[̚|t�'������;[O��_W��"w��~:���9$�H���0�S���ww�=����x��p�)M��]C�5{������UkBU8�"Ӊ������p`�ʾj��K��M�5d�@��6��_+x
�a��o��V7�=��'��ڰ����\A�n)��"j��-�����A�u�����$�"-�[��>�+u����-��l�y��Wit������ {�#��__5��RH�x���o�,2pˏSA��p���a,�ap6�c^'�_���kz iE���e}m�g1����%8�����!Y{76+�'V�!����/�lJ#���i���a�</�WP�?z�ƒ"��M=l���@/�D1���˚|�G\����;G�@�i�_�К�E�3/�^�̏�`���%uz��p�I���|�å7�����/c�T�I"c�>?~O�%s������g��oHPeav�te�+��o���Y�m�b*���DA*oI�o7�O�M9��߿q�=�����ѡ���� KP��@r��xV	��C� ���u	Z�S��W`p�5�vƎ�-ܕm�:4��'9G�b�///))���{ï��N#���m)����:���u!X�~���s��K��6)"c��(&�{��w�n���d�NuhY�`O�lħ 7c.@-=�(ė�����%��ml*�Lˍ����!#���G�g���]�=�#}�����m��e'��?ʄξ�B�Y.�����>v��<�n/[-�<M�M{t���T�z����dJ�X�Y���U�>S
������wF\|F�vJ�nJJuTwf�	t�=�A�e~��A>�K�iT�R�}�����둨N))d���h:u�H��(9�l�O8�E���揅�3�/A9����S��06,l`x,wX���؞����G&�&U��LR�Z�
�o�ƣ���r��O~�ju ��K`�k�ִ�A� �P���pʊ�zM�G�h�p.���#���=a�Rux�A9��|� ���n�	s���]i��q�OHڪ��i�%{x�n%eG�[�k��=���3< m���a�e`�6fx�r?C!D��d�5x�D���.��'��R�Vat�aC���w�"_HZ��KZ�w}�c=k����y?���L�{���?���q��;ow��B_U���@��O�Ν��@ޒ�����
��c���OQ��#�c3=�~�S	]�G��8�6�-1]f@�?��CV�M-T��; S7a�hy@8d�JL�<�{�,���ʦ��m�2�)b�#�E[� C��G�e�1M���sS�+R���c�r@� _�4�]�	���?Ӹ���Fp�Z�"����g�R
�08���ɰ,���Ԣ��8��K���>��2��J�1��!������E����c�h	�D�ƛ���5�+��6č~VR'?w�ᓩ���lVs����џ#�����"������?��Z;|}���n���= W�G[�9�ļ��dܝ���G����,���gJ?'ϲ��)�	�k���3��4MkǅY�5�.��f�b��Yy�ʧ;�9����%�G�s�ru���Lg@]��eDRBAGww�ޔI��)M�+�Q8��M�������#�헸c|~��llT�
��7^�����wz�TN���p��cE��٦���ľh��i?
���_��o��m�AGo)���)�>��FF}����V�������@u��u�����7���]8�i���M_�^�T�ҿ�Ow���b~��r�xԫ�W�H�𸞭�x{�PL��{5}�
A�q;���a�ActT\����`Z�P�nF�gR�NB�V\b�ɰ�rf��?7������'��$�c�U,-����M���b���-�|W��VӜ�p��lh�`v�!'0h'��P���s`>����� �X@��%���`l0;�32�tٚ��Ls�N���c^.nw���J���d.=(�VX̭����@횔��{�{�i��u7�l�����c�V)�����������.�V�tĂ���eBp�E� �s�a�?<à����b`�?�h\�>p��Ԛ��9}J6�cp,�F���=0l���K��YP�ԯ���鈐r;On����F��鎎>����x�G?3��.���6��.��:�t�/OZh$Q-���|<���e��,+�1�=�� ߿�Kyw��b:.-�+w%�&N3ؐ��wE� 
�brnfh'��3�]��'��"�	6�<qY�Æ�q��7W�_�L���$ڝ2�?���^jfmO��6?.�U/$h�r<��3�=2i����t�zgmv��p@�#��(X��,I�"e:I�%����,1|/{���
� ��>���T��h����lB�͟EgNK�P�u��&Kcdp��[ki�)4���o��j<� �$��D,[�*hn��N�Q���i�w9J�P-	�`0�e���,VYK439x��-�&w��g��@=F�q�#z�O���m���U�V��Y^ǲ��F���+�hi���"�.���"��R ���wtn4��Е��������\}��l�*�'�jx������R��Ƥ�"�0R#���h�	�����{���׾�g�-sI`��#�!��L�����tll����EZ|4@%7{���˫�ޥ1��G9d,m8��}���q��- ��v�V�Al���I�����W��r+���.�<�r\�Ut`�.on�ׇ���n������rb���$�}ty�5J��6G�[H����B��ֶ���������+ˏַ�?�af�G�$<ʤ��V�0u�9H�F��EV��/�*�7V(;�#��'(�M��K�%������B7����j��17�i�^U7_&�S����Q�TΝU[�sI��/x����O+=\+<�=J߹��y�)h���{1=��c�,�ւk�����L�����<�;�Ϭޞ�Ya*J�c/%�:�_�kx
3;����!��91�R���b�xJ��Γ#ã8�Wnۏ��7��쑯������׻>�B`�~o:��o����L�=�ߘg���H��*u�b�l6:����˥��f��S�;��lA�筴\<��+���.��ѽ�h.u�T����2�T*F����?�g�+�ϊW�·&SH?��ҩpu��Ξ�IIgؚ����~A9��!�g�Q�VFK��a4P�L�b��϶�IZ���C�H�ި��l&�}- 
���+N����9�vQ�'�CE��!5@�&	/�#�qnW��?����g��D��D嶹&���/ðn�^سL/k��qE �8Y	��Bb=��,1G�2.8�Ã����ģY;�`��?@��R߹B[xDc��FWk���3R�+D15�G��B��4ܹ���k�7`'�BlZQ�ߋ�ˢ�_���O�u'��J#����/"��s�'}��#h���R�7���Ϗ������E��m!�o�R7�,!��"{h�l�<$�h��~�<���_�B���W�8�� ���ΛVqD��Oj����(А������z1kn	R�XhJ�a����2͋������|��aw����1�,�n�SD��]�K����!���j.�:��̶�`��:0_ߗd����\���W�Bbr��v�IU�ё�8%d�e�y�E�|��d����^ ��kmo�DDM͟�4�o�b)s�&ZV,x_��e�>j����Ctl4n�����8�����<T��x��5�Xl�r��K2�Յ���Xdn]�f��m�[��Ԉ�׻2˩�H�z��{�tN�}��?=n�Aȟ�o��9.>��T.���j
�'zQ�# �� (&#�Ns�`9yy�hx�.��k9W�(�9?G>h�k����^���s���� [��G�tL��r�yjp*-+kG[���V�k`�׸������ݛ�BY�۞	���̠�m;��K3��p2*pWC$h��0��/�r��_�I&�]�ei~㉔#�X��~���o���GŖk�λlv�X����dH�̝V�p��Ȕ�aISQ�䧍���MB��5A�??�lۿ�#��#���ѭ�E���.���hP�������h��/�ǘ�Zዿ���.����r$d�O�`,�8��_W|x���k�5J3�֘�]�݀���3���J����J�s��|Z玦��#o����RCE-�zo�����pr����G���t�1��j�R�d��f��vN��nM \��ӍQ����9cJmV���S�V�[��bw����"3���?��4�4�u#}{�$�%MGSp�6���QxV0:�?�I������R��A6R ��d�8@P��), �8G������@o�\����Y�ڨ��Z�_� ��#:��_a�Sz��=���Q%N�#��5����GϞp֓�����f�NU���N�*wzE��TW��&�*���+���+���H���Q�q�-y�a���[����|_��/�m��'�V�c6����z^��ߟ�a0�S���^��X�>�Z�Jg�%�CF�K�h�`e�B�9���$�|��o��
E��8���*H���+q��i<�)���x��g-��>l0�15�:k-�r0b37+��Y�����������4�,��	���N����n_�����p�E�M]A	ٯj�P e�n]�Nk/��W�i������/Byo|��o����u���*��y�[v��� &��R��1����Ԩa]����'<�!��%PtݴEZ`T�<V}�0�У��9�����U'�����m?uB$�e�vR�Zky�m8��y�����Z����f��P|+QD*��;���Y��ɒ����H}�y_�з�:;�����տ�%7]�!?�E-�/��Gu�%E?�U��
��w�-�)nB��2�OR�y׋ok�;�R/	��&����փ�DW���¿갏:�����(퓑?l��'_����Y��d~k����G}�tU5����v "OKEes|9�M�+�Ϸ�v��O1Ї4��u.�ԿW�p�Z�'�cm��=+ZE6Z<E� <6?B�G�A-����*@���?�3�:�@ӝ���z����z/j���slt^�>g|�􈙖��e�Y�8���g�k�����(,���c�����E���ZƜ0P)��P}Q=A���T�R)<I���D���U��Ι]RRq%���u�!SL��Ä�+8��N��m�/�3��<k�Zn��t��R��E}Μ����HZH|rJLzGF�	�����[h�UH���e� �6�6�?�s�xsp_ӆ�Ƈα.�Q-����P�I{Q�T�`T�dPߌ� �5�H�k-�nYP֌̌	��*���n�
���HBW'�� ���]�lWU��LK>BBb��ė���ӫ߽�a(!aaK���s�ۢ��*��5&����IC���Q���N�b�Nv�<�PنƮs���1��;!)L���K�VE��84�8?���ٯ���������,�2�j����|?��j����b����n��&�l��n��@���˃?kC�D!�������uJI�N�)��v�����/����yX�<�b�tH]������ԉ���l�x�X^>hE�h��N�#>F�pT?}ތ�`X,��TP�^��[%=��g�*���畟��)}ƶc�D���q�����w�Hyۋ��yﲻ�U�H{�hN���`��L$�*�o��m]-rS-n��N$��"iG�7H)[3O	;��Z�N�+R�jkM�&�����%�=����z��y��-w���K+�ţ%T7�G�S�JΝCaM�jN_T;��}ٽ���^I
鏡�rɘ����W�ҿ<^� ��	�P��
Ϳ������K�d��>\�ݿ𣧘���c�<���ҙi�飍>؅|�
T�8՟Q+3��.y�y~����4؞nt!�����8A�k�p�E|��T_���4GYw~�T��R'T\��ć=Ɲ쀐o}��Nl�����B�.uבERT�@�p��V�+x`"㟅�QI���B�tt��
IL��"���Y�{�a�D��?mU�Β,�F\iA��W����N|�^"B��
�ЗD���՗��u *rB�>/�ܰ_,��!~<E�cmZ�3=u��]�I&)��E4�zm�e
���΢S��:ַ%�m���]8���k�a������˟�v�vW�
=�'�c���m��ey�Ճ_�*e���	����k�f��\3���L`*u�<FI9�cnN	Sd�š��zƑ�m���Q/�z����Ճsҝ{���w�6%��{��Ȉ��%f� �I#�����퉮��o�k�^h��d0[��,[���r�23ɟwLr�t��������Ԛa�,&aC�z��ւY<2��H��R��i������#kݘ�I 
��:�2����d�VtH�J�w(;�������/8�}:	jh�����M'H�&T>l�;$�sD�"<2g�U60�����i"���:|k�xfH/���8�VL>~���윝���iudg��!Ùu�Ԣ�Vc�+������	��ٛ�������SB1ٛ���z��}���蘒�(;���ݫk3�È��l`e��uA&zG��4iowp�Z�T�J�(���/���������D X���L��&$�q�ߗ:�/��¾�l9���T2��$7hG Q�r������S[ф7�Sގ�g�1�?K^.�<kMC���aYQI���zV�Q&��(��j�W�7�Ea����t�s�cey�<#m�y�r�c�daX�YQ*�`�?��f ��6�g+L�60�X'g�NpMZ��C,�_D�,��Y%Uɵ��P�LQ�v]t:��zn^%^N?'*��2��f"�_mЏ?���;�T�
���{.�v_���w��pQ:#�k�5����a��hA0��d�r~�ZIMS�>U�7m1P������l֌�I�0PJ��񅶋\���O��������p���3�vU'N��f�<mo <"t��WH�x���#�&,� �#�,dOz�qe��>]�����nᵮ���\��;�����4l�"���ơ##U��ߡ���Mh���U�%��K�N�u���HԲ�c�9��|��&�%R���)�#H8%��F3.���D"GV�~�<�*C����4����4�{���<S���G� gQ�=^��4�/���0]B��o���yiڎp�G�X6y��q'���7L�i��j�1p�V,���	�'��O_�,�*�Lm�O>렫�f�6��5�F���C�^��|H��W��|���*��?*���`_���u�1kX��z��퍪eݦ��9Ú�w�o��_��A
��QZ�}��;�M60SO7��������kK�N�����"�WD����SAɳ��f�����ֲ1�-P�>���a�Ž�6� ѢڗĆ3�Ą�xO8��G��v#���"�ye�]܁Q"��j�k�wJ�D{ER&���Y%����� ��4�ʨ�=q�&=H��fk F35R�,;���j�޷��ޫ�Xα�d��P�eN/%EH*��NK(B�G���H޹[<|�����1�99��=(	<���v�yst���h%�v���2y��:S�F6�6&���i�����Og�f����'��C#Z�s`G�*Qdj�̌dM���ȟX��Em>7��306��X\}r!���|b���i�o��d�l�X���2Ζ��7~�c�N9�)7e���3��8b)�)Z��K?�ͨϙ�6�
�����s8�͑Y���qQʴ��Gӑvq�&�W���/' ���Ne���k9S'�"�^\�;���~�Ht�?H�q�v�������3H��8���<;��s>�*�FS�Pc@Is+�����m���; C�w��(�����ߊrn�x(ټJ@!���M��g��Q����ͮ��{"�t�v8�Olt#��4v2�e��ntG+"�c^����&$���ǳ�ӉAeP���kw�u�0
!����<�0���6qJz�hY�x�
β��0�:)�%$�!Ǿuc�F!��q��u�<S}�1�/(Р%����%q�P�{O([����%8�z��DTh�ۃS��QIAZ��pT&����y͛�f�4,����r�f���t�?��+*��*9������R��f�,��h��ԇ����d��7���r��(s+��@�f�2`u"�y_<IPly�N��(}�i�hs&Y��pW�aѢ�B/h���a��KE�,�鞧z�u�?/GA�)�v�K�N�pވ�w�R�
�*BsWE/�e>y���Z҆#aUo�ഠ_��dN"��퉘�k�k�+ݗ����n��w�������8!O_Ƣ#*�IP�A(aa���9�I���R��yϨ\l���������;܊�#�s׍)k�K�W�]�����~��H�|@�j��ށ��k���^�>�.�AGi�jK��QV�B`m���?�p�(��j��DΑ�n�9A�+�a�,���/�0Z�?*{(�*�I,�����C��8&9��7�>'��~�,���t~9`�3��~�Ih��������rA�pf�س��A���I��~�J�όg_/���.d�7���ޞm�f���=�͸�5k��n�}{0�|[�|��xt]2�������Ri1z�����L��lW_���h|S�
:�<G��3%����}��5�3�T�{=e�W�\��(a�L��(}l�.��\�����#gk�r�ˆ��'�
��2�C�j&Y��B���'���T���G찎����y��,A��!b���-�Lً��?��\��ʈ��^�F|�	ߍ��e�v!��O�$��ƿX>'C�r�TbD�mp��!�o��}i���mu�	���s���j��A�7�������7�)
�
!��q�8^�*�
7e��W9$���ۼ�7�Y���y�Y��Uw��w��(�x��f����@���:�u�uT��f���y�E���`0Q!�s�c��6kD-=���kTNpVkX9��ݟ�5N{���Y� 1;�<�y˗�{D��h|�E�k
p���B;$�T�C�=1TΟ(�����?�B�zؓ�����&Z1���I餱���͉�o���RBY����(�!Mtv�o�g�o���Tl@J.�o�L��n6x`�����F�a���6E-�_��t���!/2|�-t����l#�mtC�_�iK@�����y��nj�P�z�j���-n���gE�0��#W>$n�� Q��Y����h�]^���v�u����n�qU�-���_A�C�x���뜑��90<�y@�C7�b������_1�JV�ꠇ(!J�D�='g�h��u{{��-b�gIIIЗ\�v��̓����Mw2~����OQ����ct0|����	 ���Z������B�oi����ht�VM�MV�P�*�6�ia��DK.�\�C{>�!E�z�C����2�&�VS�'(��,�Z9��/��1�ט��_�ɩzqqߺ�soo,�2Lqd��o*���>�����R�~ľ<IJ�x`KS��0���q􇋰lV�{=�{��x�t3���+�Bo�f.oo~2_eޞ��.����/�W,�\��Չ��4r�<隟յ�����TF	�?�?r�C�w�	����� S�?2�_����i�J��W�����`㜍9�U�z5�|��zȩ���b��wK�ރ������`�3 A�?��YbA*��+$B.�i7�)�����q�&=ecЛ�Э��7��$��;P�|ZA���x�-V������:�V��fG�+�w2f�#���Ydw*@��Gc|ٞ���zi�x����+hR@���}�|�>�P��/�d�c)��9t��&&�p����wU�6�9��KjQ�Z��p��#%*�Yxf��ǗI�����k��G�����o]�aW���$�=�&#P�?�3V��qA�g�+(�鹘=<�h�
�YW^��2�t�ArM
�7�*���'�}�*�+��8<T�=��ń��|hܱ|�a{,p�A�3��ٜ�+�8��응��=����qpb�6�1�U��G�����g��?��B���q@ҵ�t�ڙ ������|Sݯ �#�'(���zEf&�B��@���
�[��R	s�s6��X��I�U~wt��4���oǏZ�����.P�����+�!W�a¼v�Uk��>�;�.i�5�x�*$�KK	�� 1�V�������W���?��f}}QӒ!74D�	��{+���G*��-�T1�N�����Ǎ]��O�v#��c���C��ŲJ�5ԧE%�U�E�W�F�W4ƄGfΨNL}��b~���6��Am��i�S��2�}�M�FeH'��jm?���-��G'��A5+g����s��
7#��ݣE�l�WuE!/���"uS�����R��W���+}�gw|C�G��t���ꜚn�m�q������nhP��eSPh�`T��?*.NV�������Va���<������f�g���˷���i�s{)�|}�x�/{w�����o曩������ϛd�'�hi�U�qc��"	������B)�3_��|i�`� ����5�秝h�W��I���t{�i���'b������pZ)jWnS��T7�x,��Z��iM7�/�f�G[?������98f���OخL��k�f�5�}���R\����wn�;(���i'��y����c���؉��Έ�I_���u�Z���KW��~O\�!�`��iݮ�!�<��FaC��K�2Q-�>��{��[J:a�C��=��
��f- 
 p�1$!�o�d���J�;��w{����le��flw3%/�K�+ҭR���-vw�����hx<:�5}߭���TG{������v�L�1T��O����q�k�¥"9HD�k
�jS�%�=��I��(CC�1�u��D�Ga^'@(7NԤL|a(Q�P�UW��.����02���HZ�� I��8�?Z��u�mǚG�_=-���@���E���;�Ԑ.k��Č�B�Cy�XW�ߩ߹�!ȓ-�ٲ�J����)�ŧ��5!�md��k&drǁj�u"��*!�i� _$Ma3�Py|�ś��Β0�/].��)��tI��B�����=b�B��05
-�𨝚�ME.���C ��x��r���
��s��E���'��@O� ���+�4D��{�%�Kf�����V)H�n���便5�(S202<d�d�3�omnm4��퓚�;�˟����M{��՟4zqW��1������ӓ�LՋK�ՉKHLKM�������=7Io�3�����������X��O��.6�s	V01���C��+3 ����7�)��h����0)=�W��,�Q-�ʐ̴�� ߂K�k��,����f�d	�6��ء��]�BFK�ߍ�ђMA��h>�z.��++f�In~���q���#�_�X��.U���Z�X��[�(�[7W��
//�VE͌���Ы���[t������r�(�4�_U��WV{���U�~����� �Oi��M~[X`��
]1/\��6�7K�,��f������)�U�ۙ�ݵ�˫��Ao�WK�δ�����V�\�L�5���ήkR��<.�F�����#�R�Ǎ�1���R��B�5s[/5���d���'X�\+����E��.���
���`BƏ)h	��rk8��,�=���;l�h*|g���+M�������%w�kxxՉ>u��痽w�z��<��Wr��H�(��k�������3?H�A"��N�m����~z�����k�����!�>��nL9�.C,�p@���E�kA{��)E�ʲ�lL�L���R�P�A��XI��o/�Ķ&O,�Ř?������ۏ�f�x=g*��|�v	��ZttN�
Z{}~����?vH�vW��=P��4�-��/Fk:�nJ�;T�]���Ƣ�f�J�U��g'"P%4�/��hx|wR/E�JN��pU�X��rP}���)&:D��{y�y��v1�Q:r�d�Q�[_�Z�]��N:5w�pj���up�W�S�����=?V�_��y#@|@^�ARdCѴ�C{�(�Θ�Q (�������og��tm�,�ɏ&C<��V̞��EGo�a���Y�_��ѳ@�fA����|O=a�8!�b!�TJ��!�k�����7@>-1s��.�q�C[l&�Z��r��=���(��g�|P��'�5�wU-=�}��m�,HN�\K5��d_�v$W���w��Hg *$��)&�G5�3e�hec�FM�s~��{x~�Ww���\xV�ȱ����#�]Q�3��us�p�T����U�ǚ:`C� X϶�V��d�� xj�i��CIG�?`�gf ��8b���r\��`��Kr�2I�R���2I�\�fل���5���pvq-�:5���G������G�慫�sJI��� >����I
�]�al��R~b\vA.�m�c���ϻ�YE-�[�.tEH��%g�E��l-���w�wcr_�^�6��:*	:\�}{�w�1u{�R�|9z�|3�t�+�vY���P����j<�9�z�_/[��b��v_̻c�19��i=NC�؃����32�3��wMo�ب�3wl��Y�Fa��\���boY1-Gx,f��{�V�#P~<+v3�(yrt��F0�Ո���\m�I*ʳ��E�^V=�d����s4�Q�y�T�x��ֈ�����ͺ�V(��~g���r�yJQ�G\�ػ��?�;6�#�l����c�ԗ�Z�>]��\)q�q�E��J�<��!?7���FP|o� �.��y�� �!��ҎO�(&�ku�,ɱ�����A���Kd^���V�F}��.�����:'���aS��hQ'|��J�(
�	��&�+�p��_��/��u�=Qyjo.g������8=����炌�}.���6�����x�5�"1��3ި��}�m��:xi��:���m���;�ᶬd�S��f���\���d?P�K������]b�W}�9;�Z5�@�Pw�O���bi�B�(�ǃá���U1J�~H�܋����
����l�i߇���`����!0�F�������I�R7����
��R��W�m�!:KS�m{�0޵DV�^BK��m/]a�H��ϕ���R����Bd���B�qh�]U�X��� 5��<�EV��m��oO�M��N���ݎF�"O
�=zO�0�=�Y�=K*ټ8˓��b��1��J�v��ϥ�s�>P�k/����⡂;b�
�*T�/�H���?3B?��>���
's�Q $TH`�3���������α`� ��3�"�~i�{��ה�1�-�ON7�*�%��TL���a�	#f�i_��e-a�Fs���P�i[�ۏ�Y&쥕<U���8�Y��T)��ykk���l��1P�v}m�}D��U8�n�����{oo��y�{�U��5F�U�����?�3��]�נ�n2�y���R����05��g!�lj�`��u1i����J+	�W�ϥMҿ�{�}tw֏�V~��~���h�O?v�Z	�
�>�@}Ϟ��C� 74!�տ=�I��>��,d�7/R�襖��S�}�Σ���1�?L�g8\����E�� $�m&z���w#��F����轗 D/1Zt�{��?�����1oxe������k]+�*��~f�0��%�s��ؗF�Fy�p�,������q|�Z�ϙ�7��:W�}T�;��ݝ����д[��թNH�?�ᄟ�[������}�G��ԀC��Y�]9� �����92�MiE|�onn��n7�� '�xg*�]�WO�����&��e��e ��n���$m�,��lXd-Z'/�0����c�q��C�� �ޘ��[��~�S=+�&��͒uɾ���l���Ԥ���Ȧ�!p������pR���i��0kk��zɴl��u	ΖO����Mp��+�L޾��}dP@�Gx��hK�������^ܝ�V����Dne\�}��Ӛ�3Z2Ƚ��4n�5���"\�r�N��'��s?ip7������6��nfA�v�n�~.k�nK���tx��������ݝJ����ւ�K���Z��
������6z}...�̻O� w�R(������
��-|=\��+Q��@ �؀��S:����q:��lj���no�^ڸ��<��[���@dzk���������Dil��������&s}�6WP�����θT�6z3���܋ab�L:�Z��������P���4���=lF��F>�`kI+j������9������	g*�(�n�⋁x�-X	�n�W��!�K⏁~Ѳ������S�Pp`�����V	r��;�DDH��L��Q�&���H,�����f��s�wn��C��0ٜ�WS��X��L���ȸk
����6��vg>N:��F���a-c�]3��o�й���\2����:����B"�@�!�P��T�
QZ.w��5��`����}��������ThE���I]K
�-�����U��� �XTJ��פl�TS��F�7w(L�~\UA�����ڪ?M
�=���D2A�%�~����ws*Y�(]XT�~�#[&��t�Z�г�j�$�T�����}[Fc�Q�����u�2��)����o�J���J[������SH�?%i4+�����Q��4}Bx�گ�<}�OjUO�x��5¹�I��#����=�s
��|��Mq�=v��\3C�������Y�������	�J�����ó���S�ha�1�����2��C#$�}Ȁ�P��,�/�OI)w���:�����g�Uo�_���D�i5��'�ȚO2P�/�&zr�&�N�N��S̿���}�q�µk�?�]Pb4_k�̃Zj�����v��^)pԯ�ɷ`����&	_��ò��&�Uz�Y
P���:�$R������	���}����me���w�+<H�v�)I�ܝۜ���D"���kk�<�~�5�+**����OMMut`�C�jD���H�-���8�b�O&�_̌���?�,�x�|n=�P��#3C�g{g�&�K��V��ǫ��I��0B��(�q��AJ F]S���� ��7�4�b�5��-�J
P��QL�������}vYV~QZUK`����0���I��v�V����S�������u�k�͚Y��c���]��c]����[ę���tw��bW�t^��}�:��6�w�o�Cd�k#>s�s�|�\��N�!��E0�&��?���?��Y�!Y!Z��<��n�g�����?� &*�I}npUg���\FS� ���/��������I�<��D�ϰ�� �K��Q݅����BKrU�0��mX���{Ѵn���J�x0G�Z�Lâ%�+W�[_X�ț7��j�&~�b<1Ȇ�u�{0,���R+}�Hz�EK?mh'A��.��#��{�z�|�X���ǥp����u/����f)5����dE���$�Vﰌ�l�`X�"=�h��|"x"U^�O�l%�|E�b�n�����Υ-2 ����ؑs���{ �Ћy~	�L�%P��d���KLn���%���O�]�u��(���жQ�0�r&xy�o�hH�݀� �sx9Y�k	�H/��Xq��`	`�6����o�����%�Oz5Ȣ�$�Y4:�嶗�����,���Yo��n&��=е-���/m}��.U�t�4���Ou�`���D�E*q� �U��������^ ��N�-n����������J�#��b��7H%U3�J��P����7h�og���F!Dxv��&���Wݥ������@wO�ˆ������F|�0�Fx4vL�~��������.�p�Ҡ�{��;G+���_}�SDbu�^1B�F���~�� �|�1�]7%�q�~N�y\��x��J��!�s�_��sH�#����_p�	�b�db}�+�i�5��sv�=�[�Υ�. b8�OƠ�$�/�5A����x�w�%-��րyo^���������T^Cj���a��vQ_����3��Wu]SxhxnS�ty1mCVrSr�����I[Iesum^t�
��K �4 ��8~-�z:���҂t��^G��y��I%G�������A��߇��� ���-���DTT�����z������Z1���ׯ_ڣ�  iIǅ�}B
"��0OMA�r�T��+t|;4%3�{`*�i�nih��
>y�Z�[�/#��J��`��7�p�AF��@=�
ܢ�!U�>�����+����9T�/�Q�����EZG�����æ��s�͒�23c���UC���ŝ����Ͱ�u���MW������M����ε�ݍܹ�}��Q���ź�E���|�Ŧ^/C�(�.'����gTY[�YV]��\=�j��뷃����;#;3W+�I�M��������z�)�.s�B#�#�5u:��kI}�r��R}!w�����d�h��hd������ �s����Ag�4���Cg�Zq���C�ڐf�+&k7��Ǹ�.Nx��||��H@�{��9�x�~5�����s%r�@�FP�1���h��C>�H��h H#��>�5��O�9H�u�vX,�;CQ�ţ�O���,B��~�|��)-��z����oc!��M�
����ie���gќp�8���s/��MD�ګ�0p�|yZ�3P��r��h�����h�� ��U�ڣI��<�`#S�+K������?ت�|���� (6:�c�bK�"d=�b�1�����Ir+���(�A ��X���V
�*4�d�؏��wQ5��)'�tG9�	�I����C%�m��QX(ߐ鈠�,��<�l�h����*#nH�;ݼ�R$�&�u�������hB�oA2�nH��Lޡ�G`D`| ���BYF!��m1}P��������:� ����R�D��};X�tc�i���KWs��8�����3�{=Ԟ��,u3XHi�z�yb~͞�P����򯤁�h=�P�4�V��� �ʏ��3�X8z莻�{�=�⛚Қ�1!��y��H;NNN��f��/XXX��t��I���tc�1�yܮ�ߏ����D4�[i�7�����|�=4�|�ֻ�_x�*���S\�׵��yoщ��g�y�m���`���R)wvw,Kː,��=
�ʐ��������S��ϛY��Ņ�E������O
%{J�=��`���`nFJ�HO��s�����O	�>�����_|��ޠ>33ә�ϭ����yflll�M}��'�t�e�!$$$Q5���;�V��|F�X��hu�I���?�	?���~;��p�׃vˌ������%�)/�t<���tR��(5���%6?�&|��a��w�:H8�sӺ�� S�7/��X>оCt_�A�S��vtg��$��)4(��y>~,�����������t��F�#����a����MWq�}����!���vg��X�EI���ӌu'�;=�陸dJڝ�5c3+�ІrQȊ�ʪ�05����K��'��s�M^�u�� �2�M���B������Eo`�Y�����.�:��v�I����?o�b���H8�:I�%0so��0�,��٬v�ִ5�Mh��Fmۋ��Vw��^���L��Ɠǀ1���g���%�l�P'��1�A��fGh����q���Ǖ�#�|�Nk`�S"d�B��5���� �����8/�a�}��0�:'1Y������^c��qO$�6�i1d��=�z�� �i�q\�;&���q�T���-4�/�[�p�u�oO##ٿ�ojL%'8��U�Jc��n��p��(ՐI�Z$�� ��+Pj�ړ&��m%��1��'��7��U1u%$,����_��~��P@t6�VLb��]:Bm��<���Ÿ5��=��a�~O���؆�� �.7-��Q���`������cj�%�4h��9� �Ȭ��_q�|U�\���u4��Aތ��Z�^�i�A0e(�������'T���aF}�S���o
,�5�WJ\c��l�(=�F��'Q�!?��R�>�?��]�v���j4PG!�ދA�~�P�P�<bC
~�Ǆv�F=3�^�Q�y�����Y潛=@RO/O��^���)�-�&�h��N	�$����U�t�%�PNV��K�"�io���k�vN���3�%�9�����J"�N�ӷi�42�o����<���_xmn��{��y淋��,\���\�xȦ������,��f�{��v=a&�����\8�dҟI���yZ7%-1��������N	�VL|jVFlZ�쪕�!	����FE���I�ڂz������0��Wy�1#x_�p�S�X��lO��ٱ Bx��������::�r�E\#bo�]���߅���'�~�IF�6��q�H	|tT��FY��94Ua�>-�)%DP��p�2�,�A;�6�a������M
�ge�
����0�"�Q|�vz�7'���������EKkkk#[��њ�����zI�s��QL�7��a���2��룖��N��O�"��鶛\/�~��Fa��ך��*)>!8s��kG��'����VT�V�U9�W8?�gCtw��M���je����r�<Z����UJ�f�QL�o��Wg�o'O�.<�R�l��v�2(������K7Id&�[��?�U�h|- e�����Q")1���a�=@����ZNr@��Ղ͛��#W�on�+{� 7�5�e��B% /N_����{,-�pO�o���!T��e9�(���4J�x�k}���_�GkH���5!�Vil����4Qh����(���H\����n�����k���c�����t�z1��k^x���b0��Q���6u�I�ts`�r�B�1�v˦JT^Rqlm:����l�! _z
d���t3�`t� ��������~A0��U-�XT�T��C�6ӫ�O��BX�W���Y%�Q��X�X��N'���Bj�:���nui��/��GC�Ɋs0�t'�#I�?u�)�����#��F�4�.Հ��4��J3�{���[��h6~�Ǘ�C��i���wN�l�q�uˢ�'m�A�[�K�
��>q)@�A��` `�Q�!�'���y�2 �V����/�<��5^�CT#�]~���r�ٵ3��H�(� ��+R��yi��m�I{ص�Tl�J[함ڹ�q��U9���8�A����o��r��2��A0q���tM��L�0E�q��t� �AV�Ex%$ 222^^^0���.��6`3OK-�ʪ����먃�������^����g�m7se���˼.Bn��nV\�w�}���oJ�}�����-/�|�!jF�G�&�{
a����뵜iGUcPC���.4����ks�3���7��h��J[~C��M�9�s]l#L�EkoiH<8�( �/*�a#��T�e1ef9�<hnH���P �F8�������Q#�/O৥P�M�c�������l�[q}����Hd��U��<B�ڂL���� �U�z�y옅�
Oé&���,���"�%�o~������5o���HS؉�k,�t��͘|�B�Ó�M��1J�t��|�L,��\�,'��H����L�Sji�S�R5��c�����E5�с������{�T������]g�BlZj�,<�=auyA��xY��g�&&�~�H-�����k`�o_���t��\DGa
��oN� �dz4��]��q��Y�dGq+>2�	�?)�8�|�&T���B��p�'�O�)q�g�3�2�xm���ߞx.��_��;�lO{1+���L�]e����K�����Z�A�N�_�ճ?���T�j^.}�jŽ�M��
�p?f��kZw!��Ef[�:ը��g�/r�k�̢,d�|n+��"�ХUk��O͛d5$� z�������3��^.Aȗ���x8e��=D
}��Fe��z�E��\/������sΥ.FS�ë�l&�r48t�_;����|AG's/�BC�A�t��ZTb-�F�3��Zn���	|(k���.�����h����35ǱᔤR���$58bOC�\b���-!���N�Y�tO��+�����8��rI}�ղ2&�;F1 ��>�7�B	�SD��>�HK���Js?S�>M�9� ������4Y=?��~I�H߮M�-��p�����wTH�����[Rt��P��������IY��31�B����a���<r���H
�4<t$C�x�C�z'���_���C�&�t��//4��0/�)�xj�Y:�T��j�~���mP>Q	�!�ӕ1V�� \a�by��g��Q)�,+j��a�(�p��j�&�@E9�׌�fff�+�{,o�9��>5y���%5��]Y�/h5;�_�ȩ�y�^v��^�������ψ��M�-\]�������*�;��[��<κ�9o�����]x�q|����	�I�r�����'��V��o�O�y����g���b�X��x�bj|����rЍ*��Aߐ�')@K�8M'���J�; �y���ݣ^G{�P	���ԗ���L�8
1����������ɨ��t�����_!�H++�MG6�ϛ7�_�kmfXT�kсm ����1�~�1��z���u\��"�������=���Ak�)�ޜ��猪*�[�wu�e^�$qǁ�Sh���B��!>�+���B����Rdx|UY>�������R۾�0�w����33�)p��S��U����4g�5�/<t�^��j��:Զ]�L���j	W~����d�5�^�'lna���cD[x`pfijif�EbXjMã/�[�+k{+[k,]���ȊޱS�lg�c�n��t%����e���BUkuFt��R��Ʈa')v$�;�܀� G
�#r/;guϷ�=l'����|����R'W�§߅��_\1Kݦ ��g���z��k�����B��{���^�P��e15���<D���)�fPA	@О���p��Pк�o;IF*й(hk$�M5K@���L�k�d���Y�L5Ks52��<�W�M�#ځ����{���^�����j�M���gTf�4���7�-Ⱦ��I0���2<h4��G �Ak�v*�Eh���VU�3<=�n�qZ� ���� ��g)�ۧ# ����O�%v�l~�_��K2�����O3�'�\�����WAS�q��B�Ӌ]w�!8m9�7}�x@�釉�'Z@���ł{��-�gS�׊�ȉ�~}�|�a��x2`[��Eh.Qd<UF��.�a���}���=�5L�6��r�bI�h����������?��=LUu���qh
�I�Q��f��N&������Yt*4<�C��D�����O*���T��p�7�_(���.�����Y·啹G�3��o-���`L�L�3 #�����ߥ����7X ��-"R���&UU������Uo��-�C��Y�J��A��ټ�,�ov�pX��]�v��i�:�v?(~�a�{�cp5�/v�^�vc�{�t���{iw0�{�����{w]����4���!�	�k��G�O�O�U�~�lr>wࡡ}���K �OK=�W�ȸP�����@���?c�	���
�=%}F��

"]�1z8�� �4V7�e��d B2��"1�}��T\��F�pǫ��OSc��c�4c4�췓�g���455W7nI��|��ލ��qݝmu~Ö�%�3��
l��0nLu��烠N۳_�(?,��):2�X��c��Ք8� q(O�h�z��x�k�
�F��i�㚤��I��ث�*6j�E�V��ӌ̈M.��ccS`��%O�B]�<Y6�W֥ E��������psǘ�=U�(II@_eP����x�T�u��kG��p�P�?��*u_����ELFdh��~�Y�����]��]���[X��;��e�-�^��@����w���w�~�hc��8��3���[Mn����_�.<ujhbn0X�G������ʊ��~�7$��
Dt�:��ьs-/,���5�2���0��b�$VD�.�C�cפ�-�_[¢j��ڱ3���O��4�$������x>�~�|�v��Vj@�v��
}���p�Ww!�a~=<�sKa;0u�1���,����.#Xϥ�(����¥��ue��Eϰ�(��SD]Y5D��d��nNi���Q#�?��?�C��뼳cy����a�\���ﺑ8�r��o-���:���am�Z�;*�9�q�&u%�mHC�-��] �ä�Q{�Oxe\@\���q%��� ��ρ5����FB�'Xn5e�G��P��ϱ�Y�'r�����[���|y?��ߌ�U>�P��2s��i��pE��I
�Q����E������G�k̸�IIK.r�u���apY���TG��R���.3��	�}S��/����T��K̝D���O%�3�v8�
��G�W<���?���??h�b�-������pҦ`,�,<��󇨅¾q��XT(��	��H�G�g��W��V+��i9�q��ٷ/WNF��x��$S�5���z�G��M��7�Hg��#@� �����/�MbZ��w�
�?��{E8@y�@�ߞ_�W����`�zZ�ٯ<�g�����-	9�=�-%�-���{���D�T��q[����4K����[�x��(¡i��<��7�0y��i���J�+�"�;~���d�ٓ�Z�;���Y�(UG�b��sx�N����K	 �{2mD'��o৅����ZF@�k]X3�tQy�*��.D}28�%��?})�͠�KHh*0s�+W��#�fHl.ŽYh��_f�򓇯���|B-+X'��m�N�""V�V��EA������k>�R;��UﴼG5���Q	 H��2��\bׯ4�.���0L�f�����d'�Yy�;�#Dg�'�f>���v�.��[�)E.�O�E�ó�]�<�С��Z����7��$_�bn�O��<��hl�n���8�~�L���V������?kL}y���M���붻K��.��ŵ�����X>��ʍ-;���*o(Q���g7G]�g�ג�'���GJ�O��c<���r��1ë�s%�C�̂����$5#L5A��!��*�����ؐF1������1�PTKو�'�R ���m'x6+�I���<�\yr�J�55��o}uuskoMƽ�������g�7J���Qu�׭3l
g�	5����3�������u�TBBSr���|���q�􆘫sy`p�����ښZ@�-�����w�L	�`�Nq�lƍ�l�msG��rv��� <�{�j�
�B�����,� ;� �(*���'.��[�d�����m�� ��`��g�ю����T��I�-1hOi��?fp|� 8q��!fU2���:?}0�D=Y�P/�ϔ�0���*5�sjd`j$�����H.�('���vM
\K��oMى�u��v�����G�җ8$���ƴ/97-���VeK88���r;:�B��S�A�n��
�;���{;�F�Gǻ��R�_ͦ��������r��~f�%c��i����n��ҥiI�Aפ�b��AH	R���g�f���'�������t	��\O�NNyU���s���9�%�����nV�/m������,���jy�j������^�Č�<]���S�T(H�%G�(T��S�r/`�����Bc�IUg'4ј�W/�j�Toul�/���Do��v|���!����o�þӆ��d�us�Ry����j�5߿�2%>�Nl�\n^K�\28T[^�E��x��Q�'��)�s-���IJ �>c*�!��ò$��M��d_�
]�5����ǎ��VxyH�0Ru�`Ce�2�;���dK��e��C�)�E�_��xχ�u�k��z�{੭�y������?���s��p(z0&�L���qiy��D���k�����@��2ҳ��/�D'���<sF�9�S�W~�g��*X�ͤ��p����e��/�{jز�(���4�T��>������A�I@��v������3ds�]�Y�T�@��::.�,���Kr'uNE�J�jZϚ�hw�,�^ɧ�����B })�Bi0��������d4=�M�L)��a5��죯��(��w����"Jx�t�R�n4�qL�Ѧ��Vx9:!�k	wd�e��F�`>`��"�Dl���\�L�� ƨ�T?r�m��[<��)����A���{���p��]��m�3���+۸�h��d�|t]�N�l��i@+!#�L`"���������������c1)������;<�<�����U�~�6��2��p�so����D�]i#T��)4�K����e�����s�n��^������_����݉��U|��Y�����.��ο��U߻m��k��U�h�텛e�3.߫ᶫ�����׶�Sb:Q_���:U�d�Q���U9��Q��2�_��k�����A�(���S2��bꅠd�/*��!,�4}#[�L���;Θa#�=��$�f2����tǼ����ŲT�� %�J$g��K ;�<�ܛ�~��gf��),���,6�0<GJc�GѶ�Q:�m��K����>;U}�j�-a�3]�{�Ɋ��0j��56HȐ[�%J䙦p�SQ�����.[q��Dpr�wv���(�	q�q4ё,	$�P	��~�@���tK��EO�jt���$`�#�Nz8�?Y��i���S�]��8`����o>�r]�nR�n9q�ճ����ލ��>�<��D*N!�'V�IIg! jK`	`�F��X2G�GH��JV+T
kc�:�nx�!��7���`sp(�y�_Q�}��tv~�-,�Y� �N��,��ﴶ��Xrr� &D�3�QC�1C䵊��DA�]L]�8���iu��[�:/����+��􇘏�j�۬}�ڏt{Qj�g������X{/ݽ������U}e�l��9NA.�F��L�R�w�%s��T;�@Q����'�v�i-o�;P����&�;W'��YQH���6)�aa� �ɢ>�^X��N)�*���%
kp�p�1��^�u{d�ӟ�O ����_��������G�_m?4��~��ˍ�*�z��+T~�tyg6c�O�`N�v��:����C�p>k۷ �r�֫7��)PI���u�
���
���
L+�]�}��!�ru���tz�����ֆ�� ��_C�$�XF�$�s�0u��o.�81H��J�B]��cY���x��bKo(��?�%ǉ�-޽�=�#��!��iX�/l�Ҹ�#<5��5@�\��L��,��̜�7��?�*0�h((�7HP��^�~����������qN�(Z�j���R���ҽ����"=,��(��P	���Fx(U�DH���w�M�G����P(`�X�߈	8�t�}�?�>>ۏ@X3�Nl&��}��)Y�xݦ�F��La_M��a�HbߥBܞW�)�/���۽��������$=�ܢ�$�@�\�&�U��'�W�x5�fz|�R�qY9��\��b]��M�����[oUH������職�t}�6����Uk�h����z���)/'3���|;A��i39qS������ym#�,$O���&g�M�s���0��9�{~~���ۃ�������`e%"���ЊUQ�rs15�J���n�V��2��`|f��������ںT������x��=�nG���nx�V�JE��u�_���
����2��v���Mb��������w���Y���-w���3v�wK۾�'*^'�m��{��ב�w���sW�sE�s�^����|��{��ޣ����Y��26J�0/3yI-#��6(������� �R�"�	����'�}X�ێ�b.�Lj��={���ۘ3�p�J��W�B>?���HޟuX�9�G�F����h��O��4�h7�(�3zo��n���x��je%��O�ow��z��7��dṇ���+����t��*�
$>� ��*�k�
�D�Ε	r�*��w��SH�m:c*��9�Op���6�2t|�H9V��K4�ݝŋ�f�Y��W1Ee���Y�����	5�����i��%�r��pPQr3~��s�93���O�U<�M~�z�	wD��m�֦�����5)	�SR��6��OD������#�o[z2�7��Ƒ���P�<]LSU`QnFh8��|���|��Y�GZҪ�>Q��z!���Ȁ��;UK�)�^�[�^ٔ���l��҂�8~�KOuX�#�/�4m3N�n�gbBan�	�E����ǀϰ����@�4x��7�֦�,]����bUl0oo9ܝ9$M�rz���^C����d���O�!�̇gH� :�!�}�C��.�qn���.�?�;KA���zL�7��^�V(��?[��ݘ��
 p���,4� ��5A��~�#4��x~ ʶ����I�1S�T��4�F���=��6�WѴ����S��Á:�7Ϣ�5}<l�'Ct��׶�&��-���)@�!ԏM��fp�P��!vg@�+͘�ot&�".3���K{�K���W�3-f$�ˉC!�جo�I�%��ָ����R0���xp,�0�ya@�cQ�z썙Ό�nL��X}����XB?�	�_Ų� ��:��׵�eiw�z;���߰F����N�Ք��S�!�V
���K��,A0�h~�O!�����A\�bj����,)Y<���rd�K�^����4��'�:�T}�R;�x__Q~�r��M��"�t�.������5U�_4�s�2������e_��I�P��N|E������Y0>7�ں��\��EQ��G�T
��;�	�Q���$?<���\]Uvsg]]sJ3�Ze��/zL�]�ŗ/,�?���I-E�<#�sZ"��3t��Dʼ��̎��a�f��:M�;/K���\ח�|}�K4|.{=�ybi;�����2��n�����*���_��:���o��i�˴��m��rv-g�Y�;�i\"_v�U�w�]ߜ�V;mo1*R�%�"�+6�W�Ȼ.���������F�M��v<� u�dN`nN)�/���@�j��%����(�]���?�n��xeT����T��\��N��̜��H�7W����MC�����!���y�Ygb������'�6.ήMk�.�q��cA�dM��2�Y����H�̓�P��ɯJ�z;���?=��b ��4	�N�0M^q�u���}�U�2��7�5�d��ߜ0w+�^_���+pzu�vg8�F����L)�㊩����z��D}�Rȟ7��U\4}�A⍖Χq�"�ҁ��`\��\�&���{fB��c������r����0���s%�p�x�'-D����G/��������J(��?�T�hj���Y�ʬ�~��sb�Q��޼����d������qh�ۡ���������o!�_���|;��Z|*ĐN.�(�hd����6w
c?>kŵ�p�X�<���"M�����`B�!p9]���'�����cu�����+<�,^�/�ҳb#��������iI"X��&.��y�ڗ{��@�Q4�8��~���5[��a>gI����-*�K2~��o��bSt:ŜB碻Qά��"T���g�Xnys��M���q�����Ԓ
$�! �/U�aQ*bl�����^qtf)�@R=����%�D�u娄R��3>0q�dr{���Y��i�RI�^�De��H�3R`	�@�Z���x�y�O�V���,X��~�P>��ך�N�i�q_�k�;1�_`�f|��i6�)�sl�Qpv�O|���;�d�hh1��(��ư�۽P'Tj@�%��kb�(�4�:�>�ĖE�b�G��y��u�!c�S=�e�rcϲ��
���U����Q��QB���p�A|�g������O[.�(˴c𱣳��*�Y7:������SJ�E�yԻ�+��8:J)~�ޜ����~kK�3�q;XQ�}��������s�$m|Z�jB���s���r)��b>����[E��pr����N�c=oX�-��bN����~�n�mT���e��Uu_ۼ�� ǛYw�e����:e7{�⭞��:�_��t��&$&c�h���ע4�ͻ~3�L�����	���~�Gz�J>�M��=���1�y�!�|Zi��L��A���6��UN,/�׬�a9����F��c�t���f�ś�D�S%�~(Ch��Hs!5[To���0ǣpG����X�o� <��� �ς��wǺ;�Zn���^>H�]Rs8���1�τ2 #�I���)5S~w12v������� f@���Ws�^��;�n�*)�+;�&"�(��������{�5�Î�;��:y?��������dL�c��"�V6��I�2AF�A̸c��0\�A��	5�u�� ����5w��f��bKa�haC�+��x�b�<ނO ǎ�7-��O�޼hA��/-�x�&��T��^�o��Ɇ6��ЫHj��/����J��p.���wᦡL�ӕ̟�!c�M&�r {����|���  X���|�М&�����R�1y���t�A&{/<��?u��s��BܐG���S��
�o�qz��q��j�!7�y��p����e�f��91'Twg��Բ�bbN妙Y0��}�#Jv�#G���H��| N��d*�����t�˿ߗ�M`�� T�M�,Ju���[j �xW�B��g��M�MJ�8dǾ���a$7ݕ�v~��&KN���8*��o�_,X�{z�#��*�c)�wq<]4kOl��/�JDV����(I:��R7'K>r:����)������$������Ab\=���?n��y��>�WL|��@1��e��C��m�J���o��#Y�-+���z�Z�B�ʉM��Ά+[/}a��Qr�V^IU>,�|�"^Jm˹u�e��59I�������4�t�K
"P��S�������x�/���A�d��2vL��u�a�S]�.��k۸~i��h�U�!N@���먝��;����	ܩ���qr�u`R"�6�	�@����?ӫ�y󉚌��I�I.��Tg�Ϫ݈�`���2��^ܧ�}�=,�O�;ƭ�w�H��T�t|�.�LTԁ��N�Z��u�~����]��ٌpq��?t�ǳ�v�w��K����˹�bn�]\b�mwgC�n���w��v7�c��G�:h�h�>;�����^]h=��`w-;]h���@� ��=1�8Q�Y����B����I��'��g+戼ה��e�r��:����q��ema�yVx��s^�s֮��o[�ފ�zO�eЦM���z_�u>~��Jt�'���͠}���ْ�:.��8�uE}�~FEu7�[���j���.)�� C�S@�f�N����Lx!��T\2��s+�'}�b�А~�6>5��Ji�c�e���Io�'qX�lc-�aq15h�&:�4�=Ds?U]!��jS���M:;D�Dd�8�D0g�����+g*�!��H(B���ǣNE�ǅ�_���Jvl$�*}�K�u���tߩ������G���2�rA��?O�mS�I`/����'��4��1�<��}�k��[9��ԒҶ���l��.m?��g}��ug�L6���د߾�����;9�:�Wg�Z_���˧4X�0�,�ASi�y�3r�z=��t���X�����Ɏ���L��hā��*e=���nj�8Mr�Lӧ�!�O��<r����&9��h��z�gn�#ى7�k��Y3���3�e� �
�1\��1ǔ;�:eJ�^k7b~#0�|����Q-�wogA˶KШ����=�An.XA�0h�;��]�Co~��%n"�&�:'���Wh�`sO3*H2ATݞ�N��n�Fp�<�F㏌E��/w,/�+�$�B;6D:+��[�q(%3=�)��S�'8员>�3�WUl_�d���yS��sHqXb�%��_�Z�B�GLe�a#�z�H+�B���$yp�y0	����c�����TWc��OZC�>�Q�g��:���Ug��?l�HwH��0�Q��N��� %����N)����Hw���y��u=/x����}���sv^���a��f���,"���&"RF�t&p�ђ�wr�Z/����5\t���i��@*�^Y����&���÷�XS�-!|i=��<�JJ{��Ҁ�����������(�|�k��@T�-%S��{����M�>�k�6r��30^�\��Gh%]M�����j�3�����۫6bJT�#�PtUg��h(LNv�&cx���~�z�U]{��r0������lsu��d���+�<��XLy��D�u�[Q��W���=\�)����l��9��w����Ӯ<R>�m��~�5~���ͷ�:7;�Rw��R�˹_OԿޟ��/���4y��s�;��z�o����X�n��M�:��+1����7\�nt�.�թ�&�˖�dF� ��cÜ�y��%ʞ�q�?�v�d=�L�F)�Zc�!C��&��'@Pd�!Rg�3����B�Y��wI�E��qn��km�Ü�㶤��U���Oƺ���U/h���e°��kF�^N_I-�����`6���ȋ��E��j0L�ڼ^�ꯍ-y"�w0<�T�w�~s�LʰNIK��&]I%f��(����{T��Т �+���k��\��ë����j��m�'��R���ڤ�z (�U_�?;�h)`{��4�o'�*�W���$j1������e?�;�J�2�#nr-`ɰ�d�,Ȭ�����|LyWFZ2�{򏖉�y�:Z�l�HH�||��{*B@ z���ߛ^��0��G��G�������(u��5�Q"�L�]�?��U�TW�I�Cn��lHIW�]��������?�Nvy�B��a�g���ʙX��1U(;���/�^����3)�����3>�o�n.+�����B���?�5���ܩ�$mwN�/�z\�)��C}A(A�����Z7�L2�>��L���m��B�|;��S+��)ēK0/�q��doȠJ�qj��^;�C��-����<��nR�1}�;]����}�M�ut�ui^��Ʃ:w��d8�,Z��?0'/b���dD'�mOd2E��	x�VF����+2,��n%�vϝ�-WL;�q	�2��ڪ��V����ߠl��P�[�?a�z��~�h�-=�@���2��C%��c^���iE|1Vu�Q�ok4i�ʐ:tO�S��i`tdsG?�#z2Ӟ1Q���Һzd�ٶ�q����/����'RN(&�_�^p��4JT���]�������m��a�v�� �P�H�Dh�gN�l�I��"U]�O)	م��79
��P���k�^泅���̣[XX���׷m�}�z>�R)ޯ~��QZ`�(C���8�)K!�%Ɠ���7��mr��W8����&�^z�c�;x��Ta�۝�҇�p)��$Iv��7_ot���26�]�##�k�q�Ѝ��������b���.ox>#�r��^��m�a[�������@�ۡ��bhG06�E�Ф��-�\6VE�|�3R{̀,-��U�]т�'��l�U[�i�i÷��e��5NOM�05>(�7����z��y����Ht�*�u/���!Ej�_���E$O8����K�$�>i��z��Bb���Ҩ�7�)f��/�z[��|��%L��`�rq�kv�wq��[������[��}m��z)'2]2���ʬC�Lǘl����3�r��69>o	rO�m
)Kz=�w�)4i<��RLo�%8�
	Y�ۙ�tۣ[�%�X�Ն�3�^N7���7Ü̓����</'4�����e�ot5���i&_\Bixw��y��J���e����R�{��oK�|��G��_F�I�%�e��p��dxuLg�~����I����#3-0���������Z g`뢃�(�W[����R�#M:�f�i�ê
}*�O��;�4�mS��8-��b�a��
�ؾ���8��(i�#8�����t���e�pP�=�o��h�s.�R�j��^��:f0�'�D'j����l�����7�!n�41�ָܸ�ט��3ރ�����I�I!���G�`�D%�V�esIv���q����d���]QR�M��a0�gHp
ZY�����@b�1!R�I�@�=��h�P������ _�ٽ#��wM�R�-L�7��Չ�(�h�W�����?����2�Ѧr۳�Z		aI��'1)�@��I1�	a,�ҭ6U@��h�@��(,{gt�/ <�����_�R���$cwqyz(�2���s6+k�4�i�� �s^ 6��&�'&�K�����2ZV �����T��7>�ô�)ͯ;To�������x����;�V���h9��\�fL������Z�d�����8�$�*�&ǻ_B	�����ߢ(�?�ߌ�����Й���������(���������5��T�ps��BD��~W��4Dʘ�K����;)ѸZfJ���Z��2�\U��Q�#�Z��GCQ�n U���ԍ���$��WF�dp��W��ˡ?+��b�®
���^_	+/k$�^�}��{ˡ������+�� L�k��B�(�jwAs��S:�SCE�a&@a3=��`��y��x>��M�C�mo���x; �U�5��9��+�!�"��1(R���H.;M�@lP[J����M�j���ݱ��7C*,���M��M�����4^rzO?�L��]�36ߞ䍑f_��K�=���|9�k��ibu��̺-M��k~ү������ �ϗ;R<�:)���N�[ֽ��1����Be||�פ ��
�yS6
>��f;3�񦲁��f.�3呍`� �go�Q��\� \u����*��,׍e�	�#�5�*����B�PM�Y_h��̨�I�]����k�{�J�����/,����_tr�W2ӭF�p�[�5�<�V�~=���QB0O���憼�_濏����%&�Z����ȓ�s�u�^e���Ӵki�C���C��b��N��B�5|��|���!���;�y8��v������L� ��)�CR���h���:��+b�|�O�e�/i���b���xZ�Fn�l��@���s�>�o����p�+N\7̅���C��_�h�q�
wJ&,}�gn�oE�D�ܡ��]1�����Wk_�v���\��s�y��L.�-tL��X�?��К+�gI׿&}u�c�7�7!�U�J��jT����8��s{#�����`ȋŉ��)^	V�"�L|��-Ks���>֎4^1��-�-���6�:�5��J��������g�t���dF���-�/��z��͞��#Zc�dj����!=�|
���]��� �R�^�j6:���yA�t��&?�M!�n8���"A���V������B�|�6��E��<�+X]���$���R�@��(������}A�>���,]����p穑�����}Q��/Sa���&�7�|��GJ�Wmb�����gm9VH<�.�]��k�Saý���̮O��4}���:�U=t�y/�`?� |AL�����4x��ٞHt?�pB��mv�`�*���c8��Ѳ��R�_׺!�2�.F	���z�L��[��:�*�������'j�����3=ϰ�&>	j���[�gM�Y,P�#"�"��Y�
v,��3^/&�LcTʰ���<oy�Ŋ9@��"yR��g�
�f؉�*8*�:�a��Q���,�����Q�nSd9){����ݢk��]��J�L�M�7x&�N!���U��~�*�l�fBc9�0y�H1 ,"�R��a��[�d���j�^�'�<A,2Z�˖��S�K��ZfZҧ�	{2�{d9w�C%Jؐ!L܅cF�3K�i�ZKl�&�G�jS��7��뫂˺�η����*�W���̏ԫ�~�w��z����W:�l ���"���^
�WV�9ӎ���N�����3��c��$�@�z�W�B�T����ɹ����
 �'��.���GX%�G�I{n�t\�2�.jxX�����[T���e�·�1ݦ/����bAoq"�3�P���c��m���'�6��u�k�;�#���C��SCF|I����Y��VD���N�k�S����W�O�[�n�o�����,$�&��e�:������C<3\��7P���&G�bH��Y߆?�K�ˋFVQ��^NKp�[�Kwi�=1H����S��N/���t�o��$�32�F�8�6���;�qK�w���p�S%�S�Hx��BC�)rr����t��տ��Y����䌊�S�0��f1�Q�tn�<�4�jl��K��<�/�c�a�B+ǽk~"��?��ڝ�[ϛ�����v�����uj�1�9.���O0���7�c
�J���]B;�qO5����6�)}T�$Dg{��:0�����H�Ҍ� �׼G/�JF�k?l���!�s$��%?�4�*v�y���	~$�LA����GUs���b���8��W����&�J=铴�{�?���?� =�M��t��\f����'4���ZԾX��&{=� _�H�0���^_������k���á��Y_pZ�V�p���������R�z5�}	��\�[���283�i[�A��ь�K}.�Ӑ�f�ۜ���Q�w����W !�l�~�:�!3Q���l�a��ɶ�g��Z.;��^�8 5f�a���/���fۮ�=�V�2-�e82l��������v�G��HU��c�����
i��[m-&��ĝ��vX��f�l�ǀ��Bn�On֊ ��;>���P�m��f���(����.%��o��G�1���-����K�E�c���1�IJ�m28�;�k���+7<�`A[
�V3�~�d����T��ytb�(�꟯��Zq����Εw�E�AӆAh�<p`pa)���zq�1�1L�}��~��1�@�p�EJ�+d}��8�R�������l�H4R��
�V���1�Ɉۨ�#V41�� 5�ѐ��� N���E:&���)�ݹdv�������Q���_&��6
�-���x��33�k�6�r;�굷6��~�fF�mu�*�$d:�ؠȏ�4B� T����ggAE����N�,�V��B䰷\�7����;��O������zQ��� {ٶ���0��;߰��o��`��~��n����ţ$��W@������߽��7v�~�iG�3�(���n����r9����_����QIZ��";8o?(�Z�9��	s��jv� ����}p�B9nGf�]8N�<�I&n�����Rk
��ٸ��:���Z���0ܙ�J����������[���<�J�n/�<.��қ�0aX�xk���>j�n�R�c�a��ǿ�i��g�����0)2w�����f����Oܿ���y�q�u]�qU�p[��V����A���U]Е�M�~�@D� ̆�O�f�9�v�9��� ㄂�x��FV+�jeM��n��$![z"Sx�K4����E��~WW�>�d�(NE�g�j5��5�rN���]':H����E��q5�Gu	�E&�H�V�4�1�x%�<�=]y�������យ6�\�Sو�,	��욵�Ӌ�,�����lHS��y����)j�,���Fc�>��S�nq0���b#sSh�o��.b��]�R����=�?W���p��k7�i���� ��[p+�;�}
x�h��ǿ^��)�.=�d� �98��f@� %Q �Kc��=$�D�m��:y�����!%EQf�^�i���-[{l�f�&�m3��L��c��{M_�L@�� ���GÅ��Q&�Ҙ�����M�b��EM3��L��zՔ @S��1��[�J��ۉ��[����ZJ4�|k���1r=(�� �_��5'e^�\��o*o���݁3�W�\�T5�I��-X����X����-L8�W,D�SC4� ~ ��bl�`^��z�<O4t����$�ի`Lb� �@>wW��Ц�]!�CV�1ic�P��Fz��0�0L�<~A�#O'*WՀ\?�r���6�NN^v���K3��s��c��b��g1븴L��Q��Mž�� 3tů��/�9�Y� �C�<�ɼ��y_��3U���`�H�J@�D��<��X�`ny~Ťp�v_���6{?�\y�|T�)3h��cMӡ�O�W��L���'��⽎iY��T�e#+�Ţ��W6�$R��[�>8..!�������Q�k�i��p�[5 ���Jp�̣g���(3���87��xu_�(�$��t�
+�S�lE�(g�"�N���A�؎�W�G����'V��f�`z%k�zJd�x�&̽� H�t��N;��1�5�O�ᝪ�O�[�rs>�qR&�ԏT��`^q����n8N\d�A�t��?�Su!���Sh�����x�>HMKM��(���� KRR\l�|;�1��H�ǔ�:e2� ���ɡ8ԧ�K�/�~]tr�$��i�B�X�$,��uz�Q�h0)�*�jQ�:�������85zJؕ�y���⪡��胟��R�^�Ǆw�[��?�e�L��8��*�%�l�.��6CI����9��H����?�)-��c4.�8��@�~w�b������ *p�<]r���zѤ��������!�&E�,+&�1tU�p��AmH���U �7!���p}�z���@��zqq�a�e���c�I��r߲�Y<�vc�s��o��ͬ_��,�N,��o��N�o��s_��V��#�g�����x.��o;wai�`0Vå:_�gf�@5��3�͎��RZ�z�}�q��Vk�U�ܞQ��W����p���կsּF2+�s�q�ze~'�r(�z[X���a(�����J��^7ѝ$v9x:1p�N8U?5�m�2���`5�3n��v=G<O�rv's%A��hpi&�Cֿ)�<��߸�;��2�{(�b�24ca
/m"�`!ğ ��ֆ=���n���+(�m���>h\h� b�x3U@����J@>9AOyܘC��o���޸�:1O[�j�8j@s\R�E��pQ&��d�'��ĬD�����c4�� ��c� uT�X܍m�.�7���X��'�LIQ=P �ح�ft��L4 Fo[L�����e���%�9j,�~(t�+:@p��m��au� ��ۜ�d�����>�MW�jb5I�q;�I�qS!n��ɤ��OQX���L0^H�ͅ�v��
	Aw�d���a�v��^3b�:I=
/�%F���I�Cx�d񗹤���~J�~y�	�w�]����d��]T��t5�ZG��6�ƪ��41-�ڮ�������Vq��5�?%'d���B��9d;.ެ�5315��-͙��x�e.�f�en��w/mb�i��m<�\��x6D�|��|���t����d6����:�w��6���^�xV�O���?��0hż��P�5��3ȏSױ߫�@�(O�&
t����Icz�e�l���8��v�Q1FS�(��6�ɺق� E"�4E�|\W��z�Q�F	��,�� 8s;�B��=E�P��!wɪ��J��I$������5qq��k>��"P\�A$p�^[�%C���vS��K�cI zm�B	���`J�0��!���F8��;1��
���]�2!�ڣY;��X+�~��N�DpR�\�� �{'��(���\��w��]vt������P@�_��g����;?Kh�Fr��ل����Ӿt-�zo2#�9Q!b�ZL\�`�L�m�h��� U ���§�<���y=n0[����1w���>(<����T���
ZK}/9��%Z��o��vz��-�~��/�	��?�FF��!���/š�, B����*sE,�m�B�;"�_&S�<[���u����n*����#j�m�V�M�|��C��P�����u���C?�>����\���d��)%��m�˼M�K���rQ�h�G��D!xݗ���c���`�x��:p^D�'h�%� �S�B�;��@gc��?9yP��9��ĸ�AL��+6|#���H	
��>kw����[�#�ړ��'����I�A�IJ��1�x�\Dt�r�=�kC	:�3��lD�7�5��븃G��y���Ҡ��QɈ��mg#�7��i��҈^Bih���($��9��fd�����`�g��Τ��%��q�6�1=C�e�#5�ʋ��W��t�q�g���!���I
���i~�6�lt�A52=[���mި2�;1���}dY�U^��v�l�R�0�H]�"��(�B��a���b��c�J���U 3C�R��Nڙ.yY�9?�Wȍ�|.J�%����g"3�{d���Bs�mp(�����a����s�O|Y$�uqj?y���ӛi_�M�?l+F�6��`iԔN+���[)��Ji=��v�������)^	gD�T'���s�K�����Q�.�I=�`-�~��e�Y��x5�XLL,$��L�$�R��k=��3p;�½�-d�gz�Y��������f��ȥ���߇�c+lnv��^�W�JyG����ѡ託��ng���V�V�-K�똳`��r�]�(��H)�l"Z[�F^�@CLs��{��}�ڌ!�\A{��:RX:xmo'�z�2��{�O�Gt0�h��ݘ&�r�ȼ��u�J�s>���^��n�\R)��=�dK���S0r{��^�wxG���^���߼�����H{]��<"B*����k�v`��L�M�I��E��Y��:��;��r�Q��;���svf�z&^����!;B��&�l[j]Z�t����	����t��u��}ڙ�g)��0�����m�ò��`�-^��@b7���0�L�����Fz�V�t"MA�->X��������ZZY���겵r<� <@2�4�ǝP菚����g7�,X���l����Cəd&����%L��=�nL��!�"��4�q�M�he�~Q]���p���mHLu�i�̐k�����7�j�ރS�Ɂ~}pjm����yߓ]o��HEr|<�Z�G�+��g'��CXg���A,IP��������m�)W�� nV)�E�r�N�����VE�O�i���8e٨�O�&\���i^|)y��o5G>^��L��]�l����{n,�4���@��P�-�-@x�v�Z?AL?�������P�xaX= @ͪ�Ůe��Rk�[�~69*׮u=by|�����T�G*�8B��+!(����̞d������z<�ܷ�\�XXJ�n=�1_c�C+��I`!�Dʒ��F�[����
���@`����3�=[���2nj[p�E&Z����(O?#� ��g8� k�mt��s���B�z2c/���������ѲT�?�c��nc/���S���Fȭ}d:�A?^kM��Ǵz)��@d�n~\J�� �~��6@۴������lG��'lVS�^Ԥ�d���T$���O��1[���$P��^nO��/�������)<؇�Q��JӾ^�?Зł+Z�BF;�)�E��3��&��lQ$|������CJ��z��b�&f����ȟ1��B�HsJ�>اOM1���3������[����*�5ޡ�W��/���^s�TeJ/�_��;6�506_��>��8.>�3Jyo��{�"�=�}�6���!N��Z�S^ �kDI�gg
�'&$A?	nxs3K�� �Pg��M�Z��6��\�5(H���M��X�]�L/1�N��������%����T�)�5>S�C/����nπ���]rK�q�H��z�y^lV�7.pH|M�{.��/�enn���r�#l�+�=&-M� $��Ȇa�	C
Ă�z�z�8e?��T���	ݔ��-��55�@�G�!�;���%�Q�y�zk[�����G�z'`CiB���6��)B�c���05(�����)<h<�$QL�N�Y���o-X��)��TZ�Q=�G'��#����$�����V[�-ӿ�W����T�>���;WTz�Ip��,7���1ۦ��4���g���z�8�x�A�1���I��x�2!kKנNwؽ��ة���9���uG�$���ΧJ�����j&{�b�	�S�y]��1U�U�G�l;쯅y��g��^���`3���OV�,,�M�iz�3��^��v������éR�S^���Z+��-���N�T#-)z�Z�����}�;��ը��zA��NK��j7W[�(	��0k���u^UQ �D����� �H6�y�?(\���7r�.���a����S�Fw�F�����4I���Z���C|Ү���L�X�ͣ�;�����):���
�ۀ�<����/�g�f':�?g�]o��u��P4��N�q��0Tp�M�69�3
w����;��f �JOq@���z+q4�>SQ�.���m�L�8=��&����cTU�"&����/C�!���׌�7�!�&��������P�ZXm$�F����׳$� ��"��v>��%m9%��EqO�je��DqO�S��:!y�"R����[��b���>x�N(l�=)C!�7����:Bb7�-��53��ߴ���[�A|
8�d�pY@*��&J��X�J;˃A=?����]හ�t8�����*l����U���{D)3��C�� �CZ�_{n�����(���$s�[{;'FGQ�V�Ⱦ��H��Ő��wq6��3s����b ���y�PSz!ᱵ�kR{�Z��{�S���-���i�|��nL	��<J#���l�o�7�(�[�&���{9����l ��?/$��E �=�J��������x�?:��x��@�����o<��w��e�1Sd�,a��66bU��CQ�O����\�����9KT�䣤5|�wq�C��N�e�T�������勝����P��.'354S:�L��
�n�E`$�W�>AI��>���	ܾ����ѓ���f�LD�y�1�)�cô+4mĸ8ib�(��tb���
f�8��I��L�]4�nz��֊�6������,�������RϹh�+�TS��'g��y��f�9�yRJ�/c�C2�30�4�E$2�f&]-���I>u���Ԓ%�V����%��<W���Q��m�r<�az溶���R���d\ ��j����l8��>wrg�O�_�;؞����^�+!���g��BH6�bzX�c�{�=N,OJ2%g��+O1q������FI���ϟ�H =�w=v�(����v�,���ۛ��2$^�����h"�������$�x�����$�F�!���}��;,���Y|���J7��Դ�4�𙺬O{cc�*��U�/����l�4��n��ԫ�I~.�[M��Qc��������=�4�dQ�R v�}��)F>����j���I�V��d�r��u��I���Nq,�SQ�~Yh�ή�,�����.�U_�K(o��BÙ44BZQ�*�[������8=Ĵ�3\	Xi��v�`]$�ޗc���e�V[�3���Y�.�3e�\�Z�L5���q#/+5t^h��e���$^����k�
�ꐅ�`<�[�z�/v��=U�|����N�M�S�ZD���Z������=����_��~FO5����nT���9N6{���S��7�7:�S3*��0��ۭ�?R1q�(Z���&�`pz�jC;Y-@�d���$k�-pp�a�d�����6$����<��NZ�
*����a��-��F_������`V�\hŘ������xA��-��:�|H��8\N~�=h֋H�����?^����� \q�w&rLؔ�.�F�3����L`�G�o�D*^:�r�g�趦QAt�	r��f�gTnŋE���i�Typ��_���ۿw<�u���!��'U+����T��m<�^����3s�I]P���;�#ǖ N��u����|4 ;��..�%�_���;8����Xe��S���QLrV���
v8	�ml�� ���6`�S���;�F�N7+��F�"5��ڱJx�L���V�^��f M�����8Z��A�hzr��JrK���a�n��l�����ߖ��Mf໡�d�&ou:B�����tLG���P�n��~��L����$�GN�	��j[}��)���U�ёWi���VfRD�AL�nzV�)�r�H��j�!���
��~���m��ғ�����ۻÛ��2?�!��n�-�<_�N����u����O4��~�ݏl������#�
t|:;�8%-u�tZ�����!�n�z����a��e�Y�l���̈́�>%b��/�n^��f� =%Mcwo������FM#���4,�pT.k��L�5��}>J��|��� >
����g�_�`Uo[Kϛ���uk��OU0�_�Ae�r��߶�C��B��;	�//N\\����֫�ߓ�s�,6�o���)Z��[AoN���w��PSb�0/=��z>v-.\jH��RbR�t��_Z��m����H��3�ˣ����$A����5��"5@��l>��힨�q��qkS�Y���,�h+*���I��W������廨3��3����`�C��,��J�Z�fb{�L	>����7������|��q?۴��5c�v��'�=��'��΄���[���R�Ϊn0i"�`q!葜���ַ���"�,���L���=?���ө�]�0
{c,ս~穱k�t�w��V�g.e��U����<>c��m�Y���.v�@��$�l��[x��Jd�ԴO�/��0݄Z&~)\y+`�`x5`<�^��lEa�P�ʛ�drY&�o����7%:�-{�K����ާ��K��q��,$ֻ������Aa��$�v��2vj��Xe'���S��(��N����g��$6HX'�����}tAn1��e�k8�hX��y�2�s��$4�i���b�n�h��}8�E�&�&�X!�xn".,�a��ۆ>�>����C׆�����js���Le���bZ>�2տUnK�� �Ӥ��~�Ą��b�tZ�[\A@�j���$U@��N���L�rƄ�9d]�-a��'�u�ԫu�.2�g(`�r@w�3�D��oK�[�; M$�]D��H
���S��4��Na�e�g��8��k�N-k�r��oyuv�[�����g������-�r(�[7�cBC���-��x"�k��6F�hLe�dA@2�jZ�J�K�`��H8�L��q;�6��K����g��H���������R)�R��o7�03U�w�J��Q�w.M�!Fu��(��H9�zHE,�ݍB'MFG����,��@���L��O{������G�p�J:�H���Gx��",��:�+��7��Nm�8n���CPݮ^�0{XB���/���~�+J6'�"����K����t|r�pp̐R6Ŵ	D� ����:@���$�n^vS�@�J$<D�F���zj��y�M�ز������	F�#d&%j�̇@ �^L����b|�(�����gz�ep���E/���'����W�+bN21�p���[�Y��R��r�vv֘��]?��)�}��#��D�)omF�z#�39�gr��SΧ�ņ���'1�5���ے������������?9^�E�������fWL��KxԠ�P���VX�МE�%������ʱ1lP��(�$��M��fYۧ$�v�2E��՛��Y����==�����E��N9���ro���Ey��c\_�!r�:x��]�B��T'Y�/���㓡��n��c^�]�	<)sվ��-����f���BC�SD]M!ӣ�B�ETc��p\�$hK"��d�m�jd�'�s�u���H.��MUy��R@��#�	�	B(�{���&�ȃ���A�4Jh���w�Ee�Yy�QE�9�Y�؟�95���<�g��M3u��Ф�wY\�$zʾ�ݖ�@���	�Ǭ�ט��6�M�<=C�a4WK���QqhJ�k~�Jb�l�)Q���#�����+��t�g�k
8�ST_�?���w������u,�#��p.]�.N50�����ɶ1/��5��B=�M+g^,�3�\�H�=єa͂N�ߪT�L�,�4��kqG3��4�<[��Y@^�˹G�-�^l��_�7��6�D���=���'��_I�6n��wC�-Hw�k6�̓5T��	�	l��nK:���(�C���0���q:��dha7�^��`GK+M�(����F��_��&d&��Jl����,�0�ɏx�H�FSX�(�������)8`d�+XC�3�(��.4�i����<{��J9�ٕK�������_sآ�e���q5^�t��_J>�AY�b�t�Qo! �>�{��M��h����j����x�[�$r�k�˛��R�g��.ChY�qϙ	��G�4�� 7��f�g��@��2�p0]�)+j}\a��n��~����f��5��]���wD����ӴL��Z�MPV^E�5p�G��bJ0�=8 �M֌�@������6��/1�[?S��Z�{�(��o� 'M�g��&,�o�'��B��=p�8�q{�]��W`��<?�i| �B@��%�ǇA�Da�<����2�|����+������J���v?� h��F�_���q�!q����kQ������B�~a�7�?��Ꝗ�Ò�(h<xF�U#-b�Ub4���/�t\I�v)	!m���K�^�$"����D���Cv����Q�T�G�$��f���9�`Э��0�_�g``��O�ף��;/rPP��t�ն�2�0���� �S�.�ۯU��
]~����;T��4�Pwh<��Z�rM������N%QΖ�����l�4�a�_���ׇ����'?��6��ğn9 ����b~��Jc�o&=��G����2���>�oVN-�0/'�$3����H'�y�?}5 ��'Ώ�
�6]�j\|�6��£'o4�nr��(�5@VPN7:Ǯ-P���_I##4__���#�?�W8���s���/Ty��W�^��IW4�n��sRb����7:��V�߻�;ת�67�����v)��Wp�l�_[O[9ILp̧>�/d�x��Cg(��%�<��}�+��j��q#�� d�#܉�#��uP����E��� 8��xE�^| ���P�ɓ�R��Q/�n�X8���LڀH�w�N.u2���Y��w����RdDM��ByU���<���7	���,tI�L)-����4�Ԣ�Ut-w>���)�;]����=��e�����u�ߑ���u��y�1K�*�a�=�2��z�N%����{Q��7<Q�ݿd��?`���?|H"i�*LXv�G��7d�h�@&���x��T�j���:�bY@��Rz����}ݿ�Ul�����t�M9�Z����8?�Tie
�H;����u5�(����U��;��K-2h�~y���Et��(���=�rb��[�Vl��s4��n�����R'S��{h�[�AЈ��M{	����)�n��6�8�,k�v�;��A	Aׂ�P�j�o�d��rl�����zFD�f��^|��nk,��a�|� g�8Йa,+):��)��0�tk�=��ӳU�h�(q�k�L�~���))hN00���F�I�"�n2D�qG����8�TXu0f]j1�h��c;@��������HW����m��L�{���W�Q/~��B32ٸ�h�(&����J�8��'�,Q���Ɩ�b���GZ� ���4P�s�u�AT	� �\�3(ͷ��|O;��Ϙ��_��u���D�"�VT`y���|
�P'~�)6G?p�&j>]Z� �l��+�lQ!	�Z<]7 $º���*�
�2_��gX=��֛'+��w�����X����O�������F�x�Q�s���CK���^�8�Is�K��m[�ѠR�f�-��
��F�q!���89+LM ��<��1��������m��ELO�'���꯾�E�P5�����-���� 3z;�� Z����T���_��?�����K�ޏ����>O��ū�/��f_v�ɻҜ��?y�K�}��kx��K�v�mf�����>3����~#;;��ɣ�`�	�η�u^Ip;�Y�#g���zH@d1z�7f\m�l4���cw���'A����Q����W-5�ή(��o�b�v�����i�T���<���~yh�s�԰�me~#�q��T��k�ת�^�DO;�T�v-��K���Bqq1�Z�U��*T0�i���b
� �2�Z�T(8�D0YS1��GC�w�ֲ������7f�N��u^�vd��yV��O��O�_��%{��(�r>{~4�ppLq���"�Zy̍I�2���8�~����5��s�sfū�]��8��)k�7K_+�ޱ��*~����W��+�f������Z���{˨��/�/�nE
ŭ�;�@ �;�B��R�iqn������ ť����7y���_�����Ξ�7י{-5
��I�b�b�Qe��N�>y�RA��M��'P�6N>0M�M��+�)n|�	�q^�
A�*^M�mhV(��"ӹrHDT���n��sLP£)d�ă�rȊ���öY�Q9 %�JWޅ�3t7H����΃WA{���[�{r�m6Orm�:��-�/H`V�0z�v?Y[�x�̌m�>dld�8^���b��Z� F O�E����@�A���x$"M;��'���:����]��N�+���#J_��[���g_-�1I���k��$G\� :W�?9�e�Ke&�d��<�l�墀�)���!��XBV�~[��蒎�7\n>,��hXۡ�Z�4\�Fk��t����a"ݻ�$�¸��N��:�/��a�h(�E�C�'i]���˫H��b��G���	!SPzE .�EA��{w�&��p�>,�ח����Ҳ��mǭ^>��V��*�q���K�-Dwh-��g��n��� ���j�tʅ�%���6yo���d�G��mJ�	;�	��m$�P����8�]��,F	@�D̺œ�#*��5���0;�z�9E�:�`f'ן����½E������pv�\�!̩��^�	�$��_��T�6bp�Sٷ���:/���Cq��褶$;;�����	�s���<�G3RJT*���U�"�wv(�lw���r��9A�_M/PM暝W�=�iۂϲ�}���/�W}7?m��������>�b����'�~A��ݟjtݜL�v�,�4ל�uN��%M\"Q��>�10�nW������T��M;����g�D'�E
��Mn�5�!�����d\W����&�g�[����Cp�ӳ1u-�}�ir���j��&_��qg����+��(�	�}_AS'C�I4�������x k|���
4u*���&�^���t��GC	@����3:��޸5���E�
EH��\�
D���_sդ��5���H��ҵ	�) F�ˣ� �
�Q��#��:(�{Z�̑�dЂ�`�a�&'b������ӤS�W�~%�����\���ۜ��%���*����g�G�=9��Z���s�!(K+��6g�Eg��g��:%��2������i�A��d���2�W���E�����򸴘�p[n`��$c��I��)"�+b{�xv����p��3>@C�`��i���AӸ��!\ؿ�@5�$q�*��|?=%҈1h�t5�y�C�σL�`���i�	����T"����ww�/f�� s�r�3���7���ǥw�Gɗ�:��bܤ\��R1kF�����1�%���c�F��c�]R�5J|!��x��6�5)�D���T�^�k7)�'A�q̓�)�Py��$�'f���h�|-�"_�M������=K��¢HW�D��+/�b��.�4)�6m��ֲ���S�C|�n�"�V�}W^���	�?;�Eٝ����eu���Y�v[�h?�1#�Eܺ���28'Z������[�mSi��V�ZKn�[^��9	������po����緸B�g_g��P�L�ATђ�s��m}��N���u�����ޞ�'��`�V��"��1�B���{�Ѿax0Q�"�!m�D�'��Ņe�d����cn"��+<�wм,�q���f���T6@<G:��:<Wr5����}_��u��­_!<gh���q��h=�}I�Dr���q94�_�Ij	�
����tI�Z;Ț�$�ƴ����$����tz99�Z^���L��+HHH &&n�"vw:d�1����1�q.�n�QP�*��d�R��a�hJX�S�v��0��U�&�b���>2� 5�����wOjn�����p�l��7Y���9G��I�A��W�l7�(s&��tո#(�d<ҵ|vX���!�Uߺ泡3��*���W1s�6����olKlU�o�%��N��[$��H�F��e�� ���)Ї�����ɺ	Q��R*������H�>��=K�"$"�{2��k���\aǶ�߾̨����6����d���	�����+4kU�?r{DjS��d���L��H8����$܆-0�}WC���IZ�o�?Z����r�y�A�9�W�W���l/iP��AZ%3���A��0\�(�p)O����"�L����f�*AVt�Ta����w>y!��d��7S߶&��r��ƺ��.M��ffٌ�J�$r�4�:���W�<"�_�)�k�;<]p���<�|�+Eg�x�����J@�M���	���ݠ����T�;4�����ff6��eW'A���(Nb�b	�9N�J�bG����	V�s,��qy���TA�Z:����>~0�6Q��9\\��:ؤ�0�p]��.���F	��_�&E�R<�x�;����f�8��s_���%�-����q����(��b~�t�09��H:Pm,�;��䒤�z�jǋb(����8��ʆH4hPg��ӭ}q��A�>Q��b!F�@hhشX�i#~�l�r�	�3���e����|D̀u�[�����+���-n-#J���L>�mm�>�`mJ8Vd){�i��USS�i�Q;W�\[$�SV��(bLY)
8=WHg��M��@���	�*��L��ಚ9���j-G�3���xѤ�*�U����z�>y��ű��9Ǒz:�Ћ ��f����L�F�HW�
%Օ�c@����0�ϙ.~!E��:j8\&zi!@�H��Dm"�~H�E�����>M^�i鈒'�ItXD:�d!���]�Y$w�#}C��D��*6�C�Vl��7�L8=I���09��)�m��e�����]c�_t�A�axO��c��������XO�d���aP�?I4��5�v���*�RP
I(E������R@��V�V��?o��SSg�����`�����Q���f �)�M��\^^�5]κ;91ڍ66�򛢎F��n�oP2R~IO���MJ�%b�d)��yO*O*챳�,��4��ů.?r�+H���\�tR���5����������$�E����೫����E�������L���6��?%��Gh��V�ޘ-%5�-2�H~��z[<&	˚��C�w<�L$ }�r�bo!���P�|ژ���آaB������A����m"������§�D�$��&�&��Ɉ
�� �V��rq�6[�21 ��H�ٻ��٤d�uF��΋���y9�� ��:w�P�����|O��"�p�Z�C\� *��ދA���6�����*�F��v���K,��:�U�F����|ň�.YFJN�O���0��dz:e�:�^�;WW��6���pMDUű�	���ɩ��#�B�0���m�̶rWͼ�o�Rh-���1�Ѐ��@6�����+z:�;];�(��&�{�
�\b��F={��z�}��@������{��������~�7�cG��4A��ly��Rh���q��O8	+ ��j_��s(��ц���@^ ��(v����fkj�r2�� �]��ʺ���!YV&��o<[z�w�w~<vٌ��?���ۈn�����z��)�,�܊����}���V���Rj�1���a���mM�T:ɸnK4�>/ �A�,a@ڧ���D��g��f>�����
�����<�� ږ�ePB'�CfB�6ଜs��z�O)ONES� T���h9C@���\�?i�~������x@���R�5���1T5©>�EN�%����O��,=&�"�
#�bW�M��B@�7,�4�T�h���ؠHRɺ��@�y����p�G_=hi�>�a ����Q����7Ra�� �Hb�*-j,��`%�(���pa�5W�HX�c��*"�F�fW���n�e��FI�%	��G�v{d3Bu����f��+�O��{�I��08	�����Oe�N�{h]�}�V�81-+��O��=L���FjU�kR��'/�@^zҾ@0,���}p�=�}���Oa�d	�ֺL2�84y�o ����j�<6Ij+��q�4M�+� ��#���4��FL�Q�6����M�`OO���Ǆ�e'G�aĞa�x����%{�����npӊ��؟�����H ��q�&v�  ��0p5�泚�y�/�y��jcC�U韮JQ����6�lt,�$ݿ&�O�ؤ����^�*��W���
r"c��z�km-+�b�VI�=Z�K��W6g86>s���ێ���AH ��Ȅ���t�օ�>���e�R>�Q��7Y	:��4[g���h�`Y��xO��|���@p��Cfk@]:�}��»�X�L_�����_����'�mf�!�o����=���aɔ{�IEҺ6햐�����0:9��T���fS�Ib4K�����.��%�h��j�P��<��	*.0�8�� ��L����F��:2h�|�˰(�)Zi��z�(����TY��4�vu�=c�IR�}
-.q��6�������/Y�a���~�k�>��������A����:�yz���>�b�ƞ�J��Q�Ԧ��ѵ�����HBEr[��.�ӈ99,���'�c���Y��_�-���/���N0�qW����۶ہl��-|�q�sY��_?R�k�v�<R�{� A<�-����/i]ն�=Ç�����gю����-��XG�n��P)+钻�)I0�4�(�Y�'�2I;�S\}�uk<ì���&*4Wb��J*g�H�]��<��3M*"Ŏ���x�Z˪�I�ՍmY@L���q���s=D�b�2��J���$����IL`�0)ֆ~Fx�(�M��dx�v��	3{aR�������ʰ�hݴ��D���_�2x���T֜y����K ��u(:�i�P���a/�)N��	�����Q������h�B؍�i�����z�����擞�]�П-J�Q�ȅ��mW7[l�E��F�
��z��u�_Y,�2�2j�h�Z�SY�ӏk�I+�繊��Ip�A��v������$9�Hg�K\(�ҕ(��^�'3�B�������s���c�)Y-�'D@4�����w��8�-�E{���Y퇌�]Th����dh��Q>�仞ZJ^�fy&��)St�7�W:'�:8�ӧJ�q��g�L�D&��9�7A�><Bφ:���ӎ����S�-l�����D��($5���(��Q��k��R���0:�2,W|�����L2I��v5�%:����o��N����h'}��eU�[��V��Ϩ�G8��K��q�0���;��� y����X<̆�H�$y5n̖�%^��m�7-	z��_.`
O�����46��
���������������{�%y�WY]}}]"c�̡��܇L�`�>��A&�-��N���l���RR{Dkə�z��AcPk2v��MJ?G�k������P�U�ǳ��.�cB���~���ST�ڽ;���O��g�2���+�Es��=1����w̙?<h]��s!^���}���z�#����q��8��|Ff-]Z�%���Џq��W@M�IB�*�����:�3B���lJx��uf�{y�]����������żݝ6��lV3��-������(Z������$4�	�i+n��E:H�c�&�T,���S�噘�����}FW��#'^OM;��G�����&�шI����u�8���|�6*_!x��.�7y'�MdRm��@ ���e��x��j�-��{}��C��������d�xq��a
N�n�,�n���0eL]}݅�;��S<�(B�b�8���ħ�x����?{|&p��C~�R�R�@"���a���J���B�����n����6&gI��H�S���[� V�^������VN���kr$ř��%����+[��Q|�Z��H]���|i���sB�$o��TRF�N*���]�8��M�Y��EPԢҁg�
���������A���U��a)��#�����e���}V�hZߢ�\���]X��lZζ���s^XH[�����k�)�r�4�����u�͕��P��V?k�T�7U̔zo�1������m�ҬbY��bM�η<��E6�g�i;�_����y�c�$��k,L�>���~~��q�[=Ny���V;����N�"�6l�wM��D�-�k?������o���ws2�.�Ӂ�Λ�>��P��W0"I�E���3�],��l�7�r��j�� ��|�惖��]�}$_>�.�5�����y�S_ɁY�H�XL}TJzJ*H�����n:���F��Ҷ��$�=�O�۽%���J=k9����~�穈P0	�c<w�&�=��� a<���mƅ�_p���4�!U�+1�=^Uڡ&����cC���i"�Ik�qmd�9Ї�z��������6��;.:�=)�w��i
� �$�c� 	˦o(��KI��d�I��إ�)���e`������U\]q�{������!��V�(�[Q�Z�f�[C�$8+�����^�3�lv�(A卑�
��q�GlnkkJh�����@|��	����C�=Wg+�܏� ��j=Ubc�`gֲ����h�uF'&�4Mz�џ�ݕ�����RS�r�<h<�˷T����M���W�{+ӌ$F��H���]M��&����tY�,�54��3E����Y���H0>444'g��`L+K��v�G����}��po����y�I���@L�����h[L��~R��mlV��@fsg���m*w�6��_�,!�oNW���aaP�<(�=���ȼ@�����s������;�r��k�%�w�ƽ�$}�g�H��%����Ȉ�l(�.l_�?�.�2/�� ,�s�	����M�:U�JD�����Pz66SQy%T�O��C?�i�y�.�`V�f��}���Y��{��{����{_e���լ��t�f���qU��<��H��vM�������W
��ErR������n�I%����I5�5__��W���Wg�����|���yoV*V�V:��߷!?M*a,g�㬖��*ƛ]���b�cI�j�Ѿ{�]T��&�����t(��;j�E��s�^���������G�.���c�G��X��AQ	lhJ�������u�RE�;�u!�&=��lD�M�[�QZ|j����)��xA�����Q�(��8���_C�t�;]b�=�ˀ�&�rH����C���|��'2mB�A����in��'��T:���ҭT��qi�9��������˪�y�eLϭ�H4���0��A�HEͲxZ������Ѵg��Z�4���7�a���O�#=G�M+��S�f��=z�I��@�����,�d��d�M9�;�8<b����7��}Cj=ߟ:D���I9��/�:&��O-�� ���ͪsj�Z�ܬ����J�#QC��Vli*y3��}c�6���F^@�T�α;�G�R�f��0y��m�E�����{�&�E���I�im-.1
'ۙ���_����iCpƦX�̩�`��}*�&�I��&�<ʋQ
R�#t'j1����ޞ�Y�J�%�å�w��]5�Q�@DOC^�=�F�Q~~=k���(M�w/˩��=l&.������P��s��Oa�]~8c����g@J1eY�����HY~x[ J�D\>HJ;�)EZojx o����!+��eM�M�>a�f��&!���a��䳢X��޹//r��A�Ї���N���%��t]�y.��O��~���d�0>�z�Un��F�;9�<�33�����W�No��_��T���-+�"��%�kcccSS��������;�<a�����ߥ��ýuj�͚��(b��+�~ʷ��?+2LZ��w:R{:��~_8�U�I�!�;�䂘>�~<H�������y�q}ߗ.�����j*�2��yb������o����
���s���S���ռܣ�Beѿ�jG�!هK��Nϝ�<���L4we��ת���m������`>`�'��K�}*B �/����}��@{��y��� C�Q�nB�F���f/iEjN��A�O�:N굗������,�+�4W[l����i&�]��*_~��������QhK�,��QpN��7 ��?t����rKo`���G����+�ٵ�׳s�a,���ۜ��6��!GI�L��9����lf�~)��&��j	�o�����^�2��Yz1<�K�헧*����"��F��H.".���⫀T��s՟���@�W�vB���Q�J�Dy�4�]B�t¨a�J @��:�io�);���8ֆ:}��ܘ��2P	w��s�Mp��LK���HK�N��;cW6)�k X3��*u!�`����Y�1P�7�U�gj9`L��F~�ůqG#�ޕC�"y�����a��d�!�{�o���gt���'�Y���R��V[����IRgV����3�nP��d��M8��|w7'���*�*��<ذ~:���c� A�d��n���?���`��_��/�9]-"��/ޙ�4����Kг`t�Q����	��G�KH�-���l7b�ˮ���H��2Z�𱚨��S���c診�;�R��^i�뮰��B�ɗ^(ؖKX� *�I#�[�S��?s�XR��}L�������QH�@�o1͐[����z������=�"�GQ*�dv��i�9m6��O)���v�z6�m��b�	e5|˂�1)�a:�;�JtGpBCWR��RW-t��r�i
�d}�J!M �a����{DU)� �t�h�֔�-��:�	գq2T
�����P��?΅�%�N��g�H[�VF������g�D� �xբ��3���v��g�6��'E�#�����=@خu:��ͭE�Ymnz���56.��S^��bh+l��q���QZ�}b�	R���!@���W����8P���FYV�%�ՖV�:�U�j#�J��n��q)%���l;���g<ѫ,����aȠf��;`�l2�a��}�ړ��q-���$'W���¶J��S��p;#��^a5����W�yw��L��7��㋕<�Z��D����Z�j����ǋ�����}>�_���v�뿼���ծ�����V`�+c��˫lY?�����_�Js

*�Ӎ��Ĝܴ��l{!zQc�lu�*�����B�ҭ�Ѧ�tw/�&Y�aM���)2��7�����y������F��D� �5;�.9���7[*-wg�ߚW��^�L,?�8�Fqlo^���,�X�:��������'G���Ɂ���dN TȪuJ+�%=�E�bo��j���e����tX�A�r��q�f��d&hzMzF�9�D2C�WnY/m���nSH���G܇����@v��%w3�c�8��k������:VϽegcR�H��/Tbr���[Y`%BM�\��r�V
ϦLigt)��_'Y����ݛ��N��������݁�:�nl�f<4��マ�Z��hI����PQ5�����{9���l(?i��U��3�dv��ټC:���~�?��}�Ep�\m���1�����w���`G+G�ב)JK{��z��b��W���w��.[�%n`v�뽡v�}�C����=�e��YR��o���]�h}�O�U3g���<Pk��8�ٓ~ZK�|,��`��ω�k��d�;���ͅa4�nL���ޢ��(S�~����9o������y'4Q�������HM2�+}�RǪ�^��B46��WMDڢ����;�|3�D��5�|���Z�N�x�v/�]��Ie��<� �c�.�D����9�h^[��z�V5Aw	_i��1�[�p�bJ(�颕�55=:ch��]������_��{g�H{����ɈI�8�M�º��%K����4��l�H�ec�Q���F����ɴ�5�^/qL1@wȉ�ScQI����|t���7d;&�>�#����ŵ�Z��f��W��_w���4#%�WX|{�a��QM\\
�C����h�z���������O� �K����|�d�?�`�D�7�����Z����S�tUŬ� XP@�U��U4u����Th���_O*��A�9N���ߏ)���/)�{��l����%Z��w/�L~��xU�7�P)`2��Ӱ���ky8\J�楗���N�Ȏ�J��Y�Nu����ǣ9T��?�'����	�&�l��`�in?�ĝ�0)��O��ܪ��ߣtTQ��մ{������;���ŎF�3��׀*��w�m;����w0�e2����d��d�-��m";ɗ,zP<�?�V�9�τ"��D<�Tl�$$G�p�X����`� �}���~��N�&`�ⷵ<08�o��^qI}ܼ)�x��4Q���������e�۲so�E=�Tr��Q4,6v��a���u�q�Z��BX��o"���K�.Hu莶%��o�XqiT_eZ��*�n�:Q�8Q�"q�0Y�I�/�'[�4��.�}�;(#5��|<9?do�_j`��[z�5�G��{.;��J^d���kmi������YU9P�~�뛹�/�^) �R$`-��f0����Y}t�(�G�"ĭ���D U7:1��iei��x<Tߧx�=bMi��x��u������?s�����#���Z��M�V�~����=,�(�a�õL�pn
���N�����;Ç���fG�n�z������*>Φ�������*�w��J����MߚPM���p�r��%�t��ߟ����봡�/�o��-j�혈 �D�Bh��w�D���rB��Y�C�S��k
Xɶ� L*�E�/�~�H�#fk���-��)�J����XQ���1���%��Ha��Ԑ��/��f�������|PQ���2���0�o� ����)�m�8���Y��F�¦^��ڵ���(�Ӎ%�w*�.eX84���B=X~/0�zu
�m�Z?a����HkĦ*�6����o�IL�l����A
CR)}���}�ʟ8U���
ǖ���c)�ڗ�N�R� �]j?�Aa2��a��5u��F�Z!ղE��ގ��@����;��t��__�!��l��>͏����Atuñ�j�S{5��E!�?9�g�X����x��܄��Orx�+����b�Ǭ���8��^�����g�(���r֊��W�M/���7���B���S��B�&yUUÓ��tn:�7�~��]�����)+��+��..���	-���/�F�0߈��;�j�ʓ�1�G����{e�}�f�4jj#f�.ayoe�iHe[Lv#����	u\�}d����6b3٠����<Y���ծ�;sAg�Y]��V��QcKp\>ݎ<��s��D$��������/��
���q}�$��Cr�@�T��ȂgEzZ�&d����+��S���L<��"*��\�b���@�Zby��V+_C\X-���N�)��Q�m_Z��i�� E�ɉN�����ܮ�O��-:�ݼs��:�b0����#��!M\���^�������7�!��|a@"�C<��F�c�}��-��aefE�$��a���Z�X$��~b�����-�cY,&�K�ހ��:j/�Ao��Q�a<�Ïh��7�;�ґ���)"�uKs?�@c.�tz�|͋�z�,�¬3k����z@�D�3�/�J��dU�S\�I�b[�����z���������`�6�eA�h3]z"����5�P[��C�pH4�\v�`��F8���۾޿�����n	�]�c�F�n�jN?4z���״�UAM��!E���t�$2l�?R¥�~��/��l��\���3������u���{��-i-C���ފ=S������Ê�0�[�$� �=���k,�P �tc��H?�EK�kT�$΢)HE�\�!%�,����)}(	�'�˔�(�c�2+&|�|�p��� ����߅�G<,�e�+Q�~�\�ʴ�d���~�B�[XB�< ���&���$�>��'�sj,K��xp+�W���]>O�����\8N�x�k���0G�q�q���X�T;��k&�zp�����| u��띤�kCh�J�~������6KI����^/h���������c�O�x"�0�K�E޸4>d������G��m��Y��j����&^M�_=א������1wn�fJ5��FI�K'ҰT�nr�,k�L,R�W�hR/����X!Fv�n�dR�\^����X4���P��	:x
=q�%�ڢ�&��p�&��U���z��BHA��tv��Ќ�;:��x�m�XD����L�4t<�Q���%GaV''����g�`��m��ur�f*�Rqv=G3�m�K����U�V$7g��k��:��R˸F+kF]�\]Ֆ�.�F^:I��֝yg��Y��-|��o5Kw������#r��-�;�������̈́v��n�\�����M�y����͢�mnЭqП��4~WC݌���IG�8�7Z�<Y�K�`xW�;�:���tm�ӨO2�%�����g}1��� @n�K=OH�)7�P�ܤ�P;~c�m��ɚ����μ�96�r[�n6��A�E?�<.��%TN��קdfj
�ʑ�:8���.� |`]��j�OJ,+�D����ja���FG���*�o��5�ܙ0�W��ǵ�>˗�Q��mu	_'�K�ʜ0��IӋ�LZ�����l��ݫ �eW|">T��#���`��i%ȋ��z��-��8��/��:y�Z��t���"�0#����~�},����MU�1�)�a���|0.��i�"�F����y����W6 �G�_�L�@_�(��ȕ���t��R+�Rg�8�f �0?�F�����/Z���� XL��FB&��z�4���П#^�|�S�M��[���4��]��$¥8�x�"�E��~�K{�j���뭝Dr��[7�y�&��n0;Ь� i��^�ˤ��A�P�XGb���@�L�*
���"�!m�ۙ��L���}��}��L��7��//�/	m8�C����'������\Ҥ�dJ'�XX5gRRa�&�a`%U�&�9�}3x3���񷂄����{l���9�-���]�%���4��gkK?��a�jʹN,��=ʸ6�D�C��(�Q~+�!��/�>��P:W�m���r?��*��>Bh��Bўk�`����Q&�~#$'SJ	���
�c���>��朱��i�fч�i)�2�K�bTb�D�,�{�M�ߵ����m��ӔxY���T��]�gcȺ�þ��Fr�r�(9��j�e�AT.��Mg����w&����
��!!�f�.C�z�Ix��F�w������Z(Y>x�s���cn���ti�?�� ���Ǧ�gfߢ>�\1�ߙ�td�h�%��RvZ�L��d��|V��?���4��J՝���L+>ͩw����t���$�(�����������\�퇩�]8,4<������/�S;ѫ,1:���ٹ2��y)��^&/3�K^jZr���7����mG���s ;ZO�oo��ۂnG������]��?4��o. �h	��j��</(�*�߃�F����ǳ�y�ϼ��J�:N�-n/\?ޞW�t�{���t]��SiP7�
�k�+0h\��������7Jv���O�C�D�8C���?'�c���%�r��wƢz�2~�_M�������Sӗ�=���l�&c�eK��&���-���n�Dڶ��֋��Ŧʮ�ߧ�#ޮf7ڹ��z�}��H![n�ݚ�g�j�
TU�~��QQ��9���'���;�)f{�309�8���j	��u��4�K����^9u����[���w����=:_���?1~��3r�$B�X奝�DB~�#HSD��u��I�H���i(&#�b&��^H���rA*�ԁBg�˚B2�8��lIZ���tg����̍i5@D��M>���SGu�E��Q��~/��f�geF�C��%�����]EG`�'��0,�^���x�h�R'���o2�����M|jB�I�o�N5���lL~@UJ��	Jz�h\�x�i�6{97�(�I�L�H�������=���|dt7��9qY��׽�#P�_�=�S�%>�������/��l����}�a&k��~���xv�{�=��cY����(V�u5SyDM��+�W;��?�B�g��3��;�TG�j�rd�W҆�$��	g�[�y����n��eP�4)+��'����Ц�'�R��q6t�6���/N�
Sۣ۩�,��L��q�@w��pf�m��@��Ϋ��hR�7e[�v��{�Q�s����p�Ȁ�v!���f��'�|��)s��kH�g���󩴈��x,��aPa`�> ���J��U��zE\`�SXyh���Te���y�y�J� H��,�D(S�m |�l����	�3�S�����&W$�����a)���M;��;XB��ާm|g6�{)}n���6�j�1_/���{N~��9a�^(b���[�T�T�vK�=�ɗ�M*�)�Vn�.\�U!��I�'�2�̓���F��	K�c�A�g�c���k�d�wn�����sXu�=��X�,�x�\�+a_��X�&p����.�E��x�.���$�Ma�p�W1.�u{�����-�LqX�D]1��;q���h}�1�W��E
�@�|5/p5�K�W��7�}�t��p!E�I�H�L�d�Eȩr��b����� �4���vY���`c����:?��L��E������	�p�'z���Kr)y�D�϶�7י�Y�����q�tyl,�����o�6�?n/l����r6��?X�G�v~8��Z��w��Ǿo���Sykڂ]'�-:N����dY܎�>��w=���`�!ջ^}��z��{<�y��N�@���:�/g��'˘=ov2�/�TPвsk7/���'�Q/��)T���2e�0��u6���$�Et"�����uu[t���sYM�uG��ۏ�r ,_��Md����_r����sx�O
�Q0J�B
��ٔ�
{{�B��MMs��0t�����<�U&�lҪ��y�4!5u������
�����v�N^����9R=%��R� �ҽ�c�*�Փ��,��,I�u�Ӈ]�s[X�h`�����m�N7�<'�q�t������.j$&���vʧ�vxXu޾�3ki@h<�ȥ\O�<�$�w!��y"���4�y��T���g�(��鑝�%Ă�ŵ��6Nj<kw��Τ�s����������oAӠ|V1(��s�5�����8L��E���
�d������{#k��g�oJ�f���#:csb4{P��5��w��o�fK��q�K�FG𫑯1B��z%z���5�L�����Q�N ���[D����}O�;	
��Ys��#~fp�����a[���:����k�͊?���.���V���	��"�9����6]t<�	r��j��Nޡ�u�����F�#���_�Dh��}4"�$8&��th��lX���#����͡�I�#p~|����d�w��ۼ���ٰ�s�6Dེ�\x}���g��@�«���I_%�*�=FĵXXDg�fI����WK��ƫ�?�}�>ۙ�u?f+-�!�g���E�µ��[�l�} �L�L�
�~�ه��i���1�#����6�Ð@�P�"��T�r���Q�شL>�,}d�"|�/_M�|����mD՛C�K+k��12N68�|,K����%z^��U� 7��;DJ��eq���$~:S:�3�h�g��R����z�A�]j>!$%���,��j�XQ@�=ubڶR~��yī��2	0&Pi��k=��ۚ��0=��h�C���ܗ<ZU�l �:݅]�O<�C��Rs0�*�o�9�?��P��#�U�M�=;�!��WS���ctH^��B�c���EB�D� Ԍ�S*�!��Z�4O�sW$�&�n�2�}o	#��+���	�B�TmU	<U{�,V�q��+�����(UN���*���Y��!�e�ɧS��xq��2���y}k��>+�ww1���CO�2��F�b�7�pcF=�|�*`f��ZNiwT�����S킍�~5�*V��+�����VRv/�i�1�ҳ���K�G8��Ԋ5���'fv��:4,ϓl����ӳ���@�{,_i �&����͕fuދ�2L�~�u��=����]:�y�}����E��E�e�Eǿ��Տ$���߹"?�,w=m�u����H��jgn��YɄ��U���ݙ���ax��Y����M���҄�����m_�:�h�*u
**jS��/ə�iٌ5��C�9<�4U1	,����FF��+����L��H����i;�C��.1>��Sl5c! N�@^��r0��>�l�^�S������y��]^ۿ�<Y��$oW�^��#u�SX>2]��b���[�2�Ү�d���G] w;�5��^ �
?�� ��Ery�Op�*
��Ь%!c8��٨"��Xu&��.5	�T����Y+>q��E���)(�x�z�r6t�JZ�>����:��1u�QM��d�5BB��Fw*0���1Z@�J����nDB�����" "����{�s�w�vv���y>�瞻g9hZ-眛]zސ�E���5�v䎓Bz�$yC__��_���1fxKw���mhX��]��KŰ�6?��xA
%��u���s�$q%��!���U>��#�#�i]U�8Wf|П��P�23(��ֆ>�lj2��O0�bш�M�$�z��Z)R����X���URF]�(�hM5����N�LC�ydkL�`<�^&@�����>�I@<��R-��Ţ�����ÀԩY�PD&ˉB��������i[y����"�T���x��w�5˛��\අO�I.�՞jm淁�^��w>Y��.T�p�����2��Ph=\s�A���0<p|��/\���OD��	����P\��X�����M-���!xh�4!G4��y���.�C�T/pof�rĮ�(���T?h�H��9s���cr���,^��z�J��i�4�?�:�V�콇Gݐ?]gR�lkvz����.I2���b����t�ZDX?j?��϶���������d~�ؿ�q}(,1�9ᢿ�DZ����æN��F��@�z��A��ߞ{:�:��\HT�
!��E%`����g=��k17��{��E:$Y�8�z�E."�)h�8���J���*���"�Ѓ�2�%1[�����vnPi8�'L�������h�����4�c`�\y�l�_4�"ޠ�;���2~)��$R���©�o>��u�#��0��� ��[o2���:�g]�SO�������"���9�a�v"����j]?'4ڏ$3�F����EG|�����]J��9Y+"�~���������n'���u��~|y���C�!���X���{��Z���Pd�a;�)�~aQ�>���hU�����GB������=�S�@*�p�����q:��}+�5���lY׻"and�����E�F�l���]"k��Ģ}e����ټb�K��HB��pq��7�rqY)H�u�F5&&���II�_����@Ϟ��5�����<�ɓ������Q��0��qY�'[��x�Tp���̟�U��G<�cP輚F,!��͍��i#����q�H@�S/K�~^�� �[kjW�t7Q���v����4�:�x�L�_��!��=�L*�I���,��oSsbz���r]�����]dJ{9@a~��  ŉXZ�O>͎綴��)����v����|�A6y�(�St"�/q,qk�e��.��+��-�7�~G]!n,�T�^x�],�E�:�Ae\��l<�
��
E\��ᶃQ%�������ׯ8��5��.ڊ]O��tj�~�'NK�#a���u�����Vc����=W�
1.!�G�6����~"��Cd��=E�0�X:t>.ă-���vL�u[F��φi{��a,�Y��	��U� �OJ=]X�����@Lb�+В�f�㛪X�������2���Г"�x��l�Y���[.�(�J<���x���q��skB`���l��`7�H�H|=��"!�J���&�_X!py�4>������u�z��{I|k*���7�g�
<�y�r.&�"���}�݁��F�*�`zϵ���)��҆GTRU� 'R,`4�Q?;���s��ǯcG�f���×��#�6F8JKy�ŅK��Ǭn��"����$Ǝ�>��F�ne��9T����$A�`��P��Fiv���*�	�l��i@R�Ӷ�9A5A�=��oa*�%�m�"�x5N��Tp���%������7)�ܷ�t�@�j��w%R*͒��G2�a[w�.���!�jK^3�t�ڏa�U���_T��,ؽ�E�?H�}|�W��>�����T��s���_�o��|��&mn\P��T'))	�=5�r�law�|9�4���ZZZ��Q�*j�'�z���W6|����lј��j����>���B���#�,��/���/ք>�~,��9�I�����}3�eu3 ��l��$��n;�ß1��?��l�6V\`���~o�:~E�>�_��up��p�)	���g_��Ȥ.,Z�Ÿؕ�Q���H6�2и�b�g�q�y�@�pz��|%���!L�����Sg�7rM�PG����n^��r��V~�v���m����� ~cM,��q���6Vxyz�Y�|2�����>�=����v�^��6 ,����>��oRacGdde�7�����!�l�oQ�d���ޏ���o+T�*�=�Q�ڒ~����������_�}rw��v21�i�L���C$�n?L�`�P��y�d���L�B�ꌬMB"i��.5�n��7�B�ݔ+C�5����x�׼t�P��k�%�*�4.d�d��	�}��!nn�Ok��b�K���`�Ec��`��"&!� 6�Al�]l��o����$zL�XDħ8k2�6����*/������4d�+�E���TW���#�j�)6�F����]5l�D _���c�\�m�x�ڐ�����7î�Q���ב*1-)H��N��t�)߷P�bo�X%&L����+��Fڴ��\%c����Ri��l��%!�8Y�t���WS����t[/�z��Kpk5�M�t�j��4�O�.����[���B�}?�����1Hw�1weĐ�b�D��m�C��Re�2M�Qs6� �^#��nZO��.on|<D�qNs�oL��=<�(�~w*�X�d����Uق�����v�#Ό#A�C��d~�����qE[�]9��Rg��;�C2<H�����6���Ro�enF���\߱����՗X'I�e��=Pi@��R+-�W<z�ަ����~J<d"�q}!�F%I� �i��/d����� �ˤ@"�a��X�9��"��� l�q�"�����ꊇo(�?P��P�ǟ��CAo��p�R|�J�-e��?������$��!�r��T����M�@c��6T��sf���2'�ڶn�e�G3���	�7����B��MoN(L���0O� �_����9��l/�]]]������[�>�5��e �t���[/ͬ��mw�_9v�{ȇ��<�9蜑��V~�[�*��{f�nJ����/
�R
�w2_�>f��6��U���	cVpI�s�n����j@5	��q��2��RbK��� �0-7��Τ���8�E8�\���W�w�v�LLd;�ﶚ�
�KZ6�d��tZ�8R)���_��}���.N�ڐ�ǲA_V���s�
eB��,'�/[v���X�m���
��e�u7���~��˪x�*�/�����|�>L�zK�~X��&�aM+�g[rݶ�ǃ֭��{ �w��=N(E�C2��__K�Ub��Ds�a�}e�����i�]�����/���^$V�P��N����+6'��@�����H�#Y�qG��j�ďy�_��&4�>�9S}�gޑˍ��/%nX �:��8�W)�3�T,W�U�~�������f���u��9�[�6d]d���6Q��Ϡ����*��;.�ŀw�f���8N�����lj�(^�f��G��v�p(VxgF}����9{1�K�_�$��/����F�}DM=��Yo%W8��^G�TP �9,�4�&Hf���Z!�y0�G�,,�:0��G�~�O�!����䜉3!���9N��/hZM�ƪ��8��3�4x���y=���ܟ�P��V{@���\���"�)�s�w_��!��Bf/r݂���!�o>6=�Fp�S�'+�\<4mb�����	�J5��ȝ9�M�Y��"�]穨 ����V��@N"���Z��Ĕ��J���E4(��w/���e����˓׸�Z(�!'Hzݬ̹��tY�߳U&㨏�g T5�*'�}XG�Ep*N1Gf�	���2��U����\�K�s(q	#�����ȕUU��a�(��'Ֆ��5g����>�R���bY�Y0�<|�	!��B<e�Wj~��h*�q+:!Q�6Ҍ!��0�]}����ix[������!D5%�#)T'��?�&��cA.�n�O���_��w���M��=�w�C��l������d�ٳ��dNz�_Z��-"od����ء���Y�)���6�Z[C.5^JL����ZF�7ȆzF�)rW+�G��ccc##qF����.�:�xt�OW&,�q��V���,���ࡺd(ݴ����Mm��{a-u���I��g��/�d���^|mLx��E�e��u���vO�w}����z�ۨ�t|�g]|��b`�}�[�CE�㑯��a�
�Q���6�0��އN-��#�߿�]z� �Ρ1O��K�~��X��>����\A�k�}������t�ؓ;޽Q�����) �]}����}�8qѴ �@y�O��M����HKW�Q��L_����7�(l&�n E(���2��J����TE�a~�V�z^aoŋlMU��)<�C^��OA	O��^�Ҟ���U���99�wL����/J�O��Z�����E���������[��<E�����V(g��Zz�a9��SO٫�y�ޖeϧW��=�yu������9fv<��j��K�l��/(
ޤ����^,�V�;0�����m'(TK�������DS�m(6A��'X7���%��8ڵ~>�����z�'RG�r�B o�p{y=]��I�F�j�{�YLK��/�����\P���j�'gV����n��@�;3��Y�ւ���M�w0os+>b��'�J�nO������{�Z�2D����k�x����H��_�%a�B�72D�cѡZ�T���˻�ͼ�u�~��O�LY�΍"��p�*����Ab��t�>���uR: ��A��ܝ��G�P��Q�Ŭ��<qF�|_���}(��L�?͞� ��*�'�b�94+�˦0()��Ý����gu���bc�,_Á.����0��Q�$��� ��G���X&��E|C]l�p0����c�Iі�~���V�z8��o^=D?OqU ����NZU
l�E;��5"���4Y�ҋ��B/� .�&�$<P�9��]
���n�`�Ӣ���Oe��T3��#,��^r(��7R{;*΋;$uI���]�v�j��8�D!'�O�2ԢW7j �3ЫL*�(PNn*���;i޴��IN��/����0Xԫ�O�q]��ؿN�q����la~~>�����	���� A�rUFwqY�/��wjkjӻ��+*�kû��\�?�h1���B�����듧��sͭ�Y[v44�/�_�����6��1B��������I�������
���d��S���<]�qܩ��H�_,���ʀNP7��m�ᶼB5�,����y2��"�a��%���ů��pR���}(��;�M�PO�=ul�,�\�l�&�;{� G�\�����r�����,�h�����K �%ύw��M?�/jͬwݝi�u/Y�ZV�2�t�}̼��⽤�\l�Զ�Rx��a�����#�b*.(t����'I�~;W�}�h�yGM���aZ[�����n�|L�ׁ.*���j���t$�=6����U���nQ�;��E�ti�4 �b_Vn2��9FJ��4Fr��'��!�Ƹ��}5b5�j�Ҷ]����*u�|�\��h�t��a�O�ﶘ�����)�&�伏���x,�
�N��2P�c¬2�ɩd�Xz,�j:9/�F��9ni13���Bs�~:�a�t�m�a��-Ƣ�֩*�n�fM�^�=W_�g-n�����xF�^w��Y���oWBwR�fȷ�*�?��ɟ��wG�D�3��fq{�8��8��Pr��,ٸ��<���p�t���Ӥn�d^�1�����]�����$�Ԑ���}�e2Z�搭�5�'�6$p�!����������i�B�{�b��U*',p�=@
�����W�����O��������)��A�H�+��<ٸ)r�8���[��C"P�ڕ>�SK�?[�|�M�!��;V9��š>c�������
0$O֞V�m��a�K.#�J���f+"��3}�^!���Z��	/�G�J�Z����������k��	zJC�?����+�T��8t%NX2��-gJo��~��~c��H��!;��~$�D����:�����H�á0��X��t����\}N'����$�-�\��~�xR��Hr;��WY�����N*m� G�)�"\$�ؼ1�4~{�Ć.㳝��xN���6���0Vl�8-����zl��/��L�����Ӆ�O<�R=����l�8�V��lN��L�N����B�$
�FK5֝v> +q`?d(�o�\��u�kC���U���Վ2����V��ZI�8�P�Q����1p$Q3NFE���H����~F�B�O  �E��I��n7Y߯�i�������WVL������)Ph�J!+�ܐi����3�>��7d�2HpJ�����Т�5i�>h�¢L��xώFb�P�����κ,*����o���f�𨦝̉��Ej��{�t�*���qQ����?ӆr��i-����^�$�ǁ9�'pKC1��tz���&�ƕ�"��.�ޟ����j�i76o|u����c��v�P�g_�γ`�`Ƣ���xl������i�G��wȖ�䓧:Pq tJk�u!Y��U�1z�*��#���yP�#aO��b�^ΰy��R|�6bDB�g�D���f�0ƒ/��1Y��2 ?� Hn�Cp�_�_B����� �l91�2�-g��c��N�H�T�����75ٳ�+y�5���t�,m��56w?���A#k�XK$�rh��)�X%��]�Fq.0O8KgI�	�{Z�g;�mn��̣��c��lѹ��}3�t��tRB�#=�g$
���%g
@��z*��3(�
^0�q/=љ������p��ܿ�zy�h{Y23Z��}w�*����ؚ����x=�g�e���u���n,����5��,ڒzS��f�y?O��ѝ/�����Iv!����;�@�S�S �2��MfTH3�H�8g�V6�!
���u0��'E��8f4~+�J���Lu����g�=������3so�d|����.,Bӵ�oz�[�`B������'�F����O�4p^>t�I����t%!qd[���������z�'��ݳ��v&Y�N��|r�v�������ԧ�P>�Fp�㷕��`,���Č�29��u��:\�Q��v1�q�@Ű{��E��߶	)���ֆF���o ^��)uz]\]'i�(v���J�@�)�����0����܁���qY��S�<E��iXR���}�h�U5a{57�<����p5|���$�z��ov}���7Y��d�����G����L�������9䢣�k��:y�X�K��?8;�U)	�S��F00S*HA�|9�L����#���;&��@��@���n�ke�Ȋ�����x�8&��\Z�cw���(������t�.�/ϭ_l�M�Ğ��t]+�֊���+���
VJ�		�䝬�k�\>t�Z�(�o����Z�V��_"��!Kƅ&�A������[�W[Y��z�+y�rB�]��T���$�$�:B#���gn.[څ�\װ�Xx�S�H�ʋ:&�����M�|K�CEI�ygg��g;;��{��\ݲsQ��^ni><�U���gi�/��a�Ihj1�BrQS�9�Hg04W��V�e��냙�-=a#K��=֛���j�ÿmt�����h���C�Ѷ��A��/��vʚ�O�4�S���$98}4707��U�ϝS��pd�������Գ��8���gɣ�������:NfF�$/��#�����ծ�./iM���#g/������A�*�T�a���N�O�Yn��P--M����)O�uGg��|�^y�"n7��S����kfƟ�V[�>0�wʴ��Yj�2�=��+���`��3r�V���23���\�O+��}!�s�9[�~8�Q�藶��_j �U']�i��<}�z.ZB�Ot��ƕ��S�<3��Ŭ�,]A�|�O�r6Qs���6p�n_�.�-�F�F�Y����4GPw
���͜�[�#[��J�}>lV��1���A8L�|O&�~ϧ��QI^4r�U���$���C�H���xL3q4�L+�vIgL��d���Ec�X��7��~5����F�wi��l6�8�2�A0��
ƌ$B�\|R4��&���Q���)V�f�Ф�D�H��S"����CѮ<��,��z��ƶ�[?���"����,V�;�uS��60�ʂ;\�����4r\*������of]!�'_���,�\-�{Z��ٝ��m�Jx��)��;��'@}��OìJi'�
�;(�E�r����D��Fw�~�o��B'�;0�pm�O�h
S�y̺B��I�DC%z�j�bD%3�.�����8��"�#$���h��ņ�g�'���5��������T�g5p.Y�S"�%�m|�� ��~ۢ���o�?��ǑMƣ?z��Z�Fczτ�-X�@!�kKz��2����:�r����@��Ș�G����T^������������>�AsОy/ E�Kd��:��u��4/ ֹ�ښj��q��T�:�M��� �D��; 	��{���;f���~n�����w�k
���]���s� &�}C�_Q@@��xi���8rv��r2��V>�*c9�z��]���o7����DCh>�����멸�ت�G�T���8��,;�6�E��H�s�u���XX�=��P���/�$~��p��{n"�������Ѹ`��qޗJ�֞����'�6�|�o���L�CNݡ�����a�R/5��?�����>΂4~����>��3��\VWS�����Q�P�P+z���4�=35�D�KCC�"�6�vu���\�]W��9�˯�}S����Ǣ�c�]\w�;���ޜR�� �7�Tc1��7�������02�0�XX��	㐳����Ƌ,�����RGށ��\���u�)̠�*�Аs���q���ޏEH���4��l��>�Ҵ޴��֟���X��5t�I�Ac�톙���������Ϋׯ���~��������r,�L�� ����c��A���i'	�����(���E��lm�H%m苖�|�=G�-�&�0(�^�����C^�NQw��m�UL`2��P7J�w��)����w\��_)�(�r����]k��ƿ!$$��w��w�Ct�c����aE7�9[��ڦ�����E�s.�� 3���bT�c X�6������5����p^/ϗ�}r�v�1ǖ�_�1�HT�C�H��\O+1ӆ���>��F>�f_g�{8{?@`�����i��6�XJ�i���%�5���\��;�R�1`	=�'��{h���-�����l~_�����beY��Y�b�tg���
�a�`F��H������� ����+�4l�YN�nQ&���3���m�D��Ԉ�j�
��Ơ���Q�L��J��F�?���u|)�O���놋�ѵ�N�e������q�D�4Ki�*Ԥ���4N��{�z�'�W�d��8.�gb.{��e����aI=u����~䃏|�93�����1��ʸ�<� ��S��q_�{sӛ��`p�p���.�����Q�Dw���B��PT]xr0/G���c��H�e���Z��3�*&T��p�9;�qL������ΊG�6�;���m�xh����j���� Ժ�H~�P%�q&K�?�?�%	i(�u�T��s�,�P�4�m+�.�,�@8�=��d��^lsЩ�����< s����S�������3I��)���7��g؈:��9��qE	[�G���,b�$���s��/��W�V:­l?�cu��T���olw_���d���wz���2�5$yy��7o��
]������ⓒ�(L�	:�W��'p�Td�(i?+����������_�grb�����Lu���=�]�&b�I�y�OI��9�d�_�5�q�ٴ��	�k�E�`(������2���0��'��yGg��2W��a����:��dN;I�P}�L&�KKtA��~!�5ie���>k�颁AIuL�J%���������^fC�q�v4н��o)���P#3�et1�љ�ƙA�#�ӝ��2eq3YL��2=��E���%<l�
�k}��Bf�N7�ꊭ�����D�o-z�0�����e�31��OR�p�E^��)��z�'O�ō�)A�Ӧ�$%��q�U0�v�� �+�R�; ۱)��Z�;#7P&�P����
N��=������o�Ry<���x
�z����"�� ��)K�j�>�4M^:R���B�}uF�eE!U5�;o�0�V�뭘b$P���s�m�e��h�HG�� ��D6��GN���N�ǂ���F;�q���|S���tf]����6�?����s�K��3!S�KI/�N�Hܒ\[���_��$Q�@�^�Y�bd�7��.�;��|�ο�3~����5#0����(��$E7;-!+�3R���p�͋��E�\�X���ޥP��*q�.�`xH�˴�	9p���&]:��وhwp�1u�JO\K�Xz�vVU�LS�-��D�9�B��!ԴL�ti;f��L&c8��FD���>YS{d�����N�	@�-�$���u6M�hQZ�5.@
�J��BmWpjE��aJ=�D�Y�[���T�R��W�=`u>�� Lu�i���"�b�b��b�m&�á|�-���?��s�M��o4�2�8p�������y�K����\d_�8��l[��
 r����>[��'�sv�k��;%�F����R����x��2t�N�j�3a^Ѣ�|"I�D����9UAb��[��Y��(�m��Ǜ�$j��'G[�q��*eŵ��`���Wȹ!*`e?��Bx��RsV��Æ��l�ɵh�y3��ޭq���U�o��]�.F��j2@a��}��1�P�c��Z�)����4Ҁ7���0�ȍ2�%e�F(��^Q}~6;bF}[E�
;��@z�'Jج���iB��A�8%)�_\J��^�t��!"8��g���s�F�ǀ�_��"k��:��D�?�@w���?*A3ĸæ����t)r��"�ԓ�O"$�}�B} Xy��Ձ*���1��!���6tE,?��DvOn���s/�Ѵf�*�`����ם�E�S��@Gi���F��}�8�C�¢��Hs�{�s}W� h�1���բ��'_9+'ec� $��� ��-��I��
)Q��Sw�Zн̵�j�s�-9�-5�/�����Yͧ2o�=�o��Y�Sg��I㺆2}��e"��'��g�Y��G�pv�|�9�F^�O�Y1E�?��2)خg7
��m��*1�um^�CY�|��-�j�� �e�fPW`����}��t��"��tM�k���4����׿lf%�bҏ�����*O�:�x�¢�
�>���|�a	�:�n��G�c' x�|�>��[i�,P���o���;9��|�� C�>}	)m�M�d���w/{^Yt��`����-��g���7�G��a�C��������r� )�b�� oٟ_�0r��&�ֺyh����WQ���ذ��Ɋ V�J?��� ���|���A$����[��B����?VU��ؚ3�A L̝Do�*[�HduY�i�y_p�pʾ���y13�/qP8ݒ �cE�����+5D+��L璉꣋����^BQ���.9��f6AK(���"��g��>
�M����{ǸK�c�Z�u�;X1I�A�=J�.7���Rd�ρ�H
�x��k����*��x��y�x���l$b_���dlP��"D#�ګb���(�I�W�c#�RZ���v�B���qI_��H�/�}2g��8X�8r�P`��̷��_N �uzn�vo���G[W��ɭ��Y�=N�L�v��-3�Z:S�X��y��_��H䳐�u�
��9愽�Rrrr���Dj(����F��[�逮��S���\�����Έ|;�����W�٭7�
/_z*Z�m({w��n`n��8`jb�����|}D��4��\B��(E1+�����,�+�8Sz�)�|��3���[8���_u��NΠ�֕;$�;�'��H��!�9�?�f*��#3#�ZC��7�9�BVL���ć��W}A���m�w|�}�db�n��L�����^p`c԰��#���gq�x	Z5M�Ľ���4��=h/ek^�R�v�p6X�{��puS���g1/@$#����G�����[��G��������T�)��)�dw~���q]� ~ݿ��+� 0�:z�#{���s�'��*���ؾ{8�'�-ьX�u%'kD'�u�Κ�?��w2�4�����+�8�@a_t{�A�[�ao���~���L���޲x}����+�[d�pnǢ��֐�K�/&�[Ǒ���}F�.p����?�v�6���*d`pĞ��[��j>Z��qm�^�CF~
I6�����־�!T�j��_�N'z��>q��|Ra��X��+�qkx�~]DU��rG-L�&1�s��>W�y�G1���nLk$��NÌb6�`
�cd�!T�n� ����R�+��4�˽N�I,�$����/|�&��%p�Eɴ(K�u���HF�V���\PÁ���9�KV���a�����C�ɭ-�U�l�N�S��T����rRiv� ��I�@�쐉-�d��C�t6(@� ��T�Sݽ$z8F<*u6i�~WIZ�j�S�J��C�n��lյr�d`�<��fF�q/Sϖ�V��U�6Y]�������j��{�4��`��ó��xT���['�4���Z�Ϻ�� S�(B�Z�~�C"W6�%����*��k��o�}�ρ�a,p�*����Ø���޻�
�6��O���� k����%�Wl�;��Xo![��k���Fe؂���n`��|�GO*E���_��W�B�k�q�O��|�-M�EG��4 &��qZH����yKc8�VxG���@p�%G�ܩ��T%Ӵ����#��0����F�&���OY"Jj���t-d�7xlƓL�	 N�!���Eo��'W�vv\�%*�*�.p��^Yh35�/Co_�`/��Q�'zD�h�v.P��c���E�����b��r{�v B� U�U?
�/ߪ���ￗ��G��돊�P�S��`F���G+�rAn�9`���h��PVO���w�C,vd��ۃ1�H`K{9�>�{��"��0�дI���~Z�(	�;t�J��&	��s��ʍ�΃ ��u~�I�����,�8��;n�Ь��'	�'���e���ُ2���q>=M�ҹ*l��K�4�C�@�ɹ�]�!8߈zgF޶Ϩ
ct� �~���n�����|���`�����rc_��ݑ��x�ٕY��a0�5jFSh+���;ji�����6w�2䰅5�,؂(能ч�G�X���Y��d��΁�Z�E�t��]T��3\��C�5	9,�n�HC�
å{B��O.,��.սڳ��Ys��:h���o�em5C����"��}�1����S׍�7��R��0�5%��Jڀf"B�H9v���-X���qh�|�|R��T��j&�Y͌��tǩL&�>��ժ�3
�h��b���%G<�y�5%Z�WѲw����j��JKK/��׿��[|�2��=���_��N!|�h	��|d~g�y�O���ᯨU��3wh-*�qЇ���A��k(9�/&����u�`mAڀ�i���u}�ׇ�}���o��M�U�8CI��O�lI$�U�v�1��2���h\���Yk�-\J�e"�B��%T�����ܦ]$����_CoYM��dP �U6P;���A_ҹ!�Z69l���.��L5*+FТl��e�(��>�B�T��b����kґ�"f*.ł����qY
R\�ݔ7�ݛ�l��C�I@,�dq������[�{.�̳&�[��u[�X,a니��:���D�vO�v6:�6�bj��MĻC�cΥZ�2�o������%�=Pm��3��zh"w��Ga����^�b�T�Fq�%���.��v*[�6�� ���� ������wO�a��b0�'�σ�ʚ��M��'_��YĔqI@0Ѽ�����ϝ�sJߤ�~T@�U��D�b�{�\���7�\鐈��OjjX��I2Tp-g\R=�����TĨn�� �H��E����
����w?�8Q��j����6^�~q*�:0)U�	g'�5x�������,���ISY�L�
Q�J�1�C\$�a��0�頚�K1��=���F5YT��T��.̣Q>GT�H�
M�2V��-�2�{�>��5
�,$�PYq����Ȇ,B�{?�e8��_z=��~D��%77R�2��ښLa���۷���[�D�U�Θ�A\kFb|X��i��1+�9��׵�����N�����T��s|��5�g*V����%���e�q��n>y�vu�v-�hwJ6\r7�;~���9�\�ע���T��T �'ŭ��\,���w��.h6r��u<�~������ٺ
߿��w�CfΏ�!��^�:��ٜ�co��۩�'�X��~����v��[;$Ck�������*4�<5l`L��3�$��X��K'�[�����I�K=%�/�-�����^,��N���Yn{�K(Q��}�L`+���c�s�Ů�%{��$��:��H���ӿ���(��ۊ�6Ik�솃�R��K� ���_Z��]�PmMc$���aSH����މ!]���ʳ�p��h9�q�f�˅i���rD(��%ץX�+��H`�#(`�3|�����BB
s�j���6J����FK��-3��y�8@D������!,۽)�,��w��"��#I�Ѐ@����<�*��꛵�?Oe�6&��Ѹ.%�D�8�����e#��Y��a�B��y�t7Ԇ�y��v�1��5؝$�NE�y�\�כ���K1'x�pc�C:�����g�/`ҙ�̓C=�+��`>~�Cs���� X��)�JwM�'�$���ժEW��X���kT�L-��I�0/���d�>���Og[�U�1�<��t���8mQQ1�¨�]�BAC���,�q�sʳ%����>+G�G�����jW5ϻ�v\�O�ɚ��ИF=��z�co K+�	��D~9�D=�Q�������2�h\-/!%���Q ������6�g�H icߞ�*�����PӑM���"l�ꙸ(>)ҍ�y��-�*���'� AxkO����'G�/����k˨(Q1'16���t�����6(;�>���0�mv�Ũ0�sP��5Xovr�q��cI�#W���ߜCfMFbZ�Z�6�yL�w���̢H#���
N�;řk���O�����Ɯ�nmſѳ��z����8�@�7g�oTBrE���C'.  �TD�ENtI��Nb����7�8�O��fOU7w���v�ؤGAB����}�˴����Sk��'�y'���۩[g��D 9�Hw�~*K<(��0��E��t�lzգ��tw����|m����#P<z{Awk��h�̲�	t�gy��K�\9�4?E�6�܋���ɬ
2B�w�����/�Om���]z�����}��+���p@����Q��\�)!, 3!�|�`�T���9-��뺘�B�O�h�ݥr�d��$m�����xZɬ�#8�|(J���*�RҪ���������j�*BJ�n"�3<�H���W�A��W~�J/�HT�c���7�/`TW��m.�x���{���d��{ l���n	���[������M��ڵ{X?��q�N���Ҝ���|��2��n�C�������e��xmQ���{�]s�3^�/H;�q'�+�±#G�ȤF��U&�Sz;ESed�Zm�/tW�9�}+[�[쯴8'� ��{b7�K8긝UJ���n�^�v��i�;�;/e��]G�y��R����L˳0?�$��cK�y�a;)�����;^�y�n=�t�{�<���f��'�O} �0��s�������]�N�}�1rۻ��9IָX\��>��e�A��s�q:�p��T�fJP��t �ό+3�/�\l��)=�=���H���D�$ʨ⺸�F�r�9ʷ�E��P/zV�U&>a�f� ��`+�|Z��P�:1��'�=K^��7���T�lE�1��r�T�Y��-�Q�<)"HJM�_h\f��0PZ��]ޘwf�U���*�z�A�p�H\�������G��>�_22���Z5���J�?<�w<[���O�Q{�V��!1j��E����A�5�Tl5jŨQ!jS��;fj��Z�j�o�z~?�C��q]��z��9��`.����QmP����x��mi5O*8y$KG���z��|����2nn�>ށ�Z{{��`�������B{T�mjFgB8M���H���<tB�u�I�Y$ۙe̹�Y[x:95LY�D:��[!������<��������3��\����|}#��O�f��_C��r��A���-Bum�I���3�=��ʌ9�(/"X���7"?�捱�����$ir"�B���k��%��/�"I� �֗"�^j�Ƌ*,,��ey��-�RL��:�|3T��F�0��ݻw���3__����ى���ɉ��բ;�fp�В�ɚ���]-G�)���I�MI�y������a �$�����!�M�.R0��h��1�����|��!�=�<o��䓁'O�%;�6��7��WRV>�n'1��3�t\e��ɶ���|_|���#���M�hm.v�{��}���x8�@�C��-�R�����Ė�����U@@�Օ��+y�W�!-/&V�w�D���3��+��4��f�K��V��[�v��<O�Sv'�k�0��,�(D8
�r���/ҕ�0�)�Ӛ�\yZ0Y���V��^@*m����6 0SW���� 
 ���K�&/�`�	�i�ζ�{�l;{X���3�o�F�Iڱ�d��\�j�O2i>�3u��hJݝ����]�)t5}vq�z)�o�l�y���D�U�0�2s��J-V�UF晴�_��{)���l�&�gGrJ{�����ӷ��&�����.�M�6�g
�Q~��G����r؇�Z-�@(���*��ŗE�K�/-'OƘ(6BkMZD�G1�'PB�Y>ܘ����3/DF4BF�PE���/��C��p%� �~Lʏt3�}��_�9�.,T��K�/b_�6u���V�*��>�6b+�
;i2�$7�c�$0a3h���ᮗ9kEXRcw���k�� I�]e �Q=-5�z[��6�Oiyy�T�����*_�x|�n��e7�`�ԇU��VҀģ��؜[�8pu�i�5J{����t��v�9��+�S����3!�G��=����@�S��IJ�����zh�|�eNh2oeC%�,��� brE�l:Y՝����V@.X�>��v5n���%Io���������/?#o���l���$�-��8�_��HF�s#*_@�a�*��+%*���_�y�i�dLA����P��/�������)1��>u����x:�.�ݹt�S k	W�z�� ub��H!z$�&������[xy|��JJ<�'972R}���$����~����,�*��(�F��JF�F�r�7(64���8M���W���av>� ^�3�>R��i�hOgkQ��W���.��V&h��̍���<�e��Ò��0���f�T~�s�� �����Q��>���[1a�%V=65��|�0eds%:RSCM奦:F]c���55A�j�/�(� ��9��_�!�����i��V\ɏ0w���S!=V��wtqxsr����C���A2��r���s-���Ǵ+ǮtK����!��W9������ |=�S�i���
�&�w�e������=7������ʽ�u&z������7�F��7�3H�a=��t�5���g��q�t+U�΍�ցq�C��Vp�]C/��;Hdl)��N��a_�����1X���(�h\����Xo8u�
Zݤ�HF�΅�H.6��W��K+�Va�O�S'e50�hp!ÂDU����&���4D�?���ё���6���X�<��{��xP�C+Ѝ.;4�{ņ/ؔU�"6���A���"������-]6=Y�6a���1�F��il��#�����3�x�C+�Iٽ�Q5����Y*�'�4�vR��8��q5k���T��`��6���i3d҄
����>xa0��*͜��� ��Zޫ1���p �v�w�;"��{�3'w�V��:wd2�bob��@I�ݹ��
Y�*�j>ύ����[u���r���[%�y\��!"k��s$��oi�Q������^uh�Ո%�OC�d�����ۅ�����[�*'i-?��h��`�u���zw�,X�ؗ�A�t�Ԍ������
�0�9u���g�H�a�i�o3���>�	�Ci��S$g��-�c8��r+u2lH�q�Y&�{P�4���xe\)�KX���z�2ktwZ������]^4��p�'�e����h�����}��M�N�/��P��ff����8-�zDt�� wTk/������)���3����d���W2�% �i�$Ėq�wP��ȗ3��F����/�ǡPZf ���P��#�fּ�+SS3m�*T���.�{4�o��kyT� eŎv��(��Y��5	�T�����B�y�I�	�t��[�Y�Z�J���a3`�����͕"|�"^�#�A�5#��&]1[�o�
b//��>=�|v0:}����\`#��\��嘟�a�@��i�f&b&�fC9����cೇ�kw2<+�>�Mg�+�t�v�S{s��r�g�^�u�~::b(�1�^�/�g�LC�]��Ї��̜g`�d\��bJyw��pgd���Y���� ��z,>H@½�%���b�3��K���-5��.��t�J�?#'{�����ê'L�|�����z���/�H9xט�D�����Y��`i�I}P��}��!�~���'if1����wyW��aҦ���bp���R����*z/_C�wO�q������R�X#�r�"ktE���*kث�%��9����q=�܍�6�������F�+��f�(Y���}Y�KK�j��}���2%8��r �O����y@m��d���B2Ĥ�'^�������v�jX�(J�����*�D:�g���,����T��R����E2��rO����l�?�	�V��V����"6f �M�0f`�-v�+�c������a���	�F�P�̎����M���wLIߐƛNZ�nXk-k�6�mv��������	�9���LP��Rp���p�١N? ��3,�Sk�	0k�3�)�D�����P��{I��o�+���QLC���G�PI<L��3�V�}����{�-�ةn�3R�J2̿77���B��t^�Q���|/22
&24E�ut�~Ĝ�c�a�FHeZ)j	vj��c���'QlD���O�NBA>VXӐ���B�x:
69-�'��oX��q��~�#�]�ģʫE:�)�D�S��#d���	l���3�0l=�Pp;Zi����2!�ڰ6a����/D~\$�\Do���#�����bI�`J���.B���p.�p���aBB1z%|��<Ʌ�:x48���-�\-s?k��~�)���F��<X�� �P�R�'9~�K����ò���Ӌ��}���^������Px~C���ɸ�B�<�T�J�o`#ލ1�f���ŧ�#���mq<��M'�-�)�K��U��1`�ϟe�q�ſ-o��A�7�ǥ�O����WS�d�ߞ&��[�tw�+I� ;��2@�AF(ĸB5��S._�F�~�!�tn��ʊA�#�O��_�+���p&�AߧB�E�w`���.r�e�rܡu�����j7�8�.�;���-��_x��_&�Bl�������v�o����4��W�'������EcNj�Ǣzx���甅����Z���#����i�Xr�mV�Z���~�������[��z������ʎ�`��8��r��_���v$����ԅr��M�PTÑe���?!����}Q��-�8b)9�]nf%l�M�k����E��g�s�p��,\���"a7�q�VGxk�C�#�97���,;�.??(�������50m!8������/>�1�H��֪�����o#�jO��œS��+'s��̐y������B[1)�� �<���_��8s�2(�9K��(��G7��i84��%��;52(9:u�)m� P�o_#�C�Ģ����SD�]��c2҃7�G#�E�g?��!ߒm���^��E�|F�3ZZA��0������]�2��ZФ��j���5��t�=p��:T�Y�K|��AA��{��cǾny���T�?Y�������ٙ�����}V^��N�MD�7_ѯ��������"���):O�,(����'�b�`�9����o�~2�� �y5��uC��Z	۬�(g�*8��dVP�z�{�B1JGɚ��z�
�Q��Q�Mї�Y�!�����S������[�z,e2~���"�ݎAʔ�u�Ļ�W���y��z�Ucͯ��}\��;�0o?a[p�H�	g��󓠳�_nU ����C�H�]�u!��9ۤc�e�ٲ��Gdw�*6F��u���O�iI�Ce9/(Hsݹ�pRR�o���i?_s�M��B�`J�H�����5�����������xEin�!��|߹x7>�dп�;Q[����l0�
N8Y1�z�=����ۦJ�R=���MC��4��Z�}K9�3��e@%����i����y�5&AQ�T
���J�,A�b�ZTh#�<��H�TD��=ƺ&<M��5����sA�������.EIi(Ad��`L�Z&�1�d�#rR5Q ٴ�̀D4�!N���"�UvT��i9N��_Oj<H�+c*p�0���� 6���'�|��-w�7?�
�`PRX���w����0���f���`Z��|T �8��q��Ɠ��g�FN�ʊ�پ���H�klZg����g�����e� [aՆU�/s��c`L�9bk��Y魞�\G'�v������UU�7�uS��:r��J�;�\(E?lߣ�xw�׎/�ZI�Q���L�|u�#M��*�f5�S~5���ы@�'�d�hL������?4VK[��g���r�r��hk
��%[���`Z^O):7����1P�\�I�A���%F��P�G@�=W��s�V���Ty�:��zE�E9��E��P��N�ļG���yy����T�l��WL���"�������/k���� ��{��쏞	� A��8ش��g�c����\�2��ׁ��~h�@dֶ�c�a�'tm�Vo0�k�6!�Ƅ�[��3T3 ��q:\�K@�MCp���=�xj�Eb����������_�_���8���g����G�8 ۪�[���CO7q�o�eNf����{��;B��FJHؚ��v�)�#��'�c;i����1��"�7��s�Z��_*�����c8��5ڢ��S��E�im�Oo��C�ɂW����M[�'�O��Tm�9�ˆ�Z����)�v���Z��p��r'؜V����c�iWλ�b5�;F��5�=�v��`�II+3F�q�[֫�*
�Z!cHr��x��̗���k��?��z@��	%N(`g,�@"P�ME�xT�kH|����&&�qB�$�%��\�8� �j"�:�i!����Z>,�7��E㪸#g'�g.rt��2r���wc��۳� P\+L�ǂ�S7��ql�3�Ҵ�g?($�i)�v�Kڈ���	#R|��e�T+���B0�r3�כ>ċ�*�*|cᑂ����5B�74<i��v���c`�5�$���dp���J�G#L�:�ޅe5��甾^����Ҙ�~����G��P���f�+Ԭ�bE!ND:��&ɺ���#d�TT��3���AAf�2���uBd�;*�W*��=%�Զl�pZ��xp[,\��l,���OyV���S�wЙ�Y���a�jj��'����JGj�-�eP�~�G_�'���;�f�����Ю��*i�t��K���H�".������ �F܅�D�G�
Ʀk�2:5/D�R�<�R9��֣����ZJ�[8;X�H�9K{�CyXצ�?��sTXbi�5�u���^#������k+��o���A��qݐ��r�~F�1ʾ�e�~!��d��|�l6����UIL
�2�����	o<xV��ϛE~�j`�3�S��o����Mg8�U��kS�����o���r��$(T�;�	�ng[�X8��Er��8�<e���4䜲��3)Zcԏ����&h���
�4s�s��9�fOA�B�H����w ��Ziy	l��j��j�~���NG�:�c��pq���b2��-�ϱ�!�L]Y���$c
���BϜ�Ċ�=I8f�,�f�4��
G����WX_&�H@����E>��������L%ξ��G�z�H[���\S�}7���YQm��<\]���u��5�~�eBȟ�4���ӓ�`z�H�>H������������z+�� ׺a� ��ّuk�eB	�mG���	���E3�Dv��'��Y������V���K5)�.��o��3/-�	�������}{W�jQ�ܮ�>����>���67���EC	\�N�]��������0��F�	G��p��D��uKv
�{6Ŋ%L|�D��)�0V/E�w3m�zz�E��C�wݣm��6�5]�~F��t?,z�2�# }������;*�ke�!�)?��~�����L�Ԛ�s�И�苓��������E�#�%(=AW����P���|Dk%m�y�s�#�f �-Q.�W��l��K��\!��;����[��W�I�B��r$zE3ќ��6��W��x�[U�_��+�=;����J��Jp�?=x&u���E�^�s��A��b���dTi�a���mo��61T����Gϔ<�
}����_ؗ����&G�]�ʧ|����_�O���~g�O� |�($u2<p.f��r���t�"R&������I���bå͞vM���T��@��kr�����,/~&G ���l�V�\��/ZJBȊ��5����M<=�ūo�%��VJ�d����"�"�?ζ����u�<�
٥R���W�	U�Yh�=�d�I�M�x)'�5��r��WmU��~�JW�[j����9��LUnM���J��YɅd%5y�������0�"}EE���.ݡw��������:�
H�&+��(}���_���,Y8K��y��K�oW�$����܌fX:0�'�<�AO�>h��<�<}��&��Q$J�8��O�<CvX�}`�k�'�����^I﷪ߘ���G�-�"9Ԫ�W8���p���ә�G��&��)*T����xc�,����$>g6t��+�٤��C�9>AP�P�����A�%��0�.����E ��)��^N:
z���-�����?�"�F�X���i��P+u4-�;պ����%�b�>��_�F�=�$�R�����i}�U�*P��5/���x �dRR�[�Իi��K�'c8��R�G�S�7_1�^�[l�%��6�L����+����y��]�oh��i!�4x�+/���'����j���BӚ�׳�y�ܻ�l�[���Y4�hͮ�s�����ȓ�
�:.X}ao�a�ogfg����҇����qa�,Q$1i�6i�&)fX�]uV$�nm���D��aBخ#�����[???_߳���#����='�����]�k\�,��V"_�m��s>R���q�?Q?|/��~#�/���>H�\"z�=��jj��g�Z��`W׈����8��%�hj���f�<��]�bL�=�A�҈GX��eO�Uآ�lm�����~�J��3{�"d޵��ŋn�ڭ9�d>����WgLo����H�B.EL�ؾ=�S�BMcV�?% ���qC
�v!"��?M�V��8�6����/�!�Myλ����eա�cH�"�?�n���J�_!�Q�����r��a6�����5��ȯ��H�3̀v׎�iⷱ���t���,�t,�4��)T��t�YiT�T��kVnc�"9g�=$DZ�-��e�&�C�kW���G�$^�d�( ��
�"T��x�x�r-�yp�8�>��c�x��������:;�}$s�(�PdRc�`*��⧅�Oލ����p��(��43�sz*�־�n��;5=tt�ذ��7�"$�+��eG���/�Z4���D[��5���DU ����^�>��p:Q���r�$p�c岮l�i�Ȏ����a�8���"-'�w��{3��Ls8��f�����g��*�Á2�_$�Ib|���$�w2�{$�M�p��{X)�ah�lDZ��,~�#9޼��L+%�!�|Q�`5���g擌#�9�� ���� �6P�S���h�~�\N�lAL�ʗ�c�e6/��8wDX�mj_$ɩ�>K�Ձ��&t�����k�R%<��~�R�QՂb� J��L�ŧ'���zx�q,�Wt�|&�0٧2�'��_8�x����{:�2Mm�I��}$ϱ��i��Lf�I>���:� �T9Z{8��a�}@���Py�R���^��I�j���$>��n��o��|NT;���ZPQ��0a��ZT،�6,�1�h��{��y��=��7ӫ+,�\�Ho���V��,]cM`�C�H ��[��V��@��q����H� h�R�7�����H㾈eֈe�{��7R��?��!�#�v�т-WW�܄ggV�^��\\�~Ȯi�D\��a�Y&�j�"���۴4��5��/��I�`�a�!\�� �XI��K�F�WOy�Xe�V�E���^|�Y��~wҊ�j�m�b�����������%�`�ҷ�Խg3k�w?��|�0~a�P���O��"��!p�]uLWjL�i�;rق�g�b�FPB#(5c"U��5^F@5TUTc4�#D���>��\I��ܻ�`�A!��ޙ|�~�z�Ϲ���y7zZ1�&���R�:˴�ƯF��Z�s'��ZLűͼ7Q5)fW�4d"��4���C���% P3ϖ|��^�؋��(�r8}��^m*n�Tr������bX�	�D��L����Lk��A�
��s/(��VZn�dAV�/��
��t�:��k�[:	��{�;�'����Y�Z��0�M���v:<v�5d=�י@w�O)�/��e9*(�H��0����0�!�dCW��T���KaA��]9���@GCo�5nL!G/|�ffe����R��۝$��Yϥ�	�҂7U���p���Z�E�pK��N4��������x[	�:eJ�Y���� �Z��Q���
R���٤n��I����f�������j�}�v5�J���ۈ&���(�d��7Z.D܄�(� �X�P���q�(�@OT�����d�~y�|�
p[�F�HX�~����uʎ�K�<)%��i�f�N���w򈔄�2��٨��������G3/=@�S�M��n*Ob�Ν�J,;p/.
����Q��W>�*LD�3;j`xy����k<1��w�vD�:��_a�t@��5�e]��6��P%U����Y��ʥ�g���u�`̯�s�ߘ��fF��Lsχ��	��//i1��rd�L�o����2�=�f��v�*�=����t��f��g}��S����s����.��4��]i��׷4���.\Z��W�& �q:Ky�h�_wb����&�2�����ˠ��3��o�1�  `#_] 
���_�� ��)�q�FȤ_�MJ`k}�fe;�󇷁�ǌ�<]wm+!�P(�'`ԑ�e5N��h��Ch�#"��BG7�5@W��D���F'@WǊ/H��?�Ĳ���2��:��} ���؄��з�:�]Ɓ�:F�\��r^Z�A�;l_7u�0����kk,J��a�h051'��;,.9-��&4��3�7oະjk��a��<;���k.�lc*iǾd뀤�g^�gd]���3��_t���@��Y�Ը�������*�"��!��j�:½���>ku���l3�ӎb\y�J���KC����4|҇^)�'.*R�!�H���5��d �39�~n�d0[h�K�o�D��vH �� q!(��ҟ���^�������m>�y����XNvw�*k4�N�W�yh����?)N��ي�ʭo�?U������ݝ�jr׶�$���c,���y��Qk��>��������%v��B��E�#R=I�WWֈ.�9�W������>ċW��5�\:�J�G 7?4�O�1yˠʰ�3��_RI����mQ��s8ϱ'�a/�A�QlQD�{�r6'>P;�%���L!�����7�����@��(ӕ	���ʹ��G�����6L6*�P���N���YӯO~�L��vc!�p1��t��ms�5nA�Q��J2
�}U����Kh��+�7i��� 
��s��Q�"@�5Y�}?����C��������P�������u��U������|���4R랼��^��Z͇��_���4�*bcc�z�T�|�du�Tr>���DI��Foj~~֐[����!17nu��?�5�mā�]+3��Ý�.�E�B ��n����������-�R7�Ѕ�J2\�ϒ8?u��v�� Z5 �pժ����o�<w������UV�"y�O-#�kD����Cf4��i��z���{3A�����zP��k:2�������wb�F'��,5�F����h�}E��+����f�X�Ň��ħ�YG)���!M�^����;���o�gd[�;��M��gEEm�	-���{�l�B1)7S;�Y���\tB�۪7>9�Hx����L��p���(@����Ҕ\c���kd��xs7����ro��i,_��_�S��_/��A�nH���{��w.Ir�k}.k���5�á�����������ΩӐ�&�J����/��cS�ԗ9���i᜝��~����8G5������+u	F��'Ȉ[�Z=f�n����h~FXN�6�zm<�@!���c�9�ߩ�6��:d-K��B�qquᝠ������$��Ǧ��~�����K��ᑝʨ�J�H���2�tЅ�߮R��N�h��~{�Q`0׆z�QQq�T ,�H-�;xI�ff�X��B�0Cѡ���a��Γ�������u,E�`^Pӭ7
�u��~��e�G9�p���[�q�G�$���dӑ(���q�$rX�xΘ���gC��\/�@C��{i���A�~��q+&%K4���^j'!>8��C��ȃ�X$6.��F2!�>'dߩ8�J�J�4:�h@���"H!�g���ݜ3����������RZ�߿~��Z�T	��"��U�����
X-�a�Y��\DPދ$#?9����D��U֑�����Z��4��%>7�B�C���F��xP�:�����P�ǃ��viĜ&+���mp��J�sv��d����l��[��|_��M�����&��g���-�W��[�?OmpN�3��&�鞄M�Y_�"��f��f�H@�'���<�s}aS�i�be�`b�"@��������� +� uu���gi�=gCK6@kU��u��q�mo�JXG��;&ςpSy��Y:� ���=Q)�,A�εV�M�m����puU�Z_ zb���({W��w�u��Q���(��8Y��RG��&:���0lL΍�Ʊ^{�>�KVH�)�־����zn��i���`���үŀ��J�٥�O���-^(,�-��<O;x�=[f���B\���PQtr��Y���̩(���i�Ѫ>�xt 9���iz�u2$إ��?�=Q�/�9�����i8y0)5�E{�T��Z��tq�l����|��(*OW�a� +#��yڝ�����R�?��r+�Oh-���y�ƭ�8j�v�"�D
���?l2���+v��V��i���0P3	����gB�"_.�:n��rKm/Z��+F'�0�F��1� EɃ%����p>���t���V�Ak�bT���Lz��)��@W�$�r��D|�&6s���RBuG&���:���4sL��S0F��i~������ѯ���_|��Yҗ�D.&��e~+��~��ӆ��x�a���t�qȼyP�ث���v��6��]Ϟ����$��UYx����𒓃aI)�2������'�f�Q�����!�u#�����ꛟ��#���w~W�Ng[����нGc\�8]���444�7���*Z��
G�t�O��7� v@�ή��鑔��x��/����yV��I�x��	;�{ݍ��[��I�S��7F��rrx���x��yz�	%�L�0F�ŷ�F�*�Vkx����}�ZGէ���y���A�?��?0����?��?4������T(��Py�5�D"x����O\堡�K��NL\�}�J�B�Z>9rcb7���(�c�j��J��:�C��}sK>kM|n�*@��F�o���bT#��kk�e�M��o.3W���f�׽��.C����G5%�L�����Z�n�tdƓ���%�3o�z�4 ��KA��h�`��;qF;���6oJ��\�5�_��������ń.��	8�U���o��Q�����zW�.($xA�[�q(Q��^/�HZ�����>L1�a9����^�^h��;��ݒ�y��8���[�"�����a1�L�Lk��C�O��0h:��4�J7)��|A�ԭ�t�'#r�Ob���9k�j:j����xs�ؤi�3Ц���4���i*�IT&��ŭ�$��R/�G�$p=p>��:C�F��,�$W�~`��
iQ��-�CS�|��I��D���hȘ*��np	rh���C=X0T֜�RY�}'�G�>pv�o|W>����PD�M�^v����턅8��=�|���v���`� f'�=����3�A�Sؖ�"9�-��Q,�����%+�/����M-6�ؘ�S3�������+}��.��-U��{�ŵeE355�Ǚ�`�F�Q�?R�yKx��Vl�2��Q\P�g�{Z*ҌK��w���E�Z&���.Ay`{&Cx�ٝ�X���DjJ7>1����mo�ճ�}��1��`���n�v`�+<�YAmYYqcmUqcs�Њ�4�ׁ^�AUU��(�?�"��ّ���1�\�Ϥ�G�ă!��a��̴uL��I>A8�;pGJ�P���f+.��M�3g���h@3,�^?�����ƞ]^����|Tb��*���삼�V�Epd�6;*y�t ��C����1X'Qz����3ʒ��%�+*���$��|�T$׿�p|�Oq��J���q ��^]%GY���p/�j����[��j�/m� 9vp7�9�;�ߏQ��j(� 
��ڹ���Ф��N�"�>�����V�mNy�ա�j��`HP�<S�>2;�8�� U��a����6p�Za���.$]2�ʹ,�+�Jb.��ͯ�-�6��V��T�0(i`�Dǰ�-�r�O|�p����C���^��]�&���hS����?돊H��a�mY(w{x�c�~�{`J�v���%+��T�T��lb��N��?��s$B6�� �!�*R;$rҖಡ�
ß]�	�>RR�#�=��k=��N�'&���S<3@�����9J�.�O�Q�6؟��Iǻ�P�xq"F�[�^�RQ��ӣH�j��ɋ�Ng��"� �V�8H�\��t����O���2e��nsu��RBe�y��G�F�S��r��n
���M>��pJLo0�r1��Y����� `��2�+����*a?^vnJ���`�4���%��(�� T�����ҙ���X�K@���%U�}R޷�n�5��|��:ǊGTk�����wV��$\R��CO |z	rQ�D�����Rp)?�fN��b7�yڼ���񦼤L���G���- ����[�"��R�_@��)��B���:��?Ϲ«��a�e���[*v6zfFjf������!���,��h�Bwo�c����OP\�_
��H�)n�rB~$ø��.i�B��e�ZYS�ݰ��F����ޏl-^��#�v�G���xs6z#M��{���2�1��Ԩ��A�E{�������[�<o��Z�٭�F�Dx���DA�N$��@�U��=oA3wg��ɣ�S�<yR��Un�p���t�Aaa'a��_̎O����;e�71q1Q��L�h�tT?�lm��J=��U��_} ]É_�R)D):=������ѡb~�+��9q�d�,)�
�LG�z��������\da�D��=Y@�#�x]�o�����Ɗp�q��Ĥ&�h�pvG~�$*�L1�;8�Rk���w6tLO�Q	�s9����eG�;�h�x5������:�+ً��P���g��S�����P�2�"N�5�}�%	0����|FϪ�]^_�%�t�|y��|<Q�Y%*�L
ɰ_w~���BB��a�fG�l8ܛO`5_󯠾NY��)��\�؇NqiU��u^�31u^�%*���ٱՕﲐ;�M����#�~��,�S�M�m)ݖ�(Eo��ו�4�{�&9s*� l��e9�䩽"
��Yl��{�f���0��t��N����L�Ѡ#��x+�_" ^�пO� ���ɕ���U���T?�����}n��BJF��>9�����eM��A4q�2hO�ݭ��s~MȻ�]p*��6�L�F��n!����ʡJ��y1�`^+�mר�(��vW@%����	�����D�������DzD�Ost, Ɩ����@	˘�í=t�︤n��t��y0m�|�Wɨ��X���
m&���2�����b�9]"yA�Q�hm��0򞴥��9�����h(�@�=ߪK#q���N��p�e�7:�:@�o�z��=�u�>���QӸ�<9"f�����}����Fٞn���5R�_��[m�%��"�}m޷�X|��B=��=����u}U�N?�a�^2���Ұœ29�yã��ڋnH���J�&�sߞ�c5N�WGL�7�5��rw����z�[�*�ڦ�6hILhs+������XEE7��GB�?M�ն�1:z8���m���B!t�[#�@+̃н�/�#v����[���ĕ�i?�r�؈lh-'��+v����8��qS��d��p�p׼z[/��N��ت�/�&��vgy�Ԝ�7F�h����,�nn@q��ｴ;��E�L2w��&��f
���Q�Tq��eK�ī^�Mϻ$�ظz�]���+eYq�-�h�{��Hq�0��\ʫs�Y�:�����#e��������F섙v�+���>O�p���K(�,������iH���U�y��2mE�^Z~�����\}�B.�*���i��ӓL�B麒z���T?�D�sI����&}�V�������W��o��G�.̾� ��뽛~d�2�>po?�~�;�����Yʗv[���^�|0u��<M����0��W;���+�m�j)M�v{��(�2��1�Z7�����zEF���J�,����o�_�(Vլ��A��Ժ�-޳����GO�^��`n
@� P��>��O��N��<�$Aʼ��q���ģ�x>���:���UG0�CU��"+I�@8���"��-n����=|n���	���S���ܻ#-���j5�ݺG��y����a���/ԙ�@`q����ahgn����5B\tltL�VJ:��p���� %#��𠷉"���$��$��T���:��&��:��:��F�&IY�̯R��ES�����x�Ҧ\�'	�%�1�d����[��k��/��"�뺌�x�Vbh��s��_"��7��w�p�~�3��N-�[AϖjӶp�0xdxd����f�ל������x�;�{�������p�Ӥggc�g���
�	&g�au�)���&{�����e��mH�~�-C���2�����'f&6&p���4,,���2����-�B��f2�<�:ۚ��Wmݹ��s�i�A�
�k��9q�wG�(C"�-�7Y�=r���L8sNL0��������y�~�ZTC���'�E#�,�}��4W�o+J/g9��L�L���M���섕��/O#�.��wN9��\3<�B�k�\&kE��!;]�馈�t?��릭�i�[l�b����J�%DC�$��\��|4�k/���c;����칖��ӓ�1�kL�O��B�7��~+�,%C�[�@�>�TS�����'fM?�����5���V:X�N	_����"���zB����iw���GwkVh��e�i?�[� �	q�L���F\�(�7����׼�v���e|���V!oH�A
c5��o���������GDx��~� ���,�w6�B����X�HͰ��SI���!O�/,,V�P�ߎ?б�w��'6���x��>~�!��MA����z�ya�~���O	Eܙ���4O�������z߷���hz� 
�y�Ŝ�n4�7$�6�U�l`�
h��z��J�E�}a5I�p?�Q4�d��P<O�ஸ�7!d5{�����@B 
 �����5�R���c�-��~߸mAI�*
J�@Z�T���L�AA��*=���C鑣�Fw<��{��u���縎�u��y& ��ܚfy�]�y?GQfz���M���+�W�P�t�4��$R���m4�%}�W���n�PJ�CW�D�ON���f���F�yL�{gswb�;?��]O��6����K�E�#�O}��>t��W�p6K���"�	DdQ-�Î����n����\��K�V�Fh��Ó��=\�t�)�"3��!PU��#�U%S-SB)5�+N�g�(Y05#5q���;�x~~�֭�)�m�3��������k�/8�;��i#Ć7�US�$����bB��P�ծ��/xS��sN�w����-t>�C{��a����Y�Ю����韸��bܕ�����5�l��E{�\���Ǳ&׉��rk��eԂcJhсt�t�P�����$�2*�g�S9�;�U ��R�����| ,˦nT�S��<�d�䂆zxy�Z��Ϣ4�i�a�m��Ƴjl���13h<�t�&9'�z�c�K�Ό��F�͍���]L�IS��|�=͙�Y�>���gdZfZ�$�a�>�[��#�1�py����#ތc��lXp�E<��>N7=n��+d���������y>�.���,�M��T�d| C��8�~�ʺ~�ߡ|e.���1'�a*#=�b"���R�/�^X5��34�i��ك�jWՄ`�fX}��ǚ�3�b���3{M{^ncoV:���`;�ˀ7�@��[r��JO����|�T�ŵ�����9J�!��lZZ?���˯��� Iv�g9��G�fwz�E�G�ˊƭ���b�q��&H��s��΍���B�	�¹������mmPk[B��%ٸ��j��-��@@UeK�h3Z"���e�4(�o��b�c��6��6����0�i�q�x�q�jU�8�w;��=�4�u[j�b��-��صs��k�_�88l��`
��CZN�
�ԝ6�6�l�H�Ǡ�ے�t�V���ɼG�u���;+^E�]HJ:<�F�L�L�����49���aÖ��\�tk
Y�7.&+!/�{#��6���@���7�a��4����k�/0b��z�g�����w���x��휐�N��P�󢝇��>�s��IާX�g�~�����/h)�h�����"5�k<r�#��~��ٵ���ף�5�棗}���@�xo�.�,�p ��m��]��4R�l�'��NH��0d:�jto���N�
%+��a���3�.y���Ԡ�/�P�(��^��� �@VlO�e�+�@,Q���}�sa����Z'�
�fG�RW-�#ϖD�O$����m *��� i�0�:n>%�gdָ�	���k�BTݢp��X2�}� o��22�J�å��u���E�kܴ��/SFL?Gie��UF<A�C���=[��s�x�~�����3��$AA�&*��J�i���\oa�l���䂣��A�1(J`�0*I��b�/ܮ��ɰҢo�p�ظ7�bJ������&��j�^绞�h:���{|O梒�����s/�7[�|���t���;_X����ܟ]D�]�^��h����wogc��"�]&���j��Mv�E���� ����T�ʁ9��Xk�1G��v:z��a��E�����$F׼� XWT2lqy��w<3k`"���g0b,T`�s�qt �A�������f�S��#��W����\������r}�(I3a�3w3��0]��8I�*�Oc1w�o��^�z�[0*��%(*��&���L�c�C�z�#���m�,�*ăL�#�����ޭ^����6�}H<�Ҽ"z��5ʈ★��r23mRMTT���@�E���N���ǁ]�^eSXI��SIܧ�_����<n�+^ ;ܶ7��v'X�[�q`n�3n�T2��@�����*5�<�Cf�[��4_d�~v����h<JD.H����ȴA1wl��Ya
cd|�l�@a`��(J`���8"-� ����ˁ��D$]���������<f�m]���N�(�>bv��B�ډz{;����'he$��Ǌ"_�`fc(�w<.wt���"]��lp�I�ӗ�G�]����О+�д$�B>y�o����&��+��4���j,�gTE�ڷ���b�%�]�b����*�����d	]���+��b~d����1��"����������CXK,		��Li�my5=������q���ql)ͯ���E�?L!�x�Y<��u������?��i�x�4z�I@�d4Y�)$�|C_��4��A`�����.kX�Y�s��2���k�tg��j�^��3�L��i��2p�&]�<˙�d�m5�d�e�w�"T�|�Yq���gJi��F�^r�p�BXL$�'����n5�bw0�t"���s���$��>��Fb$ �?��T�T>Sk��L���Ϙ��D�1:��%��^rĠ�����l٭�&�Vd�z,Ь6��W@��Q�ɕσb"pe-��M����Ą��@���Aػro�޵��*����$����ӽ{����z��2�v��t��#4c�Eѽv)u%ٶ8�?(|2�����kr⟘r�TO�S�ٳ���ֹK4+����r�w2v�Fn|�9��`�;�4�n;]u��-E���5�晌��N�]�2�?ܛ�N�O���f���36c��D�j�wz�� ���6�����bh9x��yғ3��V�[�+���-6�U:�L�P�^�� �K�HgTo�eY���4Qi{�Ed܉��nC����3�<�_��a��1��񮶪 ���o[�YUF��6���|��d��&��t[9��m�  #���mn��h,u���E�`N��f�Tve�+7W�s��eܧ4��Z!��O05���uʽ�#��c�w�#��}	k[�>j�h�V��(�o�7Z�&��~�/��Z�^��J������+x�H�8��oA����y��Ei�_���x+�#��M��n���Z�$ÕR}���+�w(�o���kT�M4Ue�ܴl�\��Ž4��U\Şbzjm!�a�#� �"썵b�K�����%��>JBk���r�_��1�����;ϕ�y&�Mwf�C�N�����>�%J�|�C)g��IJtvk���3��T�{d_���9q�S�����\��W�mS�����eki��u�d�>�����k�,��IJZ8��Ǽ02L݊���������Nk�M�G;�7�f�	�}U���v�Tr�������[��y<�XP@p`a�Qr'i9׺�)����y�e�Bq�Y>��Ę 8��Y�:_�.�$_��^X#>\���� �y�����f��+�_R����{��s�hJd.����j���uD��y7\R�5�e���&��lc{h��r2�'��\����t���f�(�g!`�&\���������'�����T7�LqS�ȥ��޴���h� q�v�W}�1��R��^��Ɉ��[o�p��Ԃ�� \�X`t�h,��y7�=YxJ�_b*b�;��Z�h�������XM��5��+�����/Yٿ�3kǉ!Ԋ�c�n�	\t}F�N��Z��nӕ��k_�E�R���
��N1�2����;3|�Q��g	NW��M��|�~�v2W�ŗ�������W��������9���5V�z����X�e����t���T[��߰ᝓ��
Ǒ�	���О�X;z�5��A@G�:���C>��e��wE�E�*\�0폒D�M��i�L��m��6{/�	n��+��wP�rHGr�}jҌV9��o�2Zd}>�C̘�B�]�	b	UG?S��;ܶIC���=����D�T����������33|c���ȹ͞�;����#%�q�\��[5����&x{���r�5�XYԣ�w����֏#*H�Σ[�^3��"��چй�m��>i�Ŝ�.�~����|�=n�i�耝!8�W��%�k�yfc�&k�Xjt�/�Jc���ʫ��<<����S�������$�(�d؟
��f���������þ��4?����!���(�b>]�V�w�̫��[NN���9Й�+��w�?��'��sQ�q���UvYq2�±����[)Է�;0ĔH>� (1w!MG����̟,���·ɷ��dև���׹��08IX/��)6*�t�1�Џ��@$@}���WY�j�F�/Dzg�m��uD܍��F����c�Ƽ�w�wI@��9���I��1w�5���'K"(D~� ��	M՛YA�c�����|޻���8GQ������d& ����K瑰���f)��˔��]�-�|2(�SL��<"�DiF�p}�P�^{g���*��ɭ��?dRI�m�r4tO%J���� @V�����ĚTq
�o�}�}<�ϕ�׶�RjS夈��o%]B�~���k-�d4q��	��ΐ�4U g�=(��N�^q�& ��Z��j*���l ��q���v���z�ˆP�¯��7�6��6$��46n>~8���%�RL��E��G?F�&
-/�1������N ]�nʷ�W��A=�"���k�l	�4K��x�B�}i/�Cj8t�ϳYAΡ�N{�������+h��ge$A��/�=TA��٠�*tȡ�����s���_B/O����c��!��l!8!�ԇX��tP�A��lۮ�Xs׏:��vz3-�Zr�b=A�	�����ΦA��TX�Dң|�]��$g��24��,f��h�j��?9��O�_oq�\,���/9]p�a��M�Q��KJ��92W�N�#��{W����{����gNwfjO��O�B9T�s�uF`�wF����~��E�L�(���i�j��5����B*�B!b@{� j+.��џ�-m;KU�x1�� �f���˥���3�ߦe}D��N	("��vH�eD�:��/i��fv��\�����e�����;�*;�R�pR+?�G���kh%����٫"'�k�J���'�ˬ��W�������--`�(Q cP��eU�����a�PzĨ� ��p����H>R`�\X\(K}�g�I��{e�S���>��'���zxu��q��ʊ����q��8�-m��U�T�*�6�'��/��޳L�Uai?��	4ү�mzr��U���������'�m|R//���E�x�9�EE:�&��l��M�7BF{���Nv/�d�JMaA$���[��1}T�*��7#�a����@Nvsv�U���̯�J�I��u�SgL�������_���8����a�ls��D ��7bgC;�6��N�˸�岲��π�̘q�(Q��*�U_��Ht���zC�|8�A�l���|�f~�
J?.v�]��P˄/P�GBI �<q��5�/ti�yi�oAD���#�t��G���I�c�'���)3����
�ِ��ou�)-��XJ�OJ˽��яpƍ�q�샴/&:��;�d2[rL+L�sLq����xla�VЃ~F�=a�O�s#`���/X~m�����Z��&��y,��C�P��]Q�܊�����m5������=��y1�D(i�"����Tn�޺!�i���Qx�$#��h�c8�)��=$�6��u�j��07s�{35K�����Ҽ��Fip�	��)!ZgJ嫚��6�(N��Ζ����[�7I) �������^�N�v�t����y�?2�v��R����L�i�ۿA�J��=�䖑TGM;eZ@��Ϝ]!E/��F=3��5��M��.H^�i	E��� ����3��p�����bc�iL)�
���� 2��<�p��Ls͸�>;��WҔW�]�7����)����|o�����@�ٺ��`w�S��f�w��d��ia��B�տ��bܲ���YO��Zq������N�l�����M�Wû��x
)��I��p;7$�6nvɿ0;'?ʏ�w��h�Z�,[��h�����W����^��/H��ЃeڙVO
H�+d|4��=��MPf��1����'أ�$O*���Wr� :�Y[���E��������u�z��=ۧu�V�u%�g�VzD��7��<;Fy
{b��!�n��ZO]}=�G������{�a6 ?����$$�w~����eV�,��\�/�
b�bڒ K��
�na/�3�gW!�%P���7���j�40@ 3�/�0�۪�@Bj�Գ5sYgo��!��T�.�]w�?p��� ��x�t�+e��w}*����]m��V�����\��J ��{y����QP��E�ݏ ;�:���Ag���U��@9�3�gh������I~�FvO�b���!�nA"_�Vf	:q;T�w��˵�SI".�w���{
�� ��H��
I��2�������ҁ�� ӫ�O�~P�G#4r7j:]��tL�w���2av����q�sM~�TPɛ���͝������������A���ڷ��;:�*�Urp|��S~C���ܜ�����cHz�/ۆ�}��:s<������ؚ ���9�<�rR�2<,9h��S���|7��!��6�����/��j�k��w��wۜ�ʿ��V�	�i�y&�i�h�%�Lu���=Ij!8_����ױ�J��}��e�v�46��:&_3*Y��?��^�-��Ep�&J��zW������T�R��'��v
3�x��V�9SW�7{������t̐vo������S� Ł�����RW+�7}����Cl�sC��zB���b�ѧ���B2��Ȯ��N���cy��_��u&|Q�T.��_E;ߒ����@!k���z1�ޜ#���6�-xz �L���#���fai�b:�m+v�Ô���*��v���AS\�� ��c�_�JVF�rM�`s���,�ݻo�G���L�I�@�PH,��nm�%�L�i���t���M*.°���js�j�Tl�q��6��{L���{�w��3w�~ve쳂�9��Aa�56����j���p�s���.\O��U���_c�m	��⫿N�W����;���7�N���?�5 &χp�[���0iLE�:8��2��+ i���e�M22ʈ�Dx3=�D�kD0/w�f:B���s� ����Muf�˓�y,c�2}���a[V��7V]8Q��~�8Z�4S���y.֭5�ENU�S�+V���))a�g�2�j(��<�c�t<��i�;t�^�Vr�V�'�ł�D8G'�4�̬d��ˡ��ar<�^#>Y{�;��%��2zZ���N��r�ò�s�qz���8��g�/d��rKz5v>Yd���ݹDB����,��;S����@�s'��6���7=Y�vBF�m{��N��qL���Dj<A>���d��{����q"t��g�k]����Hx`��>!9֔���7��j�<!�I�L�S��I�C",�&���� 8
;�Qҵ�;?I��JU(��٦�Q>1Og���%�s
0t�*�1ج�V2�d�;�U�S�۲���u��Pb
��On�:aJ�;�z��F�TQ����.~/���\�������ĀxԈ�q{]~�5��C7-Ѹw��0��Nf�#f
��9���.����_H(��9����ʶ1~�y��J�kz-��L� �)@A%�#�b��	��D�=��u����������Q��땿�g���g ��/;�`B}��怣{�T��T�V_E�=&��}�7A���f��{�hr�'�H������D�b4}��,��u�����+P��yPu�r-(8Vw�L��[@u��fԑʑ}d���i���LaS;��W����`-���T��D% �[k��?pŴ��Oxf��B���px�~���:rԮE�%��[?o��{����D(Sw_�_�׊��g�����,�����!��1䃅7���X�3��I��[^�&"��F��X@�"
�K˶�Sa�D���C�5�~�_�I��z�H�W1���������{Me�f~v5u�M��n�3�W�YXl�6�zֈ�{����~���<�䚶�H��7��L�I]!�b���
���y�%���?Q�Sw�ϸiQ@E[jIX�W�i u�N�[~��Q���M���jrd<�)�8���U��J�������R��S{5���M�>�aV_N�:Dg�ǿ�u�я�dJ������MՂ|�Qm7���g�Z��'��s3zu	Х��SӋx�jWjr;���F �m�yKu�zB]C��Èe��""C���?z��������)r->>�*��~8���֨���	�]��#��� ��c��m���u�F6T��r��q.����L����H��L�>Vm�rhW�����|��?�t���o��I�a�p�L�g=͸~��}��1���9���������h=�|=y}��w~�Y���3�|V�eN�/ܽ��w�E�X'=GZB���W��b��JK��Q��2w�LN�!l�������RI-4b�$k�a�U��O�n�Z�8j��D����I:���%�
e����L?zZ����^WJ
WF0�����D��T��F(���x�+�{��|
;��'H��T��`<�#�^�h<�k���L�0M���8:��x��N��~*dl
K��/�Qf`��$����v36+����%)i1� c�wq�Ӵ�?�w}I�!�荖O� �k�@6CWH^���a�XG(�Om豫TӅ,���Jރ���E�e�Ф�}�*�ߔv��ߒ̎Ď�Ws39���Iت��[l��ߣ�kv{l+�Tq4�ގ�~�.�E�?55�rRc���C��Zx�O��/e��������[ݖ1��jo�gX`]<
���.؊�[?������M=�����Q���ŧ���Wb�f�O���vF�ZAwT�ӭ��rCW��rYh���Jqc�>��)Ɂʡ��SVh�cc�?���@&�Ǆ�Të4)�����A��5�.~X��o��D 0��ʵ�)`mC�S$���>��K�j���)�����Lg��u�Ο�Q��f�U�Ku��ܛ���A�C�9�1o��MY��ӑD��W���s�k��� ̆����5���x���;�S���}�K.p�{q�*~!��;E��sg �	Fm��(��T�j̄ ������nug��a$�ԓRrI��$�h��v$�kܕ��j��	�0��Tڭ!d��^��%'��� �@
���K�\�o���A�	���Y�m߷~V1��wU�{ f�ަ+B.�0G'�����E��0��%��@���-!� ǖ���.�k2e,���
p>L���L��y}��pT`��_+�g���+�Z*�.֐�|8@�x3 d�W�����E����"8k����ef$ bk��0g���2�We/��l_��4^�[Y��h�L����	��`���T�̿4L\����`���Å��4��[�$�UiS����C�g ��� ��u��ꖬDzEG�>K��H䗬vhl �A�<�z,�id���æ��D�0��w"!<�ZT+yV]<<�m�����G<<j�1eg���a�{;k6	� ���Ϸ�����1|�F�%�!b@ʕl��wL��b3UJ���.�<�¦��֭��_��d~Ӏ�b'MMME/��*�[|3��ꔛ(��AO�t��*�&�.%ƈz�6%��W�Z��d.�����|v���:�/��1w�2�؉{�X��z۟j~��:��a�c���;���dp���	��kT3w}��|��;���yϨ���z�����Z��2�u��h��(�;aj����t(ʎ�K�Q��V̊�	���"�R[�k_�Y�^A��OQ���ܶ����}�]c���x����k�*��ED��l�>T��FW�y팇��.b3��3���d��|wP�_�f�r�[A�İ>l;�Ȼ�a#~l�@��ɐ�1v .������l���f�G��i����z��R�Ћ|٧�W��
���`����xQ���o�3̰*e�
�ʺ���8��r41����-rڇ���z��c�@5X�m�J��UPK�=�o���)M�t�V���K�5�w��H�l��Zo�6�!�l��G~D��(T)�c��1��[�
�_ǎ;�^`�2ݫ����jޣ$O���uJˉ�|������>#��ϱ{���gr�ƽ���0jO���W8�q�꤄�JQ��f|�x2���.S���d=��{w�u3�Vx"�b���b@^j����>I	=�ZП�!|o꺤M$�?Fn�f3% ��Fp��W��N���$m7\?� +
�EzV�o�\)���r���s�������̌&���N� x��ю2�d��]\gg�I�N�H�5P"�hA���K�"-/o��4�<J6'P���{�]������/[��A�1�����%	+8�p�E�D"�/��KΒ�Z����F(�ݹ�e�Y9�Z���[�?��X�e{K���N���^�\b�WbP���2CD��qG�p���*�C��}B���p*�<��� C�ǐ���6��[���>T��J��A�	����o|�*���j�(���mn�����"��|��i{M=B�V,�5@Q�r�L�DX��à3���Y��l��,$�^1��;7gb�&
h�u��φ�\��c�6��һ�[�Qng�F��u��+�u)���$s�s`j,�{�_g�M �*ΰ���)��|?>P�H�o�9�������]��`��T-�8p��{���d5��(��?�`dg�3Z���ԛ�x�v\!5�� �4�ؠ�F�o�MUo���1mV�|� �V��ʓ?_�1�:q�E/f�*|e�MM��Љ��%����{YNTt@�dc��2^�SP�2�Y�̨��1Q�222��!�^lm��/���rY��EF��u�Q�?�C�j��r���Zʘ�b��FJ�����v���E�ާ�)j2��{HV�
��х�����2������_�%�Wj���X'�������3y,���?,��Gl���7��p�2WC92�>;���Ý��{�[ޟ�`�A\P���2[��U5��2��X�ٲ}�^���}����b:�	%�(ZC��W�0������&�p����C��E��z���n�D�Q����QP0�^&?���zO7�;�V�J����o�`�Vs3lr(E2OW�>Lz�۾��6baa�#�IȊb��F����P�lX����A�rAr�p�OSBQ5� O#��BċªW�U/���|O��z�p�v��`����� ~,�ZZD ���]�zMcC���;hMCK7N~�'�]� �`q7y�[p���\._���o��@8�󸒴V���r���-[��Z(��^��������$$�|^�Y-T������g�R��7<���ּom��ݕl�b��_�0��nVg��x����w@B�M����������em�2�>^�ĳ(9���뎞^���JS�V}\L��&.���2 }^a�J��*V��F���r�*ʦ��P���u�I ���EB��P�\TN�&øV	�~����N�,��q��t1ڷ��~��jo�����!D���ܭCzz�|�8Ki��ىh�8�$�����"
\���|��g��Y�y@���7%s�S�b=�>O�
S�����!�@���SD�7�2��f�5��D�0>��Y0�'��j!��o(;_���J�����,�	�|�Xd-�B��r�^2�����I��$؊bq0�X^UkS��n��5i�J�g�K�{J����7Q�G`��@��Z�` ����p�*י&�Q�������B��j=���*���^�)SmQoZ3&���hcqD��7� D�	�3l�W.����)�Q�PR����ΰ�l�J������-(�\3�}�#i9F��w����1�p���b���۟�r늴���2�[;@j첍Q=�� d�Do�w�d<�v���; ������)A�w�����%O��\<�+��w��??���9�u��IR�+5��{UTL���V*���yf�>h�hI:����1��O����:X5YTy<�6{j��|2露h������%��&�Ȇ��.�SUQ����R�\+�Kc|����{��yj��lȭ�7_�_������=2R��Ǐ>|pT�N�b���BΡ��w�aOS�����|�]�L�� ���y�S�iܹ��i��U�M��Φ^�	O5<��]e:�_���c�Wc�8T3>�__��a�S�/X��q�������w6u��z�@?�}Ux���}8�͗*Y��=J���~��*���lr�Z�!���|s��w^ߔ��ZYO�\����xK,�V������J������?�^^�{�Y�W�?��y���E6	��u�.�#S"nuN�+�ֳ>ۘ�w��&�U���"c"ߙ�"#q�-R{������9 dW�j���Ҷ��PV�yG�Ǽ=,=�/]��R��2�MXUq�������+��O�c��B��R��e��[�'��Nº��b/�7��B���"ߏ���W˲L����� ��N^YƮ�:�gw���A�U�����4�xF�[����8���9�AG�H����P�!&��̡36=��#���Ҏ9���?,�Yܻ�ؿx����������n}W��rc0
��\�{_mEJ'x��_��O+��Ng�6����7�ɇ͈>��t5���w���'D�_�ǁ�K����?j�[{Crm��DP/MTQ���)�Iw��ځ����,E�K;��4Wg0��ȡatTbN�p��iE�����0@.�K�uv��jͮ�~��wƀ�l2�Nj~t$eJ�˨ޕ����X�t��CD"��n6v�/g�N�����%�DFi�V7��
�d��dSB�H�@�~�W0��KL}j���`���f���V��{J3�Q�[������|>����A��6e$�		3h	8����}�ۗ��I�=�RA�c��ׯ���$���U.t�n��Q�h�y��n��葝 ]�|U�xFk.�~���D���/j�qX�!�K6 0�C�˽�c~a ��+֌Ԭ℧=~ �O���{���u˳6j�;t֐�}��!͂	aa>y���G���}�#/�J�+���F�I/�S�ނ�=1亠X�4 �>�f���W�.7���b��l>*�N(^�Pn����I}�s�N�)4�lmc�e�E�w����T@f:^����YNk~�0P���|U��14�nӉ<�����q9T��!������>�(}���9(��vT�U_�ɰ9)D�C!7G?��Z���C��eIj2?�]�j!�R����₂�O��t����Q�}[�z��,$$���w]���g�˛B~/"ݴP���v)u}a���c�5�elwDv�&>�5I��7O��I�Ή^���]��]/{�'�\��5_������7�wV|}���|�S�������?0^�}�ݝ���u�3���js�7�#�(zV��+;}h�i��>γ�\pm�/��Vg�Ia���ʲ0��i�6S!؅��Y������rW��f���^��z,��g�M��J��9<��g��F�wQ�N��rW3��M��5�K����Qw�?r+��HNN��;������ܼ�"lBsV��V@�Q�Q4�(+ ���������������o��s{Ԑ=��.բ^�!��(��^��1[���^�Q��Se�%J%"�$뢔�t��p�W���N�Ihr�9&������z���i)����ȸ�i���v/��1+
 ���0�ŵi�>�+�����sbbk���ǢR�����[z�p06>��2F��s�zߍ���ϕ��~�9����棾�&,��|0��ZM�0����e���v����YX�5$�_էS�Z�}�	��=3+h{�R���JD��y'|�9� tg��ɦ�E��������*;z~N���@ ȝ����������69C`�)ن�u���TY�'}K7O����7�o��%��h}S�ު����T�nM���HV5�Շ#���׶�I��R��>=�ۀ�U"m�u��ސ���P�mZ���`��ҧ`�/l��v�E9!`����2�9�������	��v�/Ě&�����Ie�JKڟ�AA w���0�W��	^,�<�?�\�D����hAw���S���Zc3���2E�"����-ǂ�C��-T)Ռ�M�\R�)~Cm!�ɬ�s�䂤[�"�P��-o���2��[��5rR���^@X0Xc��@	�E`�Ut>)�݌夳�H����5�n��=��n�}�&�b?Q�&s�/D���>�l�'�t�$��5&��,��~U�On��WM��Q��Df���n��ڜ�qÌ�񻬕I m=��0e�x�y7�֨?B�!��¥�RQ?��J�F\�ͽծ�z��1X�A�p�ݥ����yH�u��(Z��ݎ1�G�����x0� Ǥ�UÅ��Ѵ�\�\~�bA����sX�Xif��<��mcX�B[K0����;	�~�v0T7�jᴖ�5�A����+)))$��~��	�S0abff���ceM���W\�_g����"/��h1T8�#����p})t8�zS��d�{Qjӄ/n�qGM�檒��~�j���A�n�� ���U�s�泮�노9l���%^�X/S��v�.qS�ס���9�ӹ�u��0n�sj|�|'�cuo��';(ek�����&+8��llDR���s�q���.�p�bt^w��b�/����2m��{�O�#��7�W}t/����׽Z)�����:eI�*eK��d���Zuv��|�I�e���D������%Κ�jg�\M;�x�7���'H[�Vd�}/1�1U�Yh��cO`USS�>$u���>Ƌ�T�c����Ѷ�����|�Oe��5	r���U�pd�s!��5	�Ѩ����eV�/��I���~�@B꧍$ �'&��Y�rA����ˇC��Qy����Q���6���|�[���8xh�oe�3:6*�]E�o�w95$Wq>o:�%'~�%��ij�7k��\���K)�gNҢvz#�Ʌ�WG�c|ͮ'1'�J|�&>�q��4w�&s��s�~��a|�wL�"Ƚ��@�Ew�ﰃ-��L�����frzxV�Y2�k��jBx�m�D�����ڷ7�.��5L�WXY�����(���Mv(Ƚc��I����a�O�p԰��-��*�kF9b����f�N5�����8�h�t�`�����Q�E>x�|-� C3����ժ����(v�89�a�K7��-lU����C7�V����@f�j>������[�`3+mw�Ρo�4����%j*g<eW��xK=���K H#�oRC�<��G(R�Gp@~���v�����%m�y�7�<~��eZ�_��8R��"$a��ZX�d%�v�J�T�Bߍ����L���m��q�O�`/�V<Iy�Xb�KH��{����Э��SuYS���N�Bq*.x���@Š}�� 1KeJ�
N����?6쾠� �i���l��s	�����=֐ ś2����Wͥ� 90��g.�
�,��=>B1뇝n���7 jP}X}��M�?��.Q[�=yP�2\�h���M�����1��'H��B�O�Ͱ��by��z�e1�X�D}��w�s���2L� ��4c���P��>���/u�Q�5D�"��]�Q�چ�o��7&���B ˰����ڢl�c���maY9�B�Q�ב���DjX�'��`4���!Ŭ2�3��e�uڤ�=��/��&�,�@�����#��� ���91b���Q=��V.�6x{+��9T~�g�Q����Rӱ�ӥf�	�����*//��I<�ڎv<	�%��K2�[�^+��I��j�oM���K�><��Vk�����:�릟��K��so����w��|�/�~Y|�V|uF/�=��^�����?��:�>8�Ǻ�\��\��\��_]�D��9�� +n�>��RM�����c��N�l�]5w��ڂ4a��!��K�\�̎�Xs�]O[]dy���[�+Dx�m���[dP�ǆ8Ș�Zd����?4sy �|�1�ɛ4U� ����*ㅑ����K�+�=�r��Z�>���+<ei��b-��9�� 	�9q�K������c���ccQ.��?� ��:��$���_>�;$�ל��
($ݶ�C<7��^5MT���O�G%jF%X*s�Ef"_���|O��^�j)˸|m��5�F��Ϸ��q��F�F������ߟ;������P���Z0��$�]]-���z^ Hd�4�����: $W����1������!I_ӤU��M�S���u��z!>6��q9�Q�$V�&�zv��9.�^��>�r2�8����ߎ2�����]v�'��0�Oy�	�S��d�1��2s���$8�<�#Q�c ��T8[��zZv`��C@��R'N%s�杬�����:먦����#H3E��J����!��@����a��`� ��5'����o~~������9�;���{ߏ��������T:jm;�-	�V���Dn���������vߊx��ʘ����a�����v�J��^���0��Z�'a�9��]��۶l��5��=��|6m���Xkf|ٍ�����>7y�Rz�@��B�"�ok7_D�yz���Xf�}���9�<�yZl�flSp��2EL�����Ͷ�kk@! �ޓ����>����+|pE�Q�Z��G�o�1m��\v��:�8��k�|�|��[����?Nۻ��-�(v�r�p-�'�k��T�,�Jt�^�*�&7pk˳�y�~�׮4��/�xO���?�K��i"��>0�hG��ߑ� ������~��Y�_^B�@q`
^2nfG0%,��M0C�U(�F٣B@ݨ�GF�$f�IϦ֠j�kZ�G��p�S����[�_-�S���y���͗a�B�>!��8^�J�ʸ��F=�k�s����[������i�Y[�f6Nr��b�֘�0��#�`i�L�$˶�Kv�Q���G��'�O�su��0�47��lc3X�Hc1M�����Qa'B�ߤ�����o��B�����'9Da宖��4=����\b]����<�w�$�*aܿ1o>�)��e_��8*V��k�Z���f���+�]'.@�B�"N�c[�]G������i�K�ޢ^L��U��iU�;�pU��*r�,���b��t{����A�f��y(=zuA�wI �# �c���ҵ]�F&k���=Ϟ�n��X1��J'��f�o�?�������S��j��}h��|:%`�������������nl$�$:�o�8��#�{�W�W��E���=d_�tj���_�g�^K���1�8�W�6A��w�,*}x�;�g�e|��]T~e�ym�L�Jw0U��<߾u�x^t����5P��<�nT�HC;Ֆ�W_o�P�w��^�Ka����/����,j1}��8�i�+��^�Q��qD�իcg�Z��Ö�M%�����_U����	�K�ozJ_�7�/4_d�jc�է,�~�N�mu1�͖�X��8� �H��*�7i�&J%=�\�K�G��u�f���z`�5OU��qb!�/�����9{#o#w5Ww�q�TxSa�2e?w �&��|e^K���u,�h��ڥ�.��,`X��}C�}5�6ߗ�V�������<_lqb��n����BN��H�� j�~�sZ~�
��~�7�(�#~�&hV���)Ǣ�$�z9�bzuQ�Wiz;W�h^�ez����g�χ����ٷe��#-ǡ�7=?�D���_ת�ӟ+~Q��u�VK�J�Ee����~HR,�S�}�U�m�
?����~���l1�{�֔����M5j�T,���o�
d�t�����eX%����Uc��[�,b�C"�Я�,{�n�?V�:e��4�ӯ�����>���O��<ƦeTm���z�)��w�BX9y,p��Y�M�g(�Z��PK�=�2��iU�̇)���]�f0��yH�>�w*����){�gL=z<�n��ֲ#����6C�O~0�|&�%���(\ݳ?�)�%���=w�y�OP���y�{����xh��w���&�Th~sz6;��Y0͈��C�����Rs멜��\I���<�s?,rsɖ��|�u�L�Ir��^{����Yh0`VO�
���>�X�0: 2���<��c~h\��aFM[�i�j�MgT(�d������/B��G���JL��<H��$f-W 
� �-���ډ�d��;L[R+�ͺ8�M}����E�a�tH��v%��_D�G�һN��u�ν4��jԋ��|]�(6��<>�|�2$$7ϼ����h-�k6��7�S�( �Xx;��s8�Y.N`��]����r�9�,A��ׄ���d��E�A"�\�����'��푽�(�� a�ه��2Z�=��ۅڟ��q_$���LZ���$<�I�Ǘ)PU�'�J�5{1�vn��,`���K�Z���u��&58,���T�d�T$�GT=p�'��6���=�4� �iH���OgL���B��YU_v���#E�{�gt5i"u$K��:�Z�Rj�Y����(�)i�i�磽�G�nL��8� ��C��\�v��@ށ;�c�F��!��Gs9�gT7���q�HL�m������+�X2�T���5����L�ɭ�X+�3��;� �y�����.�\�N������v�[���f���9�o�VCdG4�wB�?'��q�>kW�..F���5zka�[�^�/�i�z��'��L؈A�D��rDV��qj>}���G*eDeѵ>*���/���Xb10�8B�Z��O� <n�_Ս֪ ���-��.5B7�
�CSU�cn����w�(j����z_���d��	�i�i����^k�^�������J���1���n�������Q����H��g��뇋|�����+�e�g�e�wk�/u���:���K�|�G�wd��3񰉔U��4�;缍653{�ƷQ�j��Ķ������L�^�sy�Q�S
���c��k2	�n?z�3Ũ3i�&r���g�?3B��5���� K
n��ƨ� ��7�T����yL�eg{�B���V~���:��~7������޻˧\� b�J�m{M'���pM�.rr�ݕ#Rׇ�7Ȃ,�*���|�����
끠�`K�E>^E^Z��r�کOi��>�l>K���3���~b���V��/%c_�+%�!ŵ$ޮ�Ck�$���b�c;��g�|���g[u�Eмr��R�2�����7���� Z�18���΍5��,}(�l��-m��x�O�b�w��]ӴK�8�\C� �ъv=�gv������V�@��<|%~��?t�ڬ�{H�w�|Dvc���m��^?�+�;<�����>;�'�L�|�0;`i+J�7k��ٯ���i�G�S��֏�����7�z�oX6���Q�"zoZ�Vo���ꟹl���5������׷~�y��H��e��ʵ�3%N\��ϖԬ����O��n���P��^Yu�5���G��@�*~CA;3k`e<=�����?��OqE���C�f�;���Y/_)5V 6�@�ó3I-�����Q͒��>n��Н��s�u��v�f}-�GK��K�"N{%;Ʀ5�s���FT�:�֪g5����Dݿ��I��ezD,I>�/���� ����a��{h��$�U�����>I)�L�*:81��I�xZ��wq��;K�^����;�N ֖U��
d���L�X��ǘ0�yჁ`=6�ڎ��0���T�H��rʚrH*(<D�&eN�yB �
Pɰk�1a!��@�t~lCx̀/�b]Q��uOI?�A�	Ж�=ם���L����L��b��D�9� �+J&^Y�.-�:rt�w�zq��m+�d�V�E�?&��.�9by�7=��j�8��j���Np�4�1��7���2Dϩ�]�R�H���/X���/���	��������o� oT=X�;�|����%�;�,ۮ�^:�J(���� <N�6�"�ma����*!��m�2����G|ʒ]��DU2َ�� ��s�3���P�[����������n �lԪ#`�����O�[��i�92��d��"���M�}0�ڍb�ug��3���=�~��+�`���ɗ�pwԖZe:H�z���-�s<g?<ǼFQ�c�(nRT�3�T���a��۬�g5I�b�$ݓ��G[�ۋ@�@W��`����Bo׫�����b?)�2�OEӫ�R�S�j�znB�֯�~?ӗ�5_�_��=������B��MW�L�(*�v��s��d�g=�jX��a���jf��&M,�,�o�/��˳�Hxs�g�nIu6����|���q~�N�o$�-ؔ�İ�713�����ҾR��sܸ��N5Z�Xq�N���/���ֶ_S�����Nփ]�	�Y�(����QIy�jD:����j*?8��8����18V"��<�vݜ���^h�8�:w2��v�� j��a�5��U�KT�6 �I�	�Φl�}���A�:BI��{P4��Z��_!U�8�Df��Ddգ��/h&�6{����\H4��� �(Un�J;�����]P��6�'<T�����foªA�����#(�oL�p����;��Ol����C �^53��'l�RKE��J&�^$�����Smxz�q�����gn��M�������y���}���F:2�h�̗�_���C��6Dm��:��=�l��߳�fv�Ol�l��y[Q���0��p2H!�Íg�m�Y|5���3��yz� !�ES���P��îC��sun�29>�E�;��-=��R���PMN����7`=��v�__�v������vFJ-���{������ڿJ��R�����j��U�*u��P��?�H^a�IT�� FЯ3zLՆNoO�����u�U�����#;@Ĉ�U*�0$�=O�B�c�3�Ǉ��W~�m>PWUr���F���l�J	�^��(}j�St�n�b�!�-R�]�<�#[&_�W��~-�b���(,r'��AU���\9���^@��f\x+�Ks䛁S���{0� o>M��}*c*I�s���Ϝ��Ћ�~�nwęN>)|v"h�(IKA��yJ����]�Sv�`;��1������������ٓt�����_���>�(��|!o�s����
}\
�
��v��^�C�6�ǁ5rl �P�ؠ_ ?)�yT�����%c��Ke����P.��&@^N;$��I����[�i� �Pi�|�V�����#,�6����Ž���ޣ����/�ӑ��k>-�l��]�	���})�
������:1��]�(@��n/��z/AO� @�;���B\`�׷���刃5��	��B��(�֒l��.9�1Y����vKr�k�.�pvBXC*}˟����I;(�Т�̊�R�3�WO'��;�aw�(V}#��\rYq٘��R�<C+(�*)�t��>���d�4Ϙ�y&�ڠm�$��C]��cvԨ��W��:��6�{C�t[��[/��n�[/�D�9s�h�����m�p�+��Z�������?�'[�����$v0�����������E�����;���1����qS6b��=X4έg�Sk�&iq�����ќ�J� ��C�^�Y���y�TL��$.�L�X�w����?sY}ܤ5�a�T���Ѷ]LgR�y|=�Q����c7,��e����wi�Y�M˭�)8+���~�|�֝�l����ǽ�8r>h�A)���oj�&B�<���a�.�^�<�!W�G�]��w���x��l����h"�̱����h�
�! 1E~�W@�=��P��/I9�7��J��^�b�Iٟ�G�&�ۤl��c[�o@��<P����x�p��{i�h�~�ر��q��\L��Ky�}88Yz�p-��a��5�>�U����t��\_�;�5�s�i���]�P>PT��Ah�mϖ�U��Z��ot^1:��W�W
�����E�SA�פ0,��V�N��'�. �����Ũ����K�^�sJ6������pɹ)__W���;��>C616�ψ)H�T�����k��y
���=��~C�������-#�Nj�� \��
F���1����]WɁw�o%�ފD�@�ܫ�S1���	J�S�(gB'r��/;� @�dYΗV��
��������0�a�s��kZnYy3�xN��H*�g�� s:�$���79;�@��f���bx���~�NG���s��S�����éRuB�T$)���2,'�z�-H��R�o��HY�`|g��F�QEeqN2J�S�F�( �y��PB�bh^��=|跲�~��b����:�����&����o��\��E�˜ M�^�u�G�s`x�a��,p�;�Jf���<t�.FD��~���l̉\��0,c!�T&P�.X�Ɛmr��[Kܶ9�%d���&����#,S�N�����)��'O����؋��2_sǜj���Ġ�.B�� �����}�,�~��£L%M �铏��w��O<�����G�һ�R�9�T�_.��L����hw��y_�!�͙E�R�uuu�����"x����������6��[�B��K�/��$����6S�y26�`�	�b���B�~��Z/��[/C�NMo6�[/7k�o�k��G�� ǟMo���9Z��΋������7L��W!�����2���c��f���c,�}J���ۯi��N�Gxb
7�!�*���;���c��Y�Q�ٍR4������e���ե��.Ao{�C��m?��c�܎�ߟ��b�:���R��j.8NMꦦ�����!7��僒y���F?t�ۈ�S5p�Կ.�`�~�V�|���ȳ���Ʒ��`;S�!��҉l�r��^� ����<8�?����dȸ;R@�_��eU� �B[G����v-�G��=��yOS�> �~��Wʠ%�+-�x�2QP4md����~�X�o�m�\�N)���5�S���_��
H�OJ��q�T̔?-.{��~�gߟ�T�1K��7Y����}}��j='�m{��D�O��[/Ӷ�>_��Љkb�n�\�D�r9y9z��9˫t}_le��j8�ôީD �U���p�W%�fT��ߨB�^���0@0����Ko1�k�	V�����U�+�@(�tdZY9.l��1߫/g@�����A��`�N�mr��n�J���r�ﶱ,C��vI>�2Jߩ��NO�#|�!��jE
��}6��PFK�sd�编'��lд�ʨ}��^��n6G2�qC�o� �@���/Cr	�ݤ��?����4P**�~���}$R��I5a�д5�v}���t�c���@�0T�vΧ��.i'�:sXhoG?�֭����73t�
ՙ��|fBLJ�lLo��������m)�#s�N��H���o�@�`�9��9�~	����7��q���R�7:��ϴ3P��c;y����6�Z�a�|")�	�3A�����+{�C)�;O�
课�8p8���=�t���J!��A���0Ln�	�z�WՑ~@�ѷ����-V�0���g�E2�5���r��=G����� �[�d`6t�? y�L(T
�<D�+'���H�!볡��ɂ��Cȏ|�N��o.�YE���������4_/�P'�y�z9�|�W���ਭ����MB�[B�ZI�D�9՛��x�;1�j���7L����r7e�ې)?��RD���%*n{=v���J�lᶇ��n���n���v����1;�|?�k�Q��Tv�5�p��k�;I?�;j|t�ܻp9�wX|v�n�:�>a�GM���.rٰ�UM����S¼��0/�Ϙ�ǜ�+
&F���d�2R��L��f���KW:}cI�_m�^�R"�۴ט�0�ۣe�7��30 y�s������ܜL����V� ��C��o��<TP"�r�,� gwe*(V�5;�`G+Bi�У�lLQ�B����O��Х�6 ǒ��dT!��,l��q&u1?#���;�^r�x�T�njD�
�q����F�Z� �zR�����Z�q}Ԕ��b�l�l�K�&O�p��Z)�#�R�� lƠ�bR-���~��\�g��U���=�1I��z�Q����\b*��V&�gQO�E�x�C�y̐�dF���V̓طꖮJե��]��]�Ac���J�`�<?��Z~��urE�`
�����D�9k�Wb�����4"�����$�5���{Q�d�����Yh1�3m��>s�=!sv�-�{om��J�A��xܳc�R70,�L{���M��^Vm�Ž��QS�T�V��G,����Q��,ߦ�`t�(9��|�4p*������SAL���LSs�ؿxUB�Cw,�a�q!�B�+|6��^��8`t�|6���z�[N��SrD`��Cz�R� F�5Rk��}�C�ę�$���9�4�e�Q9n,E��v��fi�n���>�؝��ܸ���kQ9I��6nդ)�l&a��	�ġA0��f?�u�����k9TUi"+��o�
��,��_`��>n
���*��a�|E�x��Eo���+�=�ec��(�k�& �f��'rЇDǡ޼2T��c�A$�Z�F^�'�$hp�y��+��`��Tx�M�_���:�� �6����12�b@�����QV��Q���5���Q�AP��0kX��\L��V��@=����ȓ|0��3F
��4?fO��������t9�������{��#�X�z�j{�m�<�#���C#M��|��seM�g����w��=�
B�yv��z����w߸��bz?^l�u:|,�7��v��=�g��p6Ns�#��B���Ӿ�c�w`���F����e ׎@�Ԓ���.�x>�-����L�[V�V&9n�6P<�{�j��8y�{G�D�rr�K�7��y�Cv<�	2�7�T��>PT�1i��f_�p|6&*Ol�G�RaW����j,h�g�����/oC�ǈ����'}�!}�G2p,8�{�\��{ 4	b qq��i)��܁k�l�*�����"�ryC�:/�l�o�v0+�4-�v��T����,�k=ْ7MD>���k��s2����uE�S-�~ґ8��������)ZZ��ͼݾ2���y�[����T��a
����y�kj}�6���_|�;�� U2ķh�v�\ʱ��&�nU�K�����j��� ��w�]Z~�M� 	�7܍�����H�C}]RS�ȫ?aZ*�������sw[�s+2O������[68��Y〒�.V*���f3��d%Ls��+�q3t�������jU�u���	���k�P���C�C�1?���N`X�{��r ���O_���0�����xa�����iԕ�������@l�M�J�Z��9��;��X�B�5�d,����z��Y�0^�1U��� ��=.E��*���r�	 2T���	�z�LO��1���`��֙<�<l��l��?�(�_��$w������rf��2׎�C4�e��j��;X��v��#�Lʞ�mʍH���2]VB�P�wO��a	Y۬_�����d!��av�/�$��唵�~�%����\sŊU:�21`�M��������阰�I�PS��B����� $h�gN�������F����L��m,�BSdVN��K�(�=+ x�/��
O��J3S����Iן	�;q�/����{�f��꘤�ƟWnY�����V��"��:�~;�X�oQJ��Q0%��T����x�J�	?$�l(��oy�!a�K�	II?ǥhp�d��;������t��w@�"^~~�VVt���}OQ�R�7��g��-�=3W�w�\��2��ስ�֛����`�۵�ם�w���ק�������o�@.��gt��$E]�6&��kަ�˳���AK�t�-�qH�T*7�d�d�%���l>��J�i^�1�(*�Û4$s�o���h��s��(��>���[M��o��-�=�i��7���oqa���1���\�Z�	��m���rA��֔m�q��؄�40��@��
�S\h�
��צl[���{c!���ɷ��Z�G��:��+��I�ǁ�Xh��I�?;��~"C���u� Idx���f��7�d���pb`Y���p�1�"��{����Ĝi#$8+Q9_��sI�D�)��BU��g8X-dZOoB.6��ʿZ���x?���;�����/�9�y����ʜ}5�U��j4v��qN��9+(�I�����Á����BQ�\bW����ԇ�v�\�v0~h���{m�d�M�tx�w�mH�0P�<2.U��T�X�WtY�qEahsb}bE�i+ :0ۜD|�ɓ��X��m�nL�՜|qo�g6��G����uiGV�WR��u����ҕ���u+�w��px���_CƟ=c�+|kW^���9�"quu��
������G�"Y��9�T��ф��=��&��4�Up��C��_gl�J*(����va�jQ@���L��N��]��X��2�IF�ԏ�!@,�{W�����;�V��k,��{u����[��2�����(��"�6Z���in3o^DX!m�<L*7]Z��t)��`q$8�|W$���RP_�D�����h*�eOUF�(Nhԋ<��KF��a�������,E��@##!8(\�����"Z�˘�����ZJξ٤C�����������F1�W�G��sm	���2N��rA��6$i���G~D���' Gz҃3�q�i��[��P�`��j�<�i�,�7g~�+�P��F�nz���m�Z<��J��t}�ʺ�)���D�C�h��)����e�*
	sË�Jh�+z��,F^�����G"C�9#�`�"�~ђi��j��?3mc����/�~C�?ޅ��]��_�1J{mG�܏^��yy���v�O���Xٱ�,���i���B�����I��Q���������ǿB�W�nv��.G5-����SN	P>���OGA%�A��C�	e~��Qv����G�M�#c��`�f6.�)�Q�U+��j&�9ϛ��`�NV_�����-�s�;8�Q��{N���q}���[���W]�-����u��4�,���Kҷ�����_h&����Q庛j�s�,���Hl��Rg���k*�¦��Q.��:Ne?�#1"����Ñ'A��T�LT��	3@D�(�$e�g�1a��O���`��"ǅ�n��"S�F"���Iɍk�z�=	����T/�U%�<��"�ta}S�����oj�*��"����žh�����pã�� �{�=���og���by���Ex�CJMaau��7 �P� C1�N���D��;�����V��L�4&ȴԻ�9��LV��b�>��5��aI^ͬU�Xx9G"Pt_� ɗ����w�6dG�e�B�.�*�@e��\Rq$�\�U��K 5�vng|b)�W��+����X�����_�<1��!�Mc����%e�z� ��W�}H�����s"� �ڄ{�aR�uGvV�p<D����%=V�=ZE-����:ٵ~z�k�
|O,A��M�@��?ϸ��2�W���{<J<yݤ~@q�+���g]ɻ���I�S�U�EQ#��S3���^YI�
��<�N��?V��?>5)��L��$c����'���=�u��7�� �(,�#�b�@E�n��4�k%�{�w�DKk�چ��V�7��1=	5�|y3q�0����� �z��є�w�c �H��]Rb�U������}:;H� bJ���J���gN%�do_�q��U��7�b����,��o��yҽ�!�W��2Y�����k��*�F�ڃ90���:/��ʤ�P�0�0�
<�=��.tyL���ѹrd;+˅��S2�f�W���KiU-)p�Fo�������ڼ����,����
��j���H�6�t&�7~^ ���e�F0�`�C�����P��*�ؕ{"�q�-O�~�&A'²���ۿ'��[�u�:	썉���i��m�h�A\v
�㰩t��s��S�Oy�6�
��`ʻd��pQi�RI),%>��!�6s퐌��`*4/r�މs׋�Ѱ<��7*b����[��]��/�[�{��<qX�Qw���3�\d`��?O�/��%4�g�2?n�����x��#	N�a�[� Z�?ތ@M}u.H���:��G�93��M^.�����z��Ņ�r�(������I�VV�`]���v���8�D����O��ƣ�����o�ӆ����UtѴ��o=˜��Q�VV�HV�uv�ٺ��݆�7S�-ǧ#��͢'�e-����s�7����'�i�Q���#vt���it�M~�[�i�ѻ�Ŗ�p�������>�w�3Z_ӌ��u�ff%delyx1�|�����&�ւ���QE�o�؇x�	:�/����>İ[p2f�M~&��v^����	jbE[zs���}���ɤ���ס�5%�����?��T�1���<������L1��dt'�f,3���u��������6��G�W���*OX;S�����?!�:�5�><�H�S�v���!�8��T�&>rX���~,N�{�]�_��!��:F�=������գ*�0�nC�wx��r8�A��1���X�Q9'�s�eC"X�1nۑ�NhD�P%��5<�Ē�Ax!&m�	�۽N����!�更F{Aܛ|-B���'D�IPyEil�&~5
ơȘU�WO¦܉k��,T�k�r��\)L��
4��
�!ƙ�u���3p���b5�}Cm�i�S8��np��݉C�]!��Ȩ�MW|O�ع�)��`�!��%ð;H�Dد7Pc��Uڇ#dӃ?��W;�s���uU�b��v����躁.�������љ��ox�Q���;�}���g�4QN���[mg�ۙ"L�ݝѫw()I�۵�l�y��댄��X\��v�������ƪgI	x�Xl͢P�	�����YGD�(�=�և�Y��'�|�^w�����z�utJ^n�k�e�R��g2e�i_��l�;�����ҝk��K!�+1������e���vN�F���nvz�.�"�o���q ?�s��S~�`F�q	J��L��M���Sɉ: 
�ċ]�?��Xw�49J쳦�>�놗�h'a��y��7L_��u4#i����b}�@���a䄘��f�b��j��Q�>��L���~�y�m���m�ЃKFuH>����Y��/j>'尧 )>ٮ#��}���; *S���1����,���&��Lb¾}m��	��u.�BX����|
9H�~P� ��k�5D[h���ch���I�y�L"�_��C^I`���P�E"x��M�b�� 
�D@aqxm0��K*/<D��9s���%Zh�	������Z�)%�w9)��6�8S5�}PcIe��:<�ɬ�4�s��	��%���(x:��JVx쳢��[�*~��[4M�ܞ�AClG��A��)&��f�����1?|@�A���uعu���5-N���Bj��t%Zz���o� ��t�Ξu���!yߞ<y"��DN�S�C.X'8HGA!�(�� ��QP�|ޯR��'�u���i�_�`926f\c�*�u�ܥR��t��p7�>=�.}7R����	ηk�oF��g���]]{�˕N����m���ڀg���JG�qB�gQ�M�BS�#ؤ;�o30yA�3=eu����X�: ��g3��d��<
F �����7r*��LD��>�n�����Y�|��ψ�Z�� �֣�9h��o��6��Z�����*$$�k�Z���KD��z����=&D����S����[�j=6��wG�o����aS�| h�S���7_��ck��w�6~���`'q	�nW{Q�oԀ���r¤��(?�<p����Խy�fE�LY�M�p4�7�1�x�o�n�R��t#�����<X鉲��;���y"�r��"'H�+��2h[���<e��B ����^�Y�4&(��d��^�颹a��23�B���"�zku��~����m[�S��wz��P{������۶H[����yG�޺Zu��P5k�~��U�
q3�N,c���­�0��)a��r�~�:�`P�%�%jg�2[[O|�If!]��8q���-R�m6�,�~F0C����������z��t6��8�O�d�_"¦�j:&d��T�cO:Hn��,)��߹&;���@ܖ�x2�x+�.��~����|X��O<[�Xs=!�V�Ĭ���M�`v�%�q�uBy%�j��-�tФ�-Ἐ&�Fο�f��C�\^�,qpy��QT�!ߖ�-�Ag�eN.w��S>�c��i ��FM9{��i'`=�A�Љ7��q\]8S�b vY�l��*7�nlnS\sB�%pu��L��	Xl��5��rcI���_�O�t�� D	"�&�0U�3U��(��_ Y�:&d�ʔ�)ќQܬ��Ѓ�2�?YTs¦p��qG5(F:p�O¦�����1�x�d��Yj��pŴ��h����\�&B��|ѩ��Iy�L��~E!���@XGP��<vr�虫-�[���O�$_�P���U5b��i�:dR�~�=S��,��ꨪm�(���MBB�C��+3=;��/R ���+
��F�5>����������=�߬S8��U�Chv���g�;�(_G��4KK������9S�[^8��L�󅻭���m�ֻvӀ����������X�o�C��!Ӏ�3ϖ��l[8ɚ7C0����Z,����۔ݟk�^�ĕ$n���	j�`��SS�Zg���Q8Z(�dU��3�}���|�Ɗ	hрJô��Τ����F�!+A��#��З|R�$��!�1���i�g]��ۢ�,���� q�*���m!H�-XE9^��_��@���u��9>s�F�0 ���?��F˝4=~(J�zy�bM�Jf�:p�j�Lա�X��	�5��-'�7]�+C(��L~�[�0�K�\?6?1Gawk���L֘X��nB��K�8N"u.:zm�<C�Tp��a���;&Em�gG�/��
��#�砱��ĳ��E�Ø��D[S�ɒxE=`>��6X�hFg��K�X�M�0��*���:5F)�f�Ef�5�B��b��"-������%�[_�s�Z�������zur8��3�:�o���y�>|���	K�5\��3�����b�Ѣ����a:��r�'t�E�#%#��P�>��5��{�L6���-K⒑�	��x�x?��z���.�I�m���\.�} ��s��߾�z�����@"�69���w"
�3"� 3C� �&1�wK�^=���ү�G�xW���[���xMpۚ�gC?)�	�m,���p��h��;@&�� �E�Ojt����	x���	�K?�E�%���{@�o1^�M��0f���"� ��Fcj�wL8ğ��z,���M�><o�g휚�ށS��(��(4U,��']��G��z~_�00�n�.�;KӨD*�
�TW��(�00q�A.����4�|EO6�K��a�6t[���'oG�C壢�*��bQ������H�����ezɃ(!�'Y���Eh��.)U���*��@�a�{�=�8x�.as��f��2aa9]y�)��g�2��/�Z�)s#�ڒx�6��tӊ��i�pb�:�4](���Xi�b��l/�Aw
�����O4�*ɼ��D&-S����%z��x!� ���S+��u<�i?*�6���>���*n@��%3������Z>�f��#:���Ҳ�ɩpӻ黃���KQ���֏����;��� ap��q�z_��&s����H����S���pu3o�W�����)��}JQ⤨�M۩������J8��J��P>� #�F=����Ud�f�d���辝����P���:�\B�(���y�(�7���V�|��cb�ř��v�5�+v�\��y�ֶ�� ���)�߂"9yyq�����0��E����=]��^1��H��#z��ц4�b4�_��i͓��^��5 ���T���?<����%&iD�[Ҟ����O�u�Bغ]���4j_�JQΏ��L4�h�}Yƾx�w���z�-\]V����V�bW��^~jq���L��ES��'����ȡ�$�w�4��]�����d���$M�$��vL��w*�ՁOs��e j��q��s�T�FB����^�kT��`�����b#����9{�I8`�Aa#gL�n�]��*ђO���Ь��������j}�?:8����x���{[�B;)y���Ĭ^ip�ۑlF�Û��s5-��=U�:�1��(a]�R+q8���Ln(4��3i��-��Z:4x��1  �������R��~��C���#�7��~�ltN&���1���&Aw�r�w�&�5M�����%DRɘ�8g��9�v�.�#�O�����@�2@����Zb�+ԙ%0�-1��V=6�D����G�'�:�%��4ދ��o,p�-����Z(��ٿ����* �ciC����L������$)O@�pH꛻Qx��B�Gȧ�ǻ0U'E�Qx7��/��C�}Q�'`U�NAp��
��P�U�iNg(tQ������]'�n}y�7�(�P "L?7L������u�6T�@[R�yQ���C���<ܬ:d�����鼣�~�����-���h=D/��^� �{'���m���=z-J�$zt����w-��3��s��>g��`�MC�6�}(�pDi�.%��I���u�(�g��%�� $R� ��Y5�BC'���][����e���������w+X�T��k�:p�������V����XEA�Q2�	8��X�T��iɞ�121����q���[�$�|��2h�b�\���>]M*y�x�<7p�Dj��Z���}�߫�2!φ�%1W����B{���<(ԫ���|��q�>�"7�~����W��� 5��ܠ�?�o��·�:���=��
��0��N1؎��������p�,lBكԶX�|�t�vǶ����T1"۳���|&L��a$�f����?gJ����pw��p!R.J�R��V,	�.����$����9�X1����
����Yn�me�BG�wTZ�R]ٳt��Y��3j3��1a���`af~��(Ҫ�2S�-w�A%L��LZlD��9H<9�Q+O,=�E��&�/Rřc	G)�eq,�=�M����o@Lۜ U1����G����Nv5��ұ�w�ƼEk��R"%TS/���^����M8C�Мy��P�N>hI���" T)�%��^����J=�/<��5��>�e�^���叜)��58jدH����nT\\1����쮛��U\ ��$�.3F.v�i�x��w����Z�3;ʹH���H�"հ+��^�-��Ou��B#Hd� X���༻=�5�*�>��z�'y�]� � �=���籏X�Җ�����/_'Q#h8?�y!I�mn� ��Fd�2Qb�'	������S����.�,Js1ߟ�k��HK�J�n��°�PaU��PG�\cr�"��'�:=����$o)C�-8L����ak�pS�J{�H׭���Nߔ͔Zt*�۝}?��KE�%M(�Oi� �_��x�9M˞C��3�t� W�%�у�C�Q����ښ���Y�J_�*���$�[CC1��]��;I������ګXW����O�ғ����R���̃6�\���"�ۘ0jk�-."�%��Ue�d N�	E)�?Hܷ�j���p�E�nί ƥP z�f��ږU�m��3T�	��L����J-G�dʡ3�K"�H�fRғ��8��R�̇��Hv\dih>xZz�T�w�Q������-��� P�&�k��|(C��(��滫*e�ؠ1U ٝ�0�]4����xW:0��$�X.7�8\2o�r�3rP����cS0���[]1:p�roҀE��#z��g+ߵ�z*S~z��UJ��et
�q�`$�z�?��J?�SAddᳮ��f��Cu����� }r*��M�"�cV~�m�v���/�Uq}cW����h`0;����w�d��K�q��'؎rկ�������f��Zͮ�����v�u�v�a�A��%`!W#��~='��N�G�A~GH�f��nV%y�(HV�H+f�W?}�{(�ǫ����wJ���z��7�A�� z��!��R�nD���%��Dj:�ʖ�+��(��k~���J>=�����Z,����e�Ϋ�~��ǡ�̒�q;&j�t�!���
�w�d��F�V�@�ͤ4]�g�"tN�h
ֻ�m�d�������{>�X�y���^x�w�ޢ���tsӭ��j�n�°҈\v��-+�c�w��!��~�hNv)��L����]XA�l�!�k�ʴ��|ZZL�CH����
�Ck���]�Ӣ\Xi�86��2�Ȕ���v��y-�+���+dm)[}C���Q�ɇ�\$
s�_��3�*��r4�֜@"o C���.�moX��T�Z[Ǳ�ԟ'�~���sm�#�_�������G���}�,j�?*����~�J�z��`g��q��b�m#��Q�D@�6�l.ݴ'	�$$��Zj�K��F�Z*	����^�{��E���mRjw��\߃�����}��!���"���'��;{R?�>h���y~��<��ވV�\E�\f�&�����u\{�v%��!��`3�Լ���͂����-��VV�֍��z$�--�k���g ���!���Ip��Qv� %y*st
a.��tXH�聨=����X��D�p9�3���`������P���a���~$�k��|�&��x9��IY0%�������=ɮrpv:�}�89�mM�v�J��o:@�w���Jh���������O��ΰ��o�Et��e7c_�Ƀ����ew�a��Q�O4�Wn1n�9�0 ��rz3�3��nF��2�I|�X]^�O����ǹ`��c�U��P,�)�h��"�`�j�@��'�h�(�g@-CI/�p��g#�^b�x���G᢫��3�7��� =5 ���2S9-8C�8����8B(���+.*+���g��A g�60q/���SP�Fx���+���7�u*�8_P��|�t{��Ǡ��� �3�x�ھ]��y�[��д���1ḵr��ӥ�έ��<����-ߙ�l����+ԗ���b������.}���>�⿳j��s�����y����.37�6���A�aW��ji�a�G�z�~���������/�r���%���
�mu	<�\�r�gq6u;AL}=Bs@}~���2rF;1[�4AG�T?+-�WGWi��.�5�6̶ �vo)����'�W����8������CΛ׍��N����J�\kJZ�*%�voڗ�'����.���;['�7����=��S���>.�^|uv��e_I(2���,�cv!����ӂ��E�"B ,	�^�Pv(%:�RQ�"��I��������l�/��0�H�F��6?X�M�jr�rXCR+�'b=�`I�����R��'$̂r3]��������Km����A�������&�$�I[Z��ek}"��i-�O����*��w�jt���1II�� ����j�W꬧^@�% �hG���b"S)T��<!%g|�4>i	јyQ���(b��a��Bľ��]Zm�+�p�E���׾�T-O8a�,�txʓDȲ�Zh@��������3���%׾����Ӷ��kCa�w�յm{�J'9�����T�R��عQᒝenH��]Нo��q�g������>b>L�������@����-m�G	ڸ*i!�(q����� ��)���w�F$0Q�"��(��r(xr����ҷ�Y�'��-���\X����vB������j��dV���L^�[v+�6��?q�e��];ſ���ݚb����)�T^u������$�w���doM�&�����	���@��ϣ��A`����4*%l@vs1	����u���n/��7�D8��	u�	R�C�>�E�6�/�����n@��m���X.b^�xv)l�i��jK��L	���Qk��Sڏ)�Y�sQe]�O�[��<���"�Z'B�C�		�r������B5����E���M�l�+u������쇐i�j�	��Q�.�H�CO�ҁ�g�.r�����H=��}����`"44K�,s�w��{�mݺ�k(�n�n�L�P��Yu��Vz��ſ��&�S߯�q˛�;�[۔R#D��B�1It\�ߦ:V~��b� !C% v�,1ĳ�N�-�~ o���Wl�_<�^���N�
sB��@x��Pf�)�<
���������5i[666FW�AA�2�a��u���\=�t&7�?ݯ9e�Ƞǐ�N�Ѳ`1G�S��mG��w��U��a;?~��eoǳ��6�^y�\�M�_���Q�z�K[�_��_�z8iʽߤ�|4�A~� y�W�~�H��&[��r�����~7�V��FO�(�h��'N\oL݂�o#tR�wm�������i'���� -��^�0Ap�{TA�u0�_�̤Ƨ��W�QԀ��:]���S��h��Ϸ��.Z�ْ��q "WR�%`��A�r�`���1�_��� Z�CXn�f!����8��=�8 X�0�`�U�SH	f.�'k�d��a�O���=iy�tEJg�}�� ܂gm8�<Ưbuά�N�'�j��:��K�s�E+��jG[^�t���1�끠�Vw�lz09�w�½�x�ޏއ��L�P��vd��X��!é�84j�e�7a[r���r�HSS��-��}�6�����&�0�ɧ�M��M�DgF6㓧t�(� j�x[�j-��{�Tc�"�8�k�V�ʓC��6?<̅�	�X��J�n���[���rY/Qm)<�&׳�F�4�����C��m=F�K����8��qz�v�d�Go
�l-*��V��lcy77+[�{˪���߬��ò�qx��������\��`�����|��~�:�
k�{[�������7n��Sv���W}ո0��9��:�9���\������t����G_[y�z�Q�IB*y9�T�p"z�d��c�zQ{�?��U��]E�,(,'Y�lG����a���܅�* ��}�a[KV���(�C�W>.�T�⧰�ض���F�q�C��5e�i��Cd����WË��,J��͟����[��Y[�����èg����X5�rw�^ �M}�gY_(�tQB0F���k��t��hY#�e��BӁmj�	�o���wg:_�G}_�`0{�G��*���}f۴rOK�&U����5kn[���/����v�m�?�D�u�Q���y%6*�l9Ox��S�r����O���E�{��)�X���tܦ.��tLY&z
��&�)
(�ng����A/��Nj�+���.c}�4;x�2��{0LqI�Ԋ�L���X�p�-���k�I��M�qj�/WU�M*�PYHs���"��y��L�x�:'�zsx��)��"b��������>��$��0��ga$Af�G��N���6���ܛ�U~Š�R���1�f��y@̕��:��_�����Giգ�W.d�]T ���.Q�~�����'h\"�X ��4<�㴷C9U�T�q�����<0��D`U�C�?(6tTqM�r��*{v�s�:���s��*]��gJp��9��XJ񘯃�\���]�(�m�Ɖ9a���󒔼O�kӷ;�j�Y�ܰ������1��5L��0���V3D~-�)	�=T���Z7}�����d��-
g��
��
Ј���=�*���4����By ��.M�J}���U�Dn!�K�q���z��!1�eY]�:�ބ���兽���s���D�ǠZv��v�y�,؄'{R�V�L��D�br��c�Tr=	-5�s**�����44�-�N��|N��4ls?�f������}8����* {��a���P�����*P5r0)��\��l��}��{�b����PT����Po�J��i����ٯ��_�7�ř��Q�l�{xh�z�U�{���-���8"7`���f��~}���`"����nm��a ��q���I����]֧�+�G(�{�vӌ�w��[vi�[[vv(��3x~4�]6��e�πdm�r�W�,�8}r��u��4��¾�d�G�:���fE:�-Vu���8���~�]��g$kC}o#�������}�V�1��|��fWM5'G<p�g٩V��||���&VZn���Wx�[}�N[F(��.7�Z��8������L+K�D���m������8\��u�4�y�$�(���������ݍ��"t�'_��6��B��S�[t��I��,�߮�U��XqŁF��H�c�K�6�I��Z�\��î�U���b8~~r�9J��Ap��ᇢ|�6)���xW�;�;uR(��.ʦBC�GhBG�KR/������as�-:�7Q�@��N�=�����V��Ͱµ񊵸�8�j�j�{(>7�<��!=���^C%�#,���*���֒M|�a��[������⯉�����0ө�N�dȶЀK�]�5��+�P�qZ��x? }����{��T~7ǈ�
<�F=꟎�7_�{UT��2s�Q��>$@d��h�@�T/+�P���Xn�� (ʠ j:gX��E�Aқ
�+��!e�e�;g��$ۡ�u�ˣi�g2��|s�S��'q��Bzt��~��q؞�G��9�v�<kǃ�^���7�6�"�7)Xղr��9�R]}���s�{�0o�����.q����@Mj`�Υ���I����K���o�/7�]�nG�g�30, �b��ܫ3?x@�Z~�Qp�w��J��]�-�8v5/e��>����t>�������f���s�H�s�XH���%b/���(�T��PHQ����ɸI�K�����5��<Vû���ۈ��73��0O�ހ׽�T�ޤ� ��)��X�����E�4������������~Ĩ=��1�gWif�v��v&gv��U�Pٖ2!�]��sߋ:��g~�Ɛ�~.2�H�w�I���r���|���L͑<~��W���=��/�@܁�|�J$�K�t���453��-\�s4�~tM���(F�F�2�tU,�M����)/��#N���BLt��u�8L��*Z���q̩����J)�P�q_�dg��\���REn�_�*u�!��uX��w�ҁ�?�aGBɠM�����9 ]����u�7jx� )k@���h"�i��6�w�/�y4��RM]��N�f�F���GO�x��a�bYǜx^ϵu�/�Q�%��nV���Mʔ�M���v�FbW\�b���s�����lis��ALԜ�PJQ�~hduS��@���t��l���*��Y�ֲlZ���/��?0��_*g�땤od��4�!�1B ���!�VL���L�==���/�$D����ů�yp�۬�s"(~���خ�D�Q�R����|�{!��  ����>ˢ`[�Uٷ�9���_�$���Yb�����N�$�-�^5u'��_�I���<�|��~���
�F��ع��.y<)��?��Z5z,|��x���t�^�pK]5%
J����=��Ml/g*Ù儯��/����l5M==�Mu}u?~[
��o�`m]<�E<>Xn�B�-C�Ls�����告�7$zZ�9Z
��؂G[�M�|��Y1�3k�"	Fg���w5X6�'k�Æ�� ������t��'ꓹ�A73����`t��`&�d�d�l-�`
����My�eY@���S�HW�~*z���tP���3(0J��[VQ�cX��!J0K����Vm$��z,q�qX�ǰ4��b���
L;���uZκ�IZT��@L�N׸D %&�K�\>qλQ�O}�ϓ)q�-�S@��l�[,x-H����p�C��'k���ף��`�dc��V_ZO��Z��W$c�8_@��>m���{eAkc>rX1��Mѡ�����a�:8��$-+�mGW.D0�.4�5�7j��Eawr��]i���R��Ci}=߬1��ʠ��T+܇H@հ�xz����f�z(L�,V�6��:4�Zގ+�G {H���t�Ƀ�؇�D_[����}�?)	e�j"�#�9�2��
"Qq�q_���^��[���"�Kf�i*.�.�/�/��F��y��A��w!|�r��4���ɑ�D)a�V8*ww�!�\D�9��F3o��1w^�d�-k!�oS�0@������'�w96?��Ňc�j���iMJ�����~�Ǻ�-a��e}��M���h���H�C�U��e>�Ԙo����ppJ��Я��zG�߯�@G�贩���j ;S�H=e��r��_�+֔-b:��q��k?��^å�\��T������=��gf�/�
�2"�_=���G0ԃ�+�n����K3���R?s�${�l�Ai5�أ<�@
]��y׽�4�z�e��~����a��(`5g�)f�������-{4D^Cm䶣��qF�@�$�Lw�`8��N�Ƞ�1��@��6�\:���ĵI�,�5������B�mf����G�1z����ў�'ysM��?�-�N�]BH!��P/9�ݗ9�`n�1�)AvN$����������t<Jh��o 4A�uM~-U��E��V��S>V.VO,s7�n9n�Jv:�ġOw���\��մc�>B\������K� ���@��`,��1�)� �S!=n��ɳ��mnN!�#�#��0���0#�qpp����֦mP�S�<�C�R����'��uc
�.(�;T~��?�hotp_�
cb�P����-��y��u7��~u��f���v�W�}�Y`�R���W���Q�K��J�Ã�K?�NH���|��>�Z�^m�p1�����n�$\a4��TL��c�ܤ���:	I�*H2��Q(�}J|�� �<I���m�y��xҴ ��Բ�篞Q���N��"B���6Q<�s�˭�!���q�9�����Ի��&�f��g.�����F��_0���^��I\�ջ�}��J�i�����{��o�v<*$l��T�aj��d�~xE"��M£v�_��mFʥb������Y�C4���
�ۚ�}����;�|����B�@*v<�q|�gfq �K�e�4��+�1H��_���8��!q�>D�������B�m��x?�I~̂����6<�V��-s(U8.��* �ŝrO\4zx��bۋ��4�1�Pͺ7ٽk|C�3�tt���f)��8������|�S�kih�QkV�ePqP>�>k�
�x����E�"K�����h�2m.�k_�^�.[.u@a��� �7���#F?|�ܫa'��;ۯ�Z���[��@� �M�C�R��y~��]�����\�D$�n�ы�&r��s�KW��@*i�Y��6�.b��_Sw� ֶ�a�M���(�������["U��s|m��ڧ8[�P��8���x��=蓢 ���h�I�/XA�&_mT��eT{�0>G�z�Y��8�Jk��70,����F��G.��H�����52j}���������]�OT�BƱu����*��&#�-����
�zr�ҝ���j.`Y���1{�e&T�����<�&��E�S|��ī!��q�[�G0�tl6&.����/���+��d
�h)��#A(��!��A�|b��ZFzʵ��b��`�9`���T}��>���V#��Y���&���m��؈��k14�	R>�|D5U6ͨW�֊C5���]�Q#z�b�~��P�{��'🀺�+$�l ,=;��,�^j���Y�������o�毓��J��np��ⵤ�~��{2�\�����eh�r�W[���W����Y@�Z�3���'�-��= ��W��yf&�]#3�F�`a_'/&����� �0Gɀ.Qa��>�?¼�E �q�bq��⠳1���L�Љ��\M����rW*�9�QE�aP4� (k/=�ӏ�<���̼���c���]H��'�
�2��2r�������F��4��ftqW?:�u7�[�pTF�Zw��Ҳ���U�U%>	�iK����^��M����:ɠ��������U᠇ޠǱ�Ǔ$+�w�_��t>f�D�ݟ_�z�z�|x8@
�=���p���|����?�>;�e��_b���G�)C�as�m�"���dҭ[����������p��1��|D�hRH1g��)-����Ds�m���`(cmO�&�8����c��)�%d\%;],pkc�#�u�'�!j4σ�LJ�̓-	Z��H!��t����a��4$0!~6�H<�&?���m� ���;g�A� (k�p7_�f8�\�JCuq��%��L�M��N�x��T��fÑ:<��-�#�y�9��Z�8]�U���E�J,���c��k�|K_Q�o�vƩ�D�4BI���_���5Y����D3k�9 _��ȏ��#��ϊ\y�o�%����2�&���I�XN�ߛT�_���-&�BN���.HoZo0>Q�Q�LeT�{���QWU�K)+�2�r��K��5���WT���+�>}F�^�'3vi�Vk�r�)���,�t6�<O=��IN"�j�����]�ϑ�_�IR�2&��m��ը���$@R�����lz�e_�d��p��K��G�F.P�J|�����[|��4��L�ǩW�����SI��}ٙ��G������܅%�f��
���	�����%r�l�����$}��Z�Mx�lt��dt�J����J���V��1�p�Wu^� 	/HE�'<�e�޸��~��c'�**���'�>`�����]jm5]����T�h��LuK!��p���\M��,U�S҇,���Qs���"h�����n����1�����Z�^S{�ֿ�}�t 2�$7WO�@a���7�p��=g2�
�ɚvc����wO総��@m�T���׎��ur�u̎��er�f0ʴ�u`͌rj�j1�>�Z��,�:x�,�ˉ\�	L?���v*F6���R�W��X�A����h�3�Ø��;��Y�z�An���Wi�ր`j�I�K�RQ�'������}�ѳ�������jg�}j�� x.ɛ��g����_]���C���6�G��E��`��?����܄A[����ҪVӎynې�:�
s\ ����O��/�2u�^�x��{_㷅���)J��L~~^~�ݥS��'��Ш���{˹�I9@ɤQG��x�{���#p�<��\���Hi.�zJ�uM�ƽg/�2lZ0US@eH�|ž��`���њ{6�xS1����ʀ��������܎�8��=#����_A�eH��]�i+��ſ��T�����lx?t�����w��G.��;�>��)����>��}_O޼nr�o�`c"3]�+���V�5���P8����J>�\A�c�A־	*Q��1����]>��C�uQ�)������T����׹��gz����N�Y�o�a����!�4�R�H*Wȯc6��'>�S'��9�$�Ӹ���g�J-=��TI�E��B �!��2���e���<Â�Bܳ���t�!PO�])�c8�����ёJ"r��:�:ag�	�j�Mן@wWK�O���_��;��oq�^��O�a���&�涩�&jY��ｭ�`$����I$s#��=�	AŌ�DOc�a���!Q&0�on���Y�-������Q�	rJpfQн����#$`T�7���͂@8N�������)S�[���L� ~r>�����3�@,;�[Q�79A
R]ed��\~��C�qA�_�A ��p(���r�-0�<�
����e�,��Ua��������K��bG��y����uU��2/��|����`�[en�o-,��a\�f�[Am�M^�������Jڠc{�X�4��f��G����@FRkGz���9&\m�
���7��6��� ���A�0��}{"�8_�Þ[��U����	��I�m b������4�F�]>�笽����~�W��թ 4�8�E�c������0npou�#Ò���V����LZ� =�������=����m�=]p:���	[8����_�p\(�r*�\���J]�U������N۠h䨃��tU٪r�-*_ՙ&��F[\C���G�p�Z̲��2~�WWc�0m�2T�?�eA��E��vy�HbD�'�`��cז����Bʵ��� ��X^�w�����J���B�Ӭ���m 0�����Z����)��;,�J�I��I\��8���\�B�4��2��TV��Q�����-IL���祝�~�5`gt^Tԋ��ȘS,Y��s�D���P@D��0T�p�$�z���:R�+t�]��H�i�]�v�8\�v�0��ߌ��?�R�Z3*�v��.B!?< �M����8"L�cH0������ݽ1vyp��X�&�.ܠ�]�A�_O�gr͎�a9�j��SH5�
O�����������a���A�\�b�~��z� ���7�ՇS���͋݇�WU�ǯ]:ê�n��ޚ=�6�ݎܜ�ح�|���z��_��e>^���o�t���^��:ޤo���i8])�Y�������x�%�jO+Oߘ�"/CU��?�x���y�ԘY�d+��7��D]�Ѐ�)�N�"!%BEA��)��i��>�N'�����W~���Z�R��6�h�<u�yt�z���lʰ(�Ti���zy�g���A[���a�u��%�!��u$'�Ҁ?�7�|�h��/M����P�]U�ݠL�Ae���Wg��S�jЫ<���pJ�J�I��{�/Ơ}�V�M�1Gd���'����B���ӧ��㞍�8�(��W��㎝Vk�ت!T$[Ĕ'�:N�u�E	D\cȬ���c�� ��7j���qi%A�[$�X��
:5-	����[���
o#�"���,{�њ���p��م����?��Ҙ��H�k�Ĩ����i<�=��8<�LȖ@H���in�2�z�ճ�,(�z	�q_ ��[�i14ҖDî;�J��j���Cd��8�f	R�-z�A~{,�mO��GI�z�s�E��\��f��t��~����ow�q�:u�n촀Շ��n��<���@UD�s����ܨ%$�U�E�qBf���[��$��1���cڌ'��X�jg��9������ĩ�^���ZE�����O�|��Б�i���8:��6c�kY���\��=���GG��B��x��v}T��՟���wH�X1�v	Ow�˸�4�0�Y�g�n*A�/W�ŭ��l�>������¾/#k�Sh7�i�-���-�Ve���B�L�o� �X��v���n���s���/�:,�E[rD��om�m������E��R�E#ƣ�j���[��u\��m�����ł��M��yqf������׳ܦ�Ͷ�tĮ�"��,H�,������z��]�H�HM�\�ȪT�*�(*ǉʕv�T���a}s?eh,VaX$�?�3t`J=7���voJ>M��J��� ��6q�� N��9��&G�(1�A_p�;�*Q�,d�� m��f����ʔO��ޤ\���Y'V�����MY�1�Q��l��6GLZ�E�喬 (>�.�i��V�E��9U�Š-�*
4�I'���y�
��@�+��(ʓD_l��DA�>�T�?����B[Fen�,���^Z�u��^��$�_��N�X98iv����|�@�Z��|�W���ɥ���`�4Dh�H��ɲ�1�?�?g+��χC7������t]�s��%>؟�F��vܵ���L)���>=^^z�^���8-��?b���x�{>����_n�ғi���d����?M��W�;.�n�G��1�Z�S������TW���h�g��)��o��d��0":�}�� �I8ƭ�/Ʉ�\�E����)���|�-"�ޯ-?|m�j'!��J<�Lb�5 ����'峝��u��zC�YJ�׬�ZCU�cb�ͧ ę��l�F���f9����]J||���ra}w�:]�i{N`�h�>Y1����샜Cu�h��"s��~��9�n�N�@5ؗ��m��yѼK�Ŋ��JϢ�����u�vJ[h�#o}k�q� �N���.�KI�
�|�Y\�67
7D�g5�Ss�`%!�ÖS`�{Vzq��T��#�.+��Q�C��'ߌ5_��xŬ:����7�׃��U�;���_?��{v�zm��n��<���Tt9�����$e�RIY!"�nz� �����&	���| ��.f����3]~�T��8r[��q�4@�A��`��@�Eû��l�;�(�إUeU�r���tZ#g�v�gԗ�z��9"���� au��<x���j簙�XE�+TF�w� ��z���/X���l���/�?z�"�`-B�o�b�'�z	�H7��
��#7'�@Hm� Z��0ўꟁ��3��/�xLS�����EHBd�<.��[DH�1�kQC�i�9V�Ӹ�T�:��>��R������0��]�����]�aX�Hk_�5�H�v��U�)��9�!)}��eW,\q���C^���v�l�
����]�P�_��<�S�����#{A'�<�N�Ͱ����~��U�I{\�Ǚܰ�hX��8�Y�Q}٦��ʍ8��:�j�F��ɷR���I��u�+p�uM�#��v��~Ze����pp�3s��b�@�C}��2~e1:�m�N ���_���|2��0��#`XxOC� 抁�'��5�@T�Ro�9yU��Y!��T�~��r>��@ei�]�.�^�`���@����"���N��mڻ''h���ayk��J���?�V�/D�e�s�z-��Ñ��t��l0�*+�U�8�V�'V|���}��]�;��.��ϸ�0*Y�ç����d9L�SmG�� ���8��H�|
e��\S��tt@rrbߠ�?oG(8�oCY>��TR*������	�6��z���4Km"����$+�('헶�����J����Ukp��b�&��v�H�yzM��P��`p�"��=��
|��;"�|���?D"�~n�٦���ʯǍ������܀�?G�v+���|N�I�/*Mt�� ��3{n��ȶ�w��`l�kt� ������u�6��0�5��M�Q�oBI9��������&��?�]u����=�6�@�����Ws�[���Y�x.�`)������?-�?S����<ݱ��]:@J)���{�ȳ��g�a��Y@S���RȮ���g<�l7RcB*�� �9���=�J��QQ��A�I�xk1y�� ��O�g�[��.�O�V�r2�\��=�@{aN	�X
����8¸X�84K�قBYsj*b2:j:��χ^�32��{��_;]#S��cYga�MP�Lrm�)Ӳ׉��F��5��P�܃f=�� ��Z�7A�H���CW��v�2��
T��h�@� �,`��U�Ҽ�g���A�\$������w2�z��,�@�I�Dc�L퀙��bJD�i� J�*�	��'�	����;ZZ�oZ;#i���	�a�ON	v��Y��+��&�l����M_�~����f�U�/�n�}���j"^ȄR��ǥ�=�ٿ�ys`�R���̚8�SA������uvv
��d�}�4��rc�7��^���nT�֌���6j�B��G�y�oŒ�\-n�"l킗g��4O�F'��3w��n?���M��
��L�)b�+;��-'a��ߖUV��14��%�8������6<�Vz���,Opl�8�ӛ*)VZޛeU��$cJV$�3�8GPn��(V8t�/�_0�Pd]!�;��m�_bH�"��x�7*��쳳/}����dW��	]��(98U��&�&҄�i�c��u�zܢ�(��Ր`U�#�Û^�|Z�B�	4�uP�*~�jEl�m�`]�w����}P�Ϳ�꾇<��PPta[�7���B;��Y��F�8��"K���BD��]�Y�{h7�T&�Fw���w��{��u�_}��*�3�ͦ����J�lv�Q��%sz;jSǕ֟m^zuF�nq�n���
=����,��g�����C]��$�Q��2kd��`���Y*�V��Ɯ�Fm���� %�滛;�&��~s�h�S����|z����յ�),5��Sn�h����G�e��;b���]\���iK��V1�S�Q�Ybz�ߴ��>���*y��I�\̃u�jX��{Uj��j���W:>�L�c��k��Et�t�)Zů����0���m\�����vt?�I��U����{���SC->���Je�m�s�'$~e�y���"[=�.�4X+�N4އpc�`�L�f��/
��MCn�n�k�5���<������X�x_��ks��放T�ړHfحtɻz�.�sƺTZ�0B�89֖�\�6����WBi����A\Q���UX�o+A��e���D���ӈ/m�g\���05DAaq�X^��%��=�+Z&�+��,�T�o� F8�dP�h��lr�*�>f�����:�r*�I[�G��`�ܷ��ܦ��̂���]`%�a��d��m���L���2�l�9g���5-A�S��'.g�\����;�{�:�������g���o�u>n��/~�<�_��e�/���ᐧS���a�gQ������r�ƣ����;����sf�e�����%痯���G�ա��U�je�h��q�i�Fa�o�c%=�"yi���^��۟�Ĉ��b�$|�6��[��N�+�j�E��������0�]q
�������{�&��xI�a�Jc��b��6�~�|%;Ż.�� �Ϧ5�6c�`���(ɝ����ܻ-6�L,�|)��������nq:��Qf������8��k7.O����Գ���{�c8g����Q§�f��1�6^{:�����HH?E���}�2�vW�}&b���+O�ɬ��.��1�%�Q������{��Ȩ>��Q$�ǻ@}v�p
 �����2���h�갦�7ꑒ�5�����F����J+�5��� !5:$G
*|_�����u���k�|�9����9����tdt$�dTT$d/�4-^���1���
��CB')?��S�t�W<��y��7R�q�H"m���r|5S�֠y�5#��4R�nW�Zl'ZSV Vq��VA]5O訒w_�ε������!޳0���Ғ��1B�WP'��W{T��^�n���������y&�kE�R�=H����!�g�o�������AR���HW�4�6Z:��$�����MiT�WDp>�;p}�f
�B �OǦz/�-�����D��jz[����+Ǜ���P|��ւѨ�ʃ�x׺��ƀo�Q��/Q-��֛Gf����S����{��LG[ٱ&H�������G�!p;F"�4�����B�y
����ܹ���h��rԠ~�:�����ܣ��Xx$�ǒ��Hτ���PE1�M˧$_X3��*˞�/����kg���Z�땆����׊���,첒��
݂�1@�R���d�g/ �tR"Y�5�M�~[_h���%���hA4Q*�㼘C���އZ��N.�)� I�$j������j������ �.�<�ϱQ�+L_d����Ǣ2���+NFMɼ- �]����v�����{��,u����������?2�n
��1I�p���s�(<WRT$<��?GI�ӲCP��q/�>v�ߴ�����ڬ��w9�+�z��xֺW��j����� �``�1�X��e[�5��9lF�y+��T��G�AN���|ۃ4����tZ��v�}���[n6�:OdRM��d�$����+[�O�>��IX� ,��mt~���9�d/fw��"\i���y���W⽍��� ���|�*���	�z�tT��p��;D&mp�)�!͗&��,����H�&Sv�S�o5�I)>h�M�C~"��[�f%l��m���>��c���4�LP�LmA��+�ӓT�c#�;����@�Gb*���ߔ�C�oؼA����2�&<� U�s���@9¶��G��'&��u[����'Ǫ,�PHm�,|�?9k��kG= �CmUR�D�������蘄�O��8�����m7s���L�_�^��O8����:nB߽L�Y4l����!��� �<�M�ܯq���຺��j�w��|����5�%�����Ư��3��EQS�=ϙ���f�_Y����w��k��w��ݜ|�|��3��4_���t�!/x g�1��c�닓�Jv�w���J���_�B>���m�F�Ds�>�:�,Ta�+�R��2B��{����i?��=j�p߿�j��(�0�觸�����1"����	��.}W��x��|������\��cKE�a�5^�*�(wKf[�4T]jD�r&4#^RFJJ�-�tC֪ўҔ��_,�$�1�Z6[L��&�?��֊�%He�����E5UgiM����?�X��!Y��qV�&6���}��,�T0x)f���PO�1�k�o�Yc1����ʃɗ���$�䣸�!��12$l�)����j`9k}c}~6fv&N�q�����y�Ckщ\���b���:���s�֫��x&��%{o'J0����K���ˍ��ev'=u��<��ߍ�	���4�~ַ�@1"�J�z��i�Nw����Ft͛��<@�Q�0xg�ܱ��aT9���I��	As6q)��n���+W!��?�M�{9h�h�4���r[B��'0jk�ɿFc<�j����{���wI�J tE�d� ��f*��0��� ~J�����&^���d�C�T*/\�&��!C����TW�[S���̶�K��;�6�X��k�Bgٝ�>���K��q?)J����Z�9�:r2jS��_
�y���hr_M����3Ou���T��6k��U�>rɲ2��اR�̞���t�Qͱg �B��TH�C�2B�=$1��"a��V������h���6�h`��{�3�_�C�)�]aK�s�[p���=h�T�
��R�Y�ǁǣQ87{��ļ�y���Q�x��F��b��6�?�/V�����n�0��������3����\"�ګυ8�w��X7�e�3߲�%�j�����Y�zB���z�᝵]�_E4���{��HĴ���"�\�`>������l*e�����)m�x���ʸ�[S�����>Qpû�]� �:�ؼ���HO<��?���8�폒C���W-����r6S����D*�J(��D� 0�t�%�7�vc[��/��nFC��;KcH4�����B�th8.h�T��PG�����ڏ��Z@��x���SD�?u�l=-lxR�Z��?O��,y���:W/��lዱG��?��V���#�N�5�_���S��ڴ1x��gD i>�낙� }q�Z���/�N4O�E����z�����:^�9Q�c>l̛HV@LK�0�3<:2<�VQQ)b��`�`��f���m6��=c��bCW!*��G�a���(�w)��ʯ3�RP�������e������q��5F��_%�\�૛�f��~geTu}���gz}�}��_�}{ߍ���ֿS�ϗ��}"]?��������zȚ�'�ar>��K��ZD�[���ܢ��d��w�v�Ccrl`SO��qaز�!�Xd�T�]����� ��)��7"JOл��/������=���������V�����k�S��E�n�����7������c��J�8�vJ|A�qs�J�U�]�ks��p_+T�ߠ�~���iXaYX3W>��Sr��%&���#���[kT�#�e;59@�#4�|{p
�ꘟH���y/U�6�S�V�	��Ǆe;�2�?K������&<[J(��F:���)�6��0朆q�"en�/�&���y�������Ν���q���Z�ۂ�� �^�����Q�l��^EDjx��^2���)b�D�s��7��\�=�)W���f�x߉��#�z�K���&}e��m�V�:>1_8�F?VY���.����.e�~_h�����F�\�� ���������Yd�hV��y�J��k�K�,�}�R�M�̧Nm�k����>"��i��V���+|v�b`�+C��{;��Կ�~���)�V�TR�|�|��<C���ܩ����P2]7��sv����ób�_%�QD82˿�S����'}sީK��P����/�� 5�������=|��&R��.4����Z��IF�c[d="+��f2�s�ٰLI�쿡}ܞ.p�
�-$��&=��R`�6�n5Fqawg��a��G\���`�rb<�P��Vқ�+[����ΠD����c7~{s����<��������I�{�����獧����� �P�!�b˵\d`���+�G9b����Mac��,e��r��D"�����F1�(:	V"U�[���?/(�6�&i�J�/ ��"u��\��n���Ο��F��-s���}��~��-g���I,��w�<��|˾��nN�<
T���c�Ep��w]��fo�ZjFŧ�rp]v*"�)a�� ��[ۤ�R�dF�G��/L�b�5eL4���s��~�uf��H����)�; \�|�4�"c �	�E���W��$k���9�0	
�!�e�_�6��"�c��`�~!�]X�� 넗GE��d�A�:Ӳ�E��rC
�jY�٤P�n]�����[�}$�E&t�I� �RΆ+�#J�-�ְ{������ ������Iwe�'�����-G���<EA��	}�J��%�s�Ǧ��W�+��W�fYr�z3`�-�[L���2�#�TTddT/F���! f撡�/��DYX�Ĩ�,��d���������/� ێ�~�l�xC��!�v�zwC�^G]������hmN�ٷ�����j���?Z�\�n���?�L�r�}��7���t��{V���Y���ߟ�kL�93
���f7KH�ĪՆ����Q]�VO�6ͧx
j	A��������Q�Gh.MM"��)���p~���>1h}=@��CB�v��OI_���D�-sȒ{j�j����fvA���0t.�ꯏ:�D���-2z�pl*&�����ƽ���֚=U߫um�S�,e%����sK�_�����ԥ�QHLll1:��%�|Q7O���>X�������a)2�Sko~1TQ�BH�`��r�����2�0GO��b����ld��Bs����Y]�#��q@-)(�ߎ��p�kuJ�ri�jRu!���C�LO�ϯ���850�V�]v+��Ϫ�r�`�,ѶN�F�*�/I��&?��.�Iu^��¢֌i���Jv��j�9X��|�~�vքw�65!�����6:�*�&6�_�`���5;���4w�N�oM��?���gC�o�	��$��d!W:��I/��?�!�<��5����}6�-*ON�fѝi��E& ����B.�s1�����x���y��տ.g�q��E�O����T��Qk;<{�b[�Z�k^&��5UA� �_Z�~���/?�����}JE(��N�g���m� ��>�}�41�g��ѱt�|ԛ��A�0���rҳf�ي�ܷ�|[��c����2Сya�#�+l��RjrL@��=�yQ�=N���	�2�,���T�`�O!�ۛ�m|U�>M�Z�Tw��Ps��[3�P��Dݚ?�=l�f+�}��͉�Q0:?�y 1`��|Ԃ*lGq{Ic��2��4���/Jf`�~d���y}aC�/�,:ϔ�k�L�40���z��=�T�'F�-: 2L�{Gμ2B<(�<�	�/
�[�yѳf�(U�f��&�]&�N���b_䂷0�B��AY����.D�ڹ6�c%�k�'�	;�4����Tq�NN�B�mKw2���Z���4{��C�49zN�5`�j�z^��!�~m�W("���Z}Β!���>?�(�y�3z~����D޵�h���*�Ta$;�nxj�lL�A���I���.�C��:�˂t��N4�����}le��Q���	q��Fٔ#��J��� �/�'�w�q.u�}�U��(�J�[��x�i���ٲ�!/,�)i�!k^c]�1��4 ��1�t*]x��8�w+\���jF]��F@s" W�C��f�)��[=����"�K�l�L;ϔ� �=�?�%~�i����!����O;@J��'Զ�+�>DA�k�.=��7��t��O�ߡ�NV6�,�I5�-Ւ�e&M����rĎ��?��K��Tb���xe��X����������������B?�rX��s�.s���˽�L:q�R���H�TM�Y�����0Lnۼu�k?������j�t�n濣�J������[�+��s�����'���)ʖ��B{dd�M#%/��W��l�Z����6�4�xY�����*��0HѰ�Ԑ}un��	!LՔx����9�ka&�'
?ϣܷYԩwp�7h�x��m�����<�z��kt����T2��	?%<ܮ���������w���	�Z}gB/a��x
����.d#U�``�߬�ѿ� ���c`�9�Ԁ���T�u7t�1�W�(W�ݛ�F�o*8 ��#.}&�Ψ��{�V�l�:uzl[��w�����#���
3.U��,%^9�l�|YĢmo�y�B%Fq�ܿ�o�S�y3�_¸1�����G>�c��j~��@U+J'�b=[D�R`�L)&�����'�i�jS=ٺ|(k�a �tN�f^�ȫ���׵�-�I,�t�fh�a/�ZJ�)��"Gk�>�T��o�C%��ɘ\jXy�Ǘ}^�ׯe�p��˃�`{2�h!�歝��W��aW���2�sR���Ⱦ)��G���Kg�_D4����"�&%V
������a7W�?�J@����\�,�`9�����QF�#.w�����?��p2ۺ��4ځ%b�?|���D#:ݛQ֢��ڽ�+m�c%��{X�j�7Χ�=,����Y�t�!K4��X�B���S�7bE�(����>+����3,�9L{B�~M@A�'�	���
F�P��X�Yi�Ք�T<�;d[��3��3���?���Q\Cי�M֌b�`�7��OG���B��!`���7.=�;ㅪ�Ҵ5Ċ�%`۝�b�_����{������KC*B�[��7t]�b~�ډ����w����>>�q#6�+;y�l�6��Ȓ/0���K�u=?�fb]E���bG �	�Y�R!'2�-��Ѿh�5�����{g�J�h3_aj!�ԟ̈́Y���l�� ɠ�����f7����I���b��3	A�T�-��ZJ�k��o��6[��ֲڵ-C#3S��]�r֌���(�\(���zRyNU�eJ�qE������f[��G����5.�K�$2{�S�S���D��D�)�@E�f�i"�/�<1��܊\xz���E��$�,s\,s����*�܇���z�˯��I�5�kEn%��mE޹Q�拰�WٗGa���&�[�
T������}�	 ����$��@�j�h�f�L�i��h���P��i<:�v�����\��!��K?I��<!W�p�����f�?�[�%U��	;������E�WOm���o�ɥ|T�y��.�u�LQ������1ֱ�O.@X*F� ��L�'�C��~��~�S���F<Ւ�)X��r#n;::VVV���Q�MF�ٶ5�[�X�2�k6Z>�dL�����cD�Z��M4s+看��u���VL�P����ݽ|��$�d�7�S;v�3[LX���
وqȚh,)�~�܏��3� �4qɜKsj��Rn�!�E��s�Qy���)�9��փ�e�6� ZB��@[�i�{�	����M%�_�H�,�0�ށ-�W%�
EV��Y*l�ݳ��2���t�T��Ts<>�ߔ\��7;'o5�<� W��Gd3��ng�(4�+���ڎ%�
֫HBFC�di�6�J5�[��|n��vjp0)h7��������)�P�|���$�Y��х�k��V���?�8�L���7!Y�<�ø�������p��0`��m�M�-o��Q�X5��^!)/�吿<�76�L0HqM�=��[#%0ʑ���kޫ�@�2Tz�D�F��
����3β�Qn^�]�.��z��C�����ֻ��V	�c+i����u����!����ݜ�̦��֮�,��q�9^��l�ܼ4�3ͺ/ ���@G�^���Y��B��M�!�2�E����!9E�I�tD� �@7GtQ�A������S�,�O��L[�{\��ܶ��W$
��	�_���J�G�4�?@Gxt>�!�4�k=�VC	�;<��Hci����kV���	���,2N���ge*�[����f�6��*�뀲��IE�C T�UA�>¢7�%�NIcowב�M�����qb(,���?}�Ga���ч��R��&�H>s�	�*��cN�ʔ\�'����-����;�b'����x"�\^�cml|�|D�`�C_��-]չ��S�A/"э�LS�g��ͷ�`$�!�r �#��\�? � q�v4���� �!L���������T(�JY��JS�'S�Mȉ�J͹��{y+D�����)�	��a釧v��wH��>B3N��2.�p�d�>)d1L�ĖEC�X1����FBD	���Л:��Nm�!Bݣ��hڿ�N�my���f^�vrє/�B�;��
�I��ZY��RR������Ō�
 ���ø��*�U��x�C�1t���!H�R�#���02g�Q�Gz�n\}	�/|.P�Y�K7��ϙ�<�}�:�M��_P���%7uX)Fܢ�CCө��S�����T$hY�И݌0IΠ֭���ڭ��Y\�6d�xG�W]�֙�\�Q���{�0j��T�(^����#�ő�H��ow�a	�0gС��_8��xO=�-�@.�;��ҁ.���v�Es9��L��=�-����BE�Q���@:�ք��Qz�Nck�a��K�����|�?�I��wa��kd�v�q^;Ut�\r�%:}��[g�KX��i���yg����ǡ���pgt��X�r�t5ti�|��p��"/6:*�>�H��F=w�-���7�!)Nj�N"&�Q/����{�*{�*�m~g��?���b���������@��>�u0ޙ����b�L-��W�=_b�..��B'�'UU�<by�K~�nw������G�	2��r�(E�<�Em_���ҧ&�?q���G4q�#�s���z�OQi����¶���.K������(_g�����WK�I{Wc���h��@�I<.|-)4Q]��\��T\����X�[n�.r�"@����"&�����H���B�W��]Ø9��,�F�_K%}��$,o5O3P�┦Lԉ2�����N��}o�e L��M,�9�B�Qz��Рe5�;+e')~^SP�����Ox��Ʃ�б���"���M�M�yڧsie4\�S64K��P��2�Mݼ3{^7�C`$^�~ז~�QnnˠՉ,׉�����By�Q�����ղ��rz#*�j�:c����dh����9�wv���M�v%��'�;
r=
�f}]u	*�x���N.B��e3���.�����������C��+�|��t�
!+�=$UH0K	<}d. �G אt��m���雾��#��6c�k��S�娉lh�������4q�|%㩕��ͦ���^��A���o��'Yp�5dMx��)�PY���,,����G��Ƒ�(�)�oW��8�]a6�������>=F�a���"�_�䑑�qa)}�U�`S9�[���SZ��|�L���\[�Q ����⭝o&��w�Gȧ��+<wqi}8	5��?	>��������O�T�ܣ�@���j�3G���?ț�������8�`%\U�B���8GӀ ���u;�����Y���G�Ơ����}���A"I2�̂��٥����Z�74�9�b���@㍊#9���"Rz~�c
:�Eܑ��Q䣺�� &f�K�ژ-*���7l�~���)tk|�{�m�NR ���}�b�NU'�K������L,�*p'����?�<���G�-v�j����^D>�U�B:���s�����Bz�i�8�l�����pw]���K���Q�e��Ήk[s�Z���\:X.�	&��M^&p�IN��=��y�ԕ�o�D�,�)��KIx�v�KW#�n��D�����t�P�76�Q�R�ELF��8�����ø�؇tM��42t�i�I��4���ꃸP���ݴ��N���,4%:Z�8B��(���i�[R�R�qt�9�t�}9�S�vFa%
=X�P��������ү$��Dl��B�rLo ���j��
�P�3���$"mΐ�W��XN5��W60}�ߜC�k�P+��k\M�ci4�bɱ���s<�Pb��[�J�'&A��a��^8�(�� G�0q:Ph�u��"[�_Phsہ{H�/k@-��B�{y����8\��#���B�:G������[�z߇�aK�⺙p��x��.I������g"�`������Z9�/�haM��OÖE����1�eX"^g만S���u\��!�&�.nCBR�c4fK*K-q�c���x��T0%]r�5Y25�@��K��]��)p�Pդ�w�m&��u�a)U����{ۘu�!ڦ���b ?J�;I�\07�Y��P�����Fn��R���^�����H��1r m�S�I<_N"o1�i{�]��&�����%���O��6�qna�S��,/�i���A��:2>10�u���������6���M\*xZ$�vG�wMo�t����f��mi����edd�����w,ZiX���J��j/�tAX�K�6Ր�&����u	�P��;8n�^3�����K���?�� -6{�=��Y4�Z��ڀ���� ���i��2��L&��q�����K��E�[��b�#>ʍ��55�ˋv4�1�&�r�i�U����<F�2�A������9�>���i��Y�A�M�]K�g�y�k8��yDj���@���V�ׯ�SO�_W�TC�OVt��C�==��l��`�����k=���F@n#��Gh[n C>�:5Y^]2Zz�8�������Ӭe݊y	o��˂�r�}ՙ8nv/��H}O�6?�/���C���9��?�� x�j���SLX�r���Q��S�ML'�ڮ����ng3�����=����5=���:���.��Q([=�:�i���w!U�`��z�n�b��X	?�\%m�P�R)�e��O�RG�����ɌH�y���!E�ۗ��~#���������} ���/9y$�}�����}~��������1¿���C���Ȝ��N������� �
���ݕy��N�A.-d���U�U��JdwI?�/���UI���No�����s��Tv��_��f�7�	e/�+0���6�[��>]�Lb|��[N�*�:sx�F��E�aV ��Xzmj�?��+�;�p��/;M�p�3L�|�ȑ>��O<�7��7I����hCH��>�F���_��j0cҍ?
�!ݫv4`��h?��^��C�E�v��J���e��e�/mf����P?�_�3$�oZw���yr@�y���w)K�V��b�oo�L	�䋪x� Q�M�
���[��Kj��exE#�QX?2$E/k��KK^�ب7d�V�*�y�e�[d����[�(�wP�rtt^��2�'��Ŕ�ˏ+�ɂ1QF�Ngڅ��O�!�Ъ�Ά8l%pP�<ÂFC�3!i�u-�j��ɚy��Z͘Yu{�K���#��󑺫A�^u��,��`�O�;v�U���y�qٕ�	�1�\y�$��X��{�s����qY��:MwQ+���Ny����F�Rﺰ�F0I��%�Á��f��r�.�A��ţ��݃ש9��25?d���ؼkj���g��(8�6X��գM�';�#��<�N�ϋï��6|�����H��U��+��U+)6>#�Ai��i=�`3G�@�޺Ƹ�Lv�i��*�������Z�=�ZɁ�����f?�2i�1�Y<���W�>�u��'����o�a��<�X���p��z�ٵ{跺�V�8�F�q��!Pb��L��`��޷���vu�w+eJ�n/B��Є�Wf'�3f�b5����� �6`�x=��3�͍�@��� ����si �tCc}�|5|�t7R�2�jz>澺��\����������b��c��#$5YK��v�ل��v�{ �h#���ޱ���0�N�]�Xwl/��J�Lg
�<�����9�Hbd�d��hf$[�����PR�Ӈ��jN��3��ea��l�C5$�ͥ
�la���r ?������Jߒ�<j��;�خ��E5ܢ�B�c����h�&�K�aQi_�vFᘷ���m}���7�ˮ&�hne6/W��L]4�k�p��F���d��(9H�g�����Y�O��,1���T�x�v��w�J���Ŗ��I2
��2�0�6d��d�BƬ@�X���P˘f�2���Y���
��L�wUB6��,��pB(��u{9��4�њ\�ط��u��Z�4Ӊq1�	qq0�����7�u}}]$���ڿg����Y޵��l�gb��[�߆�o����ܱs�Q�^pڏ݋��7w�©3r����1E{蓝}����)���m����{Z�h2��;cS?���LQ�acjss��M�.1��A���T�����2��
r�����l����;XJQrc8&t�x�H�ߡ���W���B��1$��-dɧ1����� C�|���p�?��c��a<l�~Z�[�}߷1���(L��+���M�I.�jX��@���9Uy�����Q����������T��}�ެ���d�Z����`���������h<�9kI.�s\"�h���)��H�^P�O�_PFܽ{�����EU�s����u~曵��!��{�)��
��Bw���`�~��ᬛ )��C�_��)aϺ�L7��f�B�R�8�;�@��(x[�9������W�/C�6��"�J/���1/[r�L�C���K�۔Z
�/�I���V�h��.�P����œ*ߡt*��1���-��pn(�5�N��}IS�6��<)��Zy�wr��w�(`�yY+���C�Li�t�A��la�e�'�ω�bH2�q��9
��J¸;��lPx��r_��5lyU���!:���1r̿&E��4���cP�$�,�aW��ƎAE|������e=�X`�d�nR4��a� 6�]S�(�&j���R�R��\��\���w�M7l���r��m�%~	�㗾M�/��^^�f��b[��������qz�&����N���j{>*�0W5��@6dv�c�L?�S(�z	!�c;�����4���6�&�{~5�!˫��h��+fg��@p��K2���2m�w��{�h[m_n[�G���>�C���W�j��ؼ����L)g���ٽ_�������{�w�5}������_���oo��.�~�I��P:U˨����*�CDl�� N �F\nBk����&�y�N{vA{���8�-*����"���"/���b�GT�,�H���ذC�д1�^�2�19&њgj4=-�|D��ȷ�a� #	��0�mg}�gt5�It��,O�A{ؒK��/w>�Fe�)P��l�}�:%k/���uk�^�������{�Р=kB<gD.��*˙T}I�(��u�@�w�7�:5)#*!hun��Ȉ�������㎲<��0N[#8D�������8��~2_J�����La`�h}"|�xi��h�S�b�q�@�M�
c!ʂ,lGq�6j��,o�]=��]<�j;�Z��K��}�-eE�T�wհ|4և����,��MM��ZR�;58b(=�s54�?�K��_���#�8��uΔ�h.�����W��}^ݭ��U�g�S��o?^|XoG?����':|��s	Y,WY"���3! ��;�����cĥ�R�Q�T�W���`9��z�|�G��(����I!Q C�|p�p2�?��a=��6a�N��dVTRRa�X��Ta���r�j�h��e��@%�ܥ�����-m���R��惠�)���|b�ЮN6�&vQ��F8f�Ȇ�' ��y7��U~�. �T���|x+ �V
/DH�} �&
�@������${����t_�D�������BAP!S,�	��'�#���|:�&I����5���!c��9>+��/g�&���sW�;���!Џ椒 �\Jf;�E���:D�����\ϰ��
��)��ò(�ɲp��-�2,���rڍ� ѯW�6�����,�_
Sy�1��"�������s#SD��]�:���6�}���|�����ǿ,WZR��i��E�ɑ0��D�'�QP��T!Z^q��=��/&�x
xd�O�,B��]�K����#_���I~�����c�'�>�2p�LNҞ�?�)
��#I>O�,��4F��iC�0���L|���7��prr��`������R�?X7?^���°�,�1��/�Y�qx""�?>{6W>**8��z%�a��:��-W	:�1�q�m,���*�I���S@�ң��@񠔷��b+h*����p��H���9:S�2�{�=�2�<2ZJć�����0s�$�f���(B�9�U���˓��V����qf�y������N^�%���B?��!�x	����2gLD�a��v<A�u�+��M��OZa������*� ��UǱ랔,8����_J.ت���L[��-��^0^�Xֱ;q�3�>��0�\1(�(� Ip�rM>s�R�u|��~��S uۇ(���:2��H��v���6�������m1��cIŞ����?����㍏��H���>{N����~<B�L.)�Fp&��!3��ّB3s`��0:��:��eV��>--�$����f�Ϝb��-�z714ʱ?�(���APNg��:�G��?�V $m��[�]�Y��;�6�0J��l$1�Nh��`������3K�_�����8����o7�,a(��l�g�w�+6!�HO���v(o��[Ts�Tы�#�?! 5�ԣ$�Ƈ�q��"��C*$�	@��Y��~��x���}�O�P)������L����;��X�M<X�����#��1a�8!�h�*�Ae]Kܦ�u�q���횒ˌ���͐�U�U��>Z�����W.��q֧��tj�[����N�7ixk�/�p��B��Y->���Y��p�ր_��"4���v�-Q���9��� ťB��WNnzF9vZxY���\��
gw1K�:�ʚyu�j���TÓ��y�5$����Aq��:#������ƥ�N�M���`�wf/��P]ϔ���:z;���[8uԷ"(� +U+���Mm3�\g��tr۲��cdu�J��L�u0�SR6�3�PX	(�w��A�^�� ��n@v����.He����39o\_F�|���Xrs1M�_�;M:����ȚY�J��x*�WdU0r����Z�lԬ��C�.O�@�O�ǓDg3�g3D�U(5m�u�J�Ö�$	cn:��������쓬h�/�j�8�j�w>�5z0�	q�N�-��iP�[��#����%���@pIy�mIB�BW`��b�2���g䶝]�7KՁҠ�0� ��<��x�R�BWh�kJ�Ö���$�Z)�Ihaݼ*&Wu{$�%!��c�?~���G~�}#���3$]�Ӆ���l���ZLtT���L��p���	A�*;����z�k�1	Y�E�c)��01�;����ȚЩ%�Ș�~��p�O�b弦�^&�k��&�xaUIJG�M���$U������N@�7t�ѠJ�u��=�Gɨ�1�W�W��k�p.�դs e���N6<���A���=�`�8K�i#0ad�ޛn��#�U�~���
������k zC�����cӲl��!ޢ󻠣�ӘM�I�b,p�tm �I=�ƴf:9�Ĉ�g��&Y��&ӛ����=*���������B~7�?��^��[�ϲM<i�{h^�.��	�>����	��Q�C�DH-`pK��G5Є}s����@t<�&lj�Y/i�G��L�Y����z&��gS�����38�O3X���^���ŬWiX��r,`]X��j�w�z_a�	.R��Jca�O�[Qmg�2M��Dd���;妶�FZ�d��Н�8�qv�v���'�����_�ҳ���HI�jy�<Q�cÌ�8kF	*QJ˳�F�&�5I�$<Gi,�U0qX=��Y�3�!t\1\a�>	L�)�b� ���r���&�̉���H6V�+ZP�H�ԴT�a�-[�#>�;<rNI�3=��	��M��K{/�(��)��إu�T�cNnZ�u��M��`��qi|���u��D7�3�&s����M�䶛O�?{e��	��n}��uR.�o���L��뮵�� ����3^FܛC��^�---L꺥�Xj�y].�0ٌ� &��&���4��X@2&E�F���
��m�0F�ضSj�	�Ԉ�s�i7�$��ی��J�E�W�0p&�Q�=�;���Ŕ���Wh
.���Cy|aK����g���~Xo�Ũ�����_}������ǃ�Gk�6��nڛL��X+l���G��i6[˩}r*��V:��!�KE��ڲB�PN����X$J *{x�a�oMyCq!�ˏg�_�r`_1�t��N&��2+�`�u��.e}���X$�r��Б �������{��(W-�������R��tksgS��䬔�@Ok_���������������7�n=���vlSyWWiyyK�0��lI���j���?�ъ������Vн�\��Y��I9�eEO5�f����3�{��z��3Bܑ��8�o�݉T�	�|6��+�}W�V��?�!��r�OHt�B�A�o�E�|7Js���X�ĀIJܢ�s��#2#r�eY��2MdV��ûh�oc?'s(�U_<�MY��R�tcU:Kl�aG?Y�1�@�����\�����$=�ͭ�uE�z��r����P+XF����+GTN�ʹ�K)����]��tI�BF!B_Ƙ:���\�1���E�cǼĎQ3[ |2:�
�����۶h	2�!�(���u��=Fj;�˹�!�Bn8�x"���;qlM�0n6��L�јPFI�ۯ�sPKnQ�)[�	cuJ�s�þ�����DG+�!""�~�X:�&���#%�s� %]#DB@���t�.�.Q@:F�`t#H���� ! -�o|�������}�>���:��9՘bT뿎��ߧ�e�U7��,�o��<���D�7	��cO��'%�� @�ۖ\��0��'���
c�f:�����Q^�T����7A�����/��n�Y�:�~w�H�cd����$��*�jL-�z��} ���O·����7�i	M_C;>&hO���ׅ�"��j�&��I'+��>?�Y�"� $.�׿��k�u��'�!�2�o��tۈϝ1�n̐�r��Q��`�ҋƢQ��Q�Bs���v
H�w�gJ5A���rV��r
�3Hˉ_~!����G���-�A��R��^2,��|��O�fp �����Z�\6������%w��W0�w~\b�Q�:ma!+3��3�}3�Y���8j8#��G2V�7���V!c��l5�(�+{���,�;GJ�̘�&������o��݌��7�c [rۮޓ��kp\	b!����6�٠�o�yB��ߌ8�����e5�˛B����Ŧ�:�,���d�P�HLs?�����w��n��m�w�mV�e�ſPjn͖"��q�m������b#���K�]�oN]���N�(f�ݒ㨮(7T-�~=�;��s.���H?�9>ר�)�$E�tq�];��-�u��d�dd�0��e� �G�G"��)x5�텠9�9R��4��L�8)���q��� ��#�q"]�,Q��>���$��P�ZU�h��u+ǤHR�a�6C�}��]�۷������/;*�53�A�{=&�gbt�����-��\]���K���mY}�Ю�.�E�6����VsT������E��o<��h' ��K��ӕ� 97���5/��w�r��L��K�Gg�lT������ZN�GY�l�aj�b� Y��o}a{}��]vl�]��ʹ����\�?z־��~�h��prs�w�v�tT�����R-P�z��!���� ���*������]���.LQ�3��x)�˚���\�]�\��eܕ��0�W�_���MN��!q5cF�����������������_f��p�K�h�D�GKK����A��RKg���র/`g&���>�/r+Lc�(||Վ6��]�|����������
Ŗuy��:_�$�_��k#ja���F��m��C��Ϡd�>�� oW�P�����<&U�4+y{��o�<�=>�_��£,Zu��X�IyD�B��W���||i*>��X=9�U�8�(�L��Q���&�dh	�6�	�IB����A��38<W�M���7s.����~�9���I;=�؛�,�唒=7�P�|�I�#KzZ��pn��������Be&�Ч#7 �'�3��to�|}�lg��{BZ96��u	������O�߹�����w�[YSSq�1p�X0���'���v� �ݲ+~L��7�)W��~�ѿ��I"�~��y<�Kc�盿ϊ�w�/A��r����m���Y'@6CN��x����������d��zG�����E��}�(2�H{�zj�����0�XAН��fD��a�@�H�s���(LO��ǎB��_a� ��7n��;��ʩ7�@����nz��W"������,�@V'��3΢�<5]��֋Q�D����2�-\�z�����v�����@Km-+k��r�C���0��^Nz!'��@6xp�]3W<�3�D�!]K aE�)k��D	tZQ]]X�'D���y�+�5zAۼs�*񚳍�Щ�':r;v���X�XS�XË��b��Sv�T*�O+�F�U�b㱄�V�=�'~�\��1;'��GW	l��m<��+P�@`���4\��eWr2\��R;?2]���{��!�n�ø^�z�*��B�A�'���t�'�ܔ�1�-�-�%���Y#{���ފL�iҦ��o{�q7u��i)�V�u�,���$䚩��  �83��il�\P�/��y��z[q+��/���j��{5O�梔ϓ�j}|/~�
�[>�/AN�@����l����%Զ��PԨ�S���_�!�;5��l�u�ݝ����Ln/����[U�'��}r�A��|B�>�����Z�����Ӝ���+�6�$�*Sѝ�N�W~��ƍ��BD�~�Ve�O�2p�3+��}�$�%���Z�{-����X7�6�aN��3@�ܧ#�z^d���1�
�y)��m[#�ۏ|�UiSm��z��o+o6T�b��[��6�]D�����4#�ˌuV��T"�ç�H��ik.�{9�JKB�$�-=�L���%��b��a���� �mu��t�3l�ҩD�f.�����y���$���sԮ��/�|���SH���c�>!�@7iM�tferynE�5jiuV߆��:UfEfި�"P�
Cr��O�mΜ��%�TC�~e�EŢ!ƀ�Bg|����>��V��̣�~�3���>I�f�wk*?C�@�{�J��4[f���`���X�)�xd�D��$�Tq�jN��: /z��Ŷ�n��R�U��p�+�OG �C���d<����$8��e�щ���r{���o���@�0snA�����3������ eؤ������~�A�*��@#��T��<�6Y8c(�;XƤ��F��ZU�Sl֌�(q����ز(BD��{��P(����rd{����$
��HY;gX���3�W_�;���2o�ħ��������@\�HhU1����j��p:&�v$M����� ���t�����+�J�����D�W�F$�7l����W��nZ�&���N�>�e�+���ɚ��E@,�L₠�h,�
�g�H
8�Ǉ��[/�BY?��G���|�'�?9�<KX�����{��K��]t wu���/J.�ZIUզ��Ե�D{-,о��ߋ��+ff"r��k��  8�jw�3�#�_c���.�^�7��z���g�4���D7q-�q�tV�v�vv�j��~'.:9E%���g �c�����J:i�d�d��VQh�W�;8K�O�om�.S�$�CD �Qxe?IDl��S�^����Fa�D�8�O��F�:���y6
�x�\��p�bC�b�F���%>�-o�b�g#1�-�`�㢕��(�y�^7�݃�=���;��N��<�\-�c���Y>��Z��?D�8��>�9?�ԧ�R�Goٔ+�V�/���QNB�@�	��gF?�[��@%yvZm�n8ۋ�<�[�;�A�㤼�� F�-�R#h��5*�ȏ�wғ�-SEӓ�"�-`���.vI�ƿx�Kv������˓ؾ�g�� y�����C�W� �2�P��Zi�%�Q�2Ȥ�Á�i�&��k�pl�d��Uig`��h��֮���T��2Ub|8Y�����v�Q��OV�$#�ᶨ63N������b4I������8)~�Yh�}���2pҫ���,�C{>�%����������"���ئ�K�i�3��>�Z�<�^��oe�ʲ�r?��|H.������U&�Š��w|�)~�p�W��w�pZ�fz�5�P{��E7���TO��j�'q��٘ۄp^�����љ
�,�2�:�
r�k�o�X���Ή��O�����d������w�G�I�R��w.��'��Sc�MX�মG���4�f��L��n��$*�Y���f���YȤ�Lj�m��)���@�̔,�~�ϕ�l�k�m~-2:P���l�$��ҕwzkkd�����dl��\�/J��s�
6�����8��UHH��(Hש��)��I]���x{�{5]x5��u���|����FH7�,v(���%Q�B� $}4a���-pU���$3@�Ue�acVQ��8A�_$��F\D[ �����e��d!7y���6;]ŧ�J�9[��窘�DQ�T��_KP�����\��bQݧ���'\+������/9H=���wn�"k���w/ǁ�A��� J���Y��sx�Ƙ��4zO�!�I�nX�� �8�D�^�=����W�v��ev%c�/#����}"�<��$`A�ɫ'�#LU��hb
f�L�7�g)�w}��}j�J�u���c�<.Y��Z&�>���~Q)�ϭ�˦�~�w���g|hz:�j��j�6*,p�sUR�p�T�!����Y���C O,���AvV��Y��h�'7abbjL������~�d�^.��OF-�w0��E;�O�*��X.1a����ޠ��
*���H"OW3�X�HQ�t���ٍ&ܻ�%��	�5W��裝ߛ���9��8\};�Z�O�3f��SZ����=�!ː�����ЙV�����ZġvEk�⃏��켔���a��\�k�Ɍ�&�MY�����Hie�l.Zk�]�� D�rоXě��Ҋ�����#M?�e�5:ٱ�A���\1��]'�됂�����<Ck��	^B��9��9u
:�nB8TqC=����OE�\�
aZ,I}�ɽ�5�beaP���I{�jsm�(H�I�� �k����L<njD����~�o3�������L6����P�����������������ɪ߿T�7odԪ����(��j�L}إu�Z�B�<�z�Pޥ{:m��#�_e���i��:X���#���x~p�9-"��DJ�/>T���]j� ��e���g�����'�������c�(w� c�h��[e{=�g��??�e�LE��9�}�����E��u�^T3�����]'�Z����E��p�Hv�+�ۓ�~ӎ��hb� ߚ�!��ˏ�%nH�.4��tk<1�W@&������h�i��0_���q>���(,~�,4�<�̀����1���O �Ek�6� Ch��喭�����E���|M�E�h@�{�A�dr�XFP0����S����}Eզ/bm���F{�]�WV��}���+w�E��73[.2�7C�h�_�E�[���w�g��wV7tD����hbO�&�����_2|��5l��?Jv���|�qF�y��f�������ѩ�N������.|*�UC�.5��\x�8�Ծ�����[g�$��+�"�	��ن4�23�����kQ���!�Ee��q�̲�1<'�F������J�Fg�@�Q��]v,꿯˕����7�Q7僈Ť����籣)��r|T�,&)GH����d��<Hz����y��9>H�>��00۱���Z��Es��]�G���&%j��r፜���hv��ѯ�����N��SΙD�4��q�Q�"U{�c����Ξ��5-J(Sv:���,��l�0��De45�����ؗR:�닕�����諹���Ӛ��c���J4�����0ص6�jE@���tPk]��Ǭ�U�'���L��Dn����t�m`�#NBf��	�,��qЈ�������U�U�a�ܧ�: ��!�xj��B)�C�Zf��Dq��'�aQ�d"�`�lu�@�=0��6#�;���O���u�A�[�G���W->W�V�i#�:U���'�Ǒ���4
�d��h+�=� ��-��=
��	5Cg��w8Sø���w���`���E J��1��h�~DoP�6����U�`��Α�쉉xB�{�f	��C��Z��˦�J�%�8��"Ӝ7����~2v�1����9$��S+������<�&tۇC���hh�<��d�]��INDC�L�u���UW�C,�u�h��yP�֝�|Mf=�Ib�J�4E��4�	˔�sU�(5��_^5��ĥA�Fq�������`*�pR��nl���Y����eL���s �X�i?Bfɂ��#�.%?.��>���H*���턵B~{XH��a�I�2��p�g?3qp��y;�`�r��d&b�,�pu��#�I�;;���KD<�4hP9�,���&�TT�F���S�obL
�M,�io��m�EmY�"������}���\?lDO�&Dѿ�~VJ�P�ax��c$�0���|! ر��E���'؜���UD�M/Ǯ)�&�4r3��nA��I\�K�f�l6�B{[�P�S�
ɴ�
�B��[�'=�c_ld���vjϮ-��*���6S�^xX1K��
u|\���8���b�@r�pl����t�� ]�ڣ�!|�'��	��e��n��h��S��H�m���@7��X���~�-o����X��WK0%&�];#�v���22_�\��C�Ϟ��#vO�u�p�*V1k�{Șc�X/f����U4� L��5;yr�N60mOE��S�?$�m�������RR�����a֋�s^�p����G�0g�<a��0��#ݰD���ilj���Tp�_�|�7���{�r�H��w�ī� I_˩�>����;��C�@��-) (u�J���Hz)���d�F�������+ż���kΦ�jF΢�(�|����ԝ9��w�#��m�\��V�eON-\��0xe���]�L�Qv���l,%��SE(��ܸ��Pr赓��\�+|S�RN��S5���U�ޡf�jk�P����\;Cb�!qļ����Q�Q5�1�7�n6A6�%u��llC	6��
�A��^�P^�����퍟_��[��\��������<&*��[�����������_{���c��cد_�-��/=�����vQ��^x���`�����.�KāT�/v���x�� ƾ'4��+�lYc6��8��"���	��9�6Z�?�l����'��+�N�q����qzgK?}��FC��������d�9��VN-*�e��mZ/���G埞r�S\������~����"���Y��cQC��= ��u�g���._1�d��U�_ȐQB�'�|cl�`N2��P���q
<����u�mv�R 0�0E�&�]�����$��U^��*i���c��0�I��~b�rr��7��=6�{��V)j���.B'����)�H\K�@Ze����.���,n��݃#h¾@�y�/�>-~�T���E��	���΢%��Xj�Lx�2B���d�<�p�oO!S�\�=�QźW�;����3��DE �V߆g�e6f��||���!qdO�+�Ҡse�e�q�+/-_$]����Z�O���'��pP)��͐v�
�,G��n�6Z�s�6����ך��_yM�2x��[�'`x�#���1�?�^wV:)o�
�<D�괞Sy|s%��|�%���
6w�=����r4c"����
�?4���F�r=
�{H�R���,�B+�+܇�ckdd�$K��i���A�cg�ȭo���0}�Fv3襄Z��ġm��~3��'����x<��99LMX�z~cd�~o#Xc�D �>�X�|�h�N$�!-y]����IΒ&
���v��Դ�|o�!�zݰ���0X��M;>܏�F�f���A �A�	�jݸ�\�����{+�0aecst!y.v!��b\��@���Ȳ�C����A��RF�������D��;���\�5S�O��r���qlH�.��M&�����o������^f��e�t�ɨ��J���z"o��d~���q�&��O�֨ĕ+���>�����P�@Y+̕*Ε�}҄̆�(a3@��h4 �3�J'\����_ȁ�>%! ע�@L��g뱃�z��y
�~�����;�����\�e|��F��jW�L��)Ķ��ڢ��'�c�E��1��J	�v����m�^��ܖ����mb�m���X�,�w�t�ٴA�4��4oQ�+ѹ˖Y���f���l1��MW
���׌r����Ξ�t����%�����?���Q׃f��?�G�D~0w����X�?^ӌ�?��Fa$tJ&���q�h|�-A��X�cH���hſ�ի�&b&�����T����ˈ����)��Glg������4phP�񇑖��3J��|R���V'���*vɗ"��4K^�u
�?��Җځ���AY�U{M�m���ځ�I�<���Au�w{����[tՕ6�Z����]�P-js����$1/��9�Ԯ�6N�|]��`:��e����I?�?u�'LQ���E��rYW��a��*-�`J�x�P�(	����?�U��i��~�1s+d5�E�S
ƽÂ<� h%yy�ւT�$5p���ȠX�%�ѯ@K��v1Ƈ����}�[7�/n�[�d�;���J��N8�����c�|��6��(UIS����N|�nel��*����":6�ݹ�RT������~v���>jzF�*���&J�A� ,�,����	��T&#^;����}o,Q�.o?�!+���������5~?�gvxug�qz�V~�is�78����kq.�w\`��dr�����7��c�E��e��OwWW{V/R�gJ��%揝j�ڂ�6��Z���Ŕ�TYx�MIj:��(
5�K�NEI�M�J���	�0��P�����a�`vt������˵��>�^��8�W~?0Q�Vk�V�d��]2�l��<��y"4����f����dU�U�+@��w:᷺�Zh�@� ���܅ �Jf�2AP�������9�j����.�k �����5f�y���8`�m�-���S%ap�����גe�+��J_&�卌�K��^���e�G�f�3α���jG��"�ܕ����Iw��ء�����W!pk�>.���'O<�N;��*��|xeU����l�l������/3�@S`��&����t�j��ȱP������b�tЪZ��\+j�L��s,�<�t��2��Z^'iýG�Į��'���KP+���-Hf�?)����	B�n���%OK���ߋ�K$1��s�������yTT}�x]�R�~���.�k"�g���V�
����	�W�8+b0\�\ j��/�3`���f���f��+�œ��{��{3��}[k���}��X�#�&8�?����t:�PD��,Fb���!��� Y��	y�?s�k��?�8F��B�,��W�[i:�m�����V����v��j0����֐����*{n�lU��%���k�{���X��7\�4�^�GU�B�#K-��Jd1/�-�O����Eb�.�t(O$�9�Riv�C5�0�X�0�p��J���cΤ��E6n���n�A�x����(
�B�]��#���l�9,dh���"
|aU��uap(z'3/Z5z��q��z��r��ٹ���|bj�������:�H�U�&�K���������Y2¢�c����<�wNn4A�A=��N���*/dp�w=�� [�>���*4��#�g1ܟ3=�H�z�V��� �0�\܍�bs���v���wۇ��B(6D29��V<��_���%�T�D������z���W�� J+y*�?MV�|���	���%�̬(6mr�Xulڹz�uőˣWuYRy���a��
)�6[��YU\(�����w�l���G��Th�"lf�����3& �I �����ME2U�G�'Rh��vZ��3<j�[
��/M��M�F��!�B�q�(�I�c��m^�)���g��c�'����+G���1����v��ɠn��h�,�r$�m� �ܚw(ܺ�pm2w6�s�8��Au���5W��N�|N�o@yd��0���Sgm5�4z��f���u�zv��x��u�Ptһ��X�.5N*�&���}i��݅d���0�S[��)�#��cS�+c��W�NZJ�M�8!��y;�4����|97�3���34��׻�x�M�T��ks�-�̙��ٳ�1�H��_ڒ���@�o�ė�G�.ռ�k�O��1o%���(wz+	-�� �Yi]��B���"-��K��Ԕ	���VhD�%*Q0�(H>��a�I0��O���i�'��%��5�0�hr��ug�s��^[�%S4w��^ �����62�3�؟:" O��>��I����\ F~J��J�/��a�#��Yq��t/،��^��I]��nŵn�U]����F����SG���I�ݝ��x��
���ϊ��c8��ZEōG��\���!�s�j�16jȘ��V�����$��N��u>���ox.�P�O�!�"�����J#qx���0�� ^�tV�s�M+�:_���;��D�N��9p+�S�Ͷ\������+�I�N�1/�L�׏F��o��bƞ�.�y/W�?�hG#0�b��N�y�b`מq������_��	�z��AV�Y,0R1Ռz��F���'Dic&���'��Z)˝Ug/,�դ���3)�ʢ�T��) *�aFi�by�S�T��@	QՕ?���j�eǪ�Z����	�~SZӊn������yn������2�EM}w?;9,	�@ш��P��Oƅ�Z~_k��"�qQ�4egp`���ұ��Ev�����Q|�S)ʴ������={�Y�ޡ�G�R+��������.������:ζ6OO!��*!���z/��;(L�C@�o��~fRڶEb ��T���ʳ����p�����T�;��W/�o�� 8'p�������j5�M�ϸ��Sر�9�uJ��"�K�`t��0���h�o<ՌY5����d��t}�I�J}Q�e��s�`��a/O��@}�DfFԀ/����k7�ڭ4��}>�kfO�3�����A39R3�«�b��2F�b��ֺZ_5u���ki�G�v�J7�^��SC=���2��tB�����i��jCWD3�T� ��h�e����$j��,>��^~���h1O4+�P�7�b��۸ �'�̠�a�#�X���4p!��n�@D�e�|������#�]�����W����S���зɐ�z���u앜i��'�d�:1�:1�7�_/��m��4��4f� ���_gB�k��NΚ\�b���?��}��1���,���Z�D%ɚ_m���i�UG���^�OY����QD*�O�񓤻�Si-�	�>�A�u1���{��`,ך��O�%��S�3e���#���?����xX�qe)+�ð��"(p�6��Ey{�1R�@��҇|kT����>}M�s��w�J5㧎�~�3}Xf��.��~:��;�=8}3�9o�w^{�}6ig5 �+�U�y�K��W����öVu[�2����~���qMн��^�̤륡Q����x���c���4h*F�T*v�'j�CЀ��;Q-�܆���ƫ!1���h�u*۟���$���5%ťn_-�>`?�^z�tS��񞫕r�w���@�8#� =
��T���C��߿]~U��|��o|-E�ybO�p}�]vl,J��Ä��6�U�OE���=�<�����#eո��� �t:4��i"L����
$��	t����
�N}�<9r��wD3���Cǃ�_ۮ3s'�3/�R��K��䭩�"vJ��F�w�/�X��0�$���Z���B�"3g\�#tV�?V6�Y��y �i��+(����x�9EUKW7pv|c� �7Ű,ح�:�18�7��yz����W�����E��X�������$�E�(򅩭�YB���o�N5�1FC��~���o�,�O���ۑ����48.A�.�w�!�v�٩�d���ͦ?*>!�!���8�-�����`U�#=͚��Hk#��D|)a:y���a�rw:)��8���v�o��q`�ncXv\�t��e�1�*Hgj�?M�MF�]d��~����4F���W��:�k�(O*�WV�קi��xwv��iŝ�V�W��#�:o9~H�R�P�óz*��jP*�ء%В  Og�ǖ2���2:D��}���Yknz���yI@�t{���_���)P��o����>SlP�ڷ���2=2��:V��o/g�}
(a]�b��1A��R(��m;%i��<k�g��H����x�-c�����=8��@���[WĿ�������EVW�Ws�Lr��2��n<Hg�2��ֈ���R�D�FR�2	�?��E�֥�~�!��a�E��H�1����w�n����5��e���J?�	�l��<�ʯ���]�M�E�R�DφXtp��M��\��ہ�>wKJ�n��������F�(���5耰�_�{kzT
 C���S��L.�4�My�޳W-b�-��b�/Z��[ڿ~k�3=�Z6��쒋���|¨����A��Uߔ��W�{4w��'6�[�6>!�!��+r�F�a{(�/�
V
�׫�D)$���΃��?	$��"�Z�)��@���U�)�x�k���<��h�6lJ���D���Uf����1?{-G�M�5)�[\�Hͅ�R:{��GK�b�n�[k���Ԩƛ����Z���U���T�!��W�T0D_!�B&C(�R��[�&�IB{�y��0�Y�q�v,i�Y���4�$�O�T�`�dSH��O%��!�URm�x��L4�F�#uo�����w�훫������2X6ƪ��&�� �^��ScP���G�#���D�Y6�$3�R}5��x7]*���⽖W�w�cO��za �s��:\\��K2[?�`���08�U�{d��g2J��Ʊ�u"�����_LU�R�?�v�
qeg8��3���d����=��"C�N}G-��ߗ٩���䞁6��zO=��}���m����w�G�fO����U�gfj����u�P5�W������^sU�������<�?�q�h�(*��1�2PrJm-��Q�;�R��.Jzӛ7i��ي8Ϯ<��l��'���#�#1�9����������	 @�j�S)�7��m�r@Y�{j��9�y�J�����I�}0Q�kg��n]�+a|��u�8 �c��^ � 9ۇ@���=��Y*P�VQ^6^��+�N��q����U�?Ӟ��kD_�N��Mk���M,�������X�^QS�����������^�����vN�G{~��ɻ��7��ƃ=�ׇ�/��d�� 摰=�H<�ؾ�聞on��A�"̧�)�S�n�3Q*pHH.F�o94�ף���a������ �`0b�rUو��� ��e�Eq��ڒ:C����ztM�w�%^x�l~����7�N��_�"�q{x�i*��"��[F�>�m2HܴEؠN�f�R�P�о�
�~G�"����/�NchK�֣qƲ���@\�K���q�|��{����5h&��qҧ�|V�S`�?9u��f����Ղ(}J�yC��B\=��?{�;Okj��<\������)q.}
�r�w�,�h���v���>>��-�~W��\RQi���R�߃��x�Fv����8���)������;,F�$��˰\��O3��i�7~�Pr�z�Ku3��7���_ ��MM�͑C=n��G7�?���[Z��қm~�wY�ĵ�I~)���2������g���Y��|Tq����P�ܼ�`�&�,ԃ��oJ�D:�|�l&'J1a/�Ս�k��;�*=������D�F7�=��i&��prW�F�KRdb��;�0p>���*��jB��^D�,�0�5�����^�@k}�%�#v.�>.�΀�f�����T�D��U� $�P�F6�f��KP�U�*��f �Q<D�5?;񭭬|������u�r��r���g�%;*ۓZ�/C;f�ĵ�Kn{��҂�T�#%^|'�����d"�Y+�t� �� Pw�DԘ7˺�>KY@�~2�)y+5>v1 hx��80�����2
'�(��2Jk}��}�/F�T��t.[���e�~�3�kA��22�.m.u�Ψ!�<�.���>�k��e�Mŭ��q�h,&'Q��z��΢g�S�&�Z�w�����#曔���В1�J�8�|H���6�߅I�s��|�'Ų��8��B�����!�?�^Ҕ�H�'�1�NA�b*4��i��V�L��OІ�N�OS�� P�q�Oހ�8&�,r����#t~?5M׶z�Lּ2���y�K�4h�zՈ|���q�U����Oz�H"���I��<�oILo@G���nZ%�L��6*C��g̗�iwP/<f�:yy����ٙ����IǠ��41����k����y0����v��4��|F%	�6��Y��DR'��[�+�r.����;^c�%#��q΢a�~�Ҽ>�;\����6I���k�����O��	�O�f=jv�_��Q����%C��o���#S�'ϐ�?>S.҈�c��"&�H��)(Fa���m����d��~�=���������B<��?ۃ��_L�d\�1ɛ�S�g�S�ФXæ��q!5�-��ů�$n��=f�_y�]xwm��uD�1��e��[B��ա��>��>f��g����'����@ �����F?��b���	��/�s�� ����Ex:��;-)�)%�(�"�>W������GX�+�:�}�O"UD�2�n6�6��K�^�l�8��
�Yû׉�	�
3yN{ܞ̈́d������֞�՗k�e�w��������!%mv!��%��d�����&WwB��@E�A�ׅR���3r��5����'?R��1��ٯ��V���{Ŀ/��0��ҿ��_6b�e��n�\���MW���v�V�28no�o����h6Kf4�ܯ��V�r~���e�g#Bɖg���;O3��r�z�p�
u���Bw@;���+R��s�0W{
E��"�-�(�h���f��`b�X��E�W��r��gO��V`��˯Ѵ����9>v)�P��r�՘D�=B?�{5�S���������+��%��i���Ʈ���9'�0M��>s�
�\lQ��OvY��B�	T�d�LI���L�/,ȉś0��i�!�07!{�x�G��O�ey/;o&��_�~�(�ZA'�P���`���n҄r' ��c ]�?����(�����9AMv�;gJw���x7����!�l��5�!-���ge���0'Q)l�i��V/`)_���&C2�N�[9Ҽ� ����w	�8#gS�\����+U�,Z��1�FdDc��e @����Pa0@`5We2��ݣpZd��0F�4����/�F��vZ]Yh��Z�� ��1V�"%�ȡgfu�G���3_b�S$6��~Ì ���Ac,��UpL��
n.z3Q���M�OhH�@>������d%"�胕�&>�HGy��V��|m�F_}�_���o�zq�P	B�����������2=�LC�L?[e��:�SY��� nn��Q���{�]BM9��R�ظ�A3�,�e�k�97VUW�?Ӄ�=��T}�*׽����pjk�pN�{/F�:�$�<�c��w6��~�A��
�OO^`p����S��i�yF"R>�P��<�)"ѷ��,!l�����4[�]���f}�m��Hm�/!��;�PK@!F!����̼R�_�LM�K��ʆ4��4}�Ԇ���F�JO8c�jq�4�2�ZOLT}$�p���(�M���S6�-5�4W������.��1���w�'S�%b��(���A�]�����kJ.��OUl1�Ex�g���J�OѬ\0eU���w��J�C�<�@�ٻE�;�{ɴ��mG�
�dRF?�~��d�Ŵ�9θV�o̢�s";�2��:S�y�]^�v�=w���&��A����5����m��9����-s�'��`ql���d�_\.^#Ғ�#���'�V�9�X�cX��O����	�����������p�sz�gi�&�&:��VV�UV�f��s��>Yz�͝ �s���d��T�n�&/;/'9�f�:�4�m}7�.{�$-��n�h|ؑ�DF�W�K\�b�-�����ue+ -օ!��#��$��I�ti�|�;�����5��2�n�S�pѠ��������,�Rl�$��j��=ݯ׋��s����V����)��.�X���v���umw��l�4��m�3����X#��-6����Aƈ?"$�������������:�-��|��	|~��J%�)��k!�{�������O�n�)>��Ὶ\p`P���xw��x߀���������Vv%y�� 2��B[�IX�*U���xT�)�]N�=�f|FdiO�"J*]�g���>2�??�͙F�S��.���&����&��R%����XY,C���~�Մ��
�;^o��r!�x���t�=��e����?��*u���KR����cJ���VE�|�@�1�~���!���j���r鸠�*��1]�:;W���Y�U�?2��0��SF����m)T�J�	mjC���w��%� Ҷ�=N�k
���
�x���|iU�G>"ݺ|	 �����j�뢵�oђ"�-��������N�
���Bqw�����z��~���M~$��\��{����3� -0;7)޳{y
�"z��xE`��ٹ�Yؕ���vQ�wr�s����*ф�Y��>��Wv�pL�[�K?��Я���;��_�H�ޗ���vQ�V���Y"Θ�^�+�pӡ'ҼH~+�d�Hb�Z�*��/j�	��[Ӑ�6G�;�® �ڜنK�֊����jc2�縊�.�٤1-*���5X9#-�¥8�i;!����� D~>�c1��Z��|kk��Ƥ�X�B��$u�
.��u;y�/\i���#��pl�.x%�(����̸0�e��7��R';0�B j���i
vr ą�QC B��1z� HW_q���ÑT�a��p���sԤJ_�e|��[���<�?0K!�B��׼���c��S6��5Q;wT���D�6�?QlίK_��8t��,k�Sx��5 �f0$G(�\���*��kނ�G�����X��.���^p�=��ߴ���M���Ӆ�u�wh2��디�BRȅ�7��ɴ8z��I�.�	�Y
��ڨ
�x	v�t�{S 
�&�̠��XńI;&AJ�1C�l1m��9�H%0�FV�������J���{Buާ��^�Q(o��0{�k�:�8�7f7���' ׼����g�1���o����~;����CK'�^�@�SM�Q��c|9�֧	~?g9�����+����U|��ToR�#�G�F�a�Dx%)	�ʰg�o)T����oR��R�-oFJ%�yc�y�E�T#�,�y������Y�Mw���tT�l"w���Î-םT�gO�WO�\D:��7CLC��t \�z:!!j���z��o�}�����CP��c�g*�<�2x��g��N/l�������L�|�����[�\���@�������"������mZ�˧�IU���9�+{�쥨x�9r�\;�R#�ؓU֌zJ�V]������i���^���d=�(�h��ʻ��W�1]�0؎,��@�������ZZ�l�w9�E��C^hM�\�T�@,�~��LN^Q��M�c8����߶�آE,�d*+��(��,� �n� ���_'r���/��w/�慄���H�_o��Ena�q�2�biv�v
�����&>���T�(D�4\)��-wf�o�4� 6�RB$�?��U����$���[dCb�'���l�O���b.2.�zi��X�,-cρ�Q��x���J�⧴�M�N�:�Dq-�I�
��A��-W�ʝGY�t����Ǖ,��z���1m�ŔI��y��E]��b��]z����T�W�ę��qO�Cb�ϙ�U��e�o�yB�ݩx`�/�U��Ջ^x%:���AaKpHi؉!����DrA�))�BmƲX�
�Ex�$����	oCC����Z��@R4_rU��k��~�F�C���z�"]�q�CR���2�he���0FZX�]th�_v������R��V�ZY:�ebef�zp�a	|o�HY[�F�[Q�Φ�[�E��}HW�l��Q�+���^�Ã�g#e���[��> �����y���8&�@&�i�%����K1��&�2�����$"���0����G�sHe����0�g%Y�@��7-3�'��/�~���/h�z�:jt'G�m�KI�{�j
�0g��@x71W`l�r��6��D�%��
�Z"�V<�Zr;2x���\B��Q�ż��iC���Ֆүu;���-��a�-�5�6�Rt�(�55F�'��1np��s��1���8�S6|uT�|��L�oG>����7n�e<�W�>��+���~K��+�cS�j5�IŢ��O�|Pxwv�4OF��5CF��-��|<�E^�9N`�* {"%n3��X$���*�l��R���aE	�Ӕ���鲑��=���p�{���).��n3&�G���c*��f2y�g�����'����|���"��"~�*�I T(�B��V��l<_���ii��1��ו��C0���&GIh��jV����^.�k��j���J����y� ɛ ��j1)L8S�
A�- pS�RiT����a݀�uq�`��NGy�'�l��Se�B7&O~�6j���O������ݺcBQ��&,����'�H�)�Z�]-Gڃ�T��S*ք�hf�Ԟ�q�X��|�aǿ͝s���Y&��i �_�����|4�g�Qw.��hN��|��b�쨢6�z�ؤ���˹XhD2�cGѭQ��RJ��d�}L7xCh!�I0��2�^�>
E`?֎5�μ7D���aQ�3$�@(�A�T��_�`W����|��O)���z촡m,��y�z�^�K%(r=�Ku�r�+r��t!򸶓�ט麡K&]&����f�:ү9������K������R��H�6k���f��S����6[��Iǂv���_U_�\����O�?�/-Q��NFja���|ڑ�uMd&.6MW�Y�n�[v�l����;�p�Iz�� Gi�Oe�L�pc�[�o�C���uI}�I͖?Z�;��F�!퍖�ƣ$��^R �B��k��n� -s�O N܉��t����B�KD��˩�;#1��
k�7�Z��{s����������4��%��U&�ۆ��O�(��X�cp[2��E���� �f��G)c����ɋ�o3b��f���z�2��!.��x?d�ūha)z��J��e�c�>�TW肉̆�����c���ʉR�m�+���L�_�~�:i�$eS�<]1�����,-�U�hHi�cA��±��z����iR:,�t��?"�	UƸ�����)���LR��d�H�D,Љ����~�:ko�q�_��k�Ե��M
ML�� �?��-"�&�$�<�b�@x��k
�)���(�S��E@>��yl��>���	�1�-'�Ip�V��L�"c���Sk������)��W��j�ǽΣ���p}Y��8,c��b�ĪBF��'3tO]��3!*jA�pU~���=4���M��N�|�ڙ���Ca��* �/�ݰ����Y�N�{3�Y"$�({�20���#���S "*Ҋ�63��K�iП�q��/���X�̻�����W��k`��~`OnW�iΰu�.`a��e9^M���aDTUY^'P Ma&Ж������ѱ�!���*����������`�a��R����N_�n0��* �~}��#�q��	�����Rݎ��4yԞ�C�C�s�ܽ&��ѝ��69��h�HV=���C��u�͸8k81��xWd��� 0�=<�s�:������ͅM0��b��L�ot���Wf�=7���K}n��`o�I�%��8���	�gLR���&������h~�ٛh�0��lA��tV��M�l�z.?ـx����y���+��8���e�}�eW�VA���B�ؼ$�+$������1�l������<		���'��v��U�F���|��u�՜�ES�%d�ݥ-&SG�vR�F��ng��J:�� nqJa<��h��A��A��Vx�6�NB+���۠C�)h��~C�E~e���;��\q�gM��v�.R1�Rp�h��~	����Y���TФ�@> �)¿9&�mk�O���Vf<OYH��@�AAry�	c
�\|���[�($�����0RjÊ��Z%Ȳmk��.��8Z�a%�=�)ks�1Ω����\��u�4�=���ҝ.�P��}���ۀE�=�/쭶��Gr!Oґ��v`��~-�sUkK��&�Lȫ�;A)���^���×�8<-�a�%H�{X!r�$������= �j0e҃j~G��(X�D3��d`~:���|��+��e��#����N���ZuYˏ���Ӯ0]��hP櫨���
I?��)�x|]�O�z�[?An�J�L��,iWJ���{�?Q1����a�(���@����GS�pR mTo#f ��gvN����U&�>^٬���n��B+�Fx�=�:{8��M��$Dv7/R �6����'n��J�s[�S!_����7�4E�d�N������gT!�TD2�}c�����5��RG�Ƽ�f�!�d��$�F����J[�9R�N-�ʦE����ߛ�N��`9�J�(B��)�Я(x'��tRh����X��^�;�\%8FQQ0S,/4�TW�Թ�of������ޮ�u��?n4�;�n}8O6F�6���S^��{'�/>����,�K:�6#\��D[�	�s@��J��`�LFo�~����n�r��fo�:����W�l��l:|��}#��T�{�41[�nnn�10�BCC�~���fL<�F3T�M͠Vb�:��ݟ���տ6�EI){��jm	�@AVm������ȦL�/S�v`ւ3V����L�שJE�؉�	���bY*����9�k�m���"�}K�mSʝ�%|��kعd�L�$M�`ϟ{���o2b?,�6���T�F�e3ѻE�攀�t}����.�G�3��E+Í�v*�yW.�`�������C�#�s=o��\8�� b�jX*��Q	L׆�ms��w��?��-X<��؇ړ+�B�������ơ䋑�cigD�Y?�W¢X�k]�d���4��ߺn]�b�_��-����)��S����DN�T�1N2M|VQK��JL]Ԍ�R�hW��\�����m<<,}���ͺ���d$�NCN	(G*�^��̳�7���_;�a6cpE\��W)�a���D�C&)䪗����4h�$��#?}`���6:����Z��H܍}�����%,�>*WWDQ�1�:��A��ߠH���e��6�66�mP�lm�H�B�kc^|�N�k�Ը������\���qk�ĵ�{d#u����Q��f6�������t7�r�����r���	�$jW��m�!��(`��W�����Q��T��T�cM� oa�{-�C��G��?>�/.U�ν�K7�y��7N�#���kf��b_�Y�Wc�8��}��-H���R`� m���lPrZ�H�~�O�`
9�,�Eo�~fưA p�C^G5���{B�a�����4&m{�q�"���ݜ���HR��izpT��G�w�M0��yo���S���ǧX�x��g��w.~hA���u+c���]+ٸ������������ �΄�pGoX�l�צ��5Z���%�ޝiCP��#�n>��n(�E��;���,�C
~�r�5�*I�
~������:Q��TϷye?o73��EB��;�"�H��7��^(S��u���>����S�9�E6�J�����PN�0kRSpic/I�̽�X��X�9S!��sB����E3��]��0'#�\��|�Ȅ&��}�[�,���<����z�&�D�qX�i9��͋���M!4�
9�!��z�J������OˣNX���F��BYx�[x�O��ys��F-�2���B0}�YD�R��	�ʥ?�_�����qp�e��p�n�0�Տ�.��1��W�
���b���f{���nhRJA���90�~<�Xu�}�V�Q��h���9&���k{�P���iJ���|�M�4�s�\I��y���c0�ȫj	�h�U��6>��D�����Y��[y�g�-O�(����傅���,�޸d("֜��l�0�%��򟝛�>�A��%R/��?�;m[�`x�{�T�.�CX"��"n��ˮK�Z��<#*c���ޖ���8*M�4��/��>U�)o/���@��弽WE��������N'>�0��x�]�>��>\�R	�ܯ�,���M]�mat�52�J�7�JL2HI����ك�S��{/����_�T��"׻�4��� �����|��Ϧ��I[=��[0Z���_�q)w~�ab�Ҫ�ºG�j�|a,��¼<;�r�p?��z>�1>soص��]Â ~�u�J�g�{����61�lG�p����ߠQ�7q�0[�ҰS`j����h��s��0��*g[��Q�,6re���p��O������j��j���s��מ��XYU*���Xt���u�A�*���#��e��`�Q�ϲ��beaCԊ��Y8{��?
HBLj�I����>�2Ps?tuX���a��#(��1�m���z��,�G.bO�۱��-Ѯf/S ���)W7K�+�;�Ews�{�����V�ކ.jq�>�NПnT�|�p3��;ǵ|b�-�O'�r�<��=�[>u��t�"�r��y:��\���5Ȁ���=�|y��fjmE��\�]��x�j.EF��4-��<�R �����ی���`3Dt-Iu!�N�~c
`�K
�H��� �<>�=��_>V���nnn����.:_a,:,�x��;.�!��m/~�k�[rsvC��ߍ��;[�~�d����ȇF��������g�;e��$��=���r�� �j�V�Bf9oz�!�x�?NX�jt>�|��u�j��o4puiX7�h��)�T�-�S���9���?�h��/�3tiZN1Q��z�� �;�8�+��ഝs2�2?'Am��ZT�􍽃B�Xq}�5-�^��5�%%�063:��%�ԂZ�B5����ɭ�W���@6)L��[�4�Qs��s4Q�`m����%~�o%\�c�<5j��b=���Λ,c�wC�t�+t�miG���Dh^��B�F�l�u1<2�'�2>�yKߟo\���E-t�I`����	���8�8�T����)�}D�<e#XuZ�c�M�L�d�/�{&�:-�J��)�8�@kE��`�Sčxk
S����J��Ա�W�p�e'VA�0��Aw�@f�LD��O>���?OR�썐����8`̠ �d.�B����_\zC��t��p�����(f�@`���G�p�.ꫪ6&=�)����4�"��'�|���>��vk6Tw���N̳�o�v�ʲt�ڴ�ɥ*��U� ���Y��So��h�>�0��n��|8v��u��ԛAT8���0���������A��E��"��w�³=����{� 
�AT����]!H�^:(Wr����G�DHa}�Dm=����& �|���v��K�K�v$tˉ����x_��t�O�Q=o�?֢?+��^9�$	%�[3��G�Ch"�!�+3:�"Ɓ�c�|s�6[��3�-Bv�r{ؔ��[���ΰ��2�Nfo�H��I`#K��(
��wװw*��׬����l�������}�<�J�~��_����Y���^�������~�a��Zs�RAN���Zyt��m�Ģ�Y��fJ���Vz����2���<����I݁�c�w�pb�ksx�ֺ��*!�G�M'�+~WK��l�3׬���у����h�]�05zF�4c�W��4W�Y��Ga	�q�ң)J�v�b��s�z��-���Ax�:����',�śz��N�+)X:�(��`�zGx~H�]?}}a4� ���݌X���D�������=D2�8�3�U�Kþ���n�'����LZ���[E�e�=SA�~T羕ZW�-��|f\�-��Fb6���W)��NAs�3`�#H�m7�2����i0B���^f��$�%{�;z��k��"���:p?��NOvߏ^��Ϝ�[N.�t//�0�ٻ�D��Ȃ"&�������}m\��ҩ�+X��Z�i���i�tz���z����EJV��4ǘ4pYE"���tI]���5Xz8=v�o� �9r�k>qK�"3�ġ��e@��I��H��K���R�#(�E�u-��X�HGV���[VV+qͪ�YR/���E�B���iӗI��E����]��:�,���J�م>�egWdA��ۺ��&��/�/��X"�J^��Cw�x������]��u��qL����ܾI��V�I���ɣFXB���[�B؍�/����M�"�ԃ��WC�ߊs՗f��'��oII�����f;�bx�A�l��q߯ �Da\��0~-��I�ʴ� �)�E��cV
I�C�� I�H��!�����`��ّ�"����? l )���]��vh�r����Ɂ��\��jj����{�;ѷ8�g;	h?�@D�Z�f9�g�$T����Ye�<�&\+�:�qj�1�O���x{HB�[��]+�NOm��]t��.6�
.h���RY7\g��(	4����
��e�B7�r���R��!��pn$~s�T��l������4C�w��j��ɁuͅL�&�Re텁G~>�� T�<��8LyH�I�M�Y0̜7���b��m����q���0S����:�Ԋ
�U h�����d���t�`.I�TհGI��4>��$��gu�;��ۇ:�N|���A7�9�s�g�a�3{�*�{��3msw\��No=��p�1	�%C�-B)�$��Y�W�v���("��I�1��i�x\wt��J1rV��dk�2�1J���iL�2��1��4Y_�uҟ.�] �E�/Q�e���h蓓�
2Q�J����ߍ��/�k�*��,�@�$�y�9�.���8)�q���	�sv��h��,����;�G���;21�c�3,Yo=��f$�����`4�
VY?��;�!�p��G@������ٖI�M翫����V�Ǭ����s����*�<��$�x$x5$IVa��F��O~��!;�3��a��q��7o�3��n��W��t!�^/Z��/��tҳ�؊k��m�Jޱ�ܥ�N����]�hb��K�,+a��+wB}G�����akTX�L�;'��^,�}�N���V�?>�/��˔��><���L�N�;���D9�B����|<��K`���<S���{f�.�o�4����>&i�L��j�r�������gt3�wF�΄/�ޙ�]��=�������'�S�����Q��9�f�	/t��g����Jn���|��z��������P�R��Z��Dg��g�TG�7��S�Nk��26R5�MT���o����������?y �����'��«(bH���5~��CYܺTxK�A �( ���V��ఈ����U掤�a�DJ��/����a���J29ۈ�8����6毄D�pZ�������g'ϊ�\����������ĥ����G��xp�}yz����&-�����h���r��[�/s�[�Ǩ������DmAF����ú��lfl&�����Y�w����ֶ*�ق�ِNC�0 Ō.��f�q���o^QR����<�\��<x[��uu����� L���E�]	� ��x��	�B`A����iI�0���cv(�_)(��%�v��￥��x_��ҕ�U�n)o$����~[���ʵ'�(��X��wb��V�U��z,
.2�4�kU�ڪ����m,�j���$��0ݼ�E��%U4�A
dY�W�rTik������b�̨h�'0��S��0��` ��R��ɣ�
Nh�E2��"L�2PHt̆��9�k�'7@��,&a6Ŏ
F@j�$o�T6��X#Z��<�x��b?�<͹̭_�)�jN�ѶgDB���RP�Hz����W����.#NP�@�/��X&���'�)��s��]��ĖY5�3xz���xL�5sc��t6�'��O�"�����F:rE"J%�,?>mw>]����p��&��U NaTEq	c��b5o�	���g{�T|�0\�;΍$�h��l���j��3 ��5��[/7��-��1�($��.?q5��<.�D�I,(Vj0^f-%�Ԉ��D�18}�����y�g�1'�����j�6q�\y^N�Y�ƀ��3�;W\��cT��r�3v$�:�1������[��b������I���_�n�(��-E��z
�\t�2��ȥ�j)�P3�|���C�E�mo�'� G3�������Ns�J����'�l����.uͭU5M�Bl�ӳ���R�A]��?�i�'r�Y��6���v��:��N��g\�t%G����ՠ��r���E�3��um�`�:Cxg��W	q������7��d����_'�ʥ�y���)�6v��	V��hf/8��,`3�/�f���	 �j
���R�S��Dx��m�L��4\���UG���A��Ӫ�풛�n�&���"��>שS�N}ҴM�)Z�R�XfJ��(I�K�N�Sෙڸ�4:}+2��[c�ő�'��9G�k�b�1��-	}�����]{ݨvR�E.��`�_�P�bF>�&P���4��~�u2w��b?�����6>���/�)���_�Iw�.\�:����S����'�2��I�������}��/��*��Rj1���G��,e��@!��T���*�UQ�^z��~�����������*9�j��7Abh�g�ax��[X���r
�ټ���_;�%�H�{���>�ּ��ס����a�Źe��>ߧ�9�ZT��Ƚ����S3gx�q1x�$�2}ױ�j���}]ΌM���?��0f��٩�j�+���μ�#�����L�����ѕ��a:���ɘ��dc����#*��Ϧ�e5�#I�?�+&����}�4T=+�[G�bD��*_�Rؕw���!5��`��>��9�{��A�,`�C3�f����nf���Qag��!}*醛�D"V,_^�ҟ=mV���-7g��7��8�Y�ƙv��%�8U% ϫ;F�ϯ�gW�2<|��V�+���C) ��d�4��rUT����_�Qɻ����Ԉ�%H��E�#�B)��w�O`����;�gAOq�
}�#�
�$}��b)��=�=w��g����A�����Q�c�@C��B���oF���^s�q~�Hg~�L�!N��*��4	5]5W_Ӷ;eB�k�3�C����i���p:'|�y&b��;�ф�����L�REvG�[?r��X�m$���/�%Ohq��-��7��-k��d'<~<Y2)�Uژ7w�A�Q"�m�rǄ�߲���wgN�W�nkys�������*����c�o�v�58ia�Znf;;��S)�n�<���0�Hb��G�أ�"H�������;�=�����8�����\D��5PILx���iw���tpZ��N,�,��>Z��*_��i���p�P�`,��Hs쪹ƀ�d����G�KK�7H�^U�O�x���}?���p1�S�ɺ���f.��BT>��X*n��EG�˸�\��)F?�`9�.m�u>�O��>Ŝ�Ȯa��Λ�t*���#�2�
6��R�
��m�ҡQ�]NS�9�A����$k��}p�"j��*v�?�k�涵���f5Y([�	E�":�~��5�k^���(R�hLo�"B^���}����3�����߼�����>�sKS�I�zӪО����q��F���K����^��=��<6�4��l��Y�^���&r	���ʬ~8��>�?�I��F��I���)[�r]��,mL��e��	�'�����SlX��WN����d8��;��p��R\O���vf|ꂫF[B!��hаu ����/R^'�RKL��B�?}V��A�P6���������{Nf���;Z.:�k�n����<L³�K ���A��y/Q7֗_R��6���✪�����b�n�L=�lM�7�6�-���~��.*�yYŹ/�>����V���' �B��1]3Wr�af�D�����CGҟDR�����H����#������P���kkgX�'f�2t�S�ݛaU�oW��P+���9����_)$��������]�mn��+UA��s�8���oJ
cP�7���t�_=ד��.�*߳�p*���Nc��Ǖ��ڧ뙕�ÒQ�3^c��46��Ӽ^c����+*
;����;���U~7Jo}��H��S,.¨O^?���r�::��{��y�z��RRb��gV�C��ʸ����h�����?C H�H
J!��FqO�f`��Q������U뀥��n���K����ѧu���[J�!l��i��tD܈2m�����C�{��������%����>A��;�ϕ��]�j:�rê!�cE�3���Q��ĩ���B �-��mo+�6H��0b��8D&,�0r���xB���X�dvQ �2>�O֎����>�OV��V���R�/���jk�eG~���g�!K�XQ�j�hw#�c���nw�{���[�AU����ޕ�WXVD=$cp$��{�V���,�<!:���k�����V���B�v�yX�0�_�����|�`Ȉ�K�6���#��@��>�>G6�AX|�@N������d���/�s��y��{���@¼��p}s�L*⎳:M�ʭ�!D�=>�OU"�7�4cN���=c)��4�́X>����)n��0�e�\����Q�w�n=����Dw�(a���Ɛ��X7�,����4�E��z�c�_���SK�7�D��)F*�E�����b5�OD�N/�.��Hd\��T�U���ع�UϦ�/�S�h���7��D�����`�d���_����;����UX+x��@c�P��/��&�ea�ia�1��I�i͙�e�D�L�RF���o�1�(dߋ%�H�:�����k�51aތ�z5B�04��O7^�'�gI%�����`��qA�����f��	�k����D��FW���5Q�Di㻻��z{��p���G:��m7o�Ry��ct��d#�ڌC>����ε��b�;k�=9ۋF��g�u/M��7��r����o�gtqm�'�V�P��)��XB�~H�v;�[<�����ɴ�Έ찷񔤡�������ޏw�4C�r�f� �rZc|
�/ʥ��l�SxIi�2 �9����Y�����+iu� ��@=m�o��F?�Q1�UJ���q����|mj�A(k���j��Q<�{딚���]�X�I��ο���(p'��[n�x���e�$gh����Ԋ{[��?cqq�u��U���t�!���<�S���̨Gլ�r�΃�d@\sE�%��5���;n$^(���w��$:#'e?�X���eC�r[� ��?Um�l��3.	Yb@��v�wR 6�� �c\R��M�NF~)Zo����MZD&�m����=8��U����<ڭ��o�Ĥ�a���Lsr�s�ġ^f~KT�MW n����^�h�~��	x8z�x:�m��`yؾj���x�9jy��𿘫]�=��i���ql����
8m�w�U��6i�9�p�	�M*\�׭O��݉W�H������,�ڎ�Jokd.�R~C�}Mc>�gC?�.��6>S*��q���\w�������Q����}���c����R�J����Jw�����F���P���)�hq=��V~ d�X���6��&��N�����/�)T�%΄��e��	*�����lZ��q.�ް���tɖ����ܥ�js��S���	�f���`#�w @����$���̱Tv0����&����JOQ��ŕB��#�	c(��!�,��N��,�]����+����P۝�O���dZ6�Q);ɜ�J.,%����V�����݇�����H���4�U�/��e\���N視]�Rjw�h��S.{����d~�?T����8�/�H�%�T�2���%u.7OųL!��FI��
`[����#s���@1��8��y_�C<���g/�����퉜oA�����6fA�x��oTQ�k���J!Ihm(���HXt��8=��ybƨV��zf�B
�l��ڢ"[ւgN8���x_}��D�vpb�cUVA�1I��F�q�E��ρ�9�J	�yU2�B��N#�����ء��ВD�i:3&A�HJ#D{�iz�~�{����<=`ơN ������D?Xu��9�w������:��}�Rm䥡&,vȶ�S�Nr�����(�L��}�ێX��� .��������_�����B�:#lPzc�wPҙc,��������Pf2J���U[����W��G@˺u��#g��_�4�Vٛ
5�x Vza�oM8Rю�	�-�G�e�ncA]���B쑅�<�hs����#�R8~A���O���`fE�{L�\�cVoyAgB+������i5�Q��c�dj,�~t+�ͯB@ƌ���q#�~-�~-u{����k�n��.��$�b���A��Ms-G��D�c�ݖ����ҕ�s���Ȭ�{���ѧ�(���#��%zff�w��v�*f
���
,���-,R���D -=�\V!X廅��M)��e������ ��;Z����X�ƃ�w��%����6�k!��\΀���e��L\}rY7�<r?����R��Q �3`pS?R���Ix�������|r�ByN���:fz�`��@]����Y��9*�9
�@�,l�}�Q�6�('�F�˼��Y��&����E�J�qw�@��<v�v�����8����a��ԋx���~&��z�M�x�1A����5%MW��\:&�6Ϳn@�Z�_���FvzӢ(x��V)MM���0�bb���P0%f��|�K�W�e��x���H	�6��CU�T���`��<E��W���*Bü���G�+�;*j�_.}�e�8�����K;�1�h����|��Q�&�{�z� �[9SU��a밺����Wq�xT�$�c�s�
���H�&j(�K�^l����~:�Bf���N��~3J�X��dn����� �nh��Z[e*��HT���ΐjHe.jM��@ȑ��Zݟ�t���XuV)L��=Z$�n$䑓1��?`L�$�k�J��:�6�5K"7c�{a����mr��Cj��XF�윂�>�s�Ի�� .v����wq�_��w����j��l�s��}�}g�v9le��a�������W�^��ό�7�I]Vw�o����ӷe�s�SyT2���&���Zo+��k�n���U�)�+��y�����N�n��z���x*n��y[ov���;������\唋��S���J~��u���ixʂ�}�Kԋ����ˁ��c�_�Ğ˓��X�)��V���	Ϝ}	�≳E{��<IĉK��̪��~R)t5�J���|�M�j���_l�Qӑ��(b�G�s�pd���
���m+����@��
�&����=�����k��;���`�2-�DAJ6v�W-Ru���uu���m9!!��cٍ��᳢ S{vd���;֏���ɤ_"���Z����?##�оo��Xa�ɠ�K�w~C����yu�Նߥ��<E���C�M�����%5XO1z%Op��P�ڛ�{3�T�h�1_K���Y�v�)^`�2���G���$8��ɀ����zp�`T@O�(�N>��K�(U-E�F���7j21�㊕/T�uPBS�
�~��ׯ_
�E~�ঘk*7@�E��£�S[�_�p" s�.�	L�(
�
%��Dk���H�B�כ��1:N\rS�a��SΨ�ZT$�>��Iv�aI�nWr��$�e�D��t�x��T<��=`o(}0k�e�q�ҚE��vN�ͼ~�]��a�+�N�F�(��pH"�(��)�m�>�7'!�X�˭�a�:w�Dz)�A�:������NE���� �Q {2���	MT�����$��[�1)ۣ���+&��|-�/��
��ً�!�o8��@+5�2���������(��<!N5C�?��*_��R����Ω��fe.D�
l��b�Y|a������J���-��ӝBs"�1Ip*�c�EḴ����+>k��쀾��[jl�6=4��T�8m}�V�# L[����^�M�͕R#�P/��C�ɺx�Q��j
�im��+	�0�<�?1iY3)�uj�j�}���L=m��q�x�s�].i�����d�r͇�
���ٕ��_2�t8q0�H�ҽ�,Wc��������-��1�g�M���p׊�2�����)��-E	��&z.V����������A�ʊ(��w.��|�:��ěQ�O��6Fp���F��,�ϰ�Ζ���X�3�:ZE���H�ٌ۟p]���ON���� _ �� F�������%$�M_:��7����t��Tï�����x��<K6oE�k�ep�P3�v	=���+����2���.��E�ܥ���s3�K,�� f#{i�<K��V$Ui'G�I��3 �T,W�h�H�_/��ͮ�G�ȏ}�ӱ�U�WK�KM��O����<Bˢ"`�Yu.J�,�n��&�R������R{�>��~L��e/ۗ"�4b����T�'-�%z61�����T����d+��@�kխ� ����gx�B"����-�B=}��g��Rb��Lۯ{cʅv��_� ܩ������G��k����g���7�GP�4(��=���jƊ��Jk�WQJ���fQ{���{�ڿ�?���+W�$�+�s���>����WN�g���b��A�	�J�J
%rJ�Q*�=]X80H�G�B͍�~a������M��ߪ��^o5i�����'��@൚W����т�1N)�
2vm6c�'XI��f���Љ.��������]�wBO-`��?�|�"GR�u�
*�=��FCY$	�ʑ����Є�N��ɺ|�1�?,.-�r�ojm�x�J:�=ݱ�}B�?���S2���2�w���ko��7jB�����܏�
�/�U�%�o��$��s{<u��A�����������e�c������I�����	�����q~�[�'����R��û	��f��
H(�(*����b�C���~Ǜ�)'�X�*I���t���(Zu��R���J �u��
��ަ�=kt+�����!B���ҟt�1荍UxF��/��Y�51S,=??�u=n��f�ޤ�h��L�P�$���;ptt��72�0
ZZb�����0���krbq)*���www�����@�����oQ�卓[����K�k��!>Rm���0<�Q�VBbZE�U+q�m�K��&P��У�Ζ���P�[t��ڧ�@ �Fq2Ma�'��)@��m�ǧ����M�2NH��䔲�-�ҞO�Z�@}ۦ�}��m�f�hEI�u�$��<_�**g�O���"�팝	�+����⭏�D�taf�aYQ�h�2tp��=s��l�Q�ý�u��������R��:��~�C�9]��d����i��)�J������B�HB`%��)�z�+|�\�&tɰM4�`оgb+�"uۻȭ	����ef9[_΅�ѵ~G2���q+>�
S����#d�{%�/�o��!+�e�7.~������EF-U�,v��U�A �h��Jk��\��d�J'����A��L�-aZԱX�7Or1t�E�x�;&�+3T|ޏ>�f���SI��4`��M��BL*5�4r��?�nAJPٔ�\U�.l{�!@(WR��6߈�ӗ�݋b�+A�6Z$����~A���)����k�9ٴ�8*�8Ǒ����4҂~��f�o��m��F��ъQM�� @�l������ ���EF���C'y�
ϐ�.� �ݓU�R^1�̤�~��爝S(�>��DHF9�p�&O,�:��2�r�S�vi��L�(�-�N��V��H[����ㅳ럍��]�-s���Mv�~ey���rCOR<����߇�G����3*�Ư!7~\xa�^~�/{��`W�BW�©����|o����,��H�L��B��įԧ����d�S�������5]~s~g����@����yT�ti���	�B���TT�O[�^�z���������@NAa�)��J�m�z$���z�(Gs|�/,vV�L�?{�ͥV$v�⿡_]��O��?}sX7%�l�ؙ���t/�i��D}�_@ 0�uAc1�T�8��Ho��,�f���l��8tSD�F\
�C1�N!�v$�3c�M�!�N1�t�x��)�����zo��*�`�C��xܹ�:3�x���J �N�i��Mn���CҠJ�D@@�)�/p>>���fS�+`�u�`4�+���]x�����].W��{[��N�L$�n �~DG5��W��'���ތX��@~�7�j��/���9��}$�6}:�|�����:�.[i�z���a��p/��7'4<6�N|�*����L��L� �*LG��ګQN��aj���]��(��s>�ȴ��o$F��u]�J�J���\^�U�?��@�����>���(��t��Nq������\ǁ?�j�=����6ڤ�kff���� �e�Y�hN��1���i�F�����H���z/�p=S�K�
��G��^�/�ͦ�K�VN(��8mF'#"~1f���	���^{v��t���^cD�I��\Pz�l�C;2x��7��Z|6v�}��$�5��I���-=����=�[��y�i�sx|�wx�mj��s3�]_h1hr���===���N�M����oLJ�f����$��Y�o������e� m)��bŗ�b��C{0���mG
:�����~�?�~��#�	I��`o�ۂPk�'��3��M \i��ⱇp� %oJ�?b���\3ݺ,V�m����Y�GDE�q�r��GF !߿���������%***111/�)�G��jg,�H��T%'/��];ѣ�g ��L1/�;�'T�fK�9T�����X[�<��Y��U��C��I��RL32�h�A�ª�V1�T�ަ-�[��%m�_�3^޽�����e�w�z/��m�!3ŉ�pk�wR,����N,�@+�K��3��b!O$Y?2�ݏ~kFسW������! l%�UOQ��J�j �уW��f��O���������� ��%Ԭ��~�4u�[4[t\����R8
o��D�*��yj�'�J��O�w=D�<�4u;
�Lh�οx�m��J��zs����7`Z 6�G_ГV`gha�Ľ�`���(�np�q��a�ľ~c��ċO/4�{�)1x۸w�sL�-�{x���Sˆ!���e�0s�\*��!A��;&�8�L�)���XA���5��'�;��r!���ʇs�0%m��F(Mw�lL2H�."T�������F��T)��_�g�����qJ�r���g=�I<՟���ߝ��^�nQ�� ��&8�K2�����~�Y&��4#�6����0��{sd�T
Nz68��8�x��7�4-����
h����IhI̽$��W�B��e�t���6���9�_$��Oi�L��/���73L|e-W�{7^��眅�H�FfXA���`���n�t�ag��҈:��J���8ײ��m��#[�v#��ݮB�.�[�Jr��ܴ��OX�t8�G�W�5��xǿ.�\����2d�I�甔��7�I.���i��e=�ח�Ō9��[�Å��){��+���Ǉ��=����[?{�ݖ:�*��@<�{����P������������m��ŋ222555`�3Aj�b�K!5�ש|����O�D��l}�M~s�XsI$�BUn��V$�C��~���?���!>�*C
Uc_�>轌�n�D������� �ĭ��Ǟ�7zk2;�OԖχJ��U�>~%���!ѐhuA@�$ڢzQ-'���]���_��_Ɯ��l�(.ʇk�<�/��&�1��ld�S�\�A�)H�3���0'^���ͦZL%1��������n��0�K035�z��/����~i@�� j���(�40!5W%C%�M�&gE�I�7���ad[Mְk�)���Y��q�s ���n�:�{�^{oD"��h:�/��	*8Rh2����0|Y�i�/�;�"��8:���W�����'{P�6���gyZ�[fk|����� l�0���� �^�!�%.� {X�� .��`y�?:nF%a��Q��hD��=pD��̤˚ːe��ɱp�����?ԯ��XZ1v�`�BaN�Ϭ���bP+Q~7 M��"U��`t|�M��iiT��D\�E��?ɕ��lzK�!I�)&D�6�����'����?�h>=�&�I�.��><�.��:,��W^�⹵Xw�t}�@C�r}���D��h�����ܸ�t>d����i�C��� &F�Yy�`��~��`{|�����ť:H�6��\q����e��8$�§�}J����0������}l�cM�9_|���� �Ė�z� ,τ�7���z�"��"��į��>�Ca������_� xazrav������������?|����%",,�$$D�YQY���z�8m���Y�7���W��Ԅ�P ��}��}��p^�=��B!�4�;ށ�8� ^ftxP{Y
�� "k�c��H�������g#�l!M��-�v-��Z���b)�1��&V�=�-	��+�<�6��+i�mg�-�D� ��*���b�k��_t??������*x&��E�RV��wd��c��W�)A�� ��HGr���|a���W����H�~�9��ek�NKG$�H���g�K�r�����ݒXXq�2�����#����v��n�&�n�6���˰j�21(���|Qz��b
=cp5�a��
�GHUa��0�Aq����	َ��f)�?կ1���>��}r5�{���z�:�����r��o Uc���qɞf�kF�I<��;X����dXm>]Å6D���p�9˶�jy6��V`��z��g��*}���*��iR�"��i��	��yS�5b9������O�]�s(����k���{a-1�䅙���� dd����ח>?�;43).|) �_(��Di@"D����R�Ǣ�����c�-(	S�`Ż�V�a7 �h�2W �q�m�!�f�K�p)`�����`��z��tǴ]������Ż���ǻb��M+���I�?'�q[#�{ݷ>�-���K�ꐜ�=��j&�Q���"�6ݼ��c�`5(X]m
*��q�?�\� �=,�\·�<��=n=�=>������������(��8����������'��I�u��$$$������`��H��0�[�.@����%�,;+�2v�"�6c��6�O�A�_s[��[��s:���)9�pQ���2~�#rz�#��`t�Sx3�6T�(FN	g07�Y06m<��<qZm���Ij2~��0,o:���16������Bޜ݇XyUn�$��0�����Y��[�ɴK�\�za���o�6�IO=&O�@;OӔ�ϗF>����Q��큙��t�伙6Ǯ~���c�����;�DV�(wʄ��؞�����F�e�.%��}��Fn�cG��!�N�vªՖ��ӽ���E��9S�8+�M?O��=�2<( �ғ�̘�ן��I �Z1;�6�7��[Qh4dh�e����A�G	�D
N�3�N/x��c�ص5�Oi�� ������f���=VlflD�sҬ��BM�)A���w=%���q������mk[=����k�˩�,����p0���i,�E�8��������;�x������6��x��U�s�gl�87ĳ�[���_�q%�p���y�����$������K���3z(�5��Z���z�r�{=�1�T����(��@?���l��sz��c?LM��f��c��	�8�c��N�ӡ�@�i�������}��������Zw�,w��4󡝭-ETWF�F^YɃޛc666555LLLvv�0�@����n&��vR�+2�j�J�O�b���{k@&<$'�	Y�$����h�B6=_DX�xsp��Ũ4:>�U9�f�q�f�E���U���������$s�^��T�V"�&���5����� w�lA����^���o%YߧȽx��֡s��V� �� |��Y*��B����/0Vĭـl��~=V��+�h�h�P�����T�&hmk�15��������¢��
k�z���A���S(o���}�\���Skx�*
�}��%�<��"I���hRﭒjO��p�$+br46H����)wg�D�Z=?��Z�j�$M)���+t#8dP�N<".�>��/T ��#�ݗ^C ƿ��b������j��I5ʶd��ϼUn;UJ�)�}6��-�����ҖQ0D�� M�"
D	fÎ���5j�Y5�{�E� ?؜aQ�z����?AT�TI�5����'@�{��dO� Y���Q�V�dd�J²����׃j����e�MS�n��)�bB��!h���G ��$z�x�*r9Q�6ʩpb5�w����[���ޑh���rWA�Fz(׺�����!���J���y����3��ec݆0�J�n]O�"
6a������Q˅5��bP�L҇�|�vu�d\��CZ��%���٤,�U�n�_��bG]����MƈD��}S}���m��y+���eLF*��b_���M�mY9�����Yu���$�FR�F���$i���c��H��}~wK�#�G~��-X��Y��W���s���ek�g�CCC9+�����O�,����44P(H@���-�����ɔS��$$�*m�.��.���L�d=B��W��u���K#ok�f��j���LKi���J���!t{P�Xs���g NH�Qy�Qy��$!>��|o9�ִX�h���*3f��<��{���p|bѯ�&Nʠ��-���Ұ]��e�K��0��ɥ}�H��ϲ&δ&�.�zY��Ym7��0L�Oô��C�,�J1B�z�(�bF�*�ˁa��-�"RRg�_a�t%X�ws��'���b�^`�̌J5"�R�ה/v
������~ycU�aV�]�'T��Tȿ�#��yq�U�8*�a{h+�K��i��U�M?q�]�㫯,iЏ�O��!ͥeC3�1������f)�n��(�N`h�L:��MT���*~q;�@:�ZC�t��b��uyg�љK��KL�0�M H�(C����)Pq���qU������u�8�Ʒ.�q����em�x5*"0��V�Oi�ܼ����x��=iƸ�{���}�y������]"�~�W#�w1qK.6�|+�^u$�җ��n�ͣ��R��U)������ZyV������U��z"��)�ss+�U��!��R�?�w�����:����+j/ǮDo	s�^�WO�Ԧ��~��#0��h�">��ڶ��-�-�(.|�=KMU3���c=9 B0:0$�W"�W���ss��l�n5��������������pCC��MRV=��ё��=�G��jpz�|�a����y����������Ց��i~ddd��o丰5���[���>�V�?��;沺��J�M�A��P�C��� �.�̞0���hK*�`S'7����$�@M@	�����L�iKqŝm��t&��0#S�:�b*�q	�<9e�^7�b�I�
&�e"�+��J���������̤�6��kŬ���P���RX�W	� ��c�#�Y�h[G9O}�,~5W�;[���� ǝU�n��ؘV��)`��U��1�tB7��:�f�5I\��o;57*FQ|ŀ5�����*�#=��8����3+��^��SbxRX�>�NX�Zv�	e'�8	0�C�>?!MN��יz�R����ئ��ẓcEqo��&Cy<�јz��ז�Ǿ~dQ��.�{�����>N�
c��S0 �[&���r̪>Z�}��VZ	l��Z��4�cj��� �:N� BIr~� �I,�/��q�����tܜ,�!ۚ�11NX�51���ޮ1�1��#��)��?(���
�&�q>e�-�:)L��:��'�P7�߳}	�j���1�{��w�LX7�� �ɏK�Pb�o�\{�i�\i�2.;�a_��~d[;荭���og7�M�|MM�R�J����L?�?�몤$�C_���=���O��W�'�ꉼ�N.�h��'mk�O^b*'�m�:���C�l�Ĉ�	}|$�:Ʀ@SZB�ϐ35�h���[*;�� =�[a�����#����7�bj�x��=,,,--���JUUUOOOFF��fmm��Gu���/,,�\ &�J/):����]5P�~�n�M�������(9ѫ.�6ۢ)��fk��ic��]�K~p��]�k���3���J��6JD��Y=�f�q�Zy"E�!����Ry>����
�|�YS/_G�}w����(����Z���gÏ������W����B�QxΩ<�=.��Y���T8p�S���z8_����o>R���M�a�^�nx���>!.ĝ����4��e)�`%�s��i�U~�b��W��b tM�s~l�l\��zac1?�м����:h�Z���nq^m)���	 �h&���9�s�ܹ7,�r�@��:��N���J��";S7�S��5�k�/�_��>J6��6�K8?m�[�إNU�Ȟ6�d�$K��l�"z/#����g�+(1E�V���wn��n��Bb ���W,䛜��Fi�9�BbJ"�]�|nRK�%��D�O4���Ud�-a�6�k��Ϸi6�^�=��AM�=�|L5iB���g���?ޮ�?�������4���	ϵ�=�ƫ�0��CWڇ>��t��[̛��0���O��F���݅�6��qzM�o��i��4�Tt�[`�Q��Z�RQ�4h��P:��ĩ���A?���M��.��� ��c޼(ڋ{��`@��}�^��x�G"�3�������4/j�-D�8d@K�$���Z�߿U`��,�-L��������*�������,����ܜ����c���������xxx�o�!-�˽�R���v��a�ܬ�J~Rf[ML10����&��236�Wra���0���W�W#�n9m��00�#t�]� 	������]r�)h���3�������hM���(�@F��E�L�Q�[f�X�I���xMڄ�Q�Ll�~� �
�G��_�Qǣ@%����@	�!j3�H�4�g�:Q՛�5�<՟]��<��P��ib�e��"+jw�/����ۈ�ζKux�d|š��J���\]i�@e�[e���_ɪ��!nRL�z;� >XI3�a���W S L�!#�<��s�Zx����$5��F�S��:a�ЦR�|�W���%��by}��+�J+��Q����)��o̳�9�Ֆ	���CEe��:Q�Iױ?nsRPis�y�"���O�ʼo�EE0�b!��eM2�A����t���cն^~0uh|��h���ԊO��@�}�D_�$�_��Vl,�V�ȕ5�l�6����Z8�U�h�X���c�xr������cU���$�r��Z�1�������f����`�kI�8p��x�åoӥ/��Ȟ��M�nCBJ	@nư=� �%�dqڌ���UUeBB�����0x�m�1K��	�fi�g��,�ʛ6�G9�ۨ���f�����ɛS�M�n�����%ח��C{�n���nO��f���2pX�]_�P�p0�M`�z>�ݼ�<�6�,)��|͂��[EA�.��F���Z[�6<��Jm���/PV����E��(+(���qpq}��yQ��-�ۅ��56t��sU���NV��F�i�v�G�#��ϝj&D���ݯ�����fr+��W��o�l���r���d;��O����0:Ԥ���0����a��i`�����!W8ƅ?: ��$d��k�����S����dn�d7��3�}C������I]Z!uz�E�_��5Vʇ��4�xxy!�B��g�Wg�y�+v{)\�O.i��9:�f�&ZL���+�m��C'>L"�zށv�W�&b�c��z��h���J��W�H�)ßi�����#��_8�,����4�W���ܟ����^��B�X�V\�R.6O�"e:6j�4�����Wë�N���r�Xf���Ôh��`C��q��W�rg�0�������	�F��v��#C�ͦ�~����}�L6�9��
�5�d���n�'�+�ǉe�����k':v���lJz(W�q�x����X��"�ᠰ���Ҏ���ʭA`Z1:.�Y�\�xE6I�����U��1mb���P\OK���o��4Q��q�d-�~#*?
%���V쯇ώG'��2/�C��gD��ܐ�����c�˺=����-��۵���7�S�?K-g���i"�K�7�*�^����t���YY�^���Vj�_?)�����wn�����-���^�﻿:��D.Q��y��1��'��"�S^�,1�������,+��&���4���CM��OL➯D�e�����U�{z�c�\�� 0�v3����"����"ck� #���X^m%�����긪�����ο�P��w������&����^n*RF�r�1��͑	�w������Z��z'�2��Ǉ��8(�7Ǜ]u��I6h����.�)�?��bæ�[<E|h��R�Q6�S6VKF~�� p�M`����w�7���Tq���x�&��f�6��\c �+3Ρ��&C�i��^��$�2���կ������nr��}��<���\�f�(�
1�N-I�Z��竽�Q�`���P�a_x]��ӷ�a�J������o��^<��C��BN_�Z�F���)��	� *x��y �t���#:ې�#�L
֡
��`�/��Z�2)��5a�����b*qr�<��+L�1��������ڍ�,;���ڌe�Huh�Z�to��=&I���U'��c��5w֩h*CltI�J]��?ԍ:�'�b�i�r��!%M@�k��v�je�:*;/ ��g.Q^��=�u���}j���#H�ϧ��r#�9�{l#���l7�7�+��Y�g-��r:x9�}Š�����
�v͗�/'����0*'��;\3g�3g B��ľ��L�jc�W �J����&�~�˿!ڱ}��B�y�6d��:E2υ��K	�An��'��g%���r a��'&��|�5�b�ҭf4M�8�k>=���(�`�1@��?�T�J�fz\��!̥�<l�b	B�`ÿ	,�������ܣ)vS) �h�!tA,��A}u� ���є����)�������8��Y]��^{�IIsn�Ws�B�C���ˉ������&cq?S��"��b��0[�I_5h���q5
j�4�sw�n�Y�HV҃��ۉ[W��*�aw�@K+}zb��W�H��ntzaqf5n��e�a5��&���3x��pSt�I����J����%��&r^�G�Z�Zm�����T�R?�r�D	}����3���HU䷢ϣr����X�~R�#��P\�L�'�c�;�)�������>���%�1).!	)^�@H�zGi,��)� �43��_�^��9��8V�ύ��PL�m7�����Bb�X���%�˵j�J͜��1xT˅>���ᑐ1.fP-�ը��/|՝�;��\U��_���C0[����o��e�	��]|Qjo�k�LIF�xn�<��=��9��M��5���_�٧Z�T ����!om�G���w�2�ȊN�K�7�B�$����JM� �5<���U��� 't"�4�dT�� �"��=\DD��V@�_j�`�����7�畫+fe��Q�֯�G.��ly��������߼\?�%������R�����F4��p�gؙ�<�8߸Du]��F�l�"�s"�3sU��hK9���v�א�0kw7�W��4�5�*3����EX@��w�B��]�1}顯���c�lo]�|䔒�V���b:&��~�b<4���c� :�Ȍ;>��d�>	K���q/�%��X��tx- ��\�'��NB�O8(T���)���k�7�d�aDU��H̻�F%��P��W�5�)B��v��Y<�Kf�O|�^���T�T��T��P����~�������ק���w��X�Gb���2=|Fr��I���H6-7�ӭ���ɍ�ԙ����9��Q%�X%��s��=�C���-������~�����ƽ����M���ť���ڜ�b����핸�n��5<i��ྮ���~�n7He�q��'��au�+b�g����򩠆�3K�4'�w�c�Ln�ϱ�e���e���77ߋg��߮apOwvv�����f��о�aH��9�mvF��O��OpWM�Z=t1�w^���ԓU�4q�E�\ :���X>��Xb�J�fS��܏Hv�tQW�����D3,��9&~N����ja�[�̳�*�l?��q=<�R��:�IU&���zu�f3���˪�j_T%���{��5E���c��<6S2=wYω� ϑ3hD�_��,6y�H���.lU�U3ԕRԔ�5�Q�����["
�'Ԟ�(��Υ�����(~�V$��.�Rd�Nd��ʳ%��Eۢ�ҝ`҇Մݏ&w�+������"�Ӥ��P!`kZ�z��4�$��-�N�%`�A�'�m�*�$�W�5�Ղ��=�[�k���E��ൾ�wlAk���&�@��[	��aƙ��;U)#|	�<�\�q�h9���W`�].��K>(=n5��\{��Z�����=��_Xh��2B��EeH	Ę������rِE�دɫ��b� k!����J=�����s/
�䧐6��zQ>s
w����A6�������/f�N�>_�I]H�����v��wF31���G���8���]���me�'���*���0����e�@��N�Z7�m�-'�^u��{�k��al�2�L��� A;\&�4�r����(��YTvG��L�w�*�/���ҕ6S`�wD�6�Fn�D�̾p?ʋ"��NF����������@���^�`x�o~щ�ǐn%��U�`���'�Z��qs��=h�l�𾂧H2��i��2$<1c���p�#}Cp�cmB]����	p����ݛE�����&#�^v�yE��}b��8��E>Bμ���WF<^ñ�SrVɍ!����9�K���;���I>&�J�MV�N��8li���'���E�(o0�[���F��<e��/k�_�*�wi����j�h�J曛��v�/�hk}^����|CC\P[�Y���{��fX;�ne��{��ǂs+L$$�rsi�D�*U\0<�-���RE�j
�,ȒA�����䢣J���v�3Si�MwV�C�w~E����f7�Vk��<��k,h�˶��ME�r���^��߅9��{�ڴ��L:������F��E�ϵ첗l��2���C���ڝ��v���S-���P<6��s�uˏL�a��8/��,;aP���L��&R�y���8��,a�'U�=��;�E��*�5?�񋰼�t��P���NaP߰����*N���{7��<�4u�u���MRe)���M�T�#B{�v��W��͇�!�1PQԑ�NУ�7��`5���D����|��X��s�j3U��`���(2��]����5 ���6p8�\�����8��n�n�|k��xP�ET�aպ���� ����
�b������G�2���`Y����e$M}��	O�{�:E���&+����5�Hgt�+t�N��a�I��B^d��>�b=��:V�Q��4��]�����5ol5R%@���������o�1d�mE+�XĮ$��n���GB;[c�����K�%䤠o�%�27�c��WI�Z?��8��)��0���W�7��?f�-���d�yu�P�[6�z.��������a�?��9�{������a�w$bs������iNP��Y�ܒ��Icy�����`�����FH����AJ��53�V�j�o�Y�!��B"":z)Q�8��Y�-���JJ��o����f��F4_M9uX=Ai}%9�ѸE�͵�9e��� ,:C1.{�1�70�J6]�G?��d��]�5����y�U��oT�G�pjm��K�����E�++�z��DM��z]�[X��pc�u0%��Xic�&�}ՌQ��mZ/&���C�9#�3�I�w>�V���q��X�4y����V?~��>%���<���O��Ӏ�"L�f�$�x��	�g>�;����Z� '�E�gI�C�D[aXc�T�#r�Z����H���{f��x\��[MdXW�MSbl�a��M��� F�	�'�&J�p��dU"7ϖ*�F 1��Q�B����1������iы���{��="����e�jڿ������~2�W#�ށ%X��[(�y����vVO�	��7P��RP���
1��N��o*J ��������D&�p��_JP,{!>p���f�i�k����;V�L�'P$ԍ���[K�z�v'�!G꜐�ÏWݿ��L���(�LJ8�A��B5��_�a@�M�:�q]y����M�U9*Lɯ���}1�ԸV=ů�t[���c���)�b��8��s����}�C `�?����OkJ���FJ�I+�(�ӱ��
��i��ł��~��0����,��Ц��|Mh�8�er�īMym-��)f��)A*W�)=l�x�2Z�T;���G�4u|���{8�2�N!������Y8P�B��Т���E�#Uї�\�.'��J���ό�s���)�����E���wmt��]����F��JM�9�uҖ��x���3�jksk�5GL�-�$NY�$. )�(��`|�,�5j=�Rz�1��������}wr������h��A��B�D���*d�=�c�@ht�n�T��P�QV�P6��*�����Rx��D��X�x���+�٥pDx�#��:Ckl����t�3:�*{���q�ٕ�Zᤉ�"�B�pS)�,�O�<Fh/�ن{�l��K�#Md������!%�(�=�A"Q�z��S8o��}�E�2J}�JĠ��/���n���+�Q�/7�R~��v���q�_��Hps�Uw��.{�mp(g`��9�I��vq�Q��ښm/���<�N�B�@��U��/H��ϕd�4d��@CLJ���[	�y�5\�`-�'�yh	[�
��Z`����o�
^>I�#���g�����ח%�\�O���Rs��N��'k=���FF/�H钗��[�I���V��QZ����~ԧF�d�9�1!XZ�z;�ߍ2	�Kp�d�zUU��uv̴�2$�pY���F%�p�Uj�|}�0�&���t��6���7F�N��Y����n���BZ����m��N����H��!|ǦH����mX>��V��E�C��a��#f�-��~`_�)�T��,�-�H��t  �5��r疗�?��o�)����[V�Dmm-2G��fy�����AD����寜���擕������F��'�3NT�#O�~$�M)��Lkj�|�� ,����K���W��s=�u9^������3'G�Qr2���,�"��1zk��p�FA��ݵ���c�5,]�Y��0�"�˃b�ݳ+Z�D쳩��i�#p�@��\N����[m���%_���)Aa:|(�*�9�P��)@��x���G��n��#M	�O�mvdH.�y�����
�2'���Sp�:�W�Ҁ�nCHp��Y��%#^��\�3��e%��I�c�!m�-�h�б�8�X�̵I����fGɝ���f��-��AJ]Iy|C��,�3��y3��ڹs5^3�1�7���Қ�-�[`+���)��C;Jr�~\����7h)�� K0C��n�����a I�`#!n�7�w�B�~90�Z����}q���D-?�p�*@��'�F��T�1trp�^"�[���np65WB�1�����-���Ā��,�'n����U]� >���!��8$�J ��c[������M�H���09��dDM\b�'�\<�f����)�_��`��26����_��R{�ߟ1��`\�k蘞X��{X8�4�P��l���>6&5�y�5����n*5,�z7�"�@K�)�
V��eӁ��8b��v�f@���gHeh$�gPY��2������6�a�����L�HKI�˂�y�{�I�Ǯ�Z̉��y0��բ��k�cx�������"���u��D�Rq�[�x���E�C�����ڢ9C�Kwj�l��ۚ�5�Q(�P��.Vk����t�����W�y�ɜ2Z�t��x��e�'K�' px���Ps&`���~�W�� �&���s!`� ���2V�E�xvD��؉b~:]��]��δ�	���/1R��#
aY���2��p��ū�IBkSH��ݖ���Ѷ�T���ެ#��me]똌��)6��E���/��9.��ɶ"��;u���|��C���Щ�<�ݵ�8�E��F��ȩĔ!�D�+
�* ��!����c��j��ox�?��$g� �B�á�qYB������_eI^���;���3-�U�%�F�[�ؖ��.Е�-�c���ڏ��?��3���]��n�?�/'�2�g����ώ���TĽxX�PaW�UI�[����&k��Yҏ,Cq	����&^k���2�=5��⊛�Z�L`Vl��'��W_�k*+��?	��Y;������U�Q����R�__=�5k'd�P>�H��Ax:�&���L�(;�)ɊX܋��*n��#]��V)�C�J�����Z;{��B�x�����t��������z>��5��$0-��������O~�&zThg댵��9�N�u��v4G�@9C][{zblr2߷�����А��5k�Y� ���z�`�߰�[]uC"چ�H���5�,b�D_DBt��V'�ջ�[Q�[������������3�1���D����8��u�zSݚ����ؠ�츰���ǂX��ֆ���,q� .sk��̉���_��a�@M�aGD�p�M�d2H��@@��� 0䕼 OT%�쩅K����5�$6[�@�}��ۋ�&���U&��	�!�ߋ̒��e5�e�_��������	��S�8Xª�մh��Џؓ��RҘ"��t�x�?�3�?O܃k�QC;���r��	`"�{`JFl�{UĂD�9�$�&G�T���kJ�ѿM~x�E;��Ѩ�"i��Zm������_Sf�w@!Csm��s��rL6ތ���'��>���>e@���V��w�٩u(��n�aQr�]���p�W�ƥ�l�T�SЦ�)�7�"&� ��G��3��g}Z���8�d�����]?e�|�:����3�ݹf���~��o��Һ'�i� $�KT�_��Y	ƔC eK���㓳����r҆���' 2�?5��T4�6�U�[��@Ѫ�L�v�/\U+��W���Ṽ�`l�+AX�k���'�����ڼA%O9���a "#�B����G�3c:{K�.��D^��f���o�A�'Q�#ReP�u��S���Ġn>���BD�~f��#����#q�v�v�@���]["*��E[����f./�y��S�C�z��5O��y��t-�B�?yQ���w�S'�L.:���������|HI��d#���&.�~e�V����C����e�>?{��Z������	CҿF���}\.=~*+�0څJ���zM#`�+��5��g"mo6y�s�y��f��<ׯ�}O�H�z�趸S9 B!��~4�����is�.�:�6�F2��<���i}�aU�� 7�@R�Q⟶:�V��������z�WU�:�����C	�t��T�'GTwMW���{V{��7�F��?�Βʩ,�/-���\moo�\�w}����!���2��z'����4�f�g���9�h7��[Tw���*%Z��z����I3ʮ���ꤷ�Qu�R����N���[L�������_���;u ����$F�C=�I�Zxzdw�∃���!��������Hd�$�_�y�r�R6���X7u��49�
�T�ԑ�W=>�Ə��!����1a�������ޮ��w����G���8b�nH&��w#����屭������/W��F\,��r	"���Qbԅ\�����6�7-)c��+�r�1��W��X��2K��Zd�4p�1��[�?X��Z�,���HF�������)'�U��v·����X3�$A���IXt6�1G�DL]�0�(�^�� ���0��P�`���D
5���y
J�T4?)������k��d
O7RZ�E�_EO\���m?�GI�RA`ȋ�o}���*B�A�����6]p�4E?ȓCRaڟ����ߴ��P�:�\llH��--�@\� :��#y�ʌ�H���;�GVm{����60�{���X2� L٫%��
\���	�u�״�����
@+ǿ�;�(�)^8��K �7Ĕ/���ޑz��|�<��x���z�F��TC���o��A}A����6)��6�_#�~b�e.�h �Z)-5.ʞ<�}��+��b,!�w�]Q�w��{�z�����{s��v���㲢�Ohi����u���R_�-+��U��!����=�	v6hH�躧��+oɋ�����JDy�]	t�"�z'n5�T�b�-�7��G�-�'!�|�-?�D�n�h�C����^���T���:X����%��G�Z�9������呬�+�4z47յ��n��:�Z�f���1�z��#q(�v�qR�l���}�2��깡ioi�;����m����Q�H1��؋Z�Z�l�T;����d��y���E=�!�n?�*p(�I�-�i$'��!�T���&� �m5�%plH�mi�7�0��+�����ac��b6��%�'���L�$(�G�H������J&ld/j�~�$��*c�"����j���y;���B��|гK@�\��&AG5�%�e�u@��>�q?pKPoN´�L2��7�4�&���\I6 �5e	!�~��k�k�cm���?���ZHL�����#��[󠫘T�����J�ƿ��~��6{�t5!
�/���l0V�fw3}���२��MNi�:��*&C�e}A�_[CK��AF���#������@)n��'�5��e�����i�|�ͷh���g�כ��ח���=��^fU��FՔ�\,�k[>�}-�����C����?����Ϡ�-?�J����t�'��A~�rP�%.3M���MI�:���?�A������ؠ^������q��E����I_���C�-o�f��%���`Q���;��&���0�������jj�ofF�`�iƞH��"!qyXI��;����Z��P���8k}�Pw7
��
�%�
$��iC�ߍ�
�����H�M �+�%1�1�����h���$ *{6�!2, 9JnVp�����dy.�C:1��7DH��p�f?��<�@RP 
5Δ�z�A'���YRƯ���o��l�����P���OH���=���a$2�0;�0�!G(;DR�u׽�<�ne�]X!m�gZc����"�y@��}���o�����z=���hߘ>�c����nꜤ�V��	�t��}>H����@��oj���1�E��r#(a+F�)��@�?k�6���Q�Z��`�I�U�Tqxr��D�s���{��Z �0:�k�
��!�ʈ�(>�C~&>�i��+�S��応�_�g�"������z?H�p����<����Y���=����:�l��//=�����#	�,RL#e�����`�8�1z������Q^I��|œ����񔺥��p�8����i)�E�ͮ{k�����f���ȍ=�k{~�~�����O{B��?�|!`r 0�{m�7�)��yc�uN��V\���=կ.)
�%�|�l@v������^�Sźf��)�H�R�|z�RLs�3W��;O�w�ܘA~5|ף81r�c>��?�:_���mVyM�\��T�yǈN�B1V&o3���~ny}��C�<@�Q�W��gތ̇�1G"�	��U�SѸY.�CB0�j���<�t�xڽ����u�j�8=��+Y�nś��Lx����*�[u��"[z�a�W��О �{���F�Gu���+�6УV����D����[�����!wZ5cni�Պ�I�g[":�&��
Y������8Oi������k��Z�����?ٻ��F����[~���_���
��D=�2G�
����dۥ�Ւ@O^�s6b��p�F��3%3�D�'�5Rqw?�����4��Ƒ\��E�"����s*%;��������h��5�G�&�b���\O�!8,�uW�����M}j�?$��
Ka��䂯��XK�Mw��B����u�K�||��ҵR)t,�7��L�:$ K�1Y�Cw��k����A �����?=���b�Z���;�=�ī�:Cs�Jc;	�Ӌz�	�~�Y���.#�]R�X[��!��R��EC��2֗�&�4I��t�t�������?V�=�j�1��Lt[���F=]�E��2@��׺����NLO��Y݌l�c�,U�t���ٔ:���Fb%F�J�V�u;;���J�a�8J�1T��7�umF���P��C[8A�Mb������5<mQd9%�f���ˈDɸ\A�k�9T�_J��Q� �A,5�����Ȍ�xw� A��wb0�Z	��C(�[t׭��<�N�򖀳�o���
�O g�!�sǙ��K�C���ߩ?�#�-���5L�p��(F.�s��lx2S��ϕ��=��c�Ŵ���q�ٸ��卵�/H|�#�$P,��U�{$*@�E6J~Fh��y�ؤz*��$F?�شR�D����َ���	�LA�(z��q�y����A~u*���� X\ �)��))��oxt���Wݕ��ã�J#nU}L����,bF�V|^G�i� �ȘL.t�೏�|o߁�%�	�y�������K$R�C%�r,n��Z��s�wș�ky�N�A��%��"�U�}�6'ic����?B���/����H��U�88�B���� S�&�ݫ���A�k@���w�ޱ���-HZ:�ؘ�zK��\V�( lP����cװ�ذ4xVRDF"^'����xL8L�m�ξF���V�OO��{�u��2=1'�k�v~^��O�V�����G���;2��r��
�_^e6�Toŕ��Ø{�)�/�S��)���.�z5���<���%�Ĳ��O�/�O|]Ýv���k�����|F��z�a�n�En��8�B�r p��f�#ѫ�k���tԄm/�z	�����}�&H����)�w�]�χ���/�� r��#��.<����E��ZB߳�o�R�M�;&��+FR���%]ko
JY��>�x�n�2Y�O*�$X�J>*B�:F��U����� �RC����
��k �by��z)�s������*l��acw����De�#�G�=��օW��:�!�k�%Ʃ�ă������Ӌ7�ۢͪ)����I���K�����6U���D�����R�����<�;�N��P�[{��گiխ�����a+�[��n99�aaaY����-P4�ou ����	Vi`@ضՏq�����>��^�ٍ�X�M��+I�˭Úہu�ĤTc}#DJ�l�~τ�r�k�����UGc��D�U[I4�lɏ?��Q�2?�˲B+�CcQ��u͈ȘP6������\�Hn=4Zmn�<+L]��ڨN�U?����⽹f:C|]� :D'&3��.�Ura�#��^��{�5�჆s��U�\s��I�P8	�[���*�� 4�x`H ߢ)��g�\:��F�%#�)��(I�
Pw�^��!�H�T[8�U�/LX���d"p�tm��
�����(��Q+wb�^h�*���Z�XZ;���f��'�_�	t��o����Y!IY+34�ES�xY������/L���<��Sȃ2PGo-�jo&��!	�~en0���|������ 5�%B�x��#$8wTOM�&[5�2�Р�pB~��.f�Ғ��`�c5Y&RގP�0��,��pCE����9=��(��-v�O�	�;�Y��:633&�)���ȍ�� ����Q�N�M�Oq|�O�><9G��fjJ:��.o�"�$�F���Ln|�P/�	9&n[�WR.�LkN.D����l�V�M��+<��E��$\Y�2���SF#�n.�����eI��Iϕp����9B�Z0�2�\J�\�MW���N�]��Fw��ˡbǽ�fo�\�!
����vw���v�J������2���B��o���-�**x�{9����P�y�
�C2>�}�����f�60���H�GZ�)�\I� ��v�)��i�x��TZ�G*� �F[K�Ħ�������h�����j��D��,��hV3u��{�+�y:�����LL?���Ҏ9��Rcğ��J�a�0,��U�kMDh˖�sި`��O��k�Usd����7)����h�@g���-��K�6���3�/��_�$�����X���T�]�k�y���I��Şp�;~�j� jH���#�Qh 7���l��|�S�0��� ��� �̜���U���
����r�'y�qQw���?|º�U�U^�,:�JvD�(ѧG^gJWT��RD��l�N��A��l5�֓��~��~����e����ѐZ��W�!���AAU�)5�d<^T7/
�f�ȎPH!��Ty433�^��W
 צ_=��|�����}]K�I��"��nw�B�sV^���?I��X~�z~Θ�݉'��D����Y�z�W���b�1��qp�G)6撀TzhVBx"6���6���|>����d?)�2�����B=7ya!�a{{_�[�����c}�=�]��FE
�L4�>�+
_��MÏ\�[|<��N^[]�ַ����gJe|��2�N��Ln��e?y5I~�%(SGO.4�����ߞ���_-�M�bA����CU]i�SM����ah���Ug�����o?5I�yZ1�_v��@�����)��C��]di�C0�)T!
���h��$ۍ�9x�Q�|�)7aݶAyu6mZ����-��9�-�Mz{xI3�!=��/xb�������.ıE`��[��
�i�<��jM��o0�İ���tv�^�o�����ճg|�S���X�Μ(���/�n�F��Ҍ�?�'�1�&ˁ�c
�����������XD��k��je���,��S��%%�����#jcSjɅ�.�^���H��W��u(Y2��s���&>R�@c��k�IV=N^9ȼk_|׆�\'�eZ�ڸ�
=�I���s�x6�񜿐�win��N`R���_e�r��C��w�}N�� !e�0r�c�/�Y�~���2N�x`�J����� ��<)-}Z��4�:�;mV�I  �
a�oF�������%6�%`b���<���a��ѝ\b��>S���u�Yf�Y��Fb���V��ٖ����đ��N/I��O�XH�X//�B���f�:"�w� AI��@ 9���oQ�ߒ������j�v�7����˺�����$M#|��9,%)aMt�9Y����3�2aZ��?%��	w�b��0�b�!�BX���ū���HpJ�x���i��cb���v�F���L��İ��[@�C��Q3� Cm�c�UyFx0�NB�$��s՟\Ԣ��	Y���h���}�7{�����[�;F,_<���r�Gn;��`�@�;��Q�$m0\�i�-�ȓ�~���:����P�d�N���񔺴[b�E���f�ٿ�:��o.�oR��k��\�B���j]��oޜ���]��ϕ�gﯳ������J	b�c��Ǥ�2'dPǧ�ꌾ6���~k��:6a4���q�����ԣڽF��|�V��;�������;O����M9�Yը����`�X� �mw*�F�T'�@?�����^��tƤ�r}f��<�S�O�,/4��AG�QGɷ�o���fb�3s*$z���x0+;�a���ZA"%B	��
�ᠸs�~Lk��I:���<l,�"�_��G��]!�q���揤� �r���� ن'EKD.m)�dy�N�~jH 7��Is�����\hٞ{8��=)Hu
~��H;����Ӌ�9��(�務#����`�$���=�Aa�U2(wL;���*�TT�%-�q�Đ�u�:��������d�|V�Q�p����dCV���q����|_�w��o��i�:��������7щU֛n��_hY9�����n��dm��7������K�A�B���D>#IYo_�?���G�ky��Z+��eB�4^�n��Q��6������a9G24�yR���]��UY�{��1]�@ �Al�p�)Ў|£�����wK�������r���p4{�k�����D����A1�@��>����ٝڣ���	�w�-!��$��7	+�B�>�Ts�8>�#6]@ �P J��r��v ��[	���p�'bL�F��Q�hL���1D��A/��t�x`q͞,ِ
YB����N��eJ�CB�<�_f�gS�k�`�*�Ѝ�/B���r�!-���4yd9ܸ��֥�4�fX��>�@��kJT�_�L�1x���H�;��;���9��B��7�O�@N��+k}k�أ��V	�Vp�N>׀u�>5,�rS�`���)������c�_2�`��FUQ�{���7h��k/S��� $�J$&\����䏲��b��U��~n�S3!,����?���kq]T�{����Q���wX���N�B��>#�o�
�L9��Qռ��٧x���9��?��@-�A��
��<�MK��xt��ljL)��>�,��'d��� IL�-~u+��D�0����@�2e��i�	�S�ҭ,����+;�E<~O�d_��9<8W/�m�4��Љ��4�Z�O���bw���ϣ�i�?���->΁��I�:Ū\�f#:��?5�b\w6u�(���i���8ms������7����ً�۝��z\�l�4%�4yZ��(-R�)^�%Y���%VZY�X�[�P��B�,�*��R��5;�{f �S\w�_Q�NA�z[��3���%�pژͼE�7}z7��!VEX"$,�Gn�C��ye�v�}oۿ�񧙤�F�
�Q�|ٯ����=V�+"��9�jA��[SM��[A� �tŞIA�T�ܭ�o�,�5s�9�����I�L�`$��	8����,6{�w���~0�V�����#[��7��e�Ձ>=���EB�w����DR��
���1~� V���|���H*+�)5M����tY��>������MsV.����_��T4ެ:L�ϋʐPvݺ?�a��l������5�C"$*|�@�x�'�
dM�8��o���dD�L�ϡ�KO�7�8�O�����^�}.�;����[�v��s�"4ʽ:M�j9?�[��o������e�6$�^T~�e�� &�a�~yz��O��L񝯢VYt
��Ӈ
���#�3'��p�c���G��,ᤜ6x�Ę?W"���=�}�O���c`9Ź�T�2" ��g�(��h�׹��v�6|��\vr��P)-�s(�޵af�����
z S+��}L�
a��!;���㽇KAe�4��ғ
$w��QS*-��v�%$HEƒϗY6[���(n����Q薬�:t�W:7B2,V1D�����Ӷ��0g��I���M�X�L�PD���@V��Ld��;���d�0�"K�@"g&@�q���R�~,���9��%�IC����b[��\���Bʠ�,����pXy�
S)T�%ܪH{p4۹�F+��c6�k\}?�<�͊�|�;��4�mb`n\w�S���=�R��gw��A\�p��d|�p< 7��j�
��T�k��X6L'�p�����a�.�<���1)�� |Tܸ'@��0��yb�����a4�X�#�{�Ű7��1��HJ]w,`"�ROl~G�}|��̼�޽q"o'��t}���5�Lꢲ�k*�j�VK���>4H~�$��2�̽	'�0�"(	�e�Y�=O�	xq/*���=�1�S�>y�
lT%�g y1�����!>뵂߫TD��D�5R`
ܸ_��d���_���Z�ꇾ^��F՚�aw!��Lӿ.�ZY?��]=��&���7�-����>4g��7�z�����&��V�d4���9��B�]f��b��V���8�l��ݔ��+D��?����ͩ)��BXmaqK^NaN]n9���M~��]���}�/2�LG�q�6"┟G=CZT�E d
L�Q�J�UUXu���(����܌���.W
W����%���
;xօ��U�;�@��i�1�e�_�;����);�$#��9>#��9��?5@��r��i`
 �����I���	5j�=gS��z1y�S�pK�C��P�t��[��E(
��׌�b2��I\�tB���;��٬C�lr��ؾ�p�!'d��j������
ymey��z��5��( �+ ��[���g�+�������dsd��(��C��Y�3��L�	@��hl�Q,��zcp��̱3�vgYAW�b��!h5�#�0Sݳsm�3}[���p�w n����7t쒥�,ޫ!]�o�KF#��m̷�z=ݒ����H��S��^��?��!k��3~?ϋDن���U���5��ȳ�DvzKd�>����N'dv��w����'1`Ⱦ��`���Z�0���
�������7F�aL�A��Q��=�1�kNY���Ae��#c&��&�1�K�̓��bhǍt,h5�?M�J.����	��1_ar�	��b�i���Y��^	 E���(��^�|	�=Ӵ�݄kN"���)��_m�G�ž�S�U��u�c���Gݯ%�_Fϋy2�R���-�����K���"��T�V�~E>J���%A�b$��v�qO�iN��>Wf���t�5b�C+�Pfp;N����:���q�F�J�\�`�%����O�6�ہ��#:��ƴ��4#�S�J#4a�pD΀�j�s	xeO�6 �n��\�|�P�r_���m�M��=��uC�_{ְ�����y�����?�I��%sL]�!� 0���p4�b���l��*SVC?2��0&`�0RZeo�l��T�є��e%24V���n
�l��124��?��m`W��xMg�)e(kg��+rxd��*���1�2��`��
�%�T���b�ә:��i �SJ�oFt��0��z-di�����e�2���<<C����)H*� s~���z"��3V&����OXIX	�l�;���kM\Ө�	:�n0	������}火���նjU��"��J-�˳����|c�������h6��Zw�SM����@����{���)�W�؝)m��,5i�{�[����׫�^5[���b�=x������٫_*�C_Jym�����x�py�8�
�Y�U_[�`QF�o<��u��M?-?h���֔k��`H�S[�<��GG�N�q�Jo9�^]/y����'h��fm(���9KN/���|�Y�������+�9|Ԟ�@����� >^\Y���B-.L��D�_,R�e�����UG6��!<�0�uE�<(��]�uٓ�2H��:��̀�]��F�"��?����#�����+������gT$ĂD03Rt��7uC[ި�1�=Lj	����Z�Y�&~��y�T=2�8��i��W��5B�t���Hw�K"�K�b�d���[\\�!��;]��z������l��N@oӣ�r�#;���a:��d��PD1�j�N�u�ti*�E����f����K�酵c�����`=	��弼��<$�|�db4s���] *$9&'2$�kP^a\Ce,�4/�گe�H�-R5	�3d[��, C��~&+?W���RT��&?���K���
ʈ
�ûD�ҧ�k�Cf����c�t-�m��o$+9ld�"��ub��Oϋ됯ֿ�%>`��b����Hq�|g��F?��|��B��@#�C	���f��p:�Co��
D�Q��0�^uz Q�o;�6NH3�d�+hzS �'q|��A܃��x�"#�Z�<,(�-���� !SNS̵�2��n܍�,�ְ"-�8����J�� �S���ć^��|+=��1���ir-}��.Q���+�w����Բ��FTswr�P�H�%�p���<G�����I/zi8��J�y�jM��)�����_'�m�U���g��;����A�Ǻ]�=�1�Z S�l$~&M��ݳr.�	$sdI2��c�X��x)-���ےV�%�,�~) �R?m�J�4舷��܉�t�n�t��-�"��2��̴�xH7%�����S���'Q%֡�8?����F �H5�����4/8Ӏx<���V@ �G��� kё�&���ᬪ6)i�)��A��?H��E;u��~�i%� �7�T#X)j<�]ߎ�������x�)0�5 �����[��I���_������t�4z�*S�٨�����yq���J���rt˧���$n�-Ě��F�L��G��UY�,fT>����Y�#���-���Ƣ,�Z�%X�jF66�>TW��CI�v�^{j_?��X�G����Ywww��ln����mv���o���|T�3##�~-�������4��]]��ܥ�D^����f���Ԓ�����eA�w����I!w'z���!�>��\3N���,�,��e//[�xKƂ+ y2�V������\�� ��������"A���X ��&�� �f!w�c�%��ؑ���'��Ό=�YMh�։�B:j����&,_�+�b�a
���p�s�S�g��7HFkb����8�� �b��Љ9��M:*29�#g��~�T<�sl��sDe!�]��f)|>ݑ��a��X�cw��Buܦ��)☗�HR5+����P�J�s5�[-ősՉr4�+]��7�y@��m�����~G�Mg���m2���M^7�������y�:>�ӱ�������b���R������q	qL�v�l�#�x�Rw�Ҙ��w,�A���|)ͱ"s�b9�8��7K�U�t_9���d�P�_�b�W�4�c)��'�ЩHۭ���|�E�݀�QZ��HX���h��ۥ�i���2��)lbj�N����*�rܛ�Q�_��tu��2UI�|��BPrC4�0�S=�
�7b��FbY���9Ć��!�����vA��G�b�L�Ƃ����B/pm�� �:3�.ʕ�����kZRE�8�J,z�����أ��5��A�&Nl=^�Q�# 6�����x������>;��?�,&����6�� �>�ޮC�� {i�ߙ��}�� N���N��N,��T2�P�E&yX�,�k3�C���ڦGQF�P��*� $�+ll�aX���D1r_"'8��7�?�hF�xӌDi���Zm++�L�*��O� ��J~|��t�c�mD��p�c���
G��y�_�Q�o��S%z�磲�ȩ��
R�:�H;�k%=���>���Z��]�D
�1�G�(b=�q#��;�5��N+��<��B� B�
 �ʕĝ�'S+��p�1;�ǐG\u (�<��]ԵB������{�/#�MY_��S%�泋��YϳS���k+�&~n�T�������;/6i��L�pyR�g��igjդ��/�/㤿4�k��ҭzL�FԈ����Z˗ɫO��'�;�՟�vhrm�%�̼ٚAlK̤\zKt�^e��F�9�s���$���%�{��p��+_�և���}N�\�3�>.ƻ�7����ͧG�f�:������W��V�ה�W1Z�ZR�[�=Dr4�q4B�.��D�Hi���t�Me�@�{��P�W�q	�@/ʄ����O0��	� �/n�m\D���̀ց[D�*�Jq�G��v��2S �7���bt��|��!k���(7��͇N�CVP��8�Z��d(#��Lxj�C*t7�% ]#�Nf?�tZ�|��c���
���^I��E�S�E&d�+�����Ⱥ,��ƃD����x�Mպ��0Kִ=@��	��Z�x���1�=�%�:��{���Dp���pM='ֺ{V�wɿX^^t|[�������^��~���e_�,V�N~�_�����X�
І,���2�Z�u]����HcJg��v,���~�>>s���RD�T�Ix8t�^���NM�ZdIU�m����	A�4p���/�m�@���XlY;�bt��l�Iqm1TA�tse~��On���1��.T�su��h��衳�KX�.1�;]��qs۽^=�/��������������5U}'�w=���p�*Y�Xi��{��������$чh��"-���k������~���ɠ�"}�����.��w:%6��+���ߟ��&�q�S������'~��H�E&��T��3����\����T2P����/�'�t��O��~A"Y�ғ_(�acn>ܯ��UJ"\z�|���(`�qi��	�S���Lk�i�ii��,���N�⚀cA�1X<3���o�e �'I 9J�4@���@k��k{2�YP�q����e���HX�<^��NhX:{�vCCb2�Cۀ�[�yX�J��d�
h�`*"F��*;,�X�
`Up'���1P���$D�D%��#��#`B�@ I6���=Js���V�l[M���t��ؚ�]�G�G,�!����_P��r�P����/'L!���=�Ets�*ՀGbZ����&65�R/��v/Z>*
K������4aE�t�����P|����e:>�$��NP���:�q́¨�A���mF�CI�a�lX�p�u���/��?t1տ����&,�����g�J��W�CLd%�-����7~��Z�s�wT�Px�h���R���=���f����C�nr�.�&if6¦����}zGk����,W�|�K|��;��l7�G0����:%p�m��̬;��-���sw�K���@������[���;����q�k��N��$Ll�}�ZX�C@l�޳}��C'}-���P�����*�J�`E�� :���4�ucc��1������X*{Bf��n+1���-6�`]�M�`�����?ٌF��!�y��9��B���7M��~&.��،�!�4��(���5���� ����8��,��
E�r!P�T!Hy{���?_�<Q�)���	�Gѭ~�p�tm/�}�t1�
UVr-i��Y�w�a5��̆CM͆����&����H����st3a���\��Y���l�_|^u
�*y⊗kX5�H��Veћ���1��y�W������pl�ς��Ȋ��˃�n

O'�X,��i���:n��7f2ir�z��͝1���;��t�ۤr�T�S�E���B�<~�~�4�Ǚ�d�*���ϗu�Ӥ���i�+� Bc$����`�M��R�7#bvش�-PQ0�=�)갂Kn,2s��?<7��$����)������=7ֱ�v�����:������{x=[I�/�� E���qIȵ��8��h�6'HT��"1�pT��RH?Jp�i.q���<W���7ߵ�O��q̪�����6(�wǭB��|��r��v�y^L&�Am��#����`+u��t�=�0P%�Љ����
�`ҷ� Nd�� �7z�nS̊�U��-���������h���N��A�?��|���.����;��X&��[j��:��7����2O"���I��X���'B�>��j�d�	��ܔ�.�Pbqo��x��؂����!���1�,�6�jS�vWx�ɢ�[���N��F�P���Lٽ&�t���;��|^O�Q	��1��mP����?5�l��`#���o�d�"��k��Ƣ�M��r��3�k�G������`���ܟ>�?��l���Zy{�Y���xx��	�����*L2Gu�zl�/#A򹆷���H��Ggy����� �~�v�6�Ng���W�|��D.$�wE�<��PrOf5H�C���C?��Bm�|��I�:�ɑ��^�A�c�Be�M�Gv=��,��2^X:L'z ��Ҷ��l�����`A
O�*Usz7� rJ���C_Xh���������y��2(�k����;�$f�;��2$���4�S|�K���<B��.���w�ۉJ~՘���]��bz (��Xo7t�I۱�X�t4���.��;���{�~�����7��q�I��4�giCSS1
UW����T�����l�*�/� 
U��x����o��^�HO�{���goiC	I�733�oR��OK��?|X_�[�<wr�>���r��]�S0�[Q�6�u�o4{�iY��-w�3f�.̲�ydSV����㈆>2Q6q����P��SBN�/�H�Π"��K�G����(�7��y����p��� �Fl�z�6-'��N�3�~6ʀ�Wl�'����[4�X��8w���9�&�F@�(|7��<�<�r8��8s�;A� y���X�FAh��]Bk�0V�-��J�}���w�;�/��/��ʙ�1�Ivlʕ
�9�����%О�.��jR��nA�f�C�Ȕ!,�!������ ��iP%����߶���]�EV@�z]%�ǿ�vl�k���U����~�E�x�3�u^?��T?V�6AR�}���[��o�i��S�0+ ~��C�LɒG�}XK�^I�c�!����쬀�z0����g�{ܔ�
���=�t�H\iޤ��'�סbZ��@@��~89yx�z���a��]�|q��֬��SǙ�dޙ{o��������y�,�c�G��<^5�V�&ޫ?�@rDm�~Nڂ9_�=�H�(+�����X���v~AlUB}`@�t�+�/�t\���rq=����rzq2��x�=7�WR�����'�d��|~�jo��b��ca��,������q��۟�R^nVU�
f�i.���r.�[�b3K\s���'�3�G8�Ĉo�w0[�:��<�eHF�W=QK�6�{LF�c[m�Τ�v�`W�W��&r��*��L�lq�Nw3:11a�mkkG�
�����4�`����F�S��j.���^��.��Bĥe<6g/���-�?��^�L��6¢&�[ѓ(�5�D ��z�pY�yv�y�oq�?G��9�s�����٨��������¬�Ғw�(���~Q�J�H�����|�d۟I(��O��iPZ�Hu1sbg�>CcCR��J���K���Q��Ǵ&Y��rw�o���RJ�<�<i�~��pZZ �{���o_��h�
���/O$_~�@fl9$-��C��`Ll�A��-d��i�S����=��^ X����뭂���pm܃�+R�@��V�@��
��)Z�@�"�B��;-���Kqw����f�>�ރd�	��u��Z������1�)cNMT�H��4�L�a�O�*��c1e�?��i�N���*U�f�2�5|��q~��ml�%A5um�?z�����K�r^�����n��jn�!�S,�h����*}jkaz��l"�6�����HD:�_ڝ�����o&4��]���3� "h����aWjQ�xH�x��.J4����%��60����jB���>1�)���b���q�W*d�.��u�T�Z��>���(�p��R~\��D0�����|�:��ϒ���~Bo
��s��&�TJ�%3�ޠ���Y:F/�;�TI2��|�s�{` ݇� Z/���Y�}��-5������������H�[�N�.!;��C�`���<)fp�z�m�	t���I�����|H1��U���R�3���>R�G���Q��A���ò��.k�]7�Y-����ŵx��Q��f�}�~�==;�8��W�{R[Rt�;���OJLxLp�e�z��ο'э">7����lll��
��8����@���	NN�>$"�����B��MK3[G{���u
j��d---�ؼ��Ȕ������Ԍ HDh~�Ç/))t���̼H�|_MՃ�L�1O��;ql]�����p�Fwěp�/Q�8Z�;�M��|�Y&�ױ��L�}�! ���)�_����3���y�4񇰨�y|O���$���[jE��w���xy�bh<`'%^^ ��{�g���I6P�v��C���%��h���h��ݩ��;�`M�~N��_ #p��ɡ��5#I@RV�NF �ƒR ,Y��_�1��:�ap���a��>k�����p��N,9��[��y�O9���4�J�T]>'����FXAq�A�i&�6aD��S�j ?�?99Y-K����7�O\O/�˩���9�l��Ҥ}cv��Z�����[s���缏�d���q� );&~wךc�jg��S�H�c���~�؁�H��~h)��bIQA����\o�.�[O�t%<%���Ռ6g\867�<��������NԴލ�e0��ߛoֶ�=T�,��q��l�i�8�q���c%�+�1K�����N�P�g�פR����ڈ���$�u�e川�PwJ>�CV0@�����^�/kɊm�m�g%�V�6c!J@�[�{U?���EJ~��iU�J<&a����s�_�sU�B�4X���mTv!�R��M�a��L���J���"�`��x@����]��Ah7��|����ք�M�ˤ痾B���NV�4<�-`@9*6U~қ���"�������?pJ`@(|�T����)���D���������y�(��L��9%E�e�6L�����74*�,���'��T�	N7���r�	�m��R�1�_T����	���ǡ]�Ya��a�{��m�}O n�$�:��U�菎��NQێta�$�մ��S{�[�I��-���'�M3�t�W4�j9���*�c��g	X#B�����!�E	��Ǖ���o7&�H�A���^��P��JkapWyCd0��̶��| ��)F:��R0&)Xf�i�s��N>�D��K������]+��pC"p:�E�S��A~�a�ER�	�L7R�I7�#��n��A��zy���Ɉo{��-�["<�D��|H����	]Q���}�]�54�S�s����QņI&Ԏ���լ� v���:�3�Q!��2��̙}yū��'wŐ��s��>;Cjn\�q`�*�3~�M�����8�ח�>^>�B�"3�s�3z7���WWW��>��o疖gPA#��-\����tY��뫦�fE%�������n�8��ナ8dLA�Ar�����6G	<��q�~|��Y��s(��T:p��cEC�(�����u��r�����2��-�s�U�mT6��\Ԇ�/���.s�F�_�c��x����M;�E�1���4�yr�[������lɽG��؁Ls�JSJᲦ�o+}�nXE��5e�������3/���Ϫ$L��4{�IR���
a��o1K��x��"J��)ޏ�i�'��Guz���79�ϫ�������Bɡr����qA�����,���OKz_i�.))UԍZ������bW���&���S�n`��~�p7�q]]'s<�����A�uٕ%���3��"�L�c�;v/�2k��~^o�|�.��NIޮ�N=`����_@\����ׇ�����Ms����g���*�u������wv�k&S�p������1�����I���Ew�-����@�����I�6�w��Hb��Iµ����T�0'X�89������I�2v'O=·�WP���(%�~��E��a'���4/�g {��ļ$7H@BX�������~�ڞ7�U<s���`*��khk��W��C��f*���~Ϩ�z�NW�N���l���f
��}��d<o����e��>�_���e�Ύ��[�#���mk�L�U }0�<�9��O��dw(p�[|�8-s��{�R>���̓�0\)��C��U,<�9���4�$��)��G�� �,A�+G�`�ؒ�D[��"�`�!˛C�oo�����K߅�߰gnE�����|�o�̲�4�~��W������P��BKjz��]��`a?Y�A�YG�Y�*?*�+"�m��-�Zp���\Y����r��@U�dДǿy���-5��ç�׏��7o�AUB^�&�$?�(���� ��7�(�z~/7�����-9$�3#9���S������:/f��hA�6�Pʁ>���3A���͋4����7�0��Ƞ�� �@�^Q�S���T��?���|Vة�&3X�8B�0�$�Άa��M$�cV}��-�����*2�%�|^��Z*��Z`a�n��l���b����HZ8��|�Q��6��2�y� D��yO��f�VQU^SM6��tW�z*+C</1��Y��~������~~t�􃃃�`:>r/|,eee[[[v_5AO��/hKh�u=#u�R��ʢ	�?�hP��KRH&���XR_y��Q���,��R�ԼO��o��I�8�&�����e?<bY�Sēr�F����D�&kت�]"^1+����"5�"X.ܔ��y�Ư��fw��p�6��/����F2Y�M<�C�-��Ik#0kOd�l�E~�H�1�c6s�sP��Y�~����,I����.�ۨ�)u�� ��TW�^�W�O/8�jX!�k3�v`��45q;����`<�����B����F �^�xA'��3j�rAL'V�����|w��젦�1{�b�P��� G�9�[���EWC{dRsbBCpD�չ����ȣ�ĭM�/k|UF�8X|<K���H;4���� ��;:�|��.���6g��7ɡw�9�7�ws�ͮs$����϶�e '�?���Қ넄�f�FG!O�Wq(#��)-�Uk����f��n�����uʟAñ�O\�(�ik�䀄d$~!4ko�y����&w�9I^)�;��$��8�UAၵ-;��w]ݦ�%hb³�
����%?)�,�R+m5����0Dz�vCgpp��2�5����h�f.�����|�cNS�-R���,��'.���Cԥg/g����A̘���Ep�;A�s�D'����yp��R߽hL���>��|,���\Ǧ޺�%��7��g�!�<E2���,�4q,��i�
8���3\�P��$��gឨm�4Kq�n�Uh��M����i�k�M��@P����׷����SX�UV�Q��\���<H>�x�L	wG>xPZ����R �r)�����8���%�����M��S��oIʗqrv"K~��rAa��jy�z���^P��K?�և�z��eG?��4����@ tc�� ��V�1�3�hxF1 ���� W&�|�ȍ{6�$���ex���&~�
2��^TA� E}J 4�-^��2��������yP��V��&F%L��J��0��[j��*�K���`K!c�0e{��~�/�u1ut���9GY�a���N�&��RF��R2�u��
c�Շ�-�'*(�Bs�%`�Aa��M�8b��O��
R��rrrZ[%["BCe�����Q)k���'4...+++QQQ/*<9iWBk/��lq������ʲ���"�[S3*c�j�_�ֻm���Ia�U=�C�y���v�[��<%v� &�&ѷ��@�JNd�ҝ�J���M�Y���WPxL��B�Qm6�(#śay�oo��6�&�^K~���?��P�����˵�O ^�p�pԧvրJ8��g���HH���K"��9�;�t(Z@������}_
� �4Y2��l��wJ�eЭ�C��Ղ(�N�>���x�����ڂ�o��{3-����9(�l[�HT����,������ѧB�D�����,�G��;���Yݰ܁Z�|Mt�M�9�lS��5������U������nvG������9��s�:������۽�.k�����'�wZ���ٲ-��͎��kGG_qP�uP��5;��Z�C������/Mx���9@������`��KQ|<������O�d�
Μ��t�5��s�4��2����l�f��:8oߎw���h�dvw���-�
�! !� k��H��\m~�L��A��P�p~	Qj�v&�
�mH������2�����$�����)o��-t��]�:�1��<�@`�v=�P�0��he	6)��1F��-Q�?�񪎷_p�^^��"D$oYe�v�gDР�+>��g0��J���3�T�+0Z̻�@�U�T�y:sA��G!�����'TU��ٮ���f%A�Q�)}�5�����R29����вR��J[�F/O�>�e�)1�v��C��d�eMI�T�$�Lg:��l�*l����_P��L�Y��>���J�`��������Ei_H;�m�⍍)�|;µ�HI=ln1[R��g����$C{akr���-�����ːN�N��/s=Xh(�,��'ʘL������x���"խV8�����n"��;�N�Q�"�C&8��N�G������N{�_d�]gc�Z�~�[.��4�@ifD����������VG�u��
�����mx�3�/�;���*��u�IԱk�x~�X�|�a���BSs����hhX���\XD.�����;{aUUUA+�6����P��蘘PE.5OO]��	�?�RF��y�t��<u�o�� �K�k�?K�p/�Ŀ��~ZI�1|��s=�����Q�7u�!��e�{�pQԚ�v��ڬ6-ڇ
��5��~i�+[L"8�}�w���k4㚯���� $�x��	�|n&.PB�VޡG����T��Ӕ�D�'���}�����Z8Q��ԙ��ǫ;�x%�^����0�
J�#��Kh�bc���P��X�'�9bַ\d�� ��Ph�&R/��A�]�!Q�%4�����[l��Z��ٟm���Z��%����{��E�����¸W/�55$J��\7�����ݷ�0��h�#�P:��:����i�6��y��]���D^��60<���i��.l�;�{�X؇����J֟�E��N^�9~�?~t�!լ,�,���}�c��h�J2YC*���$�/eV����I ��gqPgp��ʻ�#�ȡx��q���.��J��j�ö�ի�Y,��_�%tҏ��9���ޔ��� ��s��i�9��n��W�7*	��(SG�R�P��F�x��J�˗�s4�+Ͷ �W�^�%3�\��* q2�N��o�x$�1�Wel�|�>��^5�:ً0���l9�u��FV���rFƹ��#�z�_f�&!�!��DP9+�V�K��=�Zh�����x����V7@󫿘#R�۔�Ž��W�$����	�A�?�>�N�W��Kvi��,����]��Q|��@lo�����u$��`��l^�̀S۫���l��h0`���֖!EՌ!-��A
2ٸ�m����CD����W��9k�'�!���xv}�>�A������+"wq�{�*.����ȵ%R���ݠ�ə-��4WU'ś�������X� �g{.bKö#��ԁ-b�N��Z��8���0|b�(��t�uk����<�� ��Z��7O�$�>B�zA�|�[��k�F:�g9�˃��JO\h�Hr��e��n�=%�2H"B7�ǭ�����JV�CA~kn��0�������u7|�g�{DIڵ��� � EC�"�t�^uҿI0=U#1F��a��y0��ܵVa8Q�o�a�JY�]k��� uNږu��:��H�-����f�~������/�W�l������"��������mu�uX�[Q�Ƣ���������a�����C���W�?NN 33�_ss��!��B�.����5D'^��� Rg��s�z�X��~�+T��}�&EF�*~�G[��g�S�*zB-���B�Oyv�����c���
�M���Bv&��M C���c�(jr8=2߻ ��a�a!�d�[M-}{S�aA���������5�&�"��gFh֍�/A�$�:��([��+�=d���T7�������	3eB�^�X�޳��M�_y��bq	�|yʦx�u+́t
�rOL��Qa���yv]1��؝�[����M7�ύd��qd/6�f����P�).͵��<t����t*_���7�H̏v����`�_?.�i��-~�Wj��+w��'�(��m1�]��ߜG�.��-��]�:b=Ꞩq�/J��n���\�/>�ӹ���%��������X^Y��ۜ��jz�c@�t�Vq��wt��ȑ��0=3+������Y̔�U1�_|�#�Ȩv�j3�ϠZ*�w�0��Wr~����Hìȿ�WQ�����m�jK������2��?�����r�Őě�tWn�W��\pz)�
b��{^p:m������&�=�M���Z��f_�[��`Mm��L ԝ��눢7q��b��e!\PJ�Y�rN"�g��A���T�z�OC�����Hs�|v�U�)BA�������&29�y����1���a3x����H�
�}��v�sP�NHN4r�Gm�{�P5�|�S2���L[�N��Ag���W��Ю	S�j2�j���QT�z�C1KSe��d�%���rڇ�` �v���iw�A;�KC��&���:D���]C e	�i�����o':��c!y���p�zaM�|.3	���'����.���5�& E���A��	DG,*�����	x�"#���7��3�[讳%��1F�����P�W�i��/�,U'M� /ݕ�N�E�&N��8S��g�q��J��y�s����P�*�ǙK|D�
Q\2ֹ��8iT!�G4����@F��x�m���������:N�s9�
�����X8��п��j�, ��	�S`듬[PkT�C.2"6>INӼM�S��JY��b��o����NS)��5'���������z{{�Gҿ|A�]yJNN�����a���hj����㢥�M�G�����Q�kr�¿
!�CL/Zg��L`��dX�=�_���xջ'��x��HR{�V�f�!�W� �[	�S�dΆ�yRrۦ���a.��[�\<�#B�6��23i���!�J�IAPW���?��YK�#7~���ߏ�|��U����F|��U� �ӣR1	��6�az��/�^oC����)�0Δ����������Y+�k�q�O���l����|�����|15���8��8����:n�LҼ}�8݉��Yd�0�����O�+�I��Ǹ$��~�z���O�9OǙ�;Da`�p�^��R6�qD<cRȖ����Ƥ������ٿ��$�Ar��n�����Ȍ[@�m��p��\��e����������LD�Ҽ������O����ɈÀ���}��É�Z�����ՋV�����T��7�q~�vݭ�;C���˄�H�����Õ��4��0 �V�����/��ɤ�i�_ �m|J4ql6P�Ǖ!�G!�B)|��t��G�YAaYn^��12���~6��Y*G)��-�}�=L����L��JiiIe���#G����_0���:�vCj�m��VT��ݙ_'�����W��lf8��A�]?���/��xg�R6��=��D�ʄL���Tr�@?��X�IZ.N]���
��T�7���e嵍񘳪�Q
�G�.��ͪ-u�`��P�'�β��F�h��o8뵤<�Xo�վ
d\�|шjƈjBu�҇�g(x}�0�%>����凣��ls�l�C�z��טU�}�iЪ,Y��AdR	�e_��a���"���b��r����|�~K�ZD�O�BgR�������-����:gMĶYыX��z_4�%�v6���r�a�����y�|��+EO��'�O)��(��|K��HW:����[������#A��,F�14PƳ�b9.����Pʿ�#\��5�6��e�PcQr���R��[�� Tm���H`���|wq� `��FLi���\�݅zNw�~+FՆA�q@چ�a�4��B�a����|��*~�K�yB�7��F��5�d��o��&�\�ie�fdx��ns���5�5�D6	&O��[�L�
quGR{]҃,�M��]�U�;��[{���S=e �l�YZ���F�F�&�B$�bcb��s��>�NNN�����wt`܇S�a��s]��mk���R�e��a	��ކv�L�Y�f���4�oC��p��Q�\�����_4�q�)R��к��\xa�+R.s��0�iP�QC�0g��#y0��9�����C�BS,�yZ�Κ##�%��z��2�& <��}%�����r����O�QHY��,&�]ַ��Ԕ���fs��Z��U�\��bZ�����I9Ll�����*���T�� �##
:�Mf�ج��m���	(�_�cMZ��χ:h�Ժ,��Cz�O�9��Y������,��K�.6?��niCwZ�4�q�)/����$���+��&(V.�i�$��~�}�q�'.gK2�b5�<�:<��N7L��t�
t�Y!c/� e�g됿|�����\)��޴����D�/�v�%�+߅'�״S���������oi�>$����˗ꐜ��x��I�^��1}=f~�M���:�5��d��k�~�Ϡ�n+�~]��Dr��l��Ů��jdP����̭��'�v6֠���_s�s�����q�ɋ������ŇF	��x��R:�������6�O
�<�®e�n�毮o����E��ϖ�Oo�%.Nl��p�9T�U�<<��Ȕ��4ÕH���>Kӯ#s>���C���6?�s���_	�@p��Z�b���N��_d����w�#�һ�>ty.Ȕ���R�!3R��.~l�aų��uƝ?���\��8"�b�����Q�p������X��ↂo�
��<�Q�!7�o��#*,�Ё�CYӢ�GǄ\5����������n���i�rGI����ɧ�^��{s$�"(����yyy�b���()�^\P��cAiߨ�����>��Z�ї�x��0�5=t�Ǡl�)q��_�󶌲euYϐk��7E�^%$���1���/l��eg��E��C�1��G�X}��c�U_��<94�V����F�*��ЭG*~�-q�Q#(��Q}���*JW󥝃�P��3Sf�l�rb���k�>�eps����z�a�����k*�hB�o�L�-<��<~��BOa�>�����7��P��w�A��]�VN�UN���,X��L_Z��_�l/�"Ǽ2�<ǉ��g;�@��"���S�>��2�V�Z�׃8��y'x��Z�!|SO��(�(�*5 '�T�
0��&f��x�؟�R<a;�x��~0�4a �G�15.ӯ>�.(��F��u[�-�{:���l#�c��Y�c5����-�ipN��|+F�U���
��Z���j��0�M�5t�!�f�B�)&+��j��M�<��"�2�C�q"XF�ylՐKeD�X>7_�X_�X���H2^0X.�h���b��T����"��
~X:��3�!�L��W�O=4�0�>�����I؝x��'Q>�Ӧ�����d�א}����6�_��H#��b���YնS���Qg[����k��u}�R��
�F�K�����d�GdA����L�-�o��Z�%����[ZZ$n7��L���3l�P�Ȑ��wp@j�G��yqvt|r�����h��=9ߧ7%���K��j��1��Թ���y���Og�j��뮝y6���L��ʰ�I�	�����)�۱��^�\X���N��ҁ�A���f4�R��m��/ �|�x���sn >���Kz��J|�ޗ������s�}D���`�^F6XD�	a"0���ŕ���Ks�*�r|�Gw��wK�]}��-0��h
Z��e�F�'K�d��������:xxQ�6�g
�v�S��a����%}x%x��)OYC�e����~�����Ǹ���nkʢ7�+��u�q��VUِ���9;�I�e�x5кDΐ�k�f�{�#��Ȯ�k� �,�$�_������$畜f&w�f���zw��Q�9�hhP���'G�.Z����~75�$����������v�a��vB�v��� ��Kr"��)x�xW��r������?W��"�K����S�W���-���<�盯V�|�����VY0�����,��9�	�t_	#>;;�!�Y��T#�i- ��UJv?Bd��M� ��֘�׎Z�:�u�ܡ��LS�G�}�8�!}�+%%+�7$�����*����j��$o׏�pż�rH�>�!�(��&��Փ*�V�/C��S�*��ۻ�Jކ���c�¯��������H����(h�Lhn�az�~n�Gt�q�q������
����Z�)��
��AW�s��~�MH'�V^�H,u��2��3����^��c56xP?n_�\���#�~�+�oR!�]:\�w�ܠ��3j
��Q�\D:��,���utH����棕Y���Y�#����O?�����݁�����A�L�ˏpK�W��Y�[x{1���d�	�L��H_�>W��t��x��d`A=�|&e%D�f���ȡ�i�U�y=H��g��F��o�63A2	�fx��}� �O��M%I���:~�Lb\�!�"�!ŭ`ӠH�5s����4��h?
�V���C�����%}�<�$�?n#~`D��	/�~3V��M� ���Y�.��y��H~�ne� �E�PK�/�C�M��)92�0>����n���������h�i���}qqqhh��SS��	J!b>��9}�ו_�tu�S�g;��,:�f�
L��4@���#���Fr\>�=�VFuRo�h�_�ȶmZG��E]�Mc���/q{�Y���k���#�t,�����O�5��G�w�e�b�˨c�և��-�R/x����d�W�%��&$���#Cq>�����K WΈ�!��X(�\��cB�v>���ۀF��`��e�˹��՘�2t]/�!��d�F�S�s���H3���h�4��h3运n��@;n�����3M�*�u�@#0' 䮝RY��%켊�%U���l�Pc���]
$�o"
K�"����/��U]u���1�Ӊ�q��ۇj^��d(�:�s�׹��H>TJ^o�oO���������������kƇ�T�!������W���~Ke�<w$�'���g�����[3w�⋾M� Q�P�k:����6�"8�wX�x�+�{nA����}.[`i=^i�)K�Z
�瀿.��}Ґ5k[9n���� Y�}��0��Л�sbʯ���q5��*����e��.Е��c�C��S�b���۝
���ra	+��D��%r��c��u�d���ܶ�B$/C��@��wK��\�1`999c�l�����gF{��G����/,�3��e���t��}�$��=G��L�^�34��:�#W��g�!r�z���L*�>s ���
�� �?3�5�!,Q�+�"$�y���_��}��4U�P��?M����R�@'�h��h��-��|,����]K/��]Ć������_�C0��\�ƚ���M�A������ot^d@*E������J'߼ۇ���^���<>���
F��1>���b�c�܁�����pD���|M����u]5�����d�8�|�@�&rYT�,��I��$AIQp���5%J��"�$7�	����MPOF2/�C�t��}fC�>��3�o��B4�nS���4֪�L�+_�!!(�4��ovԈ��ZOy���%4���H5s��$�3�S^���P��9������:���Ox��K��stl\l{%����u�l�����������***...���JP%`���w���AE��>���˴ӂ:�=_��E]�$�������Ⱦ4*�;��<(��eP)��0�8׭>'g�/����<!wSRd��|r)�im�B���kOő>lҹ��:�I̈��T��b�Mb�9A٠��AD�T:��$����ޟt���c���z�u1��ki�]������|�Η�{����W- '�]��/yA��-�d�Y��&�o��$-\�>J"�w�~'w�1��pױ��pR
�Sᡛpp��]���/e�o�/o�.���>�	�~7J�ƅ�>gk{� �[���?��^6{F���բ/�j�Pi�w{�5��-#�j����o����^���f7	��Yo�v���^�<lZ=���/ݝ���^�b��K��C��ևcr���w>\�>D%��%��Q���gj(��_h}��l���s!���`)�`�����@���],	�鹫g�pU�t��iS��>g�Jl�;4����	?�{�I-�c5��V��o��D�/0 E��Ú���ɤ+t����\gq��8:,���L-��nQM���x��7ܭ��4ef<���_�^4���P��A|�K�r��L]�^�|uTU|:<�w�edd|}}}>:;�x��x���T�*���T��W�&i��B���3���?��1�Ė�Eŧ����2�������H�H���{���� �f��� G�)�6���i�@��
�b���R(S��n~�~4�},E)���6�(~ߨ�,bT-�Gа�_�׻��#h��i���|�d_�܏�%8�i=vӿu�%��{���2�|bE�J���2��$�jM�����^P	�B]q;SBI��i[i����	�4FU�����+Ӯ2�n}�^��ZMJg!I	���8~����p
��(����LP�Wi�?��.��Y�m�Y"����>�	���m�UR�։$���EvO�6*�ܬN?���t�1\�1ٗ9۱�XR��[�W5[�y�^�,��^0�U0}�U7}����'��߿iii�����ɨ 3??��ѱ���
=H��-�r]@__�@_o� \��C����ӔJ��Ԛ,�)=�u���𼖼"V���Q�������X���I����}�Xܟ��ACH�H!���Lw����و894��o�<�dF�`>���Y���鄿m�a��f���	��%���]��,}�0�]~�"�bJG���<o�hԂ�qj�KL���rxs�UO�aqm���뺐-��--.�����i�lQx/K���\����b��p�BdYeWai[����R��NF�A���Ľ�	����S�dq��}屼^�!F���v���*gԚJ�O�}�/��N:��k��p4���ѮE����V_R��u4���4d�N���'f�I<k[��Z/׌o'r~H>4���~��*:�f*��~3��O��U����q�]|�E�������������������l�r|�(������j����R�ޓh���<��:�1�w]}8l5,�J2�ިK�$��6�4���&;�#���OX0���H�8�-['O��� �F�D��c��q���"�+*kj˹y���N%/^.�4���*��

�-�-���w6^d�y]��^�[#��w���CH��
����͘���DD����0H�j;��������;Su� r k+�{{�{;v4���+�Tk�Tèsi�~���:��;:�≠ږ1r�8C;�x�<�����t�����]&0\}���!���D�z8�0�D�&�V�c�_!��n��$�w�d�)+�NᏯl������ |����|��-¢M�.�����9Z��08N�澦8�-��2眪�ј�9B�ɘ��q�ӇZ��^o���?�H\Eȿ�j?��7���h	U7it��"v6^��`:�\���?�~�ʠ�1s��* +�b��28�O�!����t`B�	j���~yj�B�)�'�)'�'?�b�����k������r
��Í��w'Hձ����L��)A�)�$ivEJ��T���zO�uf(G�)����j�����Qt9�WǢ�S�Z��:�Z�_)����(S(()�n>]���H��urr�������C�������[UiiiS������ׄPk��_�
M��dKf��<<��� �ĀS��ڪ��%�%��_��;��Y96������O`LsJW���eLܭd��V���1*��y�ۯY���U��]`����A�l�����2�K��?���P~t��s>z �{���&*���}R��������z��q�j�e��Ȏ��*��a�iߞ�<&���	�����\߃�u�7���_�œL�\	�1�tA�?o�t
᭙ƪu=��m����ZU����PugM';���Rґ$�g�K��
�k�F�R
�
�2`#9�����WV���VuraK��ǋ7�����-��(u:�X
�ڥ��ǥ5ࢢb�%e,���	�O�ļٱ��sWw�LH�`**R�:�܏�܍N^�^�e��s��3|�k|;��r�bP���M�m����mD��Z뭕�]/���V�i��m��]���U����X������.2�G{����'|Ox�䳄��g�7��%�����j>M��&��3��$�Y�-e
"�p1���M�we��>~D����ɬ�:0ݑ�����P� ����z�h��32��PWUیR�kcBsNCCa���(��0���|�;jV�H|3ĥ���9:���}M�B�xПs�h��&��	�oll��k��Q�S�M͏-K�tO+�I�5*�7��1
��B���cT���aGR��/���H�P:����'���p�)����^ HȧT��%���Wܗ� oa��،��H�O6�J�����!}OzkZ�؇	�f�z�=ͳ1ٍ��U����)������+��3*;ku�+s�(���V?�o�+����1�+���a�%J凢:-c�AsO0e�7�`�f��� �ߙY�m<�6F*NJE�A^uy"��:��Des(�xA?n_7�P� ��k�KmC����q�4���2��'���̠�^�0$I/m4�A�p���^�bȎ0A��?�|��r�.R����k����L�nw��Q�)��D�� 1t:=#I�"^�*6˪7�ul-eb��%�R�:�Y3��3����^�*�����u���f؞������Ί���&�R��===I��UQ
4<\VZjogWRVV��gMU���njjjmu�Q��ʱQ��$�ׯ���V�����фܣ_	����:�¯��ݍ�:�A:�Ae\}�jQ�'ε���S um!�g����FD�F��ՠ�	�b�����woR[�$FCa��Zո��>��/�
�e-~��$h�+`�p�	���,�'�y��̯b�)�r�����
8�A��d�˞��Š��tV���%�M@7����P��������OM�&��'�G��bO�=q�=ʤ]sE
�x�t�6�(��o�e���;����Vp����a>
�>��ޡ7����7��>"���4Z�ޤ������D�Q+�t�цl�����W�����3I��s�֢��z�����\��Q������Q��~ў��"�EB������|�b��;��a�I��-��GS��kj9�����ng\ޏ�KxVr�ܟH^�r=��^�P���2~�;:%�s��z{�+y�w&�T�f��~�Cݾ-ͮȒ�O^A�7�a��I������f�+$�b,q)A�}�[�<4�.-�f�(n)7��g8�E	���g�*z�-a�@*v+K�!|�E_��76�!�ff�����6ގ�Vf�[�:E�����j�Or�Oy�=�v&+�k^�� �
ꊬI�t1��
Ue�u)�Kr�rra�@]]]��<nT�ٰ�ق���2����mqJ�b��Np���w.�݋��@pwh�	����E
����{����0��L&����{=k'���,x�q���.�!�U�~c[�ʚo�pC-�S��/�Č�T���Q�Y�֓�Ķq���N��2a�#P E8��z�ϲ�"�.ʮf�kMj�NHT!`V��&�]~[�(��e1{�;x�;�4�u���u�9�]jnO:�jw�XQC�[�~�����+��4
uU��˗sYV�?v��F�hW$f�7��p�}V'��/���4��$���4�E�5Dx��b�tg�]��3�<��N-�5�sN�r�^�{�j�\�n�
��4�U��?]�B��ab?�3�x���q/T��|���W�~����I�� x4Ej���&�c#�a��>�`�X��﬊h��ˏ�E��M�Ւ��J�e0�R�g�s�4�"��4���iv,�������|�A��tu�������=�o3|���|K�G��1�Ɗ0n�nlk�z���<=>;��CiP�ݼ��:�b��։�)�O������fW{��g������������[��Քl*��q�+���ݔl�lq��zDT�G��%�0�ݰ�&<�0%�Tڐ_Z�Z�;���Zm!��ۇ#������Y�Uy��l������}�����"�x���צ�Cʀ�6�ڼ=���e��K#�����Of�����5 1z�s���0����׊U�auw���h`�s��>ʄLVg�kmi�V=T��dFXk��9
#�������E0!R��M��J���J+�J+�N!<�&ߤ|������������������������bcaabS�TPY]\XXZS�>x(9\��|���@qH�+Pn'��3Q�j����J
t��h��nA_���]#������u�����W;�D�X�U���K�����������F�����x�9�^��>��.N�;���;��/z7�����r�����G�xg����׾��˗?����?�JZ���8�%�[�9�e�f�w�P^���?n*����Ȅ&�-x�"00�����˗j��/u��$/3�M�G��}���G��I}@�آ#IQR����m��Wg9{���:��l�� u �6
��_����C�Z'�V�*v����9�K=�W�S[j���)/�ވ<������~�?>[n��ڝ�L�&!���.)y78�MN�]P���&���_��@�
���̌��uy�.r`;�4_9�]���97�ti}y�u�w�w�s���O�u��]�͟L��H$���� q�i��N��v�.тd�`�6�<O�����2RD����h^�\�(z���	!/@O�2�*�G��$=iNKt��T�Yu&yu#�!3�	�Mh������<���]�-ı���j1�'2{��|'UU���LLTש�U��W$+�xB���}6�Fpm彫x�⛛2�qw}E��J;�I������q�:��aW�L����LnC�0�	 W��B6H=��r�nÇ�D3/4s���8D����Y.�>��k��c!٨���!�k�[�j+�DU��Չ��.uf:�A�lV�"�]�u�mZF����!�����rx�.�傠����"M�Ve.VʉLVO�,ɴU��v�ԇU�3d&�Y�T�	�sI:UI����ц�W��%�65��-)�Ҭ��D�e�;��\��Z|� ���s�4�	�|���4Vuf`Vշ.2`9��'!׬�Е\>��[qA^{	d��`��Pߟ�8��?5 �x���J�����h�*�KZXK���9(����\��ZY��:Ny(S;8���=�3~�iL����{:Wm���1_=ѩQu:[^���f}M�������i��KgCG������;̱q~n���J��9=LD_L:4�?���}@_Y1tp�VaC��7?�Y������hj��N%-}�-��]ۢ>��67���C|�����p\nQ���f����q ������r
U6~P��v�h�9)2��S_��R�hs|_�����$�Wb$[�j�ʮ�Z�����f�!Q,9����,�wٹj�6��o>NW�Z�vXl�v;�t�츠��#��H7l��Kx�WJ����7p�;�E4*�yb
�!%���:��T3����H��i��go-J�����]9��{w3�5�طӧFL�XmY;���!Y��$L��#kZ���/K�K>�4�a�hR�%�-���-t�3QD���/��҅=��/Yk�;E�\CE����SW������^Kb.ZVoOБ¬ª~y�j������&B�B�퓴�@f����:�<Z줧k��`z4,��x�
��L{����q2��_˫��w�Pß�ã�j�3D0��)�����	�Y�
u��J��)&���j�����z2�.��n`mii%��wۣ��������Φx
��ӓ�������"""::`��y��/^i}��]�g��J
�5���0�:�9[?:!"� &"IǧJ"~�FB����2�� �����{鈜_G�@�p>�Ć��z�w}pwy�m��������Z�M������������#���
��zl��綯k��纄�Z ���Kk5~ya;'ό��������a�8zZ�
^
&
u�Ή�_�2�:+c�(^?�뷢"��&#���-x�̂O�%��W�MȋBڥ�U���:������\�]Dى�=��S���M�\�v��D������v�?�_�Λ��]�\hg�ɰzW�[k`X�i���gw�{��|�F<���bB<������P������Ǘ����֖>�û�ۛ�KKv�����g=�1L��;�a���dĂ����;WNpS��j\cnsd(�(��%�>��H&9��Yr������M<����6����ߞ�b9����U}|�bϛ��>�2��yc�ZE�݈@Y��c.��x( ����iI_}>}�}fo����uT��c;�}�6���.-}K�T,���(*��nY7+�I������&}��#��'��c9�OKP(a���?��OQ�� ��A���g_V9?�
"�]Fz[|�e���P��XIq�K�{�}4ԛ�rn>P���C�v������^G���~�^?^�+�|޻9܀Gy[,��2�#��c�A{c}Cw�3�t�Hm-Ѽ6).�$~���mpyـ�Ѿ�U#ɻ_�	�ն�/�"������6����tR9At���1�C~-`0��H�p�H*d��q
�!9{
�8*#0��mR��bw�9��"�� ]���
�q:�n9��,]EDh(�9��1�,�=W�~N巄L�/JyO�9f���pS�HcsQn�����6,����hۭ�D�h����q(�:8�pWb3L���$�~)H#R�ߧ+��3'$��oh�N�֞s�M����*�C�/\�yT��������W�=R��X�T�������e�_]X��uڛ����ܐW{8F��(~��+U��2�"�7Z\m�=g��r�+���g��7�����7QE����s���Q?i�p�G���v�/�;�Ҙ�QuIY%����ӧ���|���Z�ˮ�#'��=�%���R�k�&*��8T�5�4Od���Ok����N:O�Ί9�kBW���x���5>L�rYbXz=�z=�]�)��������� c�ɂ�=����=���],.������	�[Pd��ؾʋ�ʄ�2I��m�eC�f[�����[��I{ޔ2����Q���ԪD1�EAy��=� L�)x�E�erO9�mR7o`�*;�(��Hp~	���ي]&48y��(q�h��>�wW��r������{WG?����`��W�{';��X�c���9*;�@#''�+�䜜����o���/k���1�"gA����������L���ۿݯ�\������{��U�j�j�����S����%�&>6����|N�+�=��nN�Ns�:[�N�� ��I��t
�/}����%o�K�?����a�+�#�-JH�-���m�?'��u��X��d��th�) ����d��4���7�Ǒ.�G#��c�T���� �q���dۻ��g'3���>.Q�@rch���� ���߈���N�?���:5D����� ����ᙛ��������k�OO�d���g�c��- �nR�D�Jԙ@R+�MЉA?��ӄ�әC����ڣ�Y@�$�.���=�--�w�\�����N�Ј,� �ܳ3�� L䛎����eyJ����v�c���π���J����	���>�/���>��>�h�F!\�
����������T�/g�r����C $ߘ��S�"c�3j�N;����]-���}�?�>���	Y ��yA�����W�:[C^ARy��GLS�\-� ���#G�
�H�װ���Z��~�x��a���B�B�1."��L�Hc�Q ����{��Y]�^1j1�b0��bmgW�%��y�f"G���a!^}b<&2
e�J:���%*��n����E7W�{�s<ȏ��
u#�pܸX�I�#|�V{�s�%t����A\V$P�K��Q�Od�I�� b�E7�������V��;��Ɔ�o"���l�b��������������>��X����e���Q�����������K��\]Z�篭^��?y5�<����I�[�����]�0u���<�͐�󖔺9�W���}�M�t���������S�,R��������1�Lcv�� +�����7����!�2i��V��[��-=5Eu�lbt���E�Mc�������<`dMt���¹D�re���t���-�T����U�`0L��P��Ԙ�A��\���c�W�?�KYż�5�/o�i�	EW��.�c&9����O�x��w���߉�����}Mе����'�XR6�b�Ͼ=�.�,.ā���҅����z-�ӡ����?���]&We�����2|X�s<��u���ڕ���dT����#�t����kV�kF\�]�Wd*,l�mX�<�@�]��Ƚ�)įK�v]�X�
���:v�@"�ar�|M����zjjj���C���b�NN�ؙz0T_�ゞ��aL�;��w�C�o�>����K��՞s��1%�m��a�c�{���x����y�Q�MNE1����4�;�����$�Z���X��/<i��yr���f���KL�"3�/�f)����U�U@p��gv�<�Y2){GH�Q����S��e|ri!m���S	J�J�X��&��������b��-,�vt|HO���N�є딇��AGO���pk+��OSc�۟�'���-�:�g/�|����);3�����/^xxz�5NR����s/#`��N� ��E���UKcc�[�lp
��*SУ�l;�#�5�ش򎼀E� ���3���z��c�M:^��w�ߩ���{O��1�j~�:N���I���<*���?���\�4Z9Na�K^���[`K�T��#^�:"XaZ�	�̩ʲ�y[�sk������-��ԕ�+{�5��bp�ka�kpSf�4�4�ݡ���er-:e�E�<���Oߡo7�C����e!rx����U�|w����Ȧ@��R�6��\΂Md���匪Ã-$���S�i�bUǛC��4�h����p�ziæ�u߄d��V���x<�����,O󠞛������$c4.�+�����}�ݸ�	yF�*�%a-i!�x�,ϊ[%3k�Ho����������o8��؀��a ��ܗa}�4��f�$ְ�aj�.h/ءʁ�dXH'��+��ZZ�I�< ���+bt%Rie��K~ԏ���ju�m���`^ewY%Xz���:�����-J����o����(S��'�;��w�9;]Y��������3�����;w��{�29��VOG1��?o�����޽��9Lj���wu��C��nv^��!xչ�Z��9><.EɝN��K�˦����ʪ
v�Zƚr�Bיۻ����X���bGt�]E�b�]Er���XIy9��?��������*�I��!�#Q�Д�t��аQ���Э$fo�l�� ���
��w���bf��F4%���Ȳtw�"���+�/''X|M�� ���S�BX��<��9&���3	 u�� kpW� h��++Ǭ.AAn@�)SA������N�?ꙐJXn��|L�6({@���隦* ��w`Kz�� �N�M���b@{��<���@���d������|�����Q�������d2+�;N�]r��}ț;/o���!����`�q�f�	�5*F>��\���Fク��K6'�c����W�r��0Q�a�{+��C+��+"�����N���A��F�R��U��CggmW[��h�/�zN~JvVzR2�+*������J�q��=�I5����國FF.>f�w�"o8Yhx'1o��O�� ,��,�+��y��g��9i�E�aG��Dl���(�e��������խ�����QMI������ITG~vnueuj�RWgMkM���ɋ�3..��M�E������Q��������ut�x��s}����5�e�9SHd����j^�k��w�9@9v�7���p1S�"�Cx��}��>�r\��A�}C�+�@��S0ƶZF�m� :���%�>&��?�=�l�ɕز��(zQ��G��0d�XTe���J'�D�\[lSDl�B����c �QHi�N�(�ȝ�[��R8�����zk�p���Ʈ�	X%HB(L�o�\u�l��ߞ��* �G�������dq'���� �QK�-�NaF�-�/�'Z��`�+����i����")z�Zʭ{�8wm��v�p��G�c�����gaow_9�?�2�AJ
�PF�!�}��N��^����	�p_�8<\�.��@c�#�g,c���b����q~_@�2 7>~�݆,���9'��g/r�&?��������K}�[}���TP�Gw}%mg.oC��^�ؑ|�&��&�rKL���1��-�Lį)�zu��x�ݼ?_�����2`V��:�+�o���l�ˋ~?��n������<����������������݈���ͮ_ћC��՞���~t�C�򊎪��� �h�_,��G������9v:*�Ym��Zi���;۰��2X�KYBz�K�r���6�?�����B�s��|&���ZK!m)��A.�Q�=e�+��F3an�|E��1�J�q�E�h�	4�;���LUڔ�ܳ4��f��%�ݥ6�4�5�i�~ʍ�0\o�hΛ$�7���@�t���\R�ʓ�JE�O6K��&)0�e��qH8�������5~�#��+h�yW�k �f�K�����t�-���|b���*�ߦ��߀n��
ǵTA�7L�N'�l&�M��%���VV���2uյ�W��4�I�@��ᅹ���E�~��Ht���𔄄��Kl�9 `��ؙԸk���+���.�,n̈ɮ�NL�g��>�?�
�5<H�pH��QR���z���0YΩ�����$c�������&�R�6A�E}}�L���P��l���6a�m��~䀼<j���@wAn�~�T =�G�YGl�?[Pp�;�vؗsusm��kjnz�����)?ҧIHx��}����htt%3�meM�#���*_�M�~'$"�������hIJJ���L�������*F8��P���Tm���}������x�W&7ՙ���
���5�8-��0����f�Ldar�v^"�v���7M�wf5`O��$��@jy^2��<�w���1*�N�	��$��*mq�U���I.�zeN�c�k�(�w(����c������M�<���4�ⳟ�fp�ʟ����T�G�u#�Hct8�O�;��F�鏃�}�s��Q��o]!��W�l�gl-��/pA���S���?n�(��W�U���B9g]��x���ټ����x��J�(�$��)Q2�UCd�j sB�G�\�`K�奙����h�k������]!�!���{ TI��P�:�����h=4S������f��{�T�nRVL�惉����~���7Q��^�K�0��" ZUf*bH8�[@��5�J���^q~��A�7�����{��{�Jy��ZJ���bQ[\x�K�ӵ/͝�Gs'v�����$�:���{�n�ж�&�S[��6��}7��w��+�	��oR��./#R�^R��\���=��>��6�V�oI��b�/ �q~~ޜJ�Z��щ���L���c����i�d��vv"��^D_C㣺v�aNFR
0����Ł��M�eq��R[�k!��<���^R�,�N.�l�א�3�(x_N�*�����(�zg�2�j
k6��$�s��d�,8�79[��^�гMG�K��J���lR�2��7��bȻ�^��w��՛E '��j�l�V�YPm���
B1��R���pb����6�������Z`�p������6�]W9P���T�)�$T �~�Ęw�!I�RF�O�=&׭J�YW��=�8�h9*�yߊ��Ўqp'�${�{�V���z�?�I"ɝ��ݿa�`-��PVVF�Cy��ޡ���Ź�鑁���ab'�U9'+9~�"(����$PO������E&f����㪑�iO������ţ���9��&[�9�9���s�-���
l��c���=~Q ��?�����Or�-��zp�dT�8��^�&��nT<T학�d+B/�,.��n%�vǅ�6�c^Q�"���J�'ʦ�ǧ�$b�+��h��LfE� ����777���4����K@ ��f���O��}��N��bi�5ߡ�����Wc��ю����{V�x�.xtD����~JЯa�Kf)�!9����լ ?��j2� �ˆ�:Eǝ��PɧQ�s_�4, �A
#r���!�z�:�|>�����UI�r��;{O_.љ!LԎ�Ny>q1�R��}k�?T+d!z5�
�6��6}6�}^W�z��!	���ܫ����ܫ��#O>��y�j���y��7���ό����$k�b��w��U)��B �
�;{���z��Ӵ����w�yA��z%��E$Χa�		!=]��-ir8���ԝ��IN����j4���]�{�]�n4�V���@-B������*��6������u��l�}/��T�ͷx����t3�!}�;H����S�tm7��;4vt㰫!�2s����G`��H���s�R�����z%u2��"Zw�g���p�ct�W���:����-���d �����*qNG~�+{ �xx͸��񿹇�\j9���+F�k_�=�����6���f�O��{uո�ٲ���**V����g�c�t<��}��Pi0_������*>�P��/�M����Pl��֚�����B�+�]�R�-���-�B�w�����R�����>\fQH<<d}vq��֘�8C�l.Տ.�S�젒���Ў2Vy����|WR��ʺ��)���֙�O�`�-�
ƿ 8W�;��:��=����CRb&��qA��0��"qNb��^�*�ĩ/L>���y֨\�{�:�E1�
��@����`��	X�?-Ěqwܙ���%b���ހ�����5�q޺AdB"h�x8�Q�aa�0e2ӗa�M/eLF�~�9���!;%c��P��ҳ>HEcQ4��aK���>�;~~Y0UI�mw�ߐ��<����p(om�6~=xD����X�P�\�6oS'���wz���������L�0-��D��w��X=�2r<�b������˦�;�%];��%�jwk����j��}ᖼeNh^�j��)H���1(A�+��k���n���{�-񱦓�$�渔�k5O~���N�eCS�V��)���+��YY����e�չ�e:^8E�Q7���Ȧ����������!��}�xu~~~}}��g9�uYaaa|�7^];\r}򞡯_�N!�����dA<�v'��j3z?mҧ�z�$�/F��P_p�ƽ��PVqk���O���T�l��{<u��R�`z�9�LR�l�;K�R$�k��ۭ��Ի	Y.�~e !��v�w��g��7��鎪#�u��iI�(��۶]�-t���I$^��H���=y�]��=9��"�١B_p��3m+O~v��	�Z�^���bn�a��R�F.,�w�>^)#ZS��n�a��D{�!��~z^�.�{�${��7^��[��%�?�i�K��1�L�`����A�k#��q�%�p�^;ܯ�Y��Z���Hu��\����!T���_y֤�&=��3�V&�xO 2ifq�f�fA�Cq����~����L� 	��'1��H^���7���X<ܴ�j�g$:�Q�-J�M��0VuIۑE=O��~��DF�u��KrecG5�lU]�QM�?�& ��3j�-� G��p�#�S�ߡ~�?	Tk���.�V�}��IS�7Х��|�@����#���KF�ۑm�y�=n����Y���>������h����^��zr���s����kWU]���<>��U�	��1�RWSv��m�Ik�����Ud-����72r���h����L�����ޠ��^�qE�K	���@y9.p���#�e'�-O[��80O��P'+b��p�Y�s(�ʃa�08�;$#'�W�^&Wb%���8�޵ۆ���x|�$	ދQ���=�@	W+��Y��I�����n��h��s/� ��F��2����W�x���{ؤ������.<?�PO��C�s	B�U��C��k�!��X����:���@�w�u�e�Jd��E���#���	:ud���A=d��(���{,�P����Ci�Mhs}KJ;vQQł�OI	��Co��w3'b�!�. jqN��OM"�>�+?����� |��$�2I�X調wo�䙞�]\\~#*X��!,(����]J��'DVv6�*Lr�Ș��6,��H��CT�R��Δ���k����D����� G*a;'τĠ�&��q:Q�ױ�A���G���B�;���###;�ۧV�d�c��%�	Ư��l����3{ƪjW�llp��٢���Z�*_JQ��.� �&��6�F|��y���5!����q�a�w�>�Q�$3�������{�f����u+��XT;;��������҈�/17����T�k:Ed)Ch>Cl-�K8q�+��S�N�c�6������7�AK�W�ђ	,b4ƛ�� %8�C���}�D�6�������?U΁v/�N5�>���yh�����n����|^>�ZQ
����%��J�X}k���݇��A�.z5����?M����Ĺf��vȮ ���[.�g���ah���o�ݴe�У��μ�r���;����_�M����w��"��}�Z�N�J�8ȇɆ]�xH��%��� ��(���P?�РZ�C��΅ӫ���Z��)�cd�F�m�w�vR+mXHt�'YW��C9�y'�"�C�}�1B��A��b��zY�$K���n$q��V�%FPa��R]=^h�S���15�xA1:�����n�w�GY2�՗��R+Y�Dz/�c�k��\NC�ﺕ�ډl�6\���r�T=�d~���e�cⳀNZO�����H�~��ֳ�/���xJ�����}{*�c#C}]�!!S3�L1�Ώ�T��ŝ���Ǩt���{6��F�^{\̝��:][�����C˳��������G�VH``mb�E�$3�B��=x=� x�%g�"i���b�#�i���eac�P��X�[�����]����.=4	�RkLJo,�H��c�a*�́�QU,^�x�8��_��r�+���u��e+b�ץ����)�K���̗��/�:����J'傇&]�_1}�`������0�uy�<����[�I���#�*�fzv:Q���`�����ST�r`�,�-����� ��`R�k�l�t��ɜ:��>081���L��޷���Z&W�K�CF�a�<��%��?��k�rN�%8�6�2�Д1��w1H��+Y�+�����+崤�����S/������Tihz\S,�V�����Ɂ�˸<�k��Ow�d8����~��Gi)�a
��0�g�h��4{�+n�֙Xw��_���)�0��FQ���Cb�dȮߛ��N���sRΦ�`���ٝb�^���e�`CE�䯦��������/��kQ4�4�j��j�cE��D_����:�Z�s^��k���z�M�����X�#��e�3L�--�M-MmM��-�`s #�����4��RvAHOM^aOp=-���MAao߮ѝ+��e��f�	9�ᨙV�V]��_����L�M'o��YJ*�?�}ړ�����Xg�>I���Qս��1ddlT���V����T�,�������]4�����e�'n�+]�g��T�Pa��gL��xp�����Pҙc�ck��tM@���UJ��p�֧+��tj:�/�=;^���9t<��.�Uz�I�ll���S����������t�e�6G7�W֕��՚��J�|�6+�wM4�,ph���5H�'�\�%�ooG�VP������R��(�H�����ù;�*p�KWr$��J�!/6l\0��ɂF�_K����{h���e�4|z�K�O����ߙMF��������{�S���pX����VF<��آ�1~]7 f��b�&��M����U,�Y�vMg�ȁDu ��J!Jh���E�_]�����d.7�Y��y	Y�Jm�Y"��8BE���H4X�R��J։J��^:QޗD�L�@����L�ʬ*ݬ
�����n����mwfֽ&�S}{'i�%�FW��"�^�E
�C�:t��f�ǾN_<��X6t\0�
�<k�M!��&R����
#��keV���C�L�]j㤟�Z��3���Ae�L�B�-��:�
ᴺ�9�ع8i����U���6!��,+aF*���$`A�:��)mӔ�a�෴��?4�^�c���/��\K~��b�_B#�Jo8���L<��	8.p�Y���*����X!B�`x����ͩg:8�t��n�����h���W_{X;�L����%Y*L�6؇���Y�p�|�΢�ÓO�b�8��F��������c�R�%q]��lVc{�6��x���T��R�蔗#�G#`�2_�9+����Z<۶��ԫ+u��AܨBaR�XPY���"�a)����`P��{�f�p�֕�gK-o-��z�\�U�ͥ�Kqcices=��퍸(��[-������������N�v�=x�:��X�d�M�� ���\XX�M$��]�m��������#�P�\����o��J@��Q�+*�2o)G�js���8�'C����I�gg��,;\IU  9���������(�Gd�V��C����:�]0��q�_��X5�g��dV	�(�<`�L��A	9��}��˼�!;&}#u�Qh������I!�{	�Y�}0k����-ⓨ�KJF7�v���m>\*|:�x/�c�+�!� ��!��"�l"�i��c	y��Z�W�#�ûQ����d?e�x��`X9.4]nНش��kL�;'��c\;濁�����jxii!���x��,M�M�G���s, �/Q@�,vn���<�sve���~3w�}�L�u�i;L�Q��C� ��Ƭ��*�$a)�^xl�����_�u�p�����������<\�25$+<ZåK�?G���;�6���<���j�n���?�a�.���q���L��� ;��v����W��$��$��w��_�טy&�n`^���%]�p\O��DT��D���C�y�t��M���>Z��;��< J̧+���eXЈ,誔������i�NA]���x�:	#/(�*if��jV���X�Z�򎇅��p�<FՌ"��<���)t�����Y���i��*�~�><)y���hF�f�`�Q����*<����h^s2{�w+L���8���`��;2m���Uka?�m�o(n�ǳ���'�E����vMvYUĩ�T�A�ɰH&0�)nO���������30���s��#Bp�8�(��ӣ�|���h���]�B� #+���*i�g��8���ι6�>���j5���z<C.%Ql[�n2�[n&��]	,*���4~EN�hxR(W��XQ2����4Bx��L���,*q88�hO5u��c��,g+�#n`0�4��#���c��q_�KY��׏n��9�H�]��h�c���	��� �MB��6Rs�vz�M�l�e���:��K�`أʉ��h����A�.�����|J����pD���S#L�'�S�����"��nת�_����s�k�K]-�֞G(=Q�?�_Su�	���V��>5~���.�W��\�e���6�|�!��q*�Z�aJ'���X�l���o�j��<)I��j\|��>���}*̏�W�PPU�M
Ǽ��i� ��c'H*���@M���M�������M&+�����FG���9@�������TwzO����;�,�,M},��^Mɽ��9W��'�7!|�<�����1�Bx2�Y��sF�v?^�v���gv��8n��#U�3�p� SpCgU��3&�"#g���n��s
K�����l�]���R�[�����eԿ������_A��	����9������~m�_X�2NX��c�Ǣ���MUU��I���8�ݐ��Ô�Gx�`I�(R�204d[ZZB ��!Ņqz��_-  ��ψR��������[A�bU�_��^ߞ[Z]�RM�a��}��&(��b��omb;SiiO%�頚8%���/e�6�+��ѯd$����������,�I2t�!�#;��$�|��u�{&''�?'rvf~njk�z�!�s�Կb[��9)�LR*��+<#/f��A=�-�TI�S��O��K����ޡ��vIm-i��M��o2��o��XD�	d��%#('U0P%(N���n��A_I�\ a�,��"�/X˾�7��@�S1_�cM2��<��"eM~��^dC���7��_d}��?�ݖ�;������o��2����mC�����[�B�z3���W��X�ʈ�Z[p��7�3�rH��K�����i�`'?�x�oä�<"
eTح��TU�VQ����x`Iv��In�Q(��fg��c���y{;@QI~���H�:�2�K�$�Dq'S�B!�:��А$a�7��л@��BΈ)��-�(� 	��ù�d�x��Y�w�����|O؜��,���fԵ����E�V	cYďu��OBe_�u����xET����:���"������2c��Ɗbp��8��Yat0^.Ja?�2ɦ*yu�c"�lz�^�2�$�R^��.��b��?���z;DOI�Q�ſ�4�8�1d��D �����&ǿ�\פ����\ܓ�v���:7;���u0��	M��/s��}ص�6N_���[l���>�ݜ+�O-�����嗻s���˅Г\�J;�t�OWi��l3CQ������⾏��ԁ���~(6��V|�4��^��le78�;���5=�������k����\�����D��m�/��Cq����yF8���0�4���_:,�����7�W�O�`�B��G2�$��Ȓ��U�)i�okm��2�"�u"�0�HD
H�LN<�e��yH4�k��_��M�>�}�?u.��d@~��v6����-
za[}�{�6w�/rH��HE���i�{�q�DM"��9�ns�����j�krI��ט�M�$Vڮ��7�}�#R�oar.� ���.�k����]*�Bn�rv˂w��"��<���AS�b�b����=F=bFM�h�CCM��Oy���������㋼pxq�eI��ڟ�W�6O���AM������ر�*Ո���c
�����\\f�!͸��`�^�)ɻ!N����Rf$$҂�Y��3s�����JԢ�;���)U��3����,*��؋����Pa�qs3'"B�~g�ۮ�yi����a����5��{9�?��ja)��,�?!K�	b�P-z\}�� �|R�g�y�K�����B9�;h�W�i� �ꡆ�H��o�ء3�L� Yw�SP���k�����D��[��Z��!M��+mG/���ů��>�t{!Pﳿ���r��+�n�&a��/��F��n����>�J���i��VE�h���k�B������o�|@�w�q����؎����08�s������8���U&�7�����c���Q��Vtj�Д�:ߖƤ�;��W�s���9�- -s��ļR����˹ɕ�ߑG�/��@�$Q����G�U����[����S4_��ؼ�N�S �y��f�����\ף��ѱ�༳{B��k�B!�7	��4B��*�h������0=�Co�aŀF&tgU�hF��]�I��}���K9g�R��i��C�{����a�5k�V�ŧ�&f)�*����b�l�Z��V��]R{��E�{��Y�����;��x��	��>��y����@�pݙ��z5�|ћ�C�s���8] %e��#%�$�^����Uxz�'�z.xʳQt�' f1	[�J�^��S�9�3Fx/�3e1[1��y�U���7��>p�f!N�b!Q�`^�Q���_]*ޘ��g~"e��,��3�l9���c��N��i����L��x�4Z��ƿ�C�7�]n�"_�KG<�N�n���\�Uo<|p�CP齱>T����]e��A�]���A..��\���P������gmg��[�]�wL���+� ��!F�o�Խ��^��,Tl vɃ#?��=联��\�Z���.]WU)�}�����ꌦ��������&��-�?�N�vn�.Umd�M�D�W8�^ ����z��#�5V�5���R�1-F�		 ��4�:�yd��������0U�B���k|��Ul�2k�Z��@B4���!���*�JJnJ��ɝ�R2=o�qB�Cy��&aqs��L	��OU��5��c>�6��q�R"�x�Ƿ��tݝ���S��q�cبF����՘
"�
��#%@y��!K!�K5��К����MZzxPp�X��!HT����FԝF� c�_C���[�?��ls�Jm���l=�~���q�P�����K���ut#w�@S���ij�������9�<��	�������U2��G޿_� "K�I�-?�p�
�7C��~�����T �RE������\�&*��Z�⸏Ǽ��7�е��iÌI��ə�<q���|��cb��w�1����ǣ�k��T���#8,QX���(x�B��[X�P�9u�������b���p�3���!�$�A���``P�����
��6�4�l�D�ø�1y`�۽a���}�����w��E�E�)�:��e9Xe�!�%�Q��hcD�g��" ��.�(-�d�P3veUz��?a�]��<7�*tp�8!��ú{�nWW)�(�
�e��g�$����=~TX�i�$t�:zI�JK����bծڲ����
�R�zQ����0(�-$m��c<]O8ya�P���p��F�~�|Śh���#��Ѷ*��$�*EB2c��%�d�yY�Ruem@����#�K����Y1J�\��3cX�5lt������4H�Mj7�e+4~@a`k��S1�=�nA?�2�/��4��U��n��jI�q��+�/��~]�UN�W�y=�1�\�8��X6`�3-�����ů����w�&.nor�n<�2�Hy������1wZ�㟥���]<�G�&F/M�(ެ��ܬ��X�	��
�kiē����}����Ǉ�b �:ѯ�=]$�`��}��o�V�7���vtOv��~x���x��yvW�L�!v�A6A�.�8�;���̖���wu�T�6&�@w&{}&�o�h��q^"�o�f����K��
s����*t�K1O����k�m~��D�Z�tx�Y�SE#����<K�E�ޤ]������O,<K�N呙���_�J�F>brbF�c3�FV��>�T=�z�ы��ݳ��yڟj��<5�l�!�תZ!��~nڐWpbG�]+�p;Z��,�-O�N��9K���{�f}=]]I��zx�R���C%yC�?*��$��'V@�X�=PA�L�沰��4��Ɗ��;0�q3�2�F�D�i�B�ӀF�u{wwO^=��㥴�Oj������W�o�
�^f����RNĺ	xn}i�5�h��;��F[�	���l���	pe���;G�ΈQYZR�z�ob� ���mծk��v��q��/8�����L��L��L�N2p��=��{N�/x���w~�я�[����j��[X���+gP,.vL.GZ��;�q��C��BȭCa�:�ɔI��u����;Q�e	Me7�]�&�	��{R�7F�2���(~���u|�7)I<�]�x��������/����M~X�7��>b0���vL�wS��2�dܵ��~����6�R��ʿ� �)ꏈ>S���]W���ǕOF������y�Bb(���L����_�Wo����U2��9�A5d��.�װ����3�4��U)j;�|�=��9�s,�w�r�!��X
F.�B�V���
���rb��Џ�2�k����Q1�\�/�ݫ��� �~;���OU}�Iд�8���DKA��p�3���;(Jn��
�^v
��"'��r��E���8�5�༔���S��`2�}�Y)2 L�Ȅ&���V���
����J����O�3�r���g/�5�%��	z�y��*���5g�����\b�:(&0^w�M_
h}}����lk�6j���,���r��Z�z0&r���ʱ�zk����4��.��;����K�����Ჩ�벥���! `�ϯ5.�,Q�?1�~uI��<=0}f� ��=[l���nB�BQh cj�+��B�2yS�zSr�$�l`��Df�\��D��W\^�L*����pl��0��P�h�;��)濞��N2���f��ZLĜi��k�1�u��K#<n��:��j6�dQ��m�}Nԕ�[��q��l��o8�1̃C��Ds)��X�p�[����A"N�����,�F��&a:pő˗)D`Y����J4��g���R!_d���cf�J`mw��/�\u3�o��Z9$/,�ີ�������y��B����wR�@(:��O㿱'jj�
W��~�Ⱥ�
�d�����N.����z����$A ��c�ё��M[m:>_��#�ZR�&$�RO�����:�����o
�z�A��������Jm�a�0m�g�C���	Z�|Fs&�׫RXc$����ɹ.s{q���Jf;P���4Ni����Ӊ��-O��OTc�͠U�����kw-�,Z�j�*!Zp�DdnC���	S�Wi�A�<��=*�N��sqvwM�qɽ2���<<� ���S��ʎJ��EA&y�0u�5�uݰ4�b���
8�;s	(�D�=���5�R��W���v�����o�s�ٮ�S��3)r�M���נρ7�
�Z\�R��ZOi�ժ�J���5� �."eӢ3<�<�Gv��Z��R�c�f=JW���)0n�Oo�ֿ���њ���˟�1���k_�0ܡ7^c�k��ѻ]���Q�Ƽ��������3^��cx���f�`<3!Wv=ˇ���~�D��*��-�+-b��E͊�e���a��uP�+�ו�k;�����9���[耍S�3W��*5%��*��߇��F���{L�h5�ц!sc��f��"�M?�LH#�Q�ޙu>]�1>��֌�F�)�&`5]��p�ᖼ:�	�{`�m�+] җ&���E\f� *q��>��WP�f����ռ\0w�\K��B��^u�-�Umە�����Q�Iϧ�=�iiǺ���&��_�Z�Wg�s����-C.�rB�a�l��M,E��N�y���m���km4��˿Ќ=���?��V�V
~���z�w묷�?�����*��-������694us-ac��[���l&�(,� ���,�/2Xf��ˢX�M3�dA�s"d&)���:������v�)�� 1��%q���8��8oĸ�{-�
�����4௡�Y �&�z�?dP c:Z�'���g~���b�y�[�p
:�uL}��W�jw��cA�#�}�{��k��	�nG���PDV��
OD�uN�z_&�V�ş�]��`=<&�b��?�iE���>���̘D��`������m��{Ტ��^��nďYǗ�=P:���х�T=��j���S�5�\�`��յ(M'`|���.��ӑ��X�s�{2J}J��/�m���Chv�5�tMǈ����ޘ���_��8��a�7���Ξ����/f_����̙�Ek�m���l�=o�25C���jX��l)Y��w6g��~EN��p�L���Kg8J=�� /�=�Qb3|'�0!�K�?�\�[�}��DuVa��3�����6V�"��5�� N�F�^ܣ<��^�:�_Zvu�rpY^ub����D&:�6����>z4��.T;w�ư��ҋMG�N��'N�,(�u�H3���zx���p��h��U&go����:���Ømܒ^��_ޓ���)zP=O����Ets,�Eҷ�t8�6��9?cH�=ۿ�
XѤ�YIQ�q�ǘ�E6/�P��#�<���:ݰ��w8��Ψl�DD@4�ɖ���{R?Z}��>�R��T�{! ���',�`���D���ߺ=l�������᭸͆W��_y�w�MrI����i���� [�'օ{%�DY�w��ԝ#G9(�_ߧU�Gp<a�� �U��h� ���z�p�Sa�<�2L<�'�3�2�M���W��9� [׳Ul_d�,ᘺ�����Qo�Ύ�]��i����Yd�ઈ+<X|��XaA�����3�+ƫ�Zf	Y>oR{�t?����'��yP��$���rz2�#r�V��+��C�L�	's��^���/�ީ�$�)	���"���fYP���}�6���&�������-6 n��N�i	����8ǧ�<����p�V�m��5�?�;�]��#��
�����~�d��kz��'H�Ϝ6�I&�[�v&�ە7e��*�b8��.�-�A�q��,+K�y���D��K%�VT��%.�����3�7o��}�1� �z6�}�nv�=�9/���[z���t�Sh���d�,�
��� �[ae���������q�Hg-�QQ#)-:Z]!^W�����^��zz���|��#ٲ���� ��,��v�yR��5���58��cvA{)$��9ޥ��HZ��.)@��}3�HÖAP�[����D0Ul���+ޅ	ϧ�mC���� �M?$�Zy⃓�p_���N�5o�㱏�hkh;���S�g_ݞ%�:�A���t=�������V؁(q���y�(�f���L�MUi�&���脰�<�]�	�	�D���ê;F#?�:(w;�;�-��xy���H=V��k����Ć�Xk@��Ed�����=n�e�M���R-��@`����U�0�H�:92�kX�yjYZ'f�y��̹)�>��H�թ��<�>�¿�������笉O��:b�ﭳ2q�|��_�>��NSzTpa�|R%�5���4����A��тL��r���`����I�ϼ!ܬ*�ޝ��49�$̙�LX��*̡D���,&�����HV�h�|�D��TXe�64�����_L�~OW3O �i��I8:z����M���d�1��DO4�1�T�q��\I+����	^�u��Ź(ӐK��1:9YWQ���YU�_SYY]UU��+���t=���U?������ �{(��}H[�Uц�ְ2�Trʵ�h��-Ok�����������~�����#��s����md�1��v��g&�Q��yϨw?���}��qޫ�7�����1qw�w�Ky�6�>���oe��[_^�[^��ތ,�?r"�d8?nK�E��}N%Y��sEw���XC�,�vO��<�x��}��32����ɦzz��KJv�6�wuO-��r�L��׆jV(�����eaI�: �,)��W�,��2��2�"B�+�Q�G^3HS�G�ϋ\Yb�|�{Ў�I�G�;�����˥��;iz{��8��
�����f�M	��8z��(�slн�J%�}��R�X.	҈��g֯���a�w+��r3>a}2�8в�.�g f� ��}�����BJ��B%F�>V���~�_�;���XlCP��JP_n���6��L��j�tٔ7��������LC�@5��R�U��<kqq��6r/gtml 0Jκ��������-�o�Y���ؚ1s��6��P˂.�|EAM�Ll�����ֵ����V7�}a���gh�JT��v��q��Q WhT��t�g��;�tG9�-'��r��p4��=*�� 9��xǔV�d�~C&��b�tz1�i���v�tn�I�ل��h=.;.�KWR )�{L/��*�T�d���BZ�	�W���R�|d󹽭�9U�>��i� ��o�ˬi�+|�TK���s���[�e�5
���*�L�:	�����k���\�"��E��aN�R��y*@������@v���xѝ����I�=��<ń"��۝�I�N=�q|���M(wwݣ�&IPIK�OQ��������-��粲2h��������DBTrB���]�[�^��+�ul�_�v��->>K�"�[V�;H<3u�M�{��|����s=�ptdk��c�@z~�S[�p�R����@;G1�����?m��,r��-�rwwf��pGh��V�fr��$���ٺo[�7�\Z�eXಬ�M��dn~9C9��o~��m~��n�A?d��,�������G��sI��������un<����s&sBOK�����W�	K��!C�YuUu��'�n���������9:
_/b��Afl�O�9|p�Y\�jEk�	x�R"�ÈL�p��2أ���%]1Ef��?(4p�m�N�7
���+j >fl� (�N���h7�S"B��}������f:X~�6���?t�7�3����qSKs��8��ߣ�p�-~�oBY��~pD������|��g�jT�d�eNF�+��Y��̝��A�7��R��J���ŗ�KF a4;T�����mt������,==�k��߶$�r���_k_��)rup�L��嗆����j��+F�˽~4pР�FFd����$(��ACJfB�c����|l�GŶ�;[����F�:��|������B��_|tI�h��uP���C+?�몪�+<+D�k���V�{Ɯxw7�|��*�B����p+t�#ec���L�f�8V|X���
���YB��b��V	��l/}ܛ�^�Hܝ�bMz8c|��.�y��S]���g��|:Nz�rb�;]�JS�d� <��T�=EA�r�Z�3P���<�\�|�?Ee��2iC;��,�sVG 	T�ŔDd?�3�yؽS(m����V��O�?���-�'Y_�����o`����?��沽Aط�6�3co�cתB�<0dY3f9N���&y�_Ծh/ec�yl��%��S� ��,��#Ş��T�V�$scq
7�6e��;A����Dg��i���I����tb͛ܓ�)H5I�>�c���Q��9�{W�^�a��7�d~Ī�G턞b>�8-�O�%���h���Nz;�q� ���/�BnK�);�t����f�(o	G�h&5�^�D�$��� L�}6�%A���u�#_�Q�<e�}>�t��f^J�}������UF���8���=��eϱx�8�+�����������4�E(�%.'�|�zi7�����̭"�<|z��,�3��u������b��ӥ�������T\d�/T������_�����U�o����w�wR�xNJK��;���^��J8g��n{����:�O˳������B'޷R/'������e	�_S�_ذ������a_�ye-t�p�#��1��X2��I�3��=��D��#QF��)U���8E	d�P�=�H�0�|ƚD�x�4��R�;���ѝ
�\���;G`HSD����~�<צ�&9�g1�g�̪�q���
��Ia����ﲽ	�ȭ��EC��u<-����ht��/� �<���V���&Y��)�fF�Haj��}p��Y��~���h�����1D~�n�P��Zow%)At`�y�}�5��[���I��LI���c� :�%QP��#��n6W�=*z��3�Y��:w!,��%�r�r��Q��#{F��x�|�E�'�S54L�~��^�ʺ����ߚ1������B�3��9�/z���i��X>2��
aPܡ�8,�
�	&$��{H�p��d���ߑ~'�VxXd��4�E&�`���z,o�r4^�����Z��`�'���dH�+�W�ޟ�NN���.]�� ����^�-da��F�?�j������)qP�r��N����U),"� ���?��?��/� 9��w������k��IZ�����\�6��ŲҢ�5�Vf�M�F�3��N2Z}]i�L�r���#
���dT%x���2������i ]����R�"���r��q�y�%
rU[�ZĎ3E��r�Ф��Q@�vkg�Y�1V�r���1t�L�_�.f{�c9N�e��u���j	�1c���a�J�QQ�,�X/��S���Oc��v\Hf�4'U&�M���s�G:�Yp��Z��D�u#�$p�:Ї�G9����Ys�m�|S53��U$�tY(�`JJ#�V/<��k�k$�%Y=gLGu���n��9��7i#��V3�B9:LfI{ ��Tq�h0`>�@%1�:jQ�iT�*N2�@��P�B�mZ'��'���E�����b��3�-��Jg�����2]�&9��V��jO��r������An�Xf�PF����ë������b���'��k�9׿�,//{C/3,�κ{�?\,��4��k��,͘q�	d���nn�i�29-);�������Ͽ�r��p5�ЀF�]���F�r�8�T�����hL�T���l�l�NV%����/[�����l�
���=r����׋
�m�v�
�lr�ݾй�3l|�Ys1�ݍ:�x�@��#ܳo�|���=���22�&%�D*�ĺ�aXx_=��Nm"���v�FEbBL/;%}(�h?� w��M��La@q'�bW�<N=�	I!ݿU%������Lt�%k��<��?�u��ڌo�������P��"����~o�*��g1�2�KW?��s~ܾ�^��H���^���b�~�ra����i&|;��x��k,�;��۠G?�p�l�C�B�ҡwE�cx5><��-�\���3����$��_{�y��G��w~�Y�t�~�_���[K�!��v��%R؃�ա�9�<䅷��k�&P/�ݿ� ��ʯb��[/�u��䐑��`n�iEAE֘�����	�l&�5�o��'j]M��()���LpV_���p�;�>�l+(���|-�X�C:t���K'��[���ԋ>��&�Y�u%*�j�Ӿ�C�����S3&��$:��V0p��pЛD�Qp��qf��!����-ǠM��w�%1
�'��J�`!�  /+�����>���Jq���s�W� ��)��pD!��~��$��q�/HQJȢ�d0	`.YCb�� .+���µ�'�V��H\4�����U�d ��|�W��� �#���Me�݌M����eN���i�A��a��K_���ttT�6
�u�� kn�Ϳ40����6t�۠�B_E���5.���Uʰ�k8^��Ч���wߙW �^��6��U �z{g�
�!�����j�T�3��M�Go�z$��x 	��v�*2g*��o'*��Ud'����J�����R�E�R�D���,��(�$�W�����w%�#o!W������ȃ����K*�R��8s�>J������w�g9�)��E(E�講;��oM#(��RѬ��-<����ؽ�9R��~ߜs4��4Fu�S8���3�`��ٛ��ꃵQt?{��Jd�%B���u+Y�
���*�O/��������H} �46h�����ؼ��+�.F<,̂<��,�F�����x�|���}������"�;:�gk�#��,����`_���9$������n|���Iy(���K��Ɠ��-2����`0G>���S9Zπ�\���hg�)���d��fg		����	B܄ ��GP��ImV��Z�^��=��d��%���S}?K��r^pj���d>I F��GX�B���R�`�sh>oi\<�n<�9hL$n�.��f�0�b���K4�/�ZK�+���߱����+S�јp�A�y��x���>�p����%�|��Nu�g\⠒ɰ ��a�x���lzu���La`�}d��9A�_�Pk~����w��"�)F9�D�4���֒
�xR6��7!�����g/�~�追�&����|ȏ/�{��.p��|��gN?톔�����4tƠb�c.�L5�C͋t�r��ۘ!�:f�w����/�~����*弎c����
	-n�Ո�u 
��~.�Q!Sk'A���d��  ��F=�q�FƜ*�I׍utB��R��1��	<�qy89}�G�޽��U;�1�:�~�@��4U�Ƒk�j��斅�!�+�7�:�dn�0)H�]%�mt������8�կB����2/ᬶ�R����Y��|��'6�<��ܺ\�����at��BH�a��7�W,ǆ���K��8'��sx�q��2����d��}4�a��.QP7݂\��3�p����N�ol�����=rSp�(h�T�{�������h�6�VD䱊)�$UbV"g2���A���Os�B�3f�.��g��D���}�� t��;ae�\��g��1�q<�^��A(�d_��d��@�a�a�p��QZ�I*0%��hr?Pƕf��۳�3�cs��y�����>�:�� �ּ�n�S��@�c�:¨����E�z�<�VL�窐��C�knTE�FCjMI���`�G�uB�6[[y�B����S�g��ғRB�s��5.ୟ(��̠7a�*�-\},��M5c#�U�Bv5hs�	�@��-��]P$�c�s���KO�fu�!��09�0j�������$��9:ΝXE,"|���b�&o���!XS��FnAR噱/�ي�er�	�}�����}E�'����#I��"�VD��s'���N�G�S��
�T�@M*��`��g�:|P{����p�$M���̑�&��<P�Ő�I�/sB�{ۮ��r~�7�~�u�/�,* ��+�-�j��iɫ��������WZBD�T����ht`(���ʓ��Y����tj)^�'���٫[IV�(��o���͍��-M�vu��.F�<�Xz@�.���ދ�u �/'�ڈe�r��/��-\",i�Q�[�Y�#�#.�l��踀�"�M$ۄ�%���<�,o
yҗr�;F�;�" ��ME�ÊJ�E���M�F�S8���ه�p#��i��p ީi[�c�>c�P0�]�mI�����c��l�yg�M����Q�v*�-^xx��A��ܻA�Ĳ����ᤢP.IP=Q�!;�}��e�C��֔=>@z/l{q�"��-�B�*a]��4e�X��+fV����s���;���&���.m���p��'D�L~�ڴb'''�_OH!��S#��i����;d�
�IPd�~���beÔ>�S��a�?�?�>=��צ��	��|�Lz���G_4�	2�@�~�wH��JJ�MMO�MM�=-8W�h�qwxa�j�o.I���|��j��/M+U�2WJ��c��-���]h¸�'x�/ޝ
o�L��WO��ƫ�Z�͞U��+k���6������t��S4��n�©�ƞ�Ir����a��k��A�M�hލ��\��1��v��=��'��|��H�
+
�2���
�1Od�w���0�u��^S�U�$PD�2s�Z8"��LFr��V��社I�j�	�[L�6�Ӎ^=^0˹�ʄ���˰w�qMJ�Y<O���@X��N��R1	"��)���!�CJ�m�1���n�ŀ�E�e+��V��E����&ܛj�uFמd��SnX�O�2N���7��eF��DA^ƌܷ��X.PA�� ���;W$�gMi��Q��`��� o�ڦ��:4W;r���I#����1�	E����=ǒBM�V%��(x���a��m*y2M��&{q���͑�8��ǣ�|��qt�}�g�E0Ё>�8yՅ;�Ɉ��``�K�q���5UmY���//Aa]��\Y�;S4� I���B����������~�� �<�s�~z�:�5��|O����l/����<���P&1�e���Qr��x�3�$1�-���Z���UԒK�����W���=FBOv�'��r7����2h��+��^����y���\]��\�oX^={��hk���Z��K��󑀐��P���LsqCk��/O��H=P����A?���h��5�5���N���F#��'��)`���<��h��8#&=#
��ؽ0�ф|�nIiy�0e�`
T�u�r�	��	1�gI$���qÕ�Я�fC�׬�����9l�ĳ�"E��|�`��QI�ƹ<Ɠ�nB���I��	�����cl�@�/O�_ƫa���N�u����2�se㴑��	��םt���̉%���ݒ�K}�ѻ���s*��p+Z��x�"CdX]ż���IE�m|���Y��'w�O�=���W�fDt�L��T��#g������B�Xt1*��$���]�U�IL�q�}��ȶ�N���?=������K�����a����q����(�l�z��"�$O#��D�ORv\D�<g���HR:����5�y>�%� u���2�2��,��ۥ*A�`���%~�k;؉m~GlIYO⢤k�P;���ծ����D?=���qF��A�M�?�������XL��l�E�`V�)��@�BB ���%S��D�1��u��:�k����
	��?g�u��N\<��k�e��{�N�	� #�k�u\�\S�Srǧ䅊cђµ�wPL>a ��Ĕ��è���
`��$_+F��lT!ar;F�?�&�?-Let����4u�}wL�]���	fi;�2	
���#�ߕ�j+{�g/�a8�e�����T�υ���J� ؎Jԕ��� �Y�?�J���q�{�����w��Sh1M^Vؗ���:�������]���������kk��߅���0���2}n��G�!^���n�fbL�_�������ê��[�=*���<��=7����q�H���D��טG7���O(Y�X5�IN��Mq�{ƴ�-�p� �D��@7^�U�,9C>X�(;)�+��}�� iYH�9�>{,ۉ��WĊ�xJv����uJBW��^���a��W�?�i���E�{֊�t~-�2yJ�!��c�ptǭ�gA���@` e�E��?*%�?£W�q�����4��$q��yB�2������ʓ���:	9?�=�p�U�ãT���po*?�.[����0�2����e���Ѓ޶������7�+���^��d�f��Ѱ1���27uWw��5�m4��w67�$&���� "bP 
tae@S&}j|&AÙ���x�uM]�i����J���aJ�''�e��˃� $/�c�:OϺ�h�������/�����ڨ��/��,� �P ;谚g�fDn�XLb��U�y2�I����Ǽ�ٶ�9,��Ӗ  	� ��_�Vg�75�����j�;W�v��\�zqJx��a���S����g�	��".���X�g�6/�I�$��Z��o����o�T�hF0Z�ݿ}�(s>D�;@%��;����yi �^��. 
�՜��{�z�����_��y����Р��p�/\w�m��O?�dF�~E���S
�7G~ք ���v?�� j Ρ�y�jP������7��&f��� dc�^�Q�����^-.E�_����L���� ����a8�HO@��/2��@p�)�	8U���l�W.��C���4�8
�Q��fZ�����"G#4��ꑷ���;��8�^Q�a��w��,h����:����(n���[P�)�hӈ���g�"��#]�H�B��mc
"ɠ�Jm��7��|��_��:��� 
�"�P�h�7Um2�Y��)	R[�*w��񷻨s<�m���Me5(Z�Yҷ��_� �2�]u��ѦQ�ܖd�Q��H���V~��R�9<_�h.�Xjl�#6�YKi�J)����tj�<u'xى#th���#\]��:Mǲ�VR/7W�k�{>����|��)�M���� �kX�&��x��po���L�=�0�����B�|]���N��������j5� ���If\�~��Y�Sc��Ȩ=RмHK�	��>�f��f������Z
�K@�Y
�-VPJ�V)�C>��3��hr��.A��9�NM�}�A�#c����n�DQ�����j���Ps��;�Ha�Gw��<� ��ׄW\�	�晫s"؆!�:�:/���h9�k�^\6�Sql�L=�7&�M�ks/�k:���ŧ���)�е�'��9�zɑ��y�����r��iK�R���㣐�.#�In�V��d$[�H����V����U]����#
H���쇻ACpf@����H��V�7�(���N{��{�x*�X):�������3O5k�qc+D�#�Y2xo�<Gi�9q��Ó2�4͟pr�_!?EDJ"�	��b{����i���ұ]~y���v�bSxF��oe����o�ߕFz�0��)��̓j�[��^2�-�f5U�ϋ��}��e�t��=_-p�ͣ��dfn~������`�G����%����<m�+#��I�7Gs-�bu��銎=�/�����$�8�m�M���r��#�i����{{��M�	Qtij�3�U�J��/�LT3*��IL�v��V��y��b��R�?��Fqq�OtQ����m$$$QQQ���_v���zգ���UK�e7��ȭy*3'�ޜ�r1u��lɱ:�n~�e)j �9��;��;�0��0PC�����N�ٞh��Q���v_�+yg
#����[>Z��=��>��i�� �ɼ�r=f<h1�p�E��di���I��vS�+����� @��W��U�~"d%��˙*������i�ʢ��2���8�7���N ��9R��C�xQ�a�����r��۝4մ��z~n�����_��\T�S�S���%$ؙ�\T���&]F���_�Ä~d5����Xc��sG5��vNӮ>H�4�����-��Ev�C�^BI�t��)� x��|ڏ=����z��KY3W4�&�a]
z�����#����s8��S?W���a��NJ�J�j�G���V1�V=�V�kŎ���ˌzv66W77g�~!�.��4111))��!���z�N��A;*9|B��X���Y��B߿?g�2Kg�`�b�r� n�45��=縔ԞY<�R�Hb?��he�7T��6�+C�jA:92W��r�/���!,C���Z��N�����
a�-�������VR_5���Ak�0���D�E=��j�˽�m�L�\R�3�8��kJ7�:)+�8B��V7�F��f?�E���P��q�/��a�93g�#����y�i�3� ��Z��S'm�p��3��л,)[��A-V�[H�5��&��Pj����,p~ja�g�����l�,�z�nɯ2䄜��y��wR}�Fϯ���ם�~��
�ZkM�:,�������.���r�_�k������\��O��tL���Xu�Nbb�'������	T��T�$M&O�1��CyT�զջ�6��<O+F�ʿ?|#�)�xvw�tO�N��R�z �N���-������;�M'�]�����꼏~<g��0.�)�ZNu�]>`a��7�bY�N��q~����i��*��{��'�o_b�[��\�j]���)�Mܺ��\��e���VJb�P����_��{�P��o܂�۪ɺ�а���>��Ct�S��g��D��Di����λY���wm�L_!�M�˱QIX�oY����>{��c` EL�q O�e0�XM��p�ۿ
�K�*X�����(�f`�\���J^��KӒ-��t#ښ��F֚n1.-����T$L.@t�\I�06p���7��/���SPN���ᢞ�E"1���H��7��B��IfF��o��B�ozs�xl������Dp�at�����V�zS��#'f�o���Jf5��l���TF��$�N�����r�Qε�:��iuO�;�\��[H��IT,�$Db�'��0�0?����ܬ�o�N��
�q���bJ�j��3���8Y޸c=nU%�,4��?A+�}s���R`��y����	2J�n�ϟA'Nq4nv��ތ�%fR�׷�1m,�Q:R&AZn:����	�}����7�&(R&0,20<��~�|GIy���ULJLBT|R������(��Pvhg5>�w�����O������˄O"""��M]]]}|���U����*AFp�W/�^�����L>��g4$&Ufg��[����R��0��uX����?taȫ����7�{X��������X��+$(`�.d��Nw�L�UT[M���Z��A��WH��R܂[����b�-\���`ť�/~��:�\%Y�ؙ���3�3C,�4<M'�C�0M�� _�	�'�o���~�]	G�y㦴��(�j�@�SKUM�fM1^���P"z���U$]��0����
��� ���E�	k���F2QzP17"�X:��l��<)TO1��GIQ���M�Y	JDmZ��6ch#B�9	��
�S����,�|�/V.z�F�}�TӺItc����:�P���������7�����j�� ��ϯ�x@|�����O��ߢ+RT�๧,�W��c��2�`v�ꉁ��ٱ������a�����ş��==}�S#cCK��ȡ��_K��c��g��:��cb��˖�W��v}qD\�`�͝0x��BCn(�\�Q�dk<:xN7>��:�H�E̥�s����<�����I�D/�=�=s���u.�b㿌E�"'���3���̻t�o搎��#D*U�7����3��O1��m��dn�/���w�>L�A[�x'�w���^?�	S�aihh   ;_77��*x?��,���c����6v��1�.�����%d߯��A��=ʽM��ʓ�x��TR�lR��-˴C˴c��WF��f�M�h��T#�d�m0R�m�X��Do�B�m�l8)A<T,A����s0�W�v��d�9r�����#������A��8Ȩ�q��H�V�q�]g�?d�m}Eq)��ZAM!+(Av����������fv_�3�@D�iaS���R��2v��j9�c��n����y��Хw�/��O�Qvy��ф,�rX{h"hQ_i�|��6�����EC��q��4�(��ե�ܒe�Jf�{i���L���`%��vm��� �t�rJ��&�d>|-O�|�0���
�w���O��P\�5"3��n�o��K�_��
��/vW�ʲ_��4T�*��(��:s�}��4���=6PJ��4*\�[a��.��QE����ٌ�p�n�O�>�˺�)�wn�����'t��p����R<��#��z��w����
�4�G���d�H�p���K�폧LF��֛X*�n�ŗV����!s�
�\Dh��q������TD�̆��e��9�;��a�j�����I��\��.��v��fҢǒݙ���������D/����]=G����h�?�9���Yo�{e'���{=;4�x�����!B=6G:�l�AZ�������%\ì�²���h��]���,���_󰃽t�����bk��b(ZR�8<���x��)�s���~>&�C�@�Rv�\����̬@���@Y!|xx����Ɋ`c/a�d�9���|^r�p��s�p�tM}ͺr���j^�D�틲���&�$擔nb+eB]F��뇌���0��E������ / 4 ��p!���h��E��m��J</'�����⪉1.s�*ՃS�;�Tl}[��P�.����qV��(U�"9+�oS��x�L`��7+�N�P���� ���]/��h�E�,�D�/�� ���ם��'��3IQ��ƹe_� A�0��{Q�@�>�k``���s>�C�:��H#7�YUq�"֞=JX�R5�B'�&��"�f��b����G)&��%=�:&ƚ��[5����_�}M�5iii������<~̀v�U�z,,�0�+t��]����Ⱥ����н��׻'���TC�� 3�3�cjS��wl���nW��E��l�*V��岇]R�9/@3dfEE�/<Z0o<C1��t�N�."%~�7�?C�m)ÅG�v�[~��ɛ�(�;/��-Q/ �[V�c���0��P�$��ÏƧΒx ����U��ntN·ER!���[F��Skh?9����b���[R�姌7XS�O��=���OOO����7�OُO_A�}��/HIx���Ø�4�a-����zh���֟n�D�0P�څ�˅�B�Őb��3,Ub�Q"��ng���G9��8��8���+g0@��Y~�4�D:������(�-1��K�3�g����?��&��Z/g*
M�=�Z@�����<��養M�TTz�������E"�L#�劭�'q%Cx��Y4������lU$�G�Ϝy�lx,���t�Z�mp�Aڎ��"t�*����zib��@wԙ^�w6�^�G^��w�vך�'���:��-���K�j!��'�&0x(�?����"b�I%`�M�F �"7�˛i���(���1��1j�Yz:И��"�{W���L���M��,��D�e�'���z�	�@f����b��B���:�S)�H�U2��D���F�����>�m"}�C.���W�g{�^9����M򲯟gNʧ�l(�ULkL6�O����C�a�L��`�z��`dr	��.
��(��ۮKc�72o��Vl?Ή.�S����(�z������%�-u$e�����E�\�`!�&M��\V�����˪Z�;I-�h�a�N�<z�	t���8=�8�`���[�+&�9�UƬR|(FX�O�	�<�2#��o�P�AhGK�i��z�ڶ�x��ni�o�Dv�/���[���==j�}C:�����Xv�WY�4����{6Y�b�V��Ֆ��uR��_%1�*E�*}P��SV T�'H��IM���RA��m���%6ψ.�Fd��x���_.-�J��"�_ϕ���3��� �������8==�����I�Ѽ�:��V�����C�Xc���]k.��M�|��ʭo��(ͅ�>Rq�&qQ_�r�}��������j��'����R��%��F��E�m�oM���5���I~Ӛ{�Q���фC���bQ����r�8ڑ1����rHOh�πqI��u	����T*S�Nꞽ���>���7R���~B���!P�>�k�����8���'Q�y_�~�4
� S�4ꭙ�od�����6�B#?gYw�5�^),:+�g�'ާg������3�a�<2)1�/L���L�7��A�В��H��ee�:�6���$8$��jH��Bu 3Q;(!@���|��pqy93�����˻���y��,��s3�r�O���� �4=���T��HEJ�VM���#��I�M��Rrbַ��$������$�����奼�������şn�:�Ό���=M����]$�x��-���2��x�E���g�x��� ���RR�5��kI�,��k�y��+?,	�o��i�F��oyo���>�����b�a.�����2�!��k���l���i.H~ey�ok�X�iъW��髆Zo��P��K�����鶉���hYG��^��)����jE� x4�D��.N�=���M3�▋\�E�F�Fߍ��|�{�;èhք|�Hg��1�I*��ߑ]teJ5�F'�-���3��Q�`��W��֖C��(�I��k[;x��f�����aM�,����o{^P��Ǝ��`���*ȅ�L���D�������9q�-Z�l&��L*�v�p������aEM���@Y�-�σN.�c�/G�Ǖ���+v��
�$f������c���b\ =��lH��1��i������Ə��o�k�;ƽ�����*�L&*&j��c5J$G�'=ۙ�Uݽ�ӊ74/�xg��t��8�"�)��R�D�)���c�O";����D���|��\�N���Gy�{"Z�ɜfѠ��0�z�%�%�sV����X�����	ƙ	�`z9����b�I��'Ƿ���ǫy�s������
�WV�U
�!��H��X�)֭7�Qᇔ�wcV�~�>�V.���'9LH6�~�H��=o(J�2�$��|L٧�~�=��S	�j?�^m��{����ްq{������+-�~�֦�CV'��&e��uɻv�e#��cќJq��X�8��r�`T�`d�@8�xL����X ��c7�
dNk:1)\
�IzN�a�]�x�eU�<�|��`mbbbd���NDE���J��U��|����?9����_X�/YBE�Q�j$f���>�Փ���Y�^�Ѹ�,��2��^TٱUs�%XeQ���V���>���wn2M���?>���d�^�U)r��;�ј�	���Z��	����ΐ�Q�P��ɨ��0�~�1���I:zS���5��R���(9���e�i�q���h �p$�p�@;+�%`yr���X6��N�������n��d��fx��� g� ����ߖ�K�2�IfU�h=jQ=��|d#���2��s�z�Y��+�ڀ���*��i��=/ӝOShE��6ή�o�)O��� �2�{+�g"�~�PH\}y�3p��2M{��'�"�-̤���tt4�
��8�Z�Ý[���C~���iBԸ�}������g�����_`���p�e�/��*(��JW�!מ�e!�2����'�sU��7o��)�����IT�f�'Ε�%���3M/fn)�������d~V�kh,ӅB��rd -�U'��@swԄ�;ӽl��x��D� �l�]:��v*��~���Ϟi�C�5�[�� ���u5C:NQ�}QG[��Ӡ����&�ς��;F^���(ﲾ���O���u��8�-�?�`���N�!��s�c |����5+*3���!&��ԓ
�t��,#�		��yX���LV�ԯT��)é���FГQ��Z�(��G�PD#��>$�1����Qג{.��~y�._w�{��5����1���q����{:�y
��p;��z�vA_�{z�C�*��4C�o��l�'������]�׹_O���/�Zr>>�81���d�_9ю�
շ�Pc�	��ur_Z��/<��@�BF�`�I�YXL6L��Ka�C�mPBs�%��q���򁊭�df�ikЎjю����a��cL��uK��6���?�]�	��
�V�JJw��h��r��y�����Ċ�Π|lj��N�e�������-��E������Ђْ��3AspN�	4�Nw�%_iԭy_��Q��A�]L+i�M�a���T�rjrӁ� �l:��ky�U�ڜȗ�"V��[l��dP<CI�|�� ��#9�����2 �c~�G�HC�P��ƴYs�MӤ� �OQzS ���:HZÑ
y������௕⡒吔C�7a\��l���`4���c��+�LW6��vPJ	a`(< rN�6�4?XV��%:��g[�1���v��V�'?�+��O��o\���Tg<1ˊ
�f&nj�tE=�B��9U!JpҶ�v���L�m��Y{Y
�rp��eQd�8�?�T]T�l�MfI��6���VwP�6�S#K�42��UG�oϐ,���@h��X :c���#�1�N�a��#�A|�h�z;���u�:K�ƌ����sC��F���F��N��w{�&��R̛Qb�j�e��丹6Q)�>�Wo��_=�*������w<�@��K��͗�+_�o�[o�֡K\���������v�l�`���������5u�M��5y�R����z|����󕳛��!���q�ê�I��(���}Ӵ�],�ʞ��a��ջ�c��e�ն��/[p߷l��l�L���
�'�Gb���J���h� ��V���w�ݫ@��F�?"aK�[=��x��A�H��������/��'�����aQ��ؚЕ�ϦG��H,e�U�[��4�O�B Jo�U�A�ލ��sm�!�i�CO�|JE����N��ϡ���x�$P7$?���Fg�c��������67����YO���_c��q��$��df�w�����#�t�ߝ�� w�ԝ�)lKy�W��)��Y��D��q���C%?���S�U}}=99���jӟ�v���$�~d��H䫃c}�;Z���'���.'�����V���_
^B�%���/+�cnFjnY�(c��ǧ��z�A+���1�$��#���u/kJ��QH��Ym\�Ց��ߋ�U�M�ʎ�#�ʢ�τ~%�u?2Y��ia,"��2T�H��&���s�i_���bau��V$����T�889Z?`&?��Ԕ~���~#��\$fb,���@�E3��Ӑi� �3�/9�)�+-6ׯ�f�I�<�O���3�w��7������i����ɿw��Eğ��Z���[��|�$�ggg'��WZ����n�_KO1g�n���б�J{�`N y���\%.T���}i�=����=�3�ېu�T]+�_+�1tP-�at��`ڹ:�aB�\���09m=���5�a��a��/�&Џ��{P��vm��`
)�r/�$%���1�{b���uz��7Ɂ�l��YJ�aY8��!�� �x������S]s�ѥ[B�LB�.T��\X.L������U��b���V�F���:�ŵ0���%�8�n�q�'���uSvcWHPDS� ����B��,�T	��2Ш�咚֒��;�9|�-�2��I8�@�ޤ2�I��0i���$
e8�%'Z	!�-�h˓�:U8�m��>g�wy�b����8���}q�sb>�G}���������4ln���{�f���۱������|BA�DG�DQѼ�D:�v@��VY�c�dS�t�ȕ@E�z�Y�1���Ň�p����l����9At��f"�%9�9sݲ	\$�RTg`���Rm���9Q])��7�+[���/��r8��~��c~��y���W�wfQ�u�r��3��9\��Y(y}������.��s{��-�88�#�;1id����1,��r!{�>��_�F<ű:l4���{22��[DKˠ=J���b-Mg9+��b�b�M�����b	T�Q��/��|��-ޫE��yv{u`��0ҳ�3:��m2>k�7�Z�� J��b=�IͿR���F}��\�G�Xr<(o��"k}�%�\ZZ���X�����#�����ё�(�V73���%��h
�N� ��/(���sT^���a\�}<*��^�����l��2X��=\����	���ҟ�"H,��]^MfVB�Z�D��ByT�E����plu:�9��K���6vd�)��|���]'�oa��jƠT��p�\{9m����i���[�%!���DG͹�	/���sU�t��]o��������ͬ��;�Z8��� o���ԧ��(�j�����T'��s�ڧ���9�Ni�� ��s�~���ז@O�4�Y���3r�V�"U`Z�������"X�>|L�q�Q���r-ͱ�􅝬u�S4-��:%�?_��*��ݱL���PT�|n�f��I��(�I��MS�ՆS�=`bq�g|xqu�qb\����T��*�������	n�]|2?5����%���CK�j��1�����糷�����}�6����HV�g2%�	+��<IQY���ږ�\���Ʒ��RZⵝ1猗�Z^6��^Ԝ�t��t�讐�m��C���|/�s�pJKg^������Rj��<F�j����{r�i�''�-�Ss����[٩O�����	,_�=�g?=�~.��Kg�~�
��FYYFF�����V�Ne��qwW��t�c�������X��#���9��N��/HC�#�[�!p_M���e��/v+�}���K�3S�3h;���e�Ԋ������@���������%-�iE��9K<u &x*V�νg�}�I	B��I�����ƚ ��7/e�W��p�3~.������x�x�/��?ҿ�Q��+v��<[g"�v�_.&�F| ��}�0�2�G��R��S�W�4��{֟4f߁��i]7���t'�K�T!�o����S|Ȃ�^�Zt�'8�b����bJt�
��yPpHj3���t�-�ɻ�p�J덀4~���f����\�|$r�&���Y�&�*׆t���&m��	i�7��E���^��͐�a6�n Ti�Ǡ$_t�v������$4�$��o<���U���	�T�Ezy��������3_�6r-�E��Z�}ui�ۓF^5�Ufϵ9����)ɗ�v�B�)�}JI^��L��񎰭1�<H�P� 7�I�l�!��M��I�;�Cs��썔 �X?�QyH1��h]���ɽ�L��y��<��z/��?x����z+)1�K�񡸦.:,��U�(,�m���lOf*�3G�qD�0��"��G��U��hۥ���HǘM�)�q��*��9<��r��u�#x�5^܌4�
���M��XGb����Y�J�7���=�ؚR:Z�Z^RO����&4*���N�ґ%������l`�_%[T�S*�ѽ"��)X/c.Γ=��*�ƒ��������<7}��V�ƛݮ��*�~��7���P����ë��������WQAAAQ1a���b��D݀ �3��̪8�����g��앣����$#?>8��o�f:��[q�{�q����e1|T��y��Y�"�,�S?��d֡_�ű ə�#�ݳf�'���C�Y`|IG�MD���I���I��%�7׻��כ{?�rQ/!��v"�v����QD�$���BB�JRT�M�:��.���~��o!;�!_Ң���6�p^v8�N�p�d�s�}���E�g�����.�`�<ǃ*ڃ>�&A1*�mK����ns�_�QPEG#�b�fl�5��aL�`g�ݓ�=�j��e݂Lϒ��J��iu͸�!'z���FP��o��ﶊ�������nB><M�
n{(
h��Z��Q�ѽ�����C_>ߤ���#xE�{�~��
-��̘�¦�Ƕ�/'Ku�]G+O���'+1�'M�+-�`����
�9*�	�2~ےS���0�¿�0��k��keu�u�����c�B���41�Y픋ڦ��Z�&�L�%��>�[��{9U��
�s������.����������q��w�����^�����u�cE�dxH{���k�0�����ӓ	I���5Z�ݷ��4vl�A��&������M��C�s�o�o�oara�k��D��O�L�L�q0O�G5.X��}sY���^8��?�����$��%_,cs57��
eY�k��9l|
�K�wh�Yi9��0^�D��j!�f�����H�<8"a������N~��Xu�6�	������8�]rf��rv����,ȉ�K�#&�������j����(t�bE :l(D�r�f{�M�����XF阎J�:^��Jh��S;eP���
��Y0s �(�p9��-�mp�����1D&� ##�m-�f��a>Z���yz��7��g=�M
� $��W,˥0����>?Hf6��X青v��U���px�{��o��ӗԉV53+TY��!���$�5]S��Y_d?�|����'F��xl���{h�+	$fQ��Y��"Z �e�D�n�઱hy�"�H❥�Y��$�<���D��3�����$��m�!��1��[������39�4��1 :�L	�fH?,��[�J��S�E��Y�w�a0	
��M����p�M���z/�K�'"��աk	��C� ��Q�G+T�}
�<�d�۷\ψzz�E���QZ����k�_���J�����]�[7�]��X�=˜4� ]?����\�י>��?�En��3�_>_�	�6�E&̦V��;�������HS��w���M�	�y͍!���`�X���A�:Ljta�$E5*�a��6k�������T�A"� �Ǩ8��	C���	1."�~x�,��������4�臗Ă�QH�u4鹆z(�X/gQ:��R<���U��H� '���7/I�5B�n*h���d���0�����O,���A?���x��Jd~7� ��H�mC�hĨ���X��X4n�.w9�So{(Dk�4���Qf�h��Xd4��]�(�«�	ZL�/w�uG�&���d�d�:n��r��;�r�/���5�8_�Ϝ�F��n �Z��K���Ҧ|���|_�%A�uR	,�W%;��	��&c�Iͬ*�s����m�N 8�D�s�����o���٧�yqvى���h��kշ֠��h���r���C���F^��o���}<�����~,��.Nmyej�W���:����F�h&x����t��[@<�4j��-��g�3n9�ڎ���Γ��_��Q^��-Ĳ^��k3���ۣ���-��\4h�M8R�<�X5�}����8��V�SK��l�X���!L�At�QqH(�H�)����#jr�F���x9|�� �����U������^��1V.��M�4��KQ7uζ>��	ۅ
Y��E�*�3�p��f�:Z�0^w0�r��jp[��&P�v\'.���ȹ��o�]b�'�۩f�S�$F['�[�)�a_��]��-�5����qy��VUx�#uk�.�?�۵����������'��P�y�eY��*BUn�E�#ǚ'=E=Khv��Ygqx牖ޘYf�<DJT�r��=Ϳ����6��oL�	�����S��0.�\�()��w�P=MJ&~23o�*:�h��b<4�{�Z}r��X�	���&&:�_%��=n�����b�D�2��c���2�[l�W��@�X_��I���?ξ�J��|�d�!ț��n3�C32���Irf�����Q��1�%��.$�v����'���}S���@<+���r��q��\�V�6%!��G�B�:bǁ�k���(i��Z�U�Rf�� ��6/�ϝ���J����}�?u_�����\��LkX��
��|�8�~�q���yR��q�rb�x:� �w}����v2�����iHPm��Z��:����ͪ:��7M�k�nBQ#�Z��7��،}qqqq����Y�k����l��m���E3Q7P^��G�����x�\�]J�s�^N��
SHӸ9R|F��f��G�:;��M~g�e��5�1��}�Y|�[�]���-I��;�t�k��6h�4�[̬
���]twh�K���˖�4$�����y��~o�55�Z��[�`k~��I�#�a�������N���a���v���6Q,�zܯ�r��R�բC؈�}�Kg~��*�E~\\\VV�i�;0��x����V��]D��tQˠ,��EV9qE�w���U�і�������^*����hƭ>�6on�ᡨ���U0��Ϥ|��$o�P�����H_���E�i��ݓ����Y�7�^����~�!�_���Il1��ϥh��溱R-����7��i��)	wb��"		����G��.'(����؉��������+M法��D'�F��'R9~VA�?�/TF)�P�f�,��C��R͢?!I;17�>�Ǯ�>�����,�O�,g��K�s�;���t�Y�\S�l��n�w�f���혃��ԛA����b�������e��1jܳs|B��U�r�J�	cPsW�z��rge4�j@�{���J5��?�N�]&S��Ks/P�
Mp�h0��������dG$�+$(�$�?�Fev��'���߬�Ra��7���p޲W�U�O+��꒜@I� �+_��dkk�(��c��z�{2�rK�)mp�����1\�����Jzܳ��.jE�"�>�
NUV�4U N�Q?`tT�*�s��X��F��P\��WO�s�y�ݭ/�
�֓���u���@���o���z)���ͷ�RϊY��
�k�|�|�b�J 8|�b zBO�����	2���&����u���ZG��UT�م��
����ެK��$/Q�@f�/�N�O���J�U�A+��H�v��m��z��#��"D��_������LÎ[�X%��^�Zi]EJ`6Nd�r�E���G�����^�tyX���V�L��SSNq���מ�STk�s�h���OĮ�X����8h�'6L�,
q�x�X���x�.:�(JEE����x	,]��{�ۮ�p��W�{��])�AK�`�b�MS�� ���m�o檭��[5���>Qgo���,9���|�T�?�%�ƲX:�`*�"6ƺߵm����A5'�w��]�ߊ�8-��\��M⁏�ѽKqO������C�ʝ�����9�ն�S��iҰ��G��q�2��r0T�m��|v�	��i�����6�_F$�y��}_5h�h7��P8a�6�:�d��3�%�O�,�`�/���a.�cG�}��΢6�W���d]��Z�F9�?�0kK7a�$�^/��9q�ۨ���������jp�q���FD��[O����]�ENp%+E��g�b�x��8�"�"��TL�Ӟ�Z�p����ԲP���2�\����.��0����c�$��^\zT��CHt2��2�F�~��e��'��5��Q�ڨ*\\e��s�f냛������8��hY|a��������H����=�ǫ�^$��tV�V�-�J�o�Vl�NS�۬��Ic*V �x9L����|���X=#��/�4v�_��i�u�v�Tw�u4��W����^�v^u����:Y��i�|=_�5����ϟ��%�.�8�IAu���9��u8�E4����e�������?^e���=K�=uڈ��puE��v�=}�~~xwbp��C!�pgc��0F���g4���t���������z�����E�׿!E���}�;5���Tok��ab|��&�����J��M�?��d|�{'d�y#��/f���BWW��*8&��L���R��;�+���$�EX�&��v���RE�ΈBvx����SX�۵,2U�%�9c���T	M�*�=Җn�i���ך.^�_۷;��^��zX㐧�̢��L:�9K�xWD��{Ǭ���S$�"..���� 3��>�7�D:\,��%�;��Z������e��q��'.3����qˉ�Z ��񲍱�1:E�*飚��	F�ձS��x]��^{�;��Z{�w��t �M%Ҝ�g������9��0`FI��2 t$�2w�J�Yp�����|
���=_70��(�3�~c� �@�e˱C�p��r�,�D����$c8?E�p����JC� W�aH�����D���a���>l�v�

����1��Oc����#���ڂ_Y);��~�+M�敮��N�c.װ��%d�R��L �A��:��/����������dȔL� lw�8d�1u���׍D���|:.=&P.Fv3�|��}t�$�e 8��w�	��<�y2�����b��&�F��ctq�:�In0.6je�-��xoV�l֨ʿDYb�5=#���Vhb)���jxLy&�
�f7���[�JR
y_X��m��d�3�z;#�/�D�g������e_a�<���r����ʤ�����=ȵ��d����:X@�``��t�r7e{���gߓ/���̦�|�����]�?��V2�ǲ^�����t�1���Ci���[�e�~��E�i�V��wDD��ͫ�V���ElXe��� x���_�ϐH����w������Ƹ-6�@�4_/���|�x&�9��-��#dP'O6��!^'x���x�e�s6�n�~�<��w�����|�]��z��D��Tz�_��CQ��ՕK凯�����	��	�D�@jr��]�6����;w�F��m��j���'
K���������<<������������鸙��M_���m����:��&��:�-JMU@���98�Ŏ[TT~OPI��|8
"ռ�� ��~��)�'��q�ᚯIڢ���*���7�??̭�)X�O���^�]���b/�����z��)�����X8�0t����t񟌤:��6�DƦ��0v{,i&׌�`�+u�H��XWF�� ��v�ir�m�����tX0�3�(fN��NlWV`��R��v�, ��ZY�|e9�kj��'G�3���g���)���OmJ�7�1�沮R��"�䳓��<��YL	��J�4Aq�'�j^<<��_9�(tz�@�i²60�c�#���� U��:�d���^���\���Ȋ��H��_��*���}�/��~���K�� �d&��`S+�DJ�)֫�5=P������_sE"��\Ŧ�F^r��"Z�d|�~+�SU'd}g��Y�r�ܞ?_��O*�9D�'�'f�ń��k��b�^{8���1\�X��x��l>�~���y��-l�k����F{�c4q�ύH��7"���4�IE}�Iu����+�}+���ق~*9�o����_2��n"�W[.r�=�Q��^?*��7y�L;�{ߝ��l$j��n?������l���5]����*�փig �����6��}d��+�jc�~���O��T��o��pu	*QJ5Pk������l����&o��%cU��x�/}r�4x<�u`z=~JWǞ�"K����2+k�Ee7P�ur���rK��g���+��Ľ�S}�*y;��-�{��=^"-�sz���n���b��x���ω_�Ͷ����hÒ3n��ڸ���b��j�_Gaaa]]݂/���n�ꐛw���!.�76�p`�6�I:C��T^?5.[�E�F�y:$��x3b�j8Y8�l�̢�7
��q<CY!��T�R��R�@u<���΄�(S�[E�In���d
}n�(�ߨ��ޒD�X�=�P�A��bC����
N�`�����8���'�7 ��1�m��`���p�f�� �%����7�P��ҾzM���myP��^])�Գ&l�_��� ������C}eC��@��a֯�ur9���@<�|hy�]��������s|*F�8`�)�]�4��ORfn�v�sQ����E}�|�:�S�U���N��e�����Dé��i������w���
4�==?'��CG��{�����~�*(���K1 <^6��3�+(��v^j�f!Y�B�������� ��pѧo��Ug��iwG,Br��Ȉ�;�s���x��1xԙov��Z��
��Ѻ?1�������� An�d��&��qw��+�^��z&q���b.�;�oE+ńn���)^S��Ehq~z�����5%� cB\Gl�KpW���K�]�'�?m��y���k��7����T��K�b��r�V�Y��
��X������[�������3�C�Jy@\Z�k�������1�ӑ�Bl�D��/N�L�S�W#�����{m����]�_~b>�,�LIU[K�9e���fc�$?ߔ�������Yk`�}w^k��F��o����%�(/ߒ���`���!P�j@���3E�����$�����=����Y��7\-�>'H�1ͦGM!��3��o*��FQ�F�y�����H��&�#	�9Q-#=�R�@��+6G��O�I�����	H$���28��>�Kmfr�0!gi�|ݮӧ�����zf!�+OM�G����2y�ojd�+q�l����V�Xk,���C�1�WM��]g�oiuu�ZL��")��W
~��e�����w0����wK	�D|U^���+w��q�����C���V�	�JTG �kщꊓ[�l�E^lo�m�����,V_��D>d< �'I���ߘ��/"�Kk\K�����'fv�*��0b��Dz8I�1��N��;�?Gb�\�ky	XBg�Z�ҐZ���!؝�Â�*��"|��_4<�=�|�_���Aqv�";���z�G૝�\�d��d~��.��J��k�Ԅ�O���k�����������'Ee����#��<��=]h����q>.��~�st��w�Fe-�r��~�h��t��A_
�r�wi�m�<y?�����o��u�c�El�a}�E�-u+����E�N�U8FOw��$������g4�U���ԭ�<��Z;%���?��]��������-�8Z��n��V?��Hn��M'BHe����aY+�+�����%D'斗'g�'+��^�B����-0��d>\��𯸭�.�/݇��?n��Q�ly��<����e�Bj���`��0Q���4A�4�#�e��Y�@\����u�#PC����<�鍣���o�l��#T5 5o�D����D M��@�g��a�.S�b�`�d� IT��2)t�i��V�,�H�Syrc�@':��	M���[����P�@W�I>J�Aݬ\�����=���!$Y��oI&�	���/8�C�)���U��?��(�[+iξ�I�� �i�4��qF_�2A��?�ƃ�J?�8���"�\{Q��`�\�T��v��˄*E��wࡉr���!�¢z߯OH	C� "  �#HÐJ)_j��n�n$i@�A�CZ���F:���=x�k����{�g��y��/�SA�NU 9�gqx
u�2�>��� � ��p��yM��r��P��ė@�7�jB6���5nմ���
�Э ,.PEX���J�s���0�@H�F�"�QRPKl1u^�\3m����b
�R"�I�I��n۝3������R�x��,'?/�����|ъ��_z����� �w��ץ�߇J�h>�Hl���=�A�yWnc�|�vB�P��ճ�rӄ]���8����H3��:0�=@6M��w�4��gϷl&�0x�{ȑ�6���W�j��]�� ��z�����u6����C�I�{MŅO;w���mG��F�/ȱ:����sy��6��i�0�,�MdB�wr�A��0
�YQ��������u�XU/0��$�����G%}.��<]�X��?��̑�?=��2z<)�A�}���vsw�ەy%|���S!y5Fv.��B�!�������	]�������vUJ��a�r-픴�-k666��@R���	��*'g]�Mͅ�q�7��9� �u]ଐu� �I��7"o�*$�������}W�~��:�"v��fv��>y̧(�G�����G��{4Z!�V)�#�2���ZE��<8c�xޔF�W��{E����	u�������`"\�Opn^ʫ�V�D%��b|Ǵ���чOts��:�L|_T�"����a�#j_�<�O�&�G������ւS׿F��&��M�P�����ףpa�|�9��~:�+�ڋn�g}���w�yn4 �Y��;���P*N�d?(��>,��o.�<6����h?6�h��V]P��<<�I�E%���Y���@��(�]���0��5��Ӏ��_Q9i?J������@�:����DSWn��-���
"�L|����̷C�W���橷F?s4�POz�Z���e(�yk�K��
�ܢ��vtK���%ψG<��x��z��-�1�7�M�	����YdQs��8��sM��KS[w��k\��PFҊ��be��J�~��ֲ��.￶�ls�,�pɿ:�`��ټ�X<ϸZ
��^yؖz��4�{�x�@��x�x��9�|�B�_w}�i��6Z[�h�L�n�@lD��賑�&7m^�*��!O�:�N5���;��L~�#�1�C�C!+�qKH3��ʯbDUu�y��X��X�\~PP֏���/����5W����y�,����lV�Q�:�<_D��C= "(�m���~������)g���u��|#��3�X��^W;���!�.}�����[Ù��sap쀡��"	1e�a����6a�P״m�x�����,`(0�|^3�8c�=��c�+7�����C7Ղ�Bq�5�7���&�X�,;��bdq8I�k8zU �ٟ����mm�ߣw����Z���
!,<��W��k���NE{��׍�I�>��y���y�tk�"�Ȼ��wl��'4|�^n���؋ń#z�,]�^�"�M��/�6������(��A��i �pF� ���,�[�����M�M��)� b���TbB�0H[�ݐ6��wc� ��ꏏ�<چT�;�D�����C��$�vT�-k�6�TQ�d˯�Q��VM�6�^e#���:Uث�a�$�r��5���v��-�rn�`.z�26�z%����0~Pw8��Yz�6�[��C.� !�=�VOhS�VE��èr9����{5&^>�±�wR]� nΪ���h��t�!���z�4d��B�'�}�׫�q 3K�築с���'5w����w���.�:���L?�{X��h��p���� v��W���[�[�[����Pn����7��Ҏ%T�j2�S������XT�z�����#巎ش�1H^�F\�z�9�	<Y�Ll����ɀ�E`0�>�vUHz���	�?�1V�|,v�䕒c"<��m�3?!w�O+g&��;@7#�O��������_@@@TT���QB�&\��א_�=�����R��D	�q��:���	WP�֢��w����զ���a��T�O��7�K�-?�*�m�2(�7���)o�)�:R{uS�xU��!�V���U۽���[/Z�� ��R�?�!5\�2K�~���@�s��L�oX0̚�S�i�e�8�Ц�L����E����1��k�����oP���e?����o?0��@��R�[bn����&���5����D��<�AϞ��HDaUP^4iɔ<]+�RUA�^�HX�+�%�������+�c��@Ȉ	�2��8 @������+æ����Ii
�H%A.bju�O���|�q/~��
��f�C��i�jw�6����s)�詨F�i,QZ����s�p��oJ��G����܄'�WJ������%�<�j���S<���o�h�* �
Lc%3���~���8��_�t�-9Uۤe�J�\������b�F*r�_${�F`Y����F�[BÛ�	U��a`^I׭3E�8�'G�WK�G�	&��1�m�[�Nm���Km��}ˁ7#z�O���ק�f�[
�F�o�E$��4�;{�ST��p,��,�!/� �$��w��2�H����B	��"�794TX8�j��jr�"U�	�����+����:�,G��
�W$�����D@!��D_��VQ�5�¶M�[_�6�V���$�h|��싖A.r`j�m��T�i�ݑ��h�Բˠj�-���'��p8�����gx��/ʯo34��y�'/�SމxP2����!�>��E��bc�ĐTA�p��+�*�W>���x  HP*Y�8e}������C��AGQ�����D��e��MO����7���M�0��:ǘ��@���R���P!U���� Xh�{)\�JG�����-����Ы���G�Tÿ�ʪX��>A���@h<�6M�~�?O������C#,�P�Ϩ�~�L���F�E��+�`�,���v�J�E$�`�������U��D��4H�	Z��;��`�����t��nq�,{#ǌ,��ͮ*���$���+�x��th̷�Y��A�.7s�R��Kl[;��g�����kEdS���H(�Sz�1Y4e(NI�ڝ~�K�xBK��{�wA��j���o�k�pa&�.MSwOօ�����`��$h�����P+zQ�!�{���ٙ�磧 -��T�U�s(���p�pH3�i%��tgV'u����bgXl��Gɸ~��M!Ǯ��.����h���N�Ќ�����Ƚ��쾭f��z��{�3a+o���	�y)�|k�Bƞ6��#�*��>�#G������@CG3�ϊ��
�L�v��H.
������f[ɛǳ�v��nu$Zq����VQ¯ۋ�+����d|2̒�/3˸E�b���!�K�&,,/���dk�7f)6{��:?ߧlt���Gv��Ŧțۿ�w���9�5.�R]�p�M����z����>"���|>c3���5��=����*ų.�D(���-��沷�L^ֱ��I�Gy'�y�"Ca_C3L�Q�ő�ߧ��{ƉC����g]�8\���Xǝ%?L�R�`|�X��E�����-���?I�;a��:TT��~{	ꏛ�;5E�9�p�����uLu����\�Z��f^@"]�K���b��x	jS�x�I4�C[Iz4���g2��CKG��2wF��H���o����؎cGh/ǳ���+�B��2�����~�e4\��s�0y"l@�ĝ|߇�(��Q�g[h�G�	�_'�w�c
ߔ����2}���%n�p
���&���ӌ{ē	����8�����r�6n��ɋ7e���JC�x�okBZ�B�!]u��j]*<�\+��PNjY�JՅ���!5.�~V�~w57��$:w���#�"Bc�/���U��2f�5�s�%�_��b�����C0��.6�쀋���,���>��k^�V�ݬ���q��b��n�_�_l8��]~X?�x|��Y�=�����&'po!ò�=)�
�j����.;��_����C��ZA�38C<�r	�er�BmИpS���o	Z1)4��c׆m��oOV{�"t��Q#��Һ��){1�G!�|��{�������+G���w�{A�FG���ʄ�7򉉁|������-lm�_��:�)�C �����{&��@G/3�gk�Ŝ׹��m�����r>- �n9K�-W�U��#8ܗ���.5���0S'@{"��v6�Kd�[PZ�]�\���@7!���* ר�?;�_�x:�^C�;��bK�1��mx�;&D����N��vl'53������S�S�-&�����}�DS����;�5.����B�N�_����k��PZ�fZR�=����!*U@�4DN�N7�ލ̅7QB,���2YC�d۷���r��<�'�A���Ҩ�eEE�v�2�ɕ2$�~z&��1�c��[S?׻Y��`��y��Z�Z�.��� ��8��$�j��MrP��.��Ge����r��h;�.�q���Y�=����>�����WJ��~W�������jᥚZߐ0x-�`x���� �'�9gLTqdL�j7�o��@��*�y�aM߇/c���ݨ�đa��3W���Z����	��k$��j��>�@��	�Z�2�lp]���`D�'
���܊�R͓;��f��MI�l|YR/�D���Q��c-6�z��!DQ�ll(�G�킑�u��*�0s����y�Kv�L�ɯI�=�(Zͅ�@0[4�}TU}EA:�L��Z�l�zEo(z� o��.opx��9<�g��y�7�g���/�����w��X��M������l$9$�н��n�/Oy\�͢�zge�� �{�lc��l���
b	v�S�� �������������;�H�C,U�Z��<<<���?�iK�}��~���O0?��I&�2��n�#v-�C �v�G&#-ao��<|f���]�)G����=�mh�J�8��3%��4����@ĚO����:\R��1L<���1d"cX�Js=���BP=A���t�02᩸xG�h	ǹ;c�.��T��^T��{t1��k�c{�5��TB���nU����W@�7�-��=��_����ִ�F����$P�tY?��_�a+B��o����?�m�dL�b�"��7i��I�{����ؠ�@n����"�������;�WZ���$t>���j�K��d�f��,��c5\��ʷ�B&~ �y0Wcg�T�󂳫^E��<� h�V�AӴM{�:��u�z/�{����u���b��R��R[�P󩾡���_�	YSd:�)p>u��C�C�۷s������ҏ�ٟ'y�@���3H�`i��ڌ���{][߽4ֻ�o����n�
����7C<y>LM��ܭ}�} J��u?�g��;���t�����a�W���0�ϋ��	E>���t���HϦ����a���2��Ef��V�,���cQx��Ÿ��\x�����n 	$dO��,����������_6?�(6��W_��G4Zx��{;A}�>�9�2�������o�(�mQZ�m��Rm�n�{�x����qo�/|��*[��/����6Aj_ �X�;����	�]��=��;�y�
.�[;�n����G�p<+S��(���r��,ȺcƊy��pX�ޮ�jMx�yl� %$W�JⓍ~�ɎWD���B�4�LW��\"��"�d;��j!��f�cn��F75FD%�)$D[��#�"�]������UYX��Ҫ�5�L��G;�� �w��z��И�f >��Rp"X(B����W� ���V�M��5�l6��L-Y�h�hg���0��ս���=�GeţS޾&	Y�DS���8��50h��W��ByS,��,�J](q����x�y8d?����E�Z�<���Y��e���!�����/�J� ��)�_`'tzb��܊�g@���?b}�3�z=g�N�/�
+Wa�果
#��{ӣR��p0(!�s����y8JwЙ��I�<���]L��ﲟ�3>%�'\�[u���q�w�0}��.�����ӗ�D�;Ks ��Lq_v�2� 8!;Ԗ��H#��D���u��m�ڠ��eew%3��/��AJ�)��f��F� F 줹��M!��a�]���=�nK[�Jzq1Q�D�/Kg%f��7hbr����Ѿ�X�@/,ϡ_���lt��s�h��[����:k�|�w�wx���#���E��h��LT���,�3lc��2�[]��"��0��m[|��T���KT�+ox���\f8��T���4�'�n��$�<	��>�i�"kFc?n�D�tR�����D��9U����vt������H65����R[h�NN�7�հ���̈́���<�)�A���Öe��[*����Ru�˕g'CU�n>*:��a��%��_2�1�K��h~�0�,-h�O͍hY�t�{i{}Զ���c���w����z>ʁ��w��"[��yu�Ɠ-��)�%@Ix~Tvd�QΥ��LDi��7�%��d#����)S���j���;Q�<B�%o��\W����hK�� ��m7UqZ�]��5������?߀�l��6k�]D�Y򳵠UEI�����Q���V�2���4�l�X�V��������,:')A����r{��R�������h�b�*���]�����e�`r'<�.j����L��[`�H��x���q�;<�a�8a4<:�Bn*�ۯ��X��r�=�;V�ɩ[�Z�ϳ��h>�s`��L�ї��P�X��t(G��a���u�������MG����Y�W���p��V��:�'�Y�ߊJW0wl_&��������бćJ4�������'Z^�Rm_���3� /�LID4h��)D��%>Nn.e��2�u�w�϶Wd,*]�0I�B��?~����A���),� �!��>y��\������b�&�/aL _�A�B'>�����K�+�t�u<�%�����I���&���m�k�>�ӗ98p�98|��R�/��U�<y����j�}�	'|?.ea�	{�S��V�������+�ذ)�l�����k�Y'�w��%�\���}2����l����φ���*ɻ;�e���+)��uu��y���;S��k���ѥ۽c����s^��0A��L�o@ ���1�5��<�ˍ���3GB��nN9 �x�Ͼ�2k���׈���� 9��� ��e��:��h��D����ؤ���5[b��gZA�Ƴ+Xe�/,�gX&���lt���';������ǳ?��1��[�;zI~p����7mYꥥI�mmT�ߏ%�g��m�b��?'L+���RY�)���$|�\���&�[b����b��֫f>]3^�?ݨ#�vl=\��O-"���o��7mg�f�Y|z�8���]��;�:�u�	�LO�8��k�Y螅2z��M�Y2�~�q���?��?�<y<k�΄I��W�{���F4�&N���ZHġ G4,�� `,�?���/�P��GS <ITO|��S��= x�����x�5��M-�;K|��A�`���"����0�^br�ė<�Ey���J��0c�P��Xv�'�Ū �?U��s'�����ЪK�a��"*Y��]��s���=��IDc��0&S����R�)ٸ!��4q�ݻ�Z3}U-S�O��լSB����VvB@8?{�b�S�݇s�x7مI��7�8�����[�օ���L����c�#�J��г-��#Ժق�Vp���Q
��^�7YC�DgU�z����L/C�B ~P�H���E�?�+�@��A�ֱD~ŜyB�0`���P���ų��f���ڒ���!�	#�/�u8�8��]����M��
㪪��`g3��������Q9�\�C.j{e�yd;#�gG�/P'�'�R��~�x��G�%�� �P���xD^�OA�j�����{Pp�~x1v�E�4M3B�_��k� #4�ר�nxs2�id�2�!�����ٻ+a��_����U�@��b���v{�;S�%�Ak����/�G��]j���$3og� 5�P�de 9FEJ����g�n�&�p�9"p�-E7�TT�1��&<��ڏ#sS�Qo0��.�P��c�|@��Η4��"0�Ә���O��k���_�9��~O�z����{z$2m��w��O��5`7�o^��{�Kg�u�A�\ukoIg�#yM]tyu��緼+ >6=��5���(M��hBjZ�+!��;��'4����l��m�af~U�U���r���~�έ�ɦ��]֊C����� m�U���e���1>�L㽛P���|��wJ�%�<�?բs�C'T�ш�AB\��&��At:o�TU	�s�u^�S��k�W������)!'���Tj7���2]qP�L��k��Qr��/�+.�̛��}F������e ٚ��X�ʻ3���w�uctи������"����2�
p�p�ܱ�D�1�$Gb=`ñ��	�[�W�pl�D̈H�L3�)P�f�tl,��[��yӣ}���1�����2Ї���F�2Oɳ������@����'�O6>��C���E��˅�m)'�*@�J[F01J4���/���(�	���1
�r����)�z�$x5����Κ�C���/b4JC�)Q��p��o���!��^�b�u>4��������[l�9��+���.�w#��L���ۘ�5V��OfF�kD/���;��Sh���J] �#r�6"���.��[�F\O��7�N�����`�7�����q�y�[�^=��b!ϕm+^�6�\�1Y�=��Xe�ލ��RW�d�e���'.G�Zu(D0a���>����FWpF)LwB���X{3&]s���SC����2.<b����7��Ћ��Z�Y[<$+����f�;i�J�>�������F��4���g|����YYYC.�ͬ�d(/�-\�=��Jd9D3y���7n�tw���;~ږz���|��$��Ď1�1�u΀�5�A��וc�O߃a�����3��t�h��h�A�q_�N=�(��l�P�.B�j��@Q���K@�s	��^*�H �K�V�%��ɓxd���Hb�.�B�W��(��̏M��jlĨ���_��cd��$�l����1*f[�I!�ڟ��Jv@������ꣽ�����[}�2�dq��/�{Z0N2��r��jx��l��"�'�0��a.?3���\,�EK�P�6��
�Z@����S�6����(�L<����׫p[��6#Е���0ǁ�װ�K3��w!�*����_����J��F,��R�SpV%C�)R�䋆�,�O�;�a�6�uR(�@�Lv���g�����׊p���Z��L�Jv��v�M�����#���,*�c��k�]QݠSV}��s\�wN�����6�I���\�`� <4Q��W��m�h�B�4��N��V�J1l���`H��3ը ���Ф�R�"�ȃ��[Bu��L2U�{_�L�B�B*]���s4\!��RJQ �U�<Q*�5�{G[�n;�+�|�����c�ѭ��&�D�H��L��	��d�_������ď�",��(�m���+���:f�c��
�1�a{�±=�gm�~�[�s% ����gӲ���G#��O��Z�}��ܝ/﷧�d=ާ�4)���
R���������4��+�Yńl}:���b����̒�}t��3Z���r�ۓ�`�L�C�����:��#u�Bc �j���������O͊�&g��?��;�5���Z���W�G�e/��̈��x�p�Z�x3_E��t��}�8<�p�쨗���a�b�K���F�e��A�V� J�f8apƎT���_N�]$�#ʎ`��Z�3kD�P���kb7
L�xst�ݪ�w%k[������&�,Qqa.�YM+#�r�Y�I�f	\Գ�ࢱ�t����a���1���l�G/�}4�''?��	<��4�U�R[:z�h��G�Om�?�}=��mT�@��A�n����hf�Le��xvAb�f�����A�@�����	��Z�	�4��6�*��*xXS��K��<M�V^a�6W�>L��t_%s`,)����¢M��l-�E:࿫�	� c+ɬ��:��j���M��ت hڛ����0`��[7���#����D�������O�P"&�9=ϿFx|2,Ka����y�!�'B��Aԍ��ѫ��D�hL�½���A*q*R�ߑl��/���x�L�����v�t2h���;�s�o��Җ���~^D��?���e�s��7�N��s~��3��<e�.\U�J��"{"���������2N�~�X���<�)e5����`��j�rU��0�0I]���p��c�ͷ�.␿��������h���v>���9��6����@�DO�gfx���޽�1���Ž����Pt��_�ӻ���uR� ?�+Jk6�m��lQ�����oG�IMMv��a����aj�) ���SͶl�4,Ꭹ�7K>突͛�Ѓ�w�(S����/I��LW9m�<�x����]��F��Y�A����rR���E)u�c��OW_�DC��f�'�41F<��4�8۷�<Vc�+<8ʗ�Ґ���1�Xs`�GGmՌ ��h����n��c�(jp�f:�5���ߩ�`/�g�ʄ��r�ҬI�g�F~�Ƅ�J:((� OH��n�:�.�a�a�1� �H�#�^�R���~r���:�~����`��Z�>6���u���U�	�a��,�;��O������L�6��A�
v7rȽ�l�W.����2��<��@m��dO��Ma/�V�)�9F���� 
�D�h��c�c�q��[�p~!�H��Z������<M�tV�u�FTa8�I$���ײ���s4VF�@��v�Zāt���11+{<O��*fԚ�]@�:L���x:�ݢ���l���b9�����;!��5&43WB-��8�u��J��օD��K��_z��k�
O}&�g<��9m��9�Y��DP��Lk�ob}Y}f����[Vq��|�+��J��ODb��}iAHJ�]���1	P��_�eLx|�sʐ�E��I?�i�N��M�ںba��(�pM_����/������[g8_Vc|�s�p(��҆ڜ@��!
w"��Ӥ��C���R%�V މ����,j�~*\t��H�|8R_n�a���n6�U,?�/n/�ތ{�H=�$��i�*:t��L�Xko4�r���@��#���,Y*����dz(I����ӈ�WYּqE�e߬��E6�e�6��&ڨ��W�PͿ�Y��Hi�5��y�b�[nj\�C]�F���eD�K�D�J㨡z9kc�l��k���j����[�\ё�D���܌+��E��K7ꏣ�,u�hn:�4��J$���k���.��d(&H�-�'�3L���w8����!��?׊h~H�Na K�_ͤ�Jc��V�/�>|�6����ڽ���U��h�}7�\$4��>*�<`'��28���Դ~O�����ccB�at3�O4?cˍb۰�߀zQA#�y��&^7I�9� Q�6���)�=��������-ԓ$L��!!X'��c��Bz9ʮ`H�,M~���M+��}�&�o"���Nm��pa�f6�1���j�i�tG_���(�ɰ��	Kňw��V���<F�	mtmj��-�+2���cZ��/F�� G�Ԙ�d�\Ҏd�lQ)������� ��}�����u��g=���LJb�y����u��%��a�&��:gw����?�@�1pl�����8��[�zT���y��~U	,tG����ȗ��5V�T�^���D��x�!َ�,Ѫ�w���S	������A�G�L��O&[�~=����{d��{[���#��x�'�)i7�-�q���r�"�(�4qs�yMÆ�\�8,�i���MFB 55�KB����i{��+��e����%s�F� �����KM��Ί&^�wQt��C���h�L%��������0��>m�\s]��}�i|.��H8��@�w��U��k#�2j;B���~:��Z�����US����tgު��OU��էK��7����duGd = ���%� ������;��Z�Y'�5k��5���Ǟ=�(��g�#�@�2��4Q/w��38.�Aע<�;����e�ʺ�V�%Y�@w�@ߕ�.2��q���@(7�^~�cK`�F�?��	� :�1GneL1��	�~ ������p���D��؍t��Ћ�V�u�!��w<�n^�ǰzn_�+�f�^���Na^J�L"(9#%P��	�g��7���#Ǭ ��LA�]5��"��'|���X���3�� Jhj/�Ʌ5��|����.!��L삩�Rtf�<�������#�0���1��򻂀�/�q��c
�"_��|���h���CB
n��%���f����ܣ�n:�eL&�k_�6��7`������N�	�^ǧ��a1ʓ|9x�Y]��?*�~Z��{��`I�i/�����w�%�)���X�Y�hRpek^YG�>���j5��a{�~�v�Ģ3L��A��夥C�R�qm�w&�E��"~�u��2.`Ȓ��7��@!"�ے����[cOt*6���9��?�
��#m�Wf�5������
��_�V���3�#1OV�X�q(B?�.�D�-�P�d�|UXMnd1�U~~}uyY(>_r�#��@O/�?���tL�ۍʷ�3���c&��숦����?�!0l��=>b]AP�.׌��﮲��Crs¨#�'�
���泊����"�����ɇ�}ӧ�I�6��3"���L)��uӶ��+S���s^S��50�����iS�i@��y�
۲��ɯ���K���#��DA|�|�"B3�Ӌ&L�xD�ۍQ��GFT��zC�+o}ϲGRy<|ߎlY����]kO�fp���}ZB}�B}�}fY�ž�˪�LW]�t.�|��fV���[���䅹�yMK,���S!:��������Z���i> x�욠k�e	��Mv.�z��w*��A��R��:}䐽KUٸP�ݠcs ����;%P�XO!�Ӻ�T!�I!�Ժ8PM.W\a�[���Y���	��������������pH��G�Ր$�пm�p�	���iޑ�k���a�:��	���F���������d��i$�!�V:z�L��m |K3%��\uI�d�>�L�xw��gOݪ����]<A=�����ᒐ�tqk<Bz��4�� ۻ\���h�	��n�{X�|X��Ϳ��[J?kS��8�W��Z��x��ٳ�s 
4H��Xl���o%{`Y���5�5TW� �%^�:�u�;�"�TC�ḍ�0g��"��F������t"��#�:͇?~����|d�tU �BWNK��f ��)�%�<��5��v��>Eӡ{����C��0�͖)ʁ���nB��y���ڮ�+l�ק�?7�W˭W���R�珛�R7��WK��jrڮO��m��rr���.�'��j��.�2��fQW�9��&�k]�EWo��G����@,ml<T {�L�/�{*��s&��R���w�w��L�	_�|�|_B�2yi��>��fE{UIUVU/��<�s���s%蜸j1��/#0L�|�A*�����]�Å���0�I��Z�Og�k�'�`�d���)mSMS��\[�3<�p֖7�-��b��6����4�b�jL�!5��0�y~x�do���^O=�4d���G�~/Q�/���	�A�T��L����a�(��A�y�ڒ;���q�}��9��-��ԏ�˨&s���nA�UT�k�H��1ٗ��v��I��=ƑH`N��;�����+U��N�G��	Q�������ҪQ_��Ҋ�:/��<�e�%Q���$��/��֗���#�ꦭ��P�:A���R:��=���F�Q�`U�!d�5,���}��(($@ �} ����r�A�������ß���[d�<a�{�y�"�����l���Hp�31��'�g$����سτ=~��/�����k����fMq��kȽ�w"�����+�!������a�g��/`\Ro�E&S�Jq��O8b6��[�"oe��;�M�4�;��(��2�؉�����6"�K���`������I�tp0Nt�ӤC�}(�Y�s)<#��vz�b��4F#�_�L
���A�P�Uj�Ȭ|�L>Ʌ��^�ڢ!�ĩ" ����aǀz$)�~
�bI-��ӊ�k˩bVl]P�콟�9R� :�������I&s˸j��h} ��/��ax�պ:@]0�u��cv�����/�?ٿK�w,���U�z˾4-�z�>�q�����RE=���4�"&jE�y����2�W�P��v��H���m�ķ���Bהݲx�T�a@�8"�h�����` ��n>��I�P0ܘ����{�������u����z/YO��n����6'�*���Iч���˽���r�s+eWwsW�@=�����Mr�)���p��F���,:�Aƿ*`Jb���eф�@'��M]�5fߠ�����!YjBltjyBgmsk��zc�|���s���'2��(ҢW�}䁆^7�_�(�~D�� g��`��j�JA����c�1��7�:��û�Kj���R��=��3=��W�5X`9�#�K12�k���RM�uB�I�[�#'88r�sߘ�$1%)�l��X��K�gs�+�}�|�5��rL����D畢��_�����<��t4eaE;�U%����pR�o���SnLP6Q�{���q��9��_����N��`>�4#1sǦ�c��M��XTqhA��tL[b���
������y`B&� ��~����zC��~#�I@^���i�����"2���c.[ߺ�"�=SWK�2,�l�w�n;réSX�{��	I�����/)6 �?Ӹ�<UQ?�R��p��WX�yd��a7���$\qT��l�K�"��+V����R� e:�A-�q�}G��@(����������ϼL�	^GC�{�V�(�
i�$U�4݈������"�п~��r�y�Y�e87���q/
���*k4;D�T6(Ϣ����4}�n^�6*�+R�<�d؛����~<���;�a����p²�Ʉ�1���Y������$0�I�AOg�tw̮�V�븺��j�~�M_�����I���myZO+hRN�yJ�TϽN��k���i���"�dЎ��o���f���'�:���b�ߕ!�)}���������=������/|��%�^4�����r>'w���'/Ml�1��3�v��XYC�-\G�(�1�	�� �r�*E|�v�6ƺl@��I���g7��\6?[Ꝛ���G��DO.���e��;W�t,�'D���Z{�^d��������K�(G���u@�y���a��F�1�s�¬5�\�@$�(bP"D������c0�{A#[�O���{��_ ld{��ZbAp��ֿO��2V�?Y�9�YP��^iL'[���d�� nW�
� 㤲�3.4���*'0w�o�:��qV��%���s� + $Apl[^|]�P7]d����m�������F!2����C ���k��|>���v�E
|���E%���b�p���K�p�j�h%R�� �dHW"�c�Դc$��C�њ��`@�д�w���I��X5���"ht(�=�Nz��Zf��	�3ُ���`�BǄibPfv��e:����4��/�ly�<�������I��vV��ܵe��a�t/�I7/�˶>���g��.x�2��y�0���1$%<�e��X��[-���(#�Y�?yDg5��L)C�@�F���c������yTP��F�Z�x�=� ��6��g8_4��ؗ�=#��vo��g�[T��2,���pl�ae1g���
p��w;%�{~E��ᗤcJ �TO��MhGhH���b�b�{�d[i4[Y<�j�3� p��|��)G%�i�G��g�q�i�@�Z�Th��?�J���g�oВ@n̨ޯR6P�R���{�
�N�f��� ��fW_{x=����Z}��*�O{G��o�����J���ؘnq�g�݌�~s�ݸw�F��O��B�
�
N�<�r������,���������H)Z�RJ��,P�=��;��R
��n%�)^����]�����CrV���g�g��l�]>��*��+���y��}ST��u�S0��vw���v��P���V�B�V}@���{�s�p�HZ�	>����j����}�릨-�����A��y1F��]_W]U]U��l��"p᥀Py:@���?f������9Z���&q�↍sR��`�-�#�����5�}�V�2��J��&n�F_�!H��;�iD�9�I�{�v�W�W��\����)E����!?n��z[7����
T�K��?��X�j&#R��{NR�ݵB�f��WD��Tlv:z���e]��O�wC�$��#��҆���>|�y���r��U��:$"�DF�H3��'��Q�w�}P:����{�!�Qu�*2,`p&�J�c��P﨩i�?�WȩhwDu�zp��v�da�p!�V�0]H�Ts7�;�^���1
��n%e�g���mzg�X��'�@��ȇ�X���?1�~���}ƪ� C�˄�}T��`�6!���U�y�r��a���'��������+|��B7�0������rdd�6���d���Q��FX�,'�P��蕒?��6���R��2��z���[��;��2�O\]�����鸕��*ߓ�َ��L�L����c���q��_�������j������&�����`i��4Xx��Vm�+�^
��Ͽ�c`�c�*�0���?d'�~�.wY-%E�!x@��OLǜV����v�(��M	!AH�:�G<�eϧ����I��'���RrOi_�ij_��x��B@G���X�^��;���|�~s|��l�&N>�ǥɰ�_С�H"�ý~W�w[��\�����-K�R����<=���Hk�&Ϳ��WƋ��+�u�߯2kbx�w������s'�1*`qn�D���ֻ��HX�zsd�3xJj���hs�0�m �?�$�Z)P���ک%)Z(�,�?�B	`~�R*U�("�	�${g9Q"�A�j�.n��&_bZ��\b�%1RO����ɷ�C)]��P7�<U���ҲR8$��Pt�[����n��A��|Q�=���Vܙ�yވ
��{͸����ԇ7��߃�e�#�z�a�;�p1B?O�Q�%��`��,H\A&`.th!�Ҍ�Q�0!@C�5� +��$�����B<�[�"� \/,�Rc�ԗ@\���?ZYB�
+m!�þ��i�OK߉�8�'��󱥴PD�B��|I��4���r��5��8Ж_�nPP�C "�rd�d;4bˈ*�P�WE�~�]Kl��"~r{�da/��wIS� b"�K��=a��`�e(c����X�V���Z�[z7���!�6���E�&y�����}׶�ީ=������k��`R�����8��:;�d����y���,M>�&J��4�(g�3��{��ߚ��v�W��J=<+�B3��Q�NخUC	�"��k��"m�_9�ʻ�z?�5|��ߜ�8�ǋ�hM������}�r򘭬E�z��R���YԾr��^8�J��XϢ�YգX���,�@9��T��+�q�-�����x=".����=�U\+ϑ%t~�<���;�Z�2m�eS��1oT⟛�������@93	޻�i�h�.%po�,��n���8�ԬXX�/v:5>ڹ�y���Z۷Wv̩�m�:�oh��73\����t1�;��N��M�m�hm�
��)���D��&��&lֿ+ ���/�@|������Y�4S(��'�-^8 �;�l�7A�]���=V�d���;���g)@��'p�"�n�)箐�o�/����I��M [�&�A/z)�m��S�(>��~قA�����|��	�t�uF���Q���~d�У�˶s�����p���!�&���%�2���ӵ�4k�6jDz���Ypc�_j��[��^[��_�Z���q�<�:�L�/ ��=��v"�����u{�wCZ;W`����[�+v�ʅ�k]k���:t^%�j��F�՗b%w��=j�	�ݑ5璻�Q>E7�+���3I����Y-Q��3�t��y������K�� �8G̝�|ѧO���׏�*�l:TS�!;U�:�КF�W����f~ 9_齙�&t>>�D�P`.SI�l���?�l�Xp�49H���bkU��z�O�������lU{����j��T�^�}�p�H�}�tZ�Ú��0����~���$�q�"S���h3w�4梞�؜��Q⧅�����_r֓�ֶ����NᲡZ6�
1���@�IjKш�@6 A���bR8���V���N���ۚ��b�z����g��]!���Oa����o���<�?ǖ7�gf����\V�y�ycl
�_��G@
1x9B�;=�7����hJ����nh�"�.�TƐ�!��^VR����o��K�z�K��OOO����x����<þw�_�z�\�Ѩ��`s�YkS���N���q&gih�� �>gȦ��2$�CXahg4��
1s�V�q"�2��J��LB��a+��(�9$���}
�x��O��k����X�)
8-�>.�2E:�����D�oP�i��sy�|7�P�^V$�)e��?
�?�+s��O���w̜��8�eN8g*-ƜD�����e�W�I0��V,����$&f��KK=wA;��3w�14R������yx
�}ĥp)b�;��(�<q	$����JE��E/u�IB?9+fs-�	�f�Pp�C�ѫ�?�k:��z-� ��3�F��٧|��H�4x*�9����q24"���%��,�\>i�;O*1Y;����HBL�����ܯ�Is�`��H���s �1Ѥ�e�(�}a5��ޒ�-P�i�9�){tB5z�vd+���]���~��������Xrl?�^�h�҇!_ ��ը��O�t �����E���kěE^.Tʞc)��.��gb���B�Tԝ��܋�\}�m���@zϢW(�����؆�l('�������}�ZQ��u�>M`�#}6b�I�W'��W�j������"
��#�@gd��~�{��íG��� ��OCb�(�'����trZ�/3�b��O�X�M�~ay�2O��`{,��5CZ1�^EA�MSY.�>�G@h�C��t��)��/��`���zJ	ě�i�IP�W�tE��<�ig��;�/�/zIA�R{2�k	�bDV6�K/sJ3$���Є�9��^w2Vw�M��}�d۵����4�qr��!(�4D]%�������zh����wO/��:��`�+Ԥ���z�-��~��p�!o ˏ�Qlh0X<�J����FtzNW�t $�|��c�F����]��[���95����ˡ�ō]s��SǨ���ȴ�"�fS��?��fn���	�f\�cbǱ�� ZegԶ�I ��*�~Nőw0v>fi�=E��z�,�ē��F������x�q)������0e��
ƊJ�����y��-�=vǿ�%��֛.��>�ۖ�N���5t|#<l��,��g_Ϯ��_ҡ��&0ȿH�{U1�
�����
1�U���5m?ܔ齉�����,R�n5�v�:�6j���S�s�����ȧA�_ܳ�cx���"U^Zל&-���fw���c�G��k�Q�έ��_��NU�$k��.6�G�o�H���B%&Y��<4���Q�$�]��y\nٴꟑ��UX9����a,�%$\甕	�:�5�N�j���i�B\��'�<�e�v��^��`1'�/
�^���/�3�f���3�0fo���q|xΧb�[���^Q[K����B�%�w{�]������܇�3
�������ݫN�:җ���a�%X\�%?�q���}�6h��-	n�x5FKh�h_������K�d�h�[���>,,IO��se;cN��~���A˿�u���sx>:��m�1���32T�Vڜ�(�$w���.��-7{�m���|[��g,�ع�����k�cvlf�seftP�G�Ջ��۳�ě(���	�ʺF�Q��8�? D[^��Lq��nw?L�T�_���+��2h?�p��}�\�ܔ���X|�&��s���D<.8Ҩ��m.	��p�ј����uji۽!r��v��lki#p�$B�Q�%ti�A?7�uu���(ml*�*+Y*�O�M�E�|
���-�c��o�;�!b!�m��i\#bډq��S��^�F2�$�;��sNф�C���YO"�l�U�f8�xk?
����t�?>��8CO�����^*���d��������������L^D�[M-p���������K�����qг�3�%G��{����F���<��z����n���f�,{�R��cF����Rv%���7��'5����1�2��'y˃
s�<��J-�Q	:I�>Щu�A�L+햏�d��EӀ.ubIkF9�)�M��jȋ a5H,m�	lf��*J�r���J��*�ߚ���w�5��_ǋJ1kb� �B�9�m��X�0Tpk�f�-�3�!h�?�)�!�z����C<��Q4f3Nۗ���ݮz֫K��X]��Q�q�5�>��<�8����P�"��',�Ɂ�:������u^!�9�nJ�*j�:��5s�w�,g�`l�%�u�����*깕�eP*5Eko�tR�CR�p=�s���rhh�I��V}���̸V^�df✼@Գ�&K�9P#����p~r-�W�I���[v�8�h3�*��Ɓ��v�߁�w�fd;��9����]c�#:�7�̒O-�.�E՜M�`	@��[kUN`V�V�
��F�e��#=��q��Rd�`e�Q�#�IU�2�F�������N�G@�F\]p�q%�h�y�!���zΎwA
b�
��͛��e!ك�B�V���
X�;g�_�9�{f"`��4�P��,xg�	t � '���+���8&�u1��*60��Fi`Ǭ���H�y�h|A�f�����4��*b�C�j��ω`��Qn50hir�����y&d�0����H�sL�1V��}�1�Tį(�hw,��Q)E��L�\�I�����1k�s�Z�5�Ern��0���w��r���qs�/1_�Y9hT�&l"��B��#�,�'�:�Xu�oQ�9�\'�ӝ�e7���z��}�z���%cc�O;	��c���^����D��`�tX�����k�٦��ѩ��{v����fzz*_� 
	����ޅQ�V��#�3~��9���-���I
[�tff!�A�Z�Y���:&��Jh�Gb&4�x�!
��X��q.�+1�����ޮ�*n%�N���3�H[����M���v�>�osb=�Jw�L���[�ׁtĸP`���]:F�I
O�3�y�DG��XeQ�#�%
� K~E�H�V+��V�ս�^X�حF�9S_���^��Uwvk=?wX1r2��(r�����Zy�Y�9dq����1Xr�
¼T����ɤ!�|$�����; �FSJ����<l�}�\��W�� *�!���b0��k+�[�*�N�VmZX�6���g�.=yy
�?�V���M��uX���A�AMm��K�Kr11�S���CX��N=ue���\�|�U ���{�����iỉ5��mƷsL��z��z��bf�z��:N�К$(��z��}珽�G@�%��~V#W������8�1$��]���U����U���w�Aߙ5�X�#�
$v���څ��J>�^�P!"�ܼ�&Ϻ�|�/�Q��`w������{�֢�����(�����Q�A$e(u������*2�� �M�Ǫq���7�>7'�O��aa�ܖ��t����4��.Q�H��r���SJZn��Q����q#�I�)�R���!c/r�4w��80�O��n�|z���G��r��d%��.�n+d��U��M*���6s!�pP0�	�Fs�@���p��aZ�(��������a-�v���Κ�>2U5���B^�?�3�k��S)�>9��"�BM�a$��Y��~�˫m��ɡdO��Е�iY�?Zp��ݷo9�{z��{`,�"O�W��Ve3 �B�#��zs���W����r}�X�:a���w��Θ</q�c_i����F��M�������T-[Sa%a�VrhP���=���r��IQ�2�P��tF���{Mh'�E��g�"�"���kW���3��k��� p�ø5Q�>cj����=�ΰ�F?��oc0�������R�]�S�ev����V��{6b`���l�_�+��<���iW���<s�)�����ET뻻t��b&>��/]��F!���LN��Zv�s#a�YE�X}���I���_3�(@G�8�����KYΙ�	0�0$p�C�t���������C(F��?���[
��ˮ�J������Q��d��|\J�$�B���.�	f�޿�s�򫃷�ô�wM	u�d���I���HW1���-��p���5;�^�`2�V%�W���PM@�[���3�j��PG��6�`:�:��;%#}�����V�O��R5���K������\���!马��N|��Cη�d����*�k���F�aD@�/]���Fy*hK>��Q�)&5��6�y4��\������s?�#���ۗ/[=.�7`O�)��"�o���}��jƾ.�k=/���| �?�+/� �l�(�ƺ�G-�[*�M��F��>v�>�;�r�Q8GN����N�]<i���l��l.Q"}KZ"Y��w�a�Z��-�i����1�d�;�6ž�ݗ��+ݎ�~/ʷ����W��}&�RH&b�#&�8�"lrPT����P�=�����-3���W�{Dp���3p�eB3\�R��Ϟ�>xz3yU\�2hX:��X�=��@?�N4e��E�N�<�5B� �g��b�G6�tf��V��Db+e�2g����S|�㳘���+�u~�[��a�b�a�)���{�exB��<��+F���2:H�U@�w�RCG������G��(4�3d�D=���F����ߥ7J��8ؐ�@į�s��#� �Ւ��PL�S5�^APwW��?hMS��c�?S��
�S�?g%uJԔ�x��fu���۾�c������ʟ�>S¿�L$��0����{M�i��as�m¡K�yP�7b�;8Y���1��b�M������	|�5�|ϝHgFp<ѕ)��& e�N%��;8S5�X��1j_��Jt��$���j�i��B����{��N���f��TP�1�����a��ͮ�G��-|����,���ρ9~��ةMB�����p������Kr��iI-`��!0t!�	¾�9�_���o/t��/>[Y���=��@���r�#�E����a��J�����w���>�#�Όۻ0X+'��^(��?�� ��':�׭'�$�SMW���
`��ߊE�ņ��A����bJȸ�6�L 5�g���������^�m��bܹ.t��C���πx���T�ߵ,�¤���A��l�6V����-�(ɴ��D�g� 8�A����AY�9�9�Y��`Ӻy��tB^O�T:'�� P\��;����*�hl�gDe�<�ͼ�5{���[&�o	�!�1ԄU ����#��"�1�!k����	�,��!��*��T�dn���d\[�c%����:���<k��疟	P%|��G�I�Q`����x?�k݃�5�zS+1�T�s�*���۵c��� ꘨��ny?WKuM�d�{dP��Z"X�fqY��?l�k�?k��<M��J�� ;�g.L�N#[z}B�����}�סּ%�;�R��f"��s�al�Q)���ב��_�4:���}��|Kɫz�W�"j Cˎ�)���V�� >�ea7c�@��Q��i�fB����.z���ɷB��B����Eu�gZ;B��õ��=�YZ�r�ݢ������ ˅x�v��s�>E�{�</�ˏ-�����Z����0�u��)'J�����&hes�i�Lw���j�k�Je�d�Yi��ۙ�+:/�� �EV�b�%<-�j#AaS�h}{��J���7"��W|'����uԳ�/�Y����K��>,u�ьz��oG�����.�Z@h@Hr/�݉�)Q�7v��rl��4��f�H�������?	�`����i��;.(��?���q��BF��\�M������0�qvI�����ol�0�wY�U�y5�)��J[��1U��������U����iG�p/�{M݄ו��/�kM�LPTŅL�[��-RC���BV�$֌�:�OI�nj����2��Q���7J�&�?���c9S��he��,C�����O�W��(��8QȑW�7f�W� ��Kf��3@���r�1#�	�Y������l�審��c:��*�z�gzV&l�BQ�8V�?4R���q�0�A��%2(��"����H�J�z#u�#�o��u�is���F�Y/���\�G����K����T*���o�S<q���I�/j��p�'m1�KÉ?7�Ŵ
�HEs)�&��Lq#d�~2]F��E��PцC)x�(f�z�M�E^��o����9�|5�������i�����7A�M�$0�V5+]ʸ|3)7;6�ьw������{.���5�Y;K��^�Jr�-�F�s�8�#q��,�HKf��i����ݩ��Ч����~�"���^���b���ͺ��:�F={�|�F'Um��'����o��I���]�0QH�IP����WN��7�����������IDzz��R����!����|�m��]������%���`j�@.V9�k	�^�ǐOo�߻��vΊ�:'B_(ߊ�{�龰_��9u[�:��2(�}�C�8��Q�8H��On����L�9�����K�m=�����9g$�@(XzO��j�2:��6v� L�h���(B(���/�	uX�=�|�Y���';�f:��p�&8,PX����.��?g��\���m��͟8a�q���w^z��r��#��#]E$���ޓ�pX���M�W�O�o{:�ԝ���l�ik5nzϮ֮Ƕص����5sˎV6�DA�-F��HZܴ�Z�Ӣ�0��˝#�r]5�5���;��l KD�T�h���Ѣ��R�R<.;P)èO���0şY���}D�s&_s�<(!�T�apY8)q��`hS���9� ^���t�w,�n7Cl�̩PPp�9.X<#;%�9�ˎ�3 ����$���^�e|�s���s�� 9�8C�m����x�ŋ�p����ۚ�9r�B�Ga׆��B܀�x����aI�z�g���N�1�kb�NuBa�sT�hELu:�5�s/b'�w�$>9}�B�+�0Zf�m�C��3�c���Q hGH��	�a��L����u����<�5�d�?��X2�x_�����yT ��GM�i��^c������"~S���~���,�-g�:N�θD���6�^5�%�|C��^W�2���(�7w��~/��q8�f�sz'��4�~��;�s��	$��*.�}z_��j�� ��?� C���Y��.c��i�2��M��ُEh墲�߾��+�l���}O\-���6�9O"8E�i�PL�T}�CgIYO�]K�\�����iHH�᫓����K�͐S4�^�j3�L�����F��1�l�J�	��/0�ٰ���g�<ˇ��ӽ��{fp��t}��Be �L�]���PFg��΀��g��i��i�}`AJÍO�Z�#;��ɼ�g�-UkK��W�\��ww��|}�DG[�^�5@��0�d,�B��/cz4�4-�z��5҇;��X�����TN�E���#ʐTR9��e�c]�����3s	�t�/��� ;�/p,f0�Ɍ���L3#��eσ�90N�wA�q���
1�0�o��Ҷ�3�7��*�B"o
�hSM�G�n�hn�N�Rr##�G��[���Lѵ7�7��D�ࢩ���^_�%)ir�K�~>�;�9�<Y�$���N��5��+�`�[y=2��� *�g�$�dG`ژ8̃5�!Z��vs������3��F�\��׏�I�[F������qύ�R�x�&��p_�A�hx|�r;���@�Μ�l�K�~�]����N����E�5�\݂�u_JI���5l����.#��&��{^�����䁲����3y_�SZ"��7^��&�u%}X%�v[T��%u����t�B����9fy&`�!:�l9�`�HJg�1ɯ���`7�Z���x˒���+6�&�1�=���9����Xo��g���j�/捬(�܈���j���h����b�(H��w�F��`�ϲY�oCj��!>��f�rV��J�o��TjT��>��&�N�V|.��m�>�c�w6���tg�'��!5 ���vs$E-�p��/��ϴ��~2\���p��� ϋ	Vy�Cx�8�#�9�'�r(ku V�xc{s����������s� �^���H?\�b��+4 $���|}&|Kw�����1���<�>
|@�ȡj��gjt0�?HާH���=A���[@�;g����~�M���!���Ž�Kmv�zUJ	Pk^���e�_o�VΡ۝�'����#�O鷍Z��#(L�Z��Z��W���{�I��d�
���M�.p�TY��. ��l}%!N����U��P#�+����11����@/�ڨ(rWa9�Q��03`�����X��Va,�AUI٤_&h���?��{�n.ȃ�XU信k�/��[mm=iP�F�ϡ�; �(�Y����Y�ۛ�����4Ljj�M�b깾� \�|���yY��3}��.��*�5K�0[�Ï������<@)H��^d�).{�2!���x���2�plHe _���|�Ǵ_w]buJ�F���8�Ƴ���f�qC���"}GlH�UAc=�$J^�g(�Y�F�ޅ����Nȉ
ċ׉b���㈽*��
�ծ:�=�4����%̒����N�ܼ���A�g5��*��4^�|�n��Ɍ����}��{5:s ��v�.&l2��{��bb<���I���=�72�O=�k�O�m�^`q�Y��@��6AU$%tC�9��w9~�ʰ� �Z̷ud��HMd���<VX:(߁��j�]��o]+�1�]y2��;�י�x�h��0���.!�
xy��F�;���s���ʮ�~����e��j������P�t���&�yG�F�<�el�4�z��O�R�[6[�|��'A���k|��9�����j�H7g�񕷯?y��8Ew鞉랊/1�a�^g����gp+*�s�����tLĬ�:0����`tT��\A��^e%�;�4�G��X���Hpʒ��c�x�c��8�Q���sR��w����:E9W�"��f��~���ΰ��u�I��$Jh�5ҳT� ^)C�(����3(5���y��� W�����JեU��Sߘ_Vf=�Q^d]���?�
�V0H��'-�u4�#By�{���J��2��d��a����O"
E��"|��6���S�����˹�r����,ڰϭ|��9��oB��@<j8�1�-	p�cM���G8��X$<���W$�����qu���ԍ0�#��%�h�k'�����r�%	P9�贏�i�,�u�5*��І0JQ{!��(ku�l{�C��c<�O^~���Ҋ �}m��Ľ3�h�bra�X��R^FA�T�u���)��Q�ߥ<�����k�8rr]̏#�m�X���o��K�'{���<D=�V��p'�$��~�8d������W&K�UX�1U��;M�� d~�>�P��:&p��L�C��P \���Z�A��}GF�0ɣ��/>�����.
`e��/=����!q�#�$^zl����6O5�iP��w��w��}㵽.n����q_���Q�������V��r�����w s�6Q��u��J����� �A[l;���S����y����ު����!��gc`R� ^�I���}�^�/R�v�h�/�7g�O��O�;����[���5n<��L�=6��w�=��R����i�՝چ�o!����3<��{:�&�J�`H��M�C����C%�9�����C�}N�0W����~�m�p�o�+eBwv�qj�e���~�n
2�~���vyj� �v����<���΄�K�Hb��VO*IUٓ��Ŀ_r��J��(������� Ɛ��w2���'���UR��˵Cjq�y2�+���<֢'h��t{���7�=�~�e�226C��ث���H���H�V0�ʛMS)�ݠ�=�i=��s�ƌ��%���~?��}�ѐ$/�r.*��Ύ�Qi���·wM��:k��7�y>b�b�h��^O[C0ڑ�Τ>֗�r����f�C+3�c;W�pO���҃�֏?�Ki��Nn߆�Y������+���3��<?��6?�ck��ȵy�>?9���	� �v�;��h̳�X����>�k?xv++�.��H-+A�[+j��xaN������Q�>�%�Q��V�����@&����"}��I�{$���߄��p/�ǿ����>��)^s��S� ����` ���s/�"$^�[5lH�-:d��h�g��Ը���2����W[�Ⲩҥx�H�a"Up1�s��G��&�`;?�����h�;HCz�2�G#���no�	���	i���Y�X �ga?_�.���� {!'4��J; ��"�j"���Vc,�mKǚhI�#g=�h�1��[�ׄ�6!���cX������x�/�i{'��8�T�~�HQǲ��u���a��ir���o��뚸$��Lu隴��ۜn �����}��nn.����+��)��g'5^}�%֤x	�������1D>����8j:�Ɓ��F��o������>/8/8�x�͛B���l��9�?��q�i���/���@���M����כW��� t��b��:�"�[>��u��NI?։�4gh�����S_`�s�U�

;��}�uSW4��'x�㗟����tP}>'A�Ky擜84��&�2]6弧jF�pGe"�$$9��D��|ԭ(�Vv�����0r��*����ն���ۈЙƔ#����TvWG��"��2M/�t�)���^�||���i��3Q��1
O���._�0��OK2��o��|��3
�-���#_����D2��I���=F��W)��0�LDr��s<mt7*�����װG�S�O���Pr��5�u9J�'?��r�byK���)Dj���]����c�2r��Ul�r	ad}b��"T��r�Q
{���o6| �jY�4��w'Rf��wߴ�_7�x��]����w6gmg�5~�;wU�H�0��.�ӗWd��e��o�/R+(�D�����>n%�������Dħ��;�o�&�!��,r���/�����e+Ř��"���lp7L�]�=�,���$�%�(��)Q��7�S�U`(��H�	��,�!�322��'~��L��Q�1��~��[ib��W��r�S�E�Y��$ɩ=r�����uWA���P7���I�'�78=�w��m��&����8����P��q�]u/���+r�%��"�4�����w"dű�t;�t���������O�����i��I4���}{dt����2|_�Bc�&��F����)$����Ȃ�<���'��:u�s�N ��Æ��d�`�@C�`�T4��T����q�]��d�������������o��b��������^&�����6�~v-M���l���f��42�
g����]�y��p=��6��⁋�*s+�~u��.�mi+n��eX~����_1���u��B�t78ۥ6�>;p�B�ZS��J���;�]}�B��������{ݼ�� ������ݴ/�ȁ��G�'Ko����lQy_����Ze��ͩ���]>�L3���	ސde0ղ:ɼ`R0�A.�����T������X�
/A��R��Yj���J��eGcjq'���x��Th�����iL�9T�Q��D ��%������m�)#H�7��_*	�]����	���3l�ԡ�R�t@*P�B��Π��.3G�d�C�+7���$~���%�����D3�����������>�83����
��bK��2�S��g�LD��qz۳��3�3x�he3��n��i��	م�G�2E�a�����^�nnU�\�^OC��8AH�H=��U�p��3�R�P���p�5����;�Z�<��tb�;{Hc��D���WN�U\��
1��7�y����\(��|�m�3���9@��ӎpaU07��v�y��ԥ���OXi^�8ɕ�ɫ�e~���g����:~_$�Ķ���d�O�f]iSփ�!`�?�?�!�R$ДƦ��*��s`�=h��!XH����e��`����{9���K�Y��sK�{����yo'y��o�r�����͙�Ť�C����J*�*Q4�rS���2g��i��S�"��e�o��K��Z��-J��W]%�r6�Sim=~��ha0�ٖ�!�T�e7m�;����9)�fj�h�Th��������g)�lT�-����c�ќX����!�uu{�����7����Fb?Z�6D��&�\Y�*o��eY�76M|�V��M`��w뒯�L���O�$s�׺-C��VL�B&;���K�[¡`�N�K��L�5�c����dm�0M��->��ui�]v��P��0®�i&���\x^��F�`�fe���&.��[��H��uݷZ�[���W3�����WY}�&����3���(b����x2qC_q� ���\�"4�9Ѫ�Έ�y�G���r��pjz_�T)������9�+�<ue7�u�$�ʊ	}_�	�CK���&8��G���Abd�PXE@؈�&B&M�Վ�D��GݏDǧ*2�k��3�X��ύ�l�x�u8���c�X0��X�*�K˧	�����Xnt�A �U$t���-�����Ox���v�߮��?�n�}Vz��G�qL������������0����"�`(s�>7�)�u�x�4zg_�q�v,���l�S��5�d�m���s���`���b:F	��n��;����}&#���-F(�)$d���zb�
�뜌'��G�]�����꣡A�(uU��������"P����v�u�h������Mue���=k�2��^Fz�^f6@W/Ƕ�mx��̟�[�������#B��{\�jPIl��*��b)��%�ѶB���^��^i=��[(�+�K��2ѵ~P'�~	�I�!o�o�9τZ���w@��e�սf*Y��O����|�!��Q�Ou0#�8��_�=N�K��B�3P�ˌS��Δ���]&��(�T�c�wZh��]LHI��M�����NV�}���nR6���ty6yR?sEշ��˿��ͬf�-�A�n 0�[��G\/1�MM�6��H���+�$��iV�����]�6f)\�����(��n0�L�	^fi�j�fgu�5�kvhH�<j�Iq�e��2�xT��C�b��R]	�D���Ѓ��^�T^��4-=S$cH���#f|��B�J�Ij�N��u�~ ���ByvB��0.�����j�K� l'i~ކ�m�jW�|��h,d��5k��)��W�e���(�,,+`���\A�-=��d4�����p��:.ʽР݌w����F^w���u���K5�92�۝���)��,��	ɦ����Og�ovM
ƣ�g�j����h�a���M`���ǋ�-��Kg6�Y�C+<~��7�ƺ�z�R�&�4��E���Q������Ě�ٚ����������w������/��������4;����>�线�|��7ˡ�P��Ro�
Hݟ[���a��	��y�x�t��F����*�����¯*�4%�R��Ĕ�����&���RH	�s�����f�CjO�r�IYح�թg<Nk!�|�����;�"��>.>f Զ�o]�oA�,�x�=�%fф_R�,��k7�a���v��Dy��6WɽBW�/S�@׍�K[eqK�'��}��d�_������Ŀ&���/}p(��{�TJ���x�<�����m�[_��lX"�G�25�8r�AjVo��Ɖ�g�\8�{S�,�v�z�J�W�Y��o�g�ڍ}�o��5&��ܪ�&�᤼�O�Y� 䥆F��Db�2(���{���D�1{J�^�2-��m�U6W3�d�=��,a@Ug��K���s�q���{Bj�_ L
K��"�}b����YA�y+�ǳ�9��������k������Q�!�HH3�ңFH��hi& �A��k0��.I�]"�ݱ{���}?;챝sv�s�|?_�u��F�����������P����\�|�c����>ZO�mɘ�nh#���~Zϔ�ˣ!��������z�o��m^y�ftqOt�tO{�t��d{%W�G�4�EZ���GKz)g7��ۻ)��Q���q��T"�4�O�zȭ���?��^E�w�@_��)d�><6cG��M���� 5��j�@X�Q㬫�)�����D˺�g!�)����E}��:�ۂ��9�B��h��[���?b,�}��
?��&�����3"�����#y��ԃt��ঁ���;��v^U��0�M�}:�sw��y�(�{n�	�L�:��8������ǝ��ؤV���G�#��[����wRl��qa]₶kɁ�J�U������^�s�������֭'E�zye�96m�͟��̞�{������7o&s��;�]�[Oj=]�M�;(�|??�9�P���c(:s���WQ#S��T�ek���4��4s��������^���)G2 �Q`DL)��oޖ;d�c.�����l�㋷S�(���J������tߙ�Br�����C	d�G�@ב���!�}�X��Sw;�Rkb�}j��|73���u�՛��6�:j	���e h{Y�[��T����E��]�y���ԕ��s��2���RdzϪ��Ç�ѱ��@7���	ƒ��ݠwi.J�Һ�e,S+��>>��>�]�	C�5�
�Ll�e~<L� p{�_ǆ�%��*�&�"��o�K?���d;P�x�\���q���>�
/Пd��u�qNT=�'�B�����(�dૂ�����	܎���,\�GuϿ=��8ے�HjFI�S���:Bg�������C�䩴��m��nІ���:�J	�R^�����ٲ�p���n�d�}��е�*Z�|b���Q�I���e�<o�~��⭨����ȣ30n���6G/���*V|ED����BYI��l��?��:)\Pk�n-=�_��zi�on!rUr�2��A��R��)��x�� ���"	�ȇ�n;#ۇG����G^��=z 1�A⅕��M �}��f�(����d�^�.(���S{!O�?�Ȍ�Ȯa�I��
��A��l?�9��� ��AfO�
婧�q�;:��f5,ʎP"""�7�Y8 ����l\��w���p=�$շ$�����h��$l+�/0������yX��Y��R�J�l�SPI�޾�n$�Jm8!��=ӼݭY�V�����U����:`)��۲�Xmc"�<-Đ�`'N��;n��K���*��O֯�Bi������/mA�۩rZ��ʘť�է����lUy�.����D�Iu
�፣M)��L액e�|.�hv���o�R��_/�h�R�m��k��f�F�8k��RD�1DD'���A3�Z缠�A��$"�{�Q����EY3���'&��Tf$�+ȪwC=�?���V T�l�����\�(���1�d��N���:t�[OOA^��."J�,o�w,�(��$��M���R�����a1�,�)��^77���6��e��
M  �f"�sH0Ȗ��o��by�1Z�N�bp�=x�ȼ�3�_[X�BBOU���8���e-m��5~��_�$D��B�α��A.G�~G�cT|=��tu��ӻ�ojp�ǧ	��y�!�{�ZY�C���gmk9������z/܆�4X.Tm5�Rn;�6:���k�ә�"7g��~�k�3c���GC�ڶ����O�"w�����B6 �s�`.����H��4�m��Յ2/��2s��O���oA�+��2_M ��}�8z��>���]_��~�"����M��z��S�@�g�Y
��i��<>}���h�W��^��@-G4�79񺖟n�B�����n�C��0#9*U�~Wg�����zF`�x"An/�߃�ZOZ���l��b
�1��Q®N2�.2a״�[�1����Oj� x;������96��_<8r�\�>Z������(�x��˟-fڋN��+uM��k�]��%�d(��g1j�C��?��ߖ�:8Z��wv�~-�Ci����
-����?M�:is܅�t��Q�~���ݣ�>S�Ղ�Ʉ'���Bm�-ͽ?b���vn�3h%�R��_K���%0�'=�6�Il����<��.螘�����c�^���uP[IcN���O�A��m������! Jd�-2%{H���.;IX)߲�̷�W�k��)Gq(}���s9x�s���홏B%V���'�$l�vP�Ow����amNݛ50�h�k��Ȍ���j���ל�,���Z'$aktS��E>DTM�UϦJT?/�Л� |I W@e��Ӽ,��d����b*�a���
%rӻ<! ���@��SI x`l{���Z����f����"����ᑠk���(	�"�G��Y�~
*�ɣ���h����8���D��+��!-2!r�`ܳ���T<�j�9�q�B�����v�]u�[ds���-�̷�*�B�2bm�z;�)x���������C���N�L�#��9�)�W"��,зy����pZ�́�8���K�պ7��2Ħw�G�D���p��c���f,&TBd/��!)����9n�pQ�G,&}<�"��bJ
�#�m�B5d������Yi���%�3��ӓ&��LSٯ�᭰�{�r��I�S�� �R!�������Jz������A˦��v�N+K��L'�]�{�����fc�V뺔;�٥3��DV+_y��Vq�)�ь2��"������;��!��'O�U2`;_jn��H�|��s�zctߤ_4�4����OyH� �q�|����?��t🬮Qq{�E�0+��O�35:R�;�=�챨6
^m�iz1t���/�\�SA�F�q��HԢ��������o@=�����s[sÅ·�����s)�c^��n���'���K�?%)�Ã�Aûn���堰��%�k�Y?�>UȘ��~* �UQ�AMUР��7�	=� Db/�T�յK�G8�W�-O�EViO�O�݌����;�%|����[̕[��7�P	^ةꚩ�!���������/����Զ'���Zlٷ��ߏڞV��>�;��M7�����F����S~����>���k�E4F�^�m������r�O�^$5|��1�L-n��s3MKaB��-+�w�u>���vF�b���j"��9���`�� j�R�hG�H��"�
�[e���:��/�F����&O�ی��lu4��Nv��Ed����"nţ~����Zԅ`<biee���NWt�Q2�u��$D�����kz]�&Q2�������re �x��f.Q/�{��g����_�6qv�q��x���M�s���Y���)i��(��UXJFŔ\�D����n�aw�W�ަ�v��7uջ�3�Y�m�8�<h=�N��?��[ஞ*3R�N>a�&� f�و��͈O�c�_�B���.��ֆ��Q#k_ENN���4d9UZ2\�f*S��1��w?|M(~�O<�W�5�y��{�8yN�hp}�n�+�Ѯ�%��\����X��x]իKb|[/|3oW_�����R��A�N75UTT|}}�Lψ�54l00̨�=�T9�VIy�Br�9@WH{��4W�YNq��P$-�@
ӳ��,���h��M �j?b����c�s�ʇ��ӣh#�b�'�\�l�J܁$D��z�A",2 d�4�X�9oP�f�0��W�@C�J�+Dp*�L̝Ҥ>(i�
��eo�9Cc�/(�������焗�O�����y�$����,M�+�2��3�\k�]s���x�s��$��d��-��"�+�L�( n�(�#�p��ta+R7QP�y��i{�J%����2�bfC%3J�U�3t����,Dj����4�� ��w�@s��@jN�4��'��>�xjJ�%Q U�rn���9�e%��7�- ��n��P���+��_�H]�����G�i�K��,p���J�Ї5h�������-�*��<R0�ѽT׾R�$U���Vu��dC[]
xO�?���,�5�w�M!K��q1�4�'x4J�������mf�FZl]�4D���4�;� ^�E<x���V�&hGǬ���<����肩��[��rdO	���%�>j�y�y��57�L���G�if����(��jR���r�x�۟-O�l���h�(���Cɞ<<�������'0���)�B��L�{E����kZH�J{��2�a�^�eY H��RE>�?��y*��?	�``}j�c7���y��y.db�xJ��ϩ��Bϰ���������)l�|�vj6 �|�9�Z�>��Z���^Lc�~����l��kY-�Q�2�
i�� ������UXp?P萞T������"6��#[C���Z��Y�x�Y�^Ro�GH,���{n�8m�g��\�@�
�D��}7��U�|C�ZC�DC�M��E,�]&S�B2[���e��!	���T��C������;���[ ^�Ę���y����}�v��3X���߰�>ܐ&�y�M�u�|�wvl�ف���l a;�\ �~<_e��.I��9x��A��.Y���5����{��T���Q!i���7�kg�G�"�Ǖ��"��]��x9H�W_/�F�L����� L�r��n��OqYL@AA� ���L���H6�n�F���8�I�$�X�w����f���A�:љ-�w�~j
����_�%Rc���F�\n��Z�|P�k{�;����r�a�}�v���X�*`��a�]n`;�0��o2�Loo�0wK������5C�;:�z����L����.凉��=��=h��]��;u�Tq4W3K����iR#V;�O84Q��V\)($�'�܃;:��;�_��)`��95B����ʶ��G;+���1���`?�Y�FHBv��s]�t�I�"���_�c!}�7h���̸�ڼ�*�[tKӼ�u�3n�`��/rn�i3n��1'���_�u����_���$�X�������VWW%�)1�@>��z����~�G�C��xD(�w�,;*��S���|I�.z Q�w�����Il*JB�@ea� [���F��Q�zSY����W$j��"n��ᡃ� o������9�m��6Qv��A�epH��_��I��۬��d���q�kyG�_ﷸ��ܧrur����kLsW�/��8��hO���T����!Hu(�9W�!΋��/��͠����FwҠ�.��SD�EB�<s�0�qA��~��3�����%�H�?}��@y?8�-�%5��>mG��!���]}4??�����;i277��t�X�X�4� K�<��0����k���B/���,����JBkx>�H�!y�k  �)괤�l������+��j����	
�6ơ��U'/��v��Nhɂ�gq�����C ���:��h������#ςs�\�����pfi�������ie3��}׳��\�J�y���6��֮uS_x*���Ofb��Ѣ�/��T|���F*�`;�w��B_;�!��l˴s���	G
��uq<P��1V�R�ڒ��ʛx����j{�П����;���i��eٷ�)�x�x��|�o+�:���\���(�cq�A��L�u�ĵ[~^����'��k���(�\��C��C��;R1�ӧ��&ȑ(rg�&��G�R<�`��_���A/Q� �� 6e���b�s��3Q��d�l�Fk�������m��*��K�!�e��
�=aw��-s��ڇ���v��Zs+J)_7�F�^��\ӕ���������������,��h�jX,�vk�y�a�ݟ�DИ�L���O��c=<�\Bz� �?tpdgt�E�ن'�#��\K��[)}�M�]�Ѽ�������]�?X�G�����U���4M�yV�\�A�vr�@]U�!�OP	3�SZ�'B31-���y[cݯ��ɔa>֡�&��:��^;��<ͭZ���(q��ə6�f˷�}-G�pg�
uX��)�@��K��R= �,��P�f�"�n���Q�Gr{D���0O$�,PL3[�Œ�J�km[$ྖ��e7�C���jU�L!^LZ񃯢GH���i�yXn��ξ�2�9��� ��[�ߦ��[�j���(���o�srl`�wh�$��u����>�����69?��P�����XfBg���{��x5��t�fz�<pY�l˼;=h��k�YW��`.�n���/Z1sKJ��w�
�&��2�M[+���~g)@���f��zj������ٹ(][`����Q\f��&�̍��LI�,[ׂ�w���kڼ�7F�,+m�*�<~��v�F1��'z+Ƭꬲ����,E<qMps����|k+��v
`?�� �-qk�?���i1�И�0y�`�4��>3c��щi۹113!�3�؋�E�[��o
�E����^��]x��|��Gr������甆�
���?�u�����$�;��2t��پR[BuuJ��`�ת�4��.۔C�,��y~/��ء��6X�f�8`R�ϲ��'��� �6'��~OX��%�N}�_LC$�n����=���ʱ�!�+%,[.�� �[�H=	o��Y���@��?��~�~o�Ψ8:�LNm�Z��YIi�����dQݾ�޾c���G�X�`l�zܴ6�2حQ\�L��Db��{�gN2�`FG�FȔ/��>�H~� &w~�QD`�`�ۃ�7����t#�(^��?#ϴ��F8�E:�Z{R�v�x`A&U�N�b�u���G�;��/�*�v[��@�H���!��!�(�A�� ���bB������ty��2_[SV1aL�W�#��P ���<��k��w<0�ǿT�?	�-���8ڒ�zku,��Bm�j6ö�I���gY48����>�]�������H�B&����m<!0N�S�:��炞��9r��Z�*�(��b;M']P�0���<�I7�����d^�����N[�0��-|I1eɶ�g�����ąoK� *���/ �t{���jE>j��*6+�~�7%b���[�®�+���ؓ޲��a�ռ"-�(�0d|V��"�{��`��C6�u�l旍�a�&�2= +����lkf������pɌ+��$=�@�?e�9��R�}8�&�R�����E�3|��7R*yK&[[��$/���!�����/���-LR&2,���2�Kqmd���H͗�-`��m?�}�;rB.J�}��<U�9��SP�nj^ `���{N�$@5�_��V�
·���/�ޥ>���E]���@����A�|��d�.�������\�x�5�"k��J�B��$�MO*�7.����$�Z;� �λւ{��*���@`QǮ��q���W�|�B}�a�d��Q��o:������3�Q�-��U�]�O�5]E�����>,���nTv_�
��x�G=�0��8i�W��?$ee�E��s��U�q�1��.�:�~-t�n�o�?8ۚE������l��d�	���r-��k���h))�X��g�dt݉\_K2�E 62oV21h.^�y�rp"�7��	51�K����B�12�Y���i�p�m�u�EX���i`�Cמ�����9�]��h=Z9���y�G/s�u�Fn�y�[�ͳ��B��⾱l�{gY������I���bvV=ZM���;�X��S�T�>,KEe���Z@�:����wk��/�I��d�Z�Q�7�la/��=t��L)Y'X���k4?�-;9��2�u�x~�1y˵šTa�Bv!-]���ۑ
���������΃���p�dw[[�ꮃC���Q�㼃�<㮟�3\5�0���:�i v:`O1��b��)��מ�Fɤ�s�s��9�>=�:�l���ڏ��ڵ�X�r�����YH��������<F�"��o,N�Z�|�Mv�}���P����Wi��`�+E�����>����L=q!�=fJ�l8���P�w�/f�I���Zv�d��뿁!U1lb��?9 �(�X��H��sQ�*�D v��)�
�Џw���f%�m���=�_��5�y���E��z�e�/��^�-v���>�`]���6�a37���{*�=��me�����m$H���j�.x˥�ũ�'T��oD��ɧ�$d�I�_5�L���b�OSkͱ����o���R�=T���������e��A�D�x���X�߱<&Cs���#�����t���1h�\uD���.�����/GQ���fʋ�h���S|dQ�H�j]��_}oP�HWz�����SE�D�&��ٷ;��Υ�LNo=��F�+"U<Qϸ)����BU� �mq#N��?<��Cjyl2�Edk�p���b�(h�*/��`��x��#!G��oﰯY'�]5���<rS	9�@
_�f���}\�-���q�:��9����BY�"����و��Ȏ/�l��Sߴ��x�]��6C�P�����,�@���/t9�"��4�Y8��s��IYP?7��8ّ���A���/��d<H�m��*���\t�۷dZ �_ߛ�|��6o�7���a��߀�������fQ��S�&��G�n.���c�q�mWf���_����Kt����7��?RkX�k�c�>��p��3rz� C����6LA��or_L	��^>r	Õ=�f߽��G_!�C�.��y�&w�;m�w_9赊a/���}�	YX��a���|�D^%)K���<{�)Um�k���w#�'��p�����R.�x��%(�F7�p$��B��y<����T����×��5W�lƔ=&�j`r{@2��e{�F�O@��������0�Ī�M���V��[V�TZ��!��k��W�/m��п���߆�k��u8��J���׻��W�n��Y��T��4:�$arNB����Bg�üίm��'k&�w�KI��ү:.�n�2��}���(1�Q�w���Aހ�)��d	��9s��o�l$I�gbn�`���~'Q���Z'�$%�k��qgS%)Z�����}7�K���x,O^���P�(�P/��#�Cl����a?����A�P�d�Z��f�;"�'i\�?��y�Xe��s�7-���z������v�䬰Ԝptai=�c�����]����7%����_�w���
�p�d��?EEE ���Ƶ�µ��sU�gϟG����^�r�X#"���?�*���|����oBC���F�֤WbZ�9%��;�p~�s> �� �U����aME4��P��C?��˖�E3�����X\�DeC\x��ʲ�?]G�4&�7����?�'��A+��OWy��?0�ʨjO�6�����S%�H~��Z�xr�0U/bxoV�jaЇ�w	 i�"M�?0�7`�֐�yߗ<�i�";v��o�,���=���8B�e'��@<��̨�1}҇��i�	�.����#$7�,�+gg��1�"�MpZ�HT��w
��&��tN�G8�&���Ux�������e�XU�eA���>c�N�0�2�L�~5�%�mWȤ=�/��{1�}ѕ~e�Ld����^'�6�2!~�ςa��Fy���1V�����F��ɮ|�
6��4
;<K�$�:a`�P*�N��� �e�ZF�,�S1���~ɫ���NZU�	7�(�2������1+g˖�Ԗ1�:��جVB����5͎B��E9A'۠�(T,D�sP�>B�8�p��Q�zjմ�O��9�s^E�S�г	5VUP.�'��A��ɌԈ��8e�SBY+�s�)�zEʋB鰅Թ�B~'�e;�%v?�`��c����c���d;!����C�u�ă�������3�>�Pş���=ou'�ϗ����d[ES0���R�0w���#�	7�L�B?!��m�彚�G�X�i��B��7��;��p@YxFaBrQxFqdl!	���Z������v@>`��2D`�s�Xȇ���~��V(��7��ꢸf��G}�����mK>J߉ذ�ɻ):2H�b��2��{��k�ɝ8�E�B/�ҿg)ߦ
~<W�Y`�n� �?������76��� ���u�[*�~N��'���L�-#)�~Œ�t(8}!�7�nÖ����V����q�@\���E�ٗ�&w�N�6[^ �������g�eԩ��"&�d�M'����,<96n(˜ZϜX}ɹ?���92�4�V��eݕO�'�-Ͽ���i�e���4�M;qǸ�>�3U;]��w�n������.��p��?U������~�.��X~�I���wb�zf�zvP�(8q�W/u�g��z��v���f�S��h��vf8�6v3c�/���n��E+u�6�r��rƂs(���ʼ;,������Srs������x�ĸ�����ˏ��43U��)�U���u�eg3�	�G�����C�DN�#i1ó�L
��;+l5�U�����/��Ϋ� �;,�-��km�'���x}�ϭ�Dr0��k��8PS��F���='�.�hi�އ<�>ecw?��|x��{O�y;P�q�~}��s��Y�������'
�-����<֟"4��Q���ʗ� ΍
m��7�Ԛ@�GiD�]��Ɉm��Y��1���v�EL��:�{���D�bNkRz����b����|���N��V%,A=�
פk�\�H�B��z�/P)����u�I��FwO��|�OhU0���s��FPYw�f�(��\��WRE�D/4V*���,��rj?�V2���,���t�����K7���u���cB��I<T=��v�ߢ/g7{��Z\
v�mH���s��1��L�<H���� ���$6�N����e3e�>.��X��u+*�z�Př�Y(g>��o��M�<"�'���9����S�4��T�.7J������#֑߳�[/���h�*G~���K�"�/dVB"N&.��^:t$�8��>�1�����IH�YT�]sd��jX��1&��c�h}P�c��l�}�;*�w��44N��Δ��D��U�EGdJ'E��G'f�)�y������:E���� ����e��������e���te$/�����J��(��b�9�d;�2����?}$$0F��y'�?ә��[R9�S�+�<�
>hxA�i�Y��׫|}��'�y�H	�K�G�(��� 3`ߺW摲�"����T�4��%I�C1my�c��~V��e-r�(]�ZJ��"��ِ۲�/���o)6L�����R�/��7���7�t�<'�Y�Q7�Q�����L	/���#�_����tO'L�M�W�6�?���0f6 �\�����gw��OY���!�U?x	6��~���,��/�%x־N�W�z���*-)��[v��� p}�Yz2�1Q n�3�m0t:���2L<�zOd�Չ��{�=Q�=Ij���u=���B����h��^��:������f��{�ߓ�������ʑ��4��d��hɉxѹX���k��~ЬuvT�=k�,<�ɮ�ߪ�|�V�S��Ŵ6n�g8|u_Q ��;��lŹf.߲B�[�.�P��;-���٨mHdՈ)6�cr��e�n�NV���E>nn�U�g�Ua�\~��;�ZN<$��>=����'��/��u������[q�ٙ���F	�ӑl�O��j{�=S��蚣�2r������KM^�A������诛�n�vJ�z�<S���;��P_G��)ݖ��m�%ة���]��q�a�T�F&�s��z{�	����
:aw�0w����a�K��a���a���n���D�>����	��fz�>w����1 �������/�$�A�y�<���?k�IC*��#���R�'	��t+l�m����#�C7g	��&�y(j�>OF��R'�?�Ԡ�R�3[б�Z��g����&�~*�[I�:}������g�Q���>�孙���{��Ս=��7Jz+�R��CbB�Y|Z�O�;���s7�7���M�*b"k�f��gPm;)���,�5�Ȱ�=aQ��_��c�a�%�̫���H��cƱ%�;ʹ���}}��U�1�m��V�TU��3� 9����#��-r���VZ\u��A�K�T|爪 �ޖ���ubk��Es�8�^��N���3cu��'� �+��T��"_�/LG����"3��8r���go�1�����Ы�*5�.R�bs�S\�i��LD?�F���X��
��*�� ��c)��>�ɴ=v����J�n뵚
�P �@%-�����J <�~{
"ٓ��]�����Jfo
4W�T��N����E_�ݒ������"����[�}�R��`	������
h*�>0hk�)��k�����^,j�#4pV�)V=-�,T+,�V~V�VUz���;��xR:7�>�g�|�[��Vt��5:[����٭����kV�u��#j�h���xڝ�ʶ)��Қ�{\>[n��I���N#9��_���C"p����Xv��P��l#�3�/f�l�qm����7u�&����y�qD��F�a��?	����f�(tC���S�`���gy�:���Y�=5��%N/[�f�y�9ރ��,Nվ��aYl9 #��m�Q(�u6�Θ��'$�fl�	���!�N�Tg��`7����%���`��Y�S��x��2�d�\$� v�l
lY�g�5K=|��@H��TS��H?K������ b�6������^�W	c�͘7F��+�~SO�T��}%ׄ���Y����b]���P�t��y�2� ��22x7r[Ws-;ψ3�L����x��vL�w�pB�ڵ�4�h�O�tV��:?��˳+zQP�+�-�M�h$�ܘnc��z9+���ZA�q�����Vͼ�� z�1���z�@�������C1yr�ܯ���'��W`~`�K|�LM:�Ykh�7�r����3��^�a�����'[i�����@���Y���ޥmVzY�`"�t�k(mnA��i���JX'�~�fz/�p�2��_a3UQ�}?-l��G�n�(�T���`Ac����8���E���W�#T�
��rF�=���1��W���Q`�r���6y�-��-���n�������ꪙ�=W2��+��oߘ��X��B�E�$�ʊT��zᶩ)�ς5g��U�K����	�&\~T�Z�5�%a6��0��~'\�x�/1�K�+�geRWK�{��\��%�q�꘍%̖���fXv�����Ψc�n�0י���p�֓n�%�����9�F�ZN�㱡�!�a۷M��x<Ɗ�~G�W���YŁ@2q M^�۹�_Xs��Vީ`�0HDd����?�HWWv���nWw��U�:�F������������7��5����F����֟���_�u����\L�0I|���ç���4ow��2�2�c��i���Q��KpI�(�Ձ�kru�vѵ�y3p��s���b�Q(Tu�U������;��=W[�P��3��K��(L},q��f�b�뚺.���M��)��!S=�nȪO��֪���#3S0�+��*y�z^�]��i2��~D�!2�,P���3�i*��ǩol��PŉYR�b�,�ua����з߭�M���M��e�/W�+��S[C�W�\�S���ߢ2�V��W�S�|n"`�8�b��i��j���*l�V��ht���K%�]�������r}qu�}"�v"�GgG�\�z��J��U��6��?�E;���$��4�8i�f�ƍv��xf���O|�ʶ a������5Oc���v��dˎ��qD��4�0�Q�a��Y+�/!��\�,��n�wbT�t�)CZ�n(Ⱦ鶏����j��F%��P�
������ؒ�n���m2�,��� ޾u�Y���2�.!>�	d��Jk��gYF�1+C@��f t��fTK=��+��d=ɒ9b��rbn�K���϶'���Yo��{ �r�O��1�D����mT}l�!  ��e!�4_�ـ��j0��:�#i7��4��h�����Vǩ�D0�C�c�&�̥G2�/�����t8����m>��*\k�M�ܸ�����wӦ�7�s]jNN��ԑA�by>�p@�(���џ�<�~�!o3�{��w��2�aN��}�|@�����?&W�?D*�V1~]W�QT�8����t��a��`V���{O'�i"�q��gm���m"�R�_��I<�;�V\ǲ�?7S�^߷^�yf�|���6�"7j0����R�k�6��*�:f��/G9�`�G���=d⿎��N����$�$zw����~[�������+V����m��ڐ�&��@+E;`�}uJ��{��$y��&���*�&9+������U{�y���U��W���.��t�e%��˟_�&��Ӟf��f_ɛ���1�����yj*bwnj�K୐��$7ǫ��z}��J��SB�������8������fg�ކ��~���:f� s����վ�]�;ɼߟ�қL���~�7�>����!�v&uӗt���lq���߾*nE����I���F\\�,OH�y�,�GO�ǂ�Q7��50\ ��*;��y-n/&����SP�kyy��n~�拯Ӳ��X^��r	������v�?|of^_;�~_���n��l���2�����|KM{O䦷{�����ւ��]屔�ri�׆�aQL��7���΃fvG�\�Ѽ�p�a;�2����`Ֆ70��Ȭ��f+U@'���3ɡ��i��j�ɚ?������C�߁�x�d{=�d����* "�D�MD]����@� B�����s���?�N�I@�c���c�{�/(�nҠP=��e�����%Ê��� Jc�dNQ�� rV����1��ʍ�㍛�8�����5�� Гv}j�v���p/�z�|w�x>����5�V�E*B�R򳿇��d*���	��E��O�<�%����Dd���`�߱��R����9>$�\���r}��|JKhW(���\�K�&��/���������|٢��Թ���Iz�_��,���)XsX5? �l{C*�B�讷Tɯ5�����,��p�x�Z֍P^�|2gg��wW��|�����)��ax��|�i�	���?M�y�%�/�rEς�u:�[˚'׼S��y� ��Bp�3i��?]��T��� |��T7�gNL���r>� ]�>�oO�"�������&�|���;z��?�r�pCxjܞ9� z,i!��qԈw�ʩ�@�}�if!1�=rd�ݑo�4�#��3�%DZ�	}��$Fn�Tj$#Rf���zBB7������"?��؅�@����u�`��U�����b���
,��{�~���o&R�'o�f����ܬ-NR��+X�U�Qiga����o:�b����܆���捻I�A��p�񖻢��g��$�w![@��O�@�}�����eٔ �Û`S�g�V����6�. f��$e���]g%ri7�~���������
f����V*��rq�5��9�(>w�[Ja�+�-�6�p��=>�q���+�:x��;F�
vr�~�ts�?[u��J��`����_����O�V�6k��K��N �莬A���ф�W���(�U����<�V(%/���J�By��;n�����mD�*K]�p��h�o��W�����	sp��[�=g�o�Z�mD8���\?[Arj��k*���%Dl�t�w��@�ީׇ���bͯۆ���m��t���.� .���KS���|�/��'-��4��ӿ���3<��6_���� +��x����=�돶Y���U%v^Yn֟l�]-<���ww�xZ��GC�;����\��

a��f?�J^�Y������'F�oL��2�W_�x��
��1�f,��B�.6�.w�N�@��P7�ŭъq��\N�eN�e�ceԠ�����9)�)��P41P4F�\kp��}��ݼ����Vu�����w\� ��NF�ň 풜��SdC��'��`��� �	oT�F k� �@yU����Q���AF���7hU��C����&	4�J���|(�*z�Ш���N��N@��q�V_5�n��ރ�n����*]Ƨ�}sC<��U���0���?�< ($����fn �R�Z�ub�(����!�|�R�*���T+�"��Vw%�k}f�l |e�^� ;n�Jw	�#�#J�z�cP1����#wU$*�	eyZ�7�-�K55c+zH��p���Ӿ�#Q�"f�%�ʾɰ���	3�2�c�dD�4�BP,|"$��d���So������� )q�H�H��������hA�c���0Z`0B�$�$��������=?�x�vv��l�������녭x�<�����֫�"��l��}m���l�x��y ~p���!�16�ͷDj��N/>I+�`}d n����7ɐ?ȩ�u���ji��o�#�w��&ip�,@�E���2Ƭ�C�O��C/�rA�-�`�֏ ; �z�o=A��8B�`D��\�����:ے���b��zJ;U���<�w�
2yT�\�{��*�����m0zPq��I8�%1t��m�oSm�0ӓI&IЧ�ޝ@�mHU�b��wU�S�D1n�0yx&"�� ���'��: �te�@t��4��'�R��O'�.��Y��һl:�����_Lо(��#4� ��#Om���i���3@j4 E�C���v,G"�Y'7���l��0�+
c���=0(�[s�ɖ�~8V���^?m̵Pl�$����Fb���[����~�k��	A���><�?��=M�<Ǉ�kK?}���ʊ��Kǫ������h�㚄���^��i o�o$[N��]$m��ssY;x3��+$Ç�Ko��UPȣ]��f>؄6����9��5��_S��u����N@7���9��+'���x���k��cҐ�uBW+�9�]B-������_�����s25uP64�8!1�ۧ^�0u��FA�3���q"߀�������[���.>��Z҂ �br����X#kZ��(:�����r>�\��0ab�A^+�j�+��0�@9m58I�����x"��-��9��1��Y�t��)'�w{!'�7+�
�Q��,��[.Ʀ�M��Ɔ�ޜ[�U&�=�6�T����W�r|����o-�Zf�x�k[TK`����[���ҖzĎK�^J?<�uI*�fmb
N}�l��T�ͨ��Pyբyp���S�~TX�.XR!%D�����8������:m��V�V��守�9���O��v�T��#w�?�[����D���N�>?�|�O�Y��+�A�U���q9:5
��h����-���_��`��>�"c��cڿ�u.<a��b�/E������ADyv��)� �ђ�)Y���/:��:�ز=oh��|��ap�Лѝ����hڟ�%�6�g�2���ち ~<���#������O���9�Q����21,�|\,e�1#/�ҁ�.y�C/~Q���4.�T�ze璼�J��N�	�;�˲S;n���WFpk���+�j��Q9S��i٧	����=�g>Ҫ��h
�FO�C����cx�^�L�x=zm2��F�o+�0K�Ha�1u����r���K�g����8S
0��{�X�wW�q�������s���ok-�&���(ꏾ��F4xNٞ��u8�^�G���|9��~�نF��F�^���]��R�~�1e��`Wj���Dj�ħ�ӭm��H�~��pU�g�R������>�.#9�p_��%m(؏�)���t�{�i�Ec�&��zs?u=*� �~}�� }�{;�ȺD�-N���`�����{@R�I"�LZ���"��(��x.J���C�:Xܽ�^��ꯘ� tN_�H�{W��#P�.�7}jՇz��h�0��P9���[Y;�gn	���/Q�0K����P�l^�YFVvvn���8=#c���o�3��_R�-�h4�p+x.���f_�g���M����=���m1��/�=9-&9�R�_䇡إ���&�bP��S����R���р���_+;��RN��v~-}�~�C�֦�?sjt�����UP�f`{~������-�6�W�{.Z�����W�Q�hm򫲎jDA}uy��Q��e!/���٭�"�~���?{��=6��HSt����t&���/x-����Թ7�{�{a����"�߂���QY���������y7�u)M��y�ƾd���GG�Z�a������-����
1�Vq_��L-�Y99�nmm��9�dIk���#���?q�U�Guk �5s�Z�c�|"��OZR�/���)C��䜀ʍ$�p�,�fK�sÑ0�a�~;����zޱg ��*��gP�:� _��L�*X/����!p�?6�ׄ���>t����(]%��H�;B2grj�I[zֆ���IR��x��I����6c�#hL�C�j���{��PkU���9��Z�����8H_��ۧ�j����߶w��;Ê� X����U� &��V�b:�q^�'��4Wđę1c5| J/�p Q.�-�@@�8�>O��
��.L�XI8Z7�
E�O�!�������}���M!>�%���93fL�ʄS(�j2��j�T����E�5ʕ�lNd�8�
�ԍ�h�Is=&��Y$"����hU�s'C|���8��u��V�q�ˁl�y��_�V�	��^v��5�粳|�{��yQ��2��������~D�a
���Ə+��Q�sfϓN�j��*�E �02l��	���QϘ}�6M%���e�s2q1��FYN3E�ւn�'�i��$[fi[�`�������~�]G,w�tK�_MH_`Pc-��˖�Ktd��;fwX���tc�7T6�Ҩ�}�W~�e��S�\��Yš�"��r���4�sL��,H�
�����d��l�G�s�� ��g��Rt���-�eO�k%�
x^7��?��

��Ϲs]�>Ļq��%U��^�!�RA ��^*m�rK��K������i/�"��B� �Zy���!���d|M��J�}2R
4�G�^��X� ��*��l�_���UUU����	�ֻ���?�@�?:�ߥ+C�=?���B'�TJ�|�k�m׷��N^���Ir>������s� u�*O͉���'ꃟrfY߿�j�x�l�
T,��]�������R�^l	��{}0;��u�+mK����Nѧ��{w���Q�����}�ܸZ�{�<��ё���D9�;�V�@J\r�����������[�ْ)�_ə�Xk���aI�����=s�ZjN|�<m^�Z��\G�a�O
%�_힜L�/��R;u�P�Nj�N�`�-�@�m俵���쳗_��O���lN?K�G>+�F��,`�t�n�o�J����u�j��Z�3]��0lO��^v�$� S~�ԥ8�'��'J�p������F�?㰖��KR�l������͵�k(x����W ��CT�ѤX��߯s�y,���>m��,<Ԅ��%$�a�S��O8�4�%�����HP[ip��1ݹe���Y]��#te�-3�Ƭќ�;�%�#p �$�L.멦u�D���	��	x����नS)�ǃ$�O��x�Q
�G�13�VZ�r,?���a��F�4`#��39ES�K�wwJ�(å�n�|��Ѱ�g����'�A)棟��7����H��S�QK��J�*O��7J[代X�S��kI�A�ر���3��0���O���M�E���������+� ?��\��7�=@�����z&ă��7����h�����<���by�0�;'5��x1x���_[�u���e�	��t���B����'�ͪ�Q[@8��`�'�����#��zv
y�������ng��N���Q�E_��O�%_֔))5~v����mK�˒xB��/��j��3�?'��m/?�9rX�j�qqq��>PdF(��	T*�g�
ɀr�������Oc�T��]`�[K�Xv�_c�J���,xe܋�2UPs��(7f3�(�-�o��O�AgE�"�yK�;1XFGl"Pw���L�5�~�������қg��O��9�x�N�~�Y�]�TF<觬��YI�y^4�%����e�,E�����uJ��!�A`kb~o���D��jb6�M$o�S����5��.?����e���ͷ��i�_f{S�9�}O��黎��tho��]{��u�?'f��|#�)��G�F:j���?����N�o���jpo鹂��(Z��=��ÍgG�ʙc�ګ*���d�G&R�8@���U�2�,[4B���`/\�L��V��ѮҎ��J���/��.0�uG�_|ۄ�~��9i��.��>�~��=e`�����umEM���ۯ��7)?[���f�nB�;�}�8�`�ov;h����^U��X��;<K���L�Z�EK�ɦ!<��8�"��*fA?�r��DގO��B��	ܸ��pZv�~�x ���@��P���<�٥8P��=}\0��T9���gj�:q-��K�.Lh�G>0Y����xds�������Mf;���y���I�J;�꛽���ی�OZ��/w���e���To-F>t���>H��gL��Q$�hK�tq:咮���8�.�gJ�Få�W*d`˪��oV� �j[�$�W*3���z6����D��P'Nc�z�mav6���fB,`�0O��f@I	Z82�9�3u������?���؏-�˥�)�'�F�EtM��S��\�M�#��1#��5��vg"��G��Ȑ�g^In� �F��w1+T(��;t��0>E!#�����l�G4ej}����0sd-e�� �.�o��s������.�ۀ�7 �=�Ba��{���D�{VE ����\R��wC,p�F�����qO_�*�m�K�=��4��s S�-�	Ѝ��EV
�E�2���Җvظ�.�]�4�aЈw�$W\w)�Ї(b5���_�v���ې���X�ݲ-{�(����e�k̠�N�� ����(�j@Q�%�S(����KE/f��B��I����/R���l �)�U��Qp!ZR*�0i��ȿ��v���T&��i1/x�,�,B�3%�*�s���Փ��.��*%;����d=���˓���H�
/�/�~W�������Wyj���I������|���=�I���N�K��%BYإ��fC�`�)��z`�0*�bHy"+����a��1,�]Z�t�Q���0_i	���:��3�'d�9@�Rļ�:�2�qԨ��߲4CVI���s(B��f��ڪu��������QJJjzz������t�fq1۠(55�]�+�5^&�s=2}�AG(A��MȘ6��611�@�f	��YX�nX����?��\�]A�9&;�C1yޣ
G!;#�Ps3C�Y}әY����l���7���h�@K�>�7���_��  J2�_�e���ʎ�@����������|��gp�,�w��w޿O #G?���gω�� �/6���3���D<[���͖h���J;�4?�4�����83���1��[�ܓ!9�:�Ĺ/��]��h���hU� ���*Is<�"�ľ{����nu��U����3������?��j�x��	�r������)O�|7R�Sم��ݖʗ;"xxx�E
{|{����m6�mW��V��P�_�6��)j����A�j���/2F>�}h��E��%gN�!����i���炷�
�W��H+�M(���$�o��o� ���;_j��_��=�y��@e��:���G����%��	դ��x��nLhg��Q�-q��w=�<r3�	�X,��8(�: ߭ԣ�\�0A�q�q��!�u?����x���v!��b�^J׭��D���-�|�����w�L[�h}��U�͞�`����ھ�,i�W�kYM��M�}CY��i���ۓ��r-�b:[��������Ͻ��L1J;�J���<iM�PjU�I�$�vaʰE���Q'��哥��)L٣��ae���Uw�2#��hE�0r�8Wp����h�"��l�(��4I�r9gw�9���~=+�Ȉ/�q�I�f%�-�,����aeT�nL���A���R���t�qS�n�4��+bk'y6hF�����GT���H���P�"���G�S
MIJD��" kU8�ӥ�`�e�2������=�t�?���f:�3|�o��Q���%7��	/���$RmӭS� �Z�����N.n;]�X���&��%g\b��s���~������d�bY�ġ�,%c��i�!R���|a@�S��F���!�J#N��]۳c[t����ĵ�1e1?`�	�gO�W1����a1�����%�&ɉ�m�e�R��u9xO���Mc����^���#w��z��ҪU�R2���ee����Я�a[�c%>��H�5$��F�2��V�0;+�g���C��F��V�󣝳3�?{��&b��<�OO���ѐ�H�H�D�@�A��!�#RG�JJ�yyI*���f�_;��T���������^�XGG����A��f��t���Cn����
g��J���҈�������.����#�ߪ�S$��4�|b(M�Q��*��r����-���H�IϘLK�J�~�;k����eCbr2�3�������O��A)�'�����t��V��d		���?��#�ϤN?}�6��MY��n�V�Zt�L��Q8��pFP��%�E����y�U�v�lZv���*��4���Ҩ��qc�9"�D4���Z@ϮX1�/����?��|��<���X�����p��|z��`�Y�j*�;ϟ�^1#0�ޣb�a�2wz���{���';tH8��=L5c��#S=����Eհ�cW?����a��a1��(xΐ�8�41�(~�v�zt�ñ���\�^��;-�X��9�ABG��llu~&��1���S'+ԣĔ���$
�'��;xdA�F2��D;��4{R*Ť�.ye�-�5����0hi �Co��ilk���Q
E.X��hܒ��󥞂Y�:�3L�w��
����2�F'�S@��c����:Q�Ha�$��6_1�>ş<_�9���V���	^�G�VN.t�C��. �����0����dA�2t*�l���+����k6 IМ���
?���.�⛫W�+�L�X��G6$��2�C޺u�f��o昊0N�,~����Vgz��yν4��ջa匿����GG���|�z; �����7��9��s�Ջ��Q�&�B�p��^�L<$���IXa3P|�@�QGs3���&�X��[E�����j���f~(8ē��Q�e�o]�D�a$F��HT��e���V^����/��߲�"v�D��O@3Bn7��O����'ܛ�to`�t�ck���l�r\���Zy�&�����ỏDyxy����o�����;�R�uQ�T��JLL�3KD��	81;i�OC�(Xyc7t�vא�HF�M�I$R�Y�j7��KFʬA-y/��0���lm������芕��J���(!������?�m蓯�� ��+VO��t<�ޭ��)#$�W�6�\��]�dm��޵�_���L�]������gez[��ݓ�ǆ��J��ڡ�v2���s�}�9�����x��%S�9�Զ���O���[ői|�X��ێ�D�di7<��`xR�;'� ����WS�1"�n��)���O�Щi&��J{��ɟw4�;�G�qʰBǫ���r/��{���I��W	���&[c�����e�!3	�)7I�	�X��J-�?��v�����Z '`����jy�<"c/��f��Јr��	�I�{�.$�I1�^ùRyT����UgV���M畜	�l?�̊Z��OƟh�h���ؙ�LZ�����]��~�{���������z�	�}���絎!�V�Ox#k�Vuwxc�U�R'߉OC<;?Н'���w}�܏0��R��D�`�{^���B/Wx�4��n��q:-]�P�Nw�w�<S|J��J��v>'������O�L��$����z�+3�B�ŋ���xT�x���g� �۸mP��E��*��?�8�����/l�NZ�s^�3���:4t�G�Y�%5�jmx��ӭ.\N@]�p�v�@E<��+����!����0\��uc��=���S(��p��_W�Z�}f�P&?��l��ij`�#6e��]1D �C�N!��p�;'�X�%�9��,�!�� ��UJ	�q�n��N\i�W�}�܋@�WE���c�a�F�/�/������m��]#���?��ȎG��i��� Rd�	�A��>C���a���9����=3K��:���K6���<��t����Ԝ-���w�\ff&���#A5V�m��$v���;��q�s�˞�3bzfz�Ș��g'2�0u�e���R�R
h@���3��<���]j[�,�έZ��YSW�R%�{G~ʒK!���R�[<ED'!ql	⋛<���$yP6$Xljp��!'������;Y:V6�{�w/��Bh��v�ѝ���(�.�T��R�ǼƷG��.���<�
��R���	�u~}�8��`�o��c�� !����셃NX����J�1�;�V��[�HZ�;�Gx���ՇZ�CxfG3�{�Ye[�Ujy�d�Xd��B��![V.[JQ��l��?��}�f�uҚ1��6uԞ%n���d��}����b-����.�8)a��ۢ9��%������b+[\蒭�^O�F*-���>"A��?�{� ��8��N Ჯu�u��t���s?��"1WÓNL\�}�����|���@Q�DM��}c��k��_�ñ��vL�k�y�9��X���X������&
��}i��5�,)����
�8i�;ȍ���~����8�s���*ͳ��k�1�(S�C����OP\����YFnG>,�c�?�G���dة���C�\ȓS@f�Z���Ť�f���(}�޶}i�hz8���-<�f�@q�g<���1djt7�'�L�5�5/$|�Q/�W`�0��	�)������d+�''�J_^l�K������|w�	s��%�20�٥�d�����
7�^���A�iU�D��XPK��I����m��Dɥ���%8�>��챷���r �(����2�6Ė��k[n%� �J(1=%��_�
�����O��*g�`@�����>7� &Ҟ�q+�/�vΐHFv��a�@�_�E��\6���<ݻQ<��!cs��㼄�E2e�Sr�չ�Q⥫�6��Ea�}�X�+��W���Eŧ��W�Z2M�d��dee��;F�T�*���o`gVN.`��Ý��c�?�:�p�C]=����VXL�c~}:)_��]:���'gp*�����ٓ��N�ڟ�����J�d|�5,o�xc��P��&�Sk�8�����R�*6N�{z���q�Tpָ�=��(�dG͏����ǆ�t� ���b9n�ٿ]O��7x��������Ԍ�����NXeMm�DMuUe���v�e�݂?��r�K�<}�-�G��ή{�-�����Ot�Tlr����"zoru�@o����R3��bcV��P.�Y�G�ݬ��]]���:��/͙_g�j}U*ڻM�O��3��2�Ꞽ������G'F{��V�"<d�=z
����yˆ�N̤*Z�H�"����	�ⷅYA��7�{�x��g�y�Q�N�"�只���C��Sy�.L�DQ|��m$�}WoO�`{
��5i�d~�Q��+�1���tDI ��A��\�
R�4T#��Tv۶H�)34��[�u�8�Q�ģ���� ~aH����E�^u�Xd?+�]Ѷ��)�Ν�{�-4�1�����JH��e�� �.���WƷ{�G��}�x�l/l����i��T�/�hy�UA��l!����Bu'����h��U�x��_�l�o� 2J
�I8W>�[áO��4d��BSx*��(wt�l��v��'�O����䖑�O�Y�>�ߢ�������8�:����#`~"fSAx���R�+!���5��y[��*9��S*u�����'�4���+ xp���y�3٣�77E�@N��;�4}%���;��2�~p71m���L�H5�d_�X`��4NC�r�@#�ۊ@����9�>�(h�P���H_4��"�x=��̰�4�h�5{����i��'�mV�u��]���� ���͍���щ������(�H���*���w�-m읚��$���{{K�ky����N��6`֙��Y���؋<�]C��j�(����]aV0k8�gl^y'�`o�	[��u``Pkмv��fB]!C���[��E�����ϙL�Y,�tl,4�� C��\��Hӻ�?%�LA�˖��<~a�X�-��z29A��d��)������_g�^���B�cȐV�T@�����*�W�w���<AV�i�Y��̋{��Sc�c��װ6)�7g��`��SV��-\�n�h���WJ`s	^"�پ�Ѯ��Ɏ����������^-;F��D;��b�(R�ר>X7�����h����.LoKQ@��du<�%\�_� wu(a�R���c�a��BN:<�NF��-8�6�W��M����j\9ςF����{:b��O�P�]�Y]��_�;&� ��M'�;�m/�<�g����.�D%�[���N��l��s?���ɧ�6�����A�S/q�鍀�����V�GK"l�V�4�'ҮM��b��OV$�1K2 �ڰ�"I�K���a����P�ۚr�I�9Uʧ���1"k7V��q�U��&X�Fm��%^F���ϙ��2�z�c��9��������
�2����u��P�)@�A���/��G7:���b#Nu��<�a[����:x�FN����&UȒ�6�Wtj
�(6?�^��"� �~a!�㐌�8���)��W��(j�J^j
������*�$��1�5ސ�ݖ5_ǥ$����*���f��6�B%��_9$i���[+��*��ɇ���<e�ұz����Յ�;fRew�y�[^�)��x�m�\A������$	��ԟa���اzH1��*H��X�K��wt��kT�g��h������/�rJ���=�E}	&j&�l:h>�������������]�<^��q��t�N��^���������c�C�\���.,e�8�t�s��u��rqt�u�y�6n�����D9[ٽ8�L� b �W���n����V~�A�e�Qy���s�~1��ɝ��Q���Cٖm}#���ت��Ml�=o��<`9���?�P�B�\����i�������FT�DM�pU�DMU]e�D����7���h*�L�*	I��*o�TW��5�|�����T{3A�[wM5(e4p0nӛ��[�o��Ջ�����fb����>���(�q�|���L��L��Kg�ϑ�l��s\��8��$vݷ(�-ר�>h�E�	i�����0H�E"�ma�VZ��Ԟ����q9J�b�]F�b!�Sv��BMz4�RI�����ukF]d_�J�B������X�v��x�Α+ࢷ��]�]�+�A�bP�w��˓��ª������Tl"�w 7{.�Vf:>td%@���]O���������0����o�Lj�*{C�y��Q��-�k���˗y�3�r�)I�`Ř\�E&I�����b�c)��`F}E�X��`ɭO�+�DF�d�x�� �5r�8��R%��g��76����~��s��J�x���k��SUm42�HG�'��+Q���Sꀋ��仛�h�1��f�l(�ۆu?wlw�U�U��R3쒸�&�&��K�mtz�:�A�өdC�3�ɐ�4"���CUe;�����w_s���ϯ����G
������q\����w�چ��\�>�kwk��wG�����(ᯥ�)�'e"�)�ӡbf�u6P聂�#�M�rx���z�*��o�K��΍����9{ʸ��q��6m�Hޔ��ە�M��wk��	���jV���EeS Kɘ�Xf0��N|i!�����p����-~���W�ٹJ�ԲeG������o�u�L�׬�b��I\�6�+�\��1,$�/)6�+�sX�fV�sد�6�h�b�}�z15>���R�/�<^��Oܷ{X�/X����L����I6�)�Ɇ7�M��m�&�Z7�
�)����x�L�/�R������Cc�+ݫ�.�i�.�p�2��s�'��g����Z��`�dop�X�������ٌ�haUH|��@��&��������ꁋ��7���E�Q�	KJ��X�z_M��5o����;
.�������lk�i68��m�s�曆7!�VObh�Ύ�12�@��������k�Xu���Վ��Ή�٢�~�5��ؓ�!��A�a�ԋcȱ�����`,���_N巨:��Y?ҍyڕ	sx����}zTq�֜���<�� A����"�a��$'������[�D�@��nZM��y�QA峘�Zb�m�}Phmӹ�1;���ؼ���+j0�p
^ �:L�^�*�案��H/�񀖇u.~+��߼�!�nc-�w����rǅxx��/T��[��Xkgݘ�p7;]CCָ��2��ZbQ���]p��jRTqX�E�ӿ8�E���b�>mEg�7h0�o�����2�h���(��wpQ.�����~:�a4��1�n����O�O�ۏX����#�f 95�/t���Z��(��.>�hx�o���҂�'p�����ˣ��;�é왿�>lu.�<�,�3�R�&��Pl����H\*��!:-�W�|�yU�j�/ŉҘ>G���w}��@m�a�}Dl�i��\X;�Mx�-8y�M(�%� oL<4n���I[�}��*a9U�9�<鈑�i9�B��$��SZ^�>'
Rͯ+��������7wM�ߞ�n�pӓ��5���-M����(ue�{�wR��mz-L��)��n���RHg��; "r��3)��q�5E�o�1�����N_z�:5j��x�8&>_�&��"��1�~������t������ N�������S���֐����_QJq�x��"7���O��)5���*O��nQO��D�l�(����r����7f��&�!�Բ�6�\�f��T9�5�G�dЅ����^Ӧ��oL/~'�?����}ۺ5��mS$�P�?�2UGc�y�v,�޼?w�C�'�5rҖ��l����lQ�����ZT��
�랢����ޮ���#+E������"-�I���JJ������{���666}��cC3?fF�G�>к�dU�V��7� ������,#.�m&T{�����>�JT>�x���F�:t�Y>]��?)_��Q:����ا9�4�X�h�6��9Y��7D'���̷�.W->�J�(~�T=Q�ѝ*.׬��s:kDz�c��v�
HH�Zq?�����z�S���F��( �#bH�}�.�L�����yY�,5���޳��枷cnp�Bz�[�s�x}y�����h%_-�M!�*2��?z),&f�9������|[U-�b���z�К�͘�U���Ϟ���_��d&��L��������yRՒ[�to��z>����bn����j���`��Gԋ�펄�g�]{IN����,���O�gy%��@6�.ˍFP�旵do�m�ߖ�g��u�vR�m��F�x�<S��~��r���j��Γqc������zNc2) ����ߩ�);�+�ϓ_(���Q�F>�ǃ�BFN�A�V��
�a�E�?�A]䑿���PFnݻ�A7�B���Α�̊��2+����i����Ԛ�w�gw�.����n�k�UP�}
jz


��e��Gr����s��%� '"	�ⳉ;���WGڕ�-����tt�X)'��ć*��xC�����!�z�(���٬�q/�9e&��3�Cj����n6���wD.]�@� ���0q4_,̀7�i	�p���I�E�=.@��� �wrTE�a|$����<�W|y[�n�lN��%�K��5�)dL��f�?&�u84��c(�vr�S���I��AyJ�TW<`�%��!F���?�Q�_n��}0� 85*�%��u����a�Y���Kdj�Sd��ˡ��#�>O
͛K�l�]ͬԡ��S<�.�_���V�9���A��D�k�G��κ�x�6[k�i��B_*=�I�Kv���]ф�9��)��_o��a��T6�g������{�(|�d�Fy��|�Bhq4�<s+�Q���Ѻ����w�BoϪ[Z�6��p=���lH���҇�m�'�>∔S�p�p� _�tWh���"��/P _�Hu�+�"�+����-+b:�>C5舭��ԇ���Xz���?%[�qj4�q|���v�#���c"��G:^M	����g�����㌖0|K5w�	����ArAO���<�װ�]Ԓ������3�9�3_�ʺ�f�����v�`���=^���U_H���wL��z!�|��O��]Hx�I���S������(0��%��^�⠺����dm�rm��T	-�m�&8�>�&���?L��|������f�2��=���[���a_L=?�B��2>v%�B���r/}ͦ�x�i��ns8��ȹ<�ř0s�ˌ��,�����C�Yn����H�ɩ��`��Em4JIbW�i��U�} �KΉ���6�WUp�$���?eMG|\�o�� ����k�-��;�3�03�;o���cKi��~ܝ�	���y^��%D�~�}o	���������^���3�z�jxd={d�-aREv��F>?�,���R{�|`0)Y��qu���(?���Q���؏uI_d�>�Π�ߕ搽�[�g$yc�u����������۩*qz���4�(������h��(%^L$p�/A5�U�^���><��F�x�u�D�H.W��9��S�R��o�۩�:�w+9ag������)�Dgg��(V�R֮�;��L��4 -֯�mJ
F�.u���nŨ��"�yC�"�aD����}�'���S�"Nv~}Ql5� ��yN�����%Z+�8�z��A���y?�G��43�~�b9�߱�%�xN��]HV1�/P�3R
�8�@�n_��G�x�c,լ$��>L��D�j\�ZA"��ؔU���ib8�:¢Y*b,��-n����HӰ='�P�־9��GO�ĬaG�%~of�bH�ŉ���HRH��p��(N�OU�+< �v�2T�?�gYL>[��j�pʦO�nV=+ƙ��':Mi�ӎZm]�� 9�TPX�	���N&�g��l\�o�W���u���~�O���G��Z�	�AE�Z�0�����v�y�A@A��k�u��P.�*�}��XN�8�v��p!Iv�X�N������@N4����e�j��>H�'A��pi]��!��K��ѫts+������r��y�Sf��S��~����Y�tWG(��'6W�'�9�wdC������y�)�l�P�Mo\PLL���SCCC@@�����Ȉ��������U�u�^�d]vfބ����wxva�!6�3�m��z�r�-a��\N�����	�I&QP��#_Uo�k:�+�61����$�*(GcK��ǡeV]��~+�[a$�=h����$QIޅ������6eu;���F5����{��Lv-:��;D�u���f�s��͍�6���R1��=�Ѿ�F������"W;^o/Te8q=�Q��� ����q?��!ܞF7��pO�Q-��p��J(�U��s�5�Lmp�m�}b�<SL��ŋ����"7�z#NP��ҝ>��p����F���tbh����%w�bD��EA��s��u�x��V���@�({F�S|�8�##g�b��\S/`�d�
�Ա�+h�qFXv����n�i@G�D;��x�����ʒG1�`|MU ����؍ᓣ�����V�N\'T���ъ��`2`&P�Tuh�Vn��7�mqF-��'­��i:�۟k�睆t!��>k
�7�����������%����n�Ot��8��$��$�2rI��#}�/c'�ju���j���qI��;�����������y+O��E�;�B�]&���²$/������z?څ���&�1$�@�l8��Vge��~E|�YG�ޤ�J��RQ,Zn���F���>�C�`<���𼩍�8Sޡ�h W��dB�wJ��o'�v=R�6z��T����{&
2>FԊ!p)U$�m���=K;�Gmwe�I:L݊�SkR"�|AP�����rV^yK�!�7���@�t�$����`��a�`��H�ޗ.pqh���$�)ڜ,��wB���{�a:F;��WZ�6�8 �R�K{o%�ǲ2ܿ��Jt��.Ro����� _###��r(3�'�'���$��[@����a��+�[-@�@�%L�Dq���F�.��1�N��s�x�'�f� *��������e&D�]��^� ,D��oXK5o;��O�t}�&��!��0��|+Y������XQ��:4"@�D�ն�0�_���:����nV��� i��*�V	�O�v�T�`	���gI����s���m>}�3�`�&���j����z%pɌB�j��}�
3�|g��Q�%/N	����T���9�����UA�:����g3l�w���kE%j�%����
jV��A�Ml*�^�(5JK� U��Z�W�����|;����%�/��_�s_׵���U���Q%k$����W_?���G�ʀ@��8�@o�b���'��+}x����U���T��,����V���l��e�L7��\5\&���Z�������H�!���<:�{,f�v��6�9K�c+B#��h|�|� ��W��~tw+��]�\����y��|���ώ�����.�xY1V�40�i�.��=������aJb��/hۂ��lޱd
s4�Ǉ�]�gs�)gh� �R!��Z����N�i���U�+r\7�Y�Bp�/yo�S��?}h�ZT��9� U
�YkN[1[������([|oF�Ǩ+�ؠ�z�G��!�L�?���KJ��`x���/�VM����-�ci��uJ�I� �)��������}��YL���qzԬ��@p��R�yF!���8;7��^��v~��{ui�"�ś?�jN�sQ���_�c����v�!	��p��V'�E�g����k��"=/�	щ����c0TR z?�sw��H1'w�j"����A0�Ȏ��Ȉ�in�ɥ�ld�O��ڹ��6@�\31*��>�q ��s��D�W���p
|ه���rv'���iz"'�K���J�b�gX	4gt�]P���d�G��Q�	>�������͞�K��Z;�����!Tu��{N����qTM��)p������Y��������װ��#���u��d2���D�^��x�����^�<�g<����H{��xP6��H�� ڄcؘU��> Zs��z���y_$!qe��5L�w+~���tJ���	}~	�ri}�2����`�n��R)����8�9�P�b������Q;�99�k��R�Z�SX�������z\Z^�<oee�+:KK���&q.�a����#����R��r���<�����y|cS��Ǽ3��%���J[�d8�,�G��k+K�m��nƭ�D�ۢ�wA̦YQ�v�t1!q�A.$�
�8cs�U�1���i��U��'Է~7����D�8��Í�s�ּ��w�ch勮g>�`�_��+��ua�9U4%��]�&c��/*j^�AMf	��Ror�r��t�y�vgg�����fw2])�������-��
����1�6�^2{�Ar�i͐��I���~�|�u�d\�������j�qo�y�`�R��r~TO��H8�|�
��^ɓ����U�6�bX���7�;��Zy2藯���t��~D'���1-H�^��z����|����	�jl,�ڍ]�3V���/Z��!<�^;�G}�[�״�w:-9SN���7vd��ӊ����O'�R��������z��Z�ɒ��*&�ͱ���C_i��x�c�%�i��|��$4�A��4F�]��+:�<�O�z��MvNNv��D��X�$����o��Bv6�Cf�����~l��a'��U�Ɗt�U���_��=yZ@��,�{�[k�/nE�#9�\�r�G��~���=���|�*y����	�_��"��p���1-.\5Q=jW'��_���	s���y)/o���ޭH�k�u�Q�T��r��Kݤ#F���,�.�q�3��7�
z�u��K{N�lVy �ѥ9���vE����W(�i��o#�NY
Q������=j�Z���eD����~�|�<�E�N'�D��X���2��ZCX�&W�Q��<!��e�
�?���1���`� �p.13�J;�jB;�0s�ZN@�'�@��[`5ܺ�'�E�G6�k�S�\��Ÿ*���=*v����z��I�^BX�}K7%h�힏�h��7�jEc_�] >߀�u����\J2k*�Ro?��
r0Yf��4o�ǘ���֪H�4~�����mF��j��t�'�o��'i�w�^���� u�\��+�p��pf7ӛʜ㣙!;r;��I�C��Ddt�wD�A�ڶ &�����&-�l�(+��uF=ާ�+A0��}$G)����녟�������V�Y��P.�U��
W'��cq0��e1�x��2�"�'����b����9�p��묨O�_������mZ�ۅ䭀��=&Z\:�\�y��2��o��w�3,�!w���	�>�47Z������ s�����m���I{F��)�ʯ+̺ڂ���xY�T��Y�p�ʲb���bkk����jn�K�9u4�-#��o5�\��M�Eǉ����mq�BH��J�3�-�5�c�˼=%���=�����.�+y?S�T�"�&%u
�q������!5kBO}:��qer\6-}C8�Is�CU-�<`�j�8-�c�v����li ����`b�ۋ]�Z����NN�.����v.O�)W�I�N|&[��U(�#�GF��� �����E�Ky_py yF��Z,"Ze�2�V�����F9�0h�!��ޝg�H�M���
�"g�!���//�?@�0y_�� V.�\�	���/��?��Y�n~��<�[1��R�m���c����%���$���r��Z_6���J���rp�:K���=��w���:ԜM�˼��&H�峷��BdgIBQ�d�ZZ׆���� 2b�l��3\����c����b9��P2I�7PB��`��,>₞%��wӠ.�Y�j�V<��̓��'�d��'����O{ӾD��R5���H(W��y7�\g@(�X��j�n ���`iH�ר.���X��I7�֡N����է��j�1T^莩�}TN�D@ ����'���=����uA/��zo.��Ta��L�%�m�q� eb�3��/j����
v:QX��㡤3�'#�c3� |������e�i��hEt)~��|9	�<�&�*�V�,��j+���Q��:�*���S��%Ѹ�xKME�	�e0+ݕ�<�)y��u��()��Y�Gٿ�pz��Z�����	'w���_�a�IGI4
�Я(Odk�ȧ./�N=d�|'���9j_�6{-�x,�7����ʞ�H�}U(Rݚ�#AR�6�컢�_�1���x&��!ub��y�Ύ��K{�1̃��3�ǧCq��7���U#(j�!����.~?:���
�Gt�NOL���.��^��p���;�� ��K�n׷4/#`�]'`�-
�>�j��sO�K��n�����EE'!��-:�lt\��;X^ǑF>����O�8ϊ��6Z���?����;��L�c���aO�!<�&���& �>o���"�g�>�`�iS��$��D�D?ہ���<�=�i؝�<0�	�7�~h�k�X�漣͎rk}�>`���G������okT�%��������FC��A�轚�����#�*����Y��e|�ݤh��C�-Ú�[�Y�7~}Va�/����#q�~rO�m�1�l;�T�1�x@����4i�&`�J@��Aߝ^Q�������$��8	�Q1���v�D"ۿ�xUt�%p
�Cgv�?30�=5pPo�c9�y���L��I����̹+F����Q��6B���gv�Ȭ)xŋI^��
Ì�Bs�\D�r�<k��Gw���?� ���r0Į�ѯ(D�����c������y��� #�l�C�@��D��R�UV:����$_�I#�� rp"���N���}��C���rQ�sr֥�i��?)�\`'�ݷ�`(c޽>ѐ���>o�l��sN�?��ґ�7*��������uoD��qܿ� E���� �#��2�4�KݿQ�!��"F���Phg`�P�ej֏d8���?��W`�4����
C�@�h�G�(�]�����x�+}M[���%r�\��mt1�ޝ��	��͛�A� sJwo�/�?�"�&Y 
`�(��1#�H�,n9���K�6��+@�R�R�@#"�}!
甽��-�|b����n�D�8QG���j; �e8Eo=<�n�+�Z�Px�,�32xO�_o�	�-��'�:�`SY�'W�� �a�L¦��&}��K(ۯ�L��>���=��/�Cy.(�E���44�O��+�l�v��6N:H����T����9ҰIS��T��98��C�/�l�JqF���;��j��v~
uX����_���Dߜ��}<�uT�f�mC��Q��#�gL�&��:&�J�+�	D��A��A����n((E���*��}w4yE�DR3������P��4mJ���-k��x����"�Sa�!��!���q&���C�7z�G�-,)��tT+�4�  R�ӫe2)�0�=�ft�mDGh&����HtI��ɾ�8�T�ܒ��fY��Z��M�������{��Հ,�_�bR� �����d߶��&�w�ث���F��w�̮+o9����or��=}�E����1s��	������ʘ�0�9��j+"c�U r^�Q
��"�.�>{�ϿƇ���������C篘�.�C`Oez5*Z6���o�_��5��aJn�2�K;�Nt�~����3�j��||cߺPj~�xc�wi��װ�3)��=CRJ����,g�t���P N��mW��!������L�s�s�g��7q��o��N8�m�\������m+��Ӷ��&P�[X`���.���(��F��9��A��?�IX���F�a{g�9�(�����������Jy���p�s�[�I}��(zt��`{�����r�>�G=\xn�X��a���ohq]G8U��ڒ�3*�l 0_���BI��$�'R���1]��b��xn%��\�QQ�B{ו��_?<�3��w�P��Z��6�̉P�n�B���2��)H�c�F��M�]�>�>�����\61�6pޖ!t13%�c�h��I�u��Oa�O�p�H��l�~[+B� 8ի5�2c�v������86$��-~"Е��*�����_ݩ0�����p�Α�X<��lϣ���7��L��#���K{D���7���[3{�ŵ�K�"�P�I��b�� [IR�g(�"9~����$,*Ɔ;�;!ݐH3���r��(@���5=��ጐF�|�~�wY�#�;�W�~~�ڔG0ƒ��K�|����Ƙތ{�����1����o��gssf&���Od�rL��%.���ݿ�$����s�t�kN���4+|ịF�m�Z�}<�uT8	t�V�[�PCD�l�����L�Ê1J���("����J���{Uc�IX0�!�`�e's��2@1����5K�i6i��.�h�g[���\B�/4�� W?�EO�z�uѾ����ܮU���_�'�{G�&z�{��G��>�Ho�ǥ�S�E�:E�Q�K��3�Xs
�� �%^�����8�1�<`��|ių�jU�/X�/xƌ𧻓%!��!�����8_�p�R�֝ ���_�S}%˂��D����Ճwݾ�u��Ȉ�*T�ua�h��N�����0j����>y�E�Ȩ��ЗH�9�����z��*X*�M*	������}:n~�V���a�\K�dy����C����E�p����L��(7JyB��ٱE�3آe;K�2�*�$	p�T���,_,	��a�6�r	*P|�-byW��/��I@��]	9qD����nt�/����,��(�s�5,B9�� �?� @��rв5�pM����ŸI�'���4�@Br���

�Me�%�^�0���|MoC'\�������[��B�,�\^+Uia/`�@�T|��0:�"�8�������K�S/�cgi��NZP�5x�o��uV�m�I��#>h�y�+Ym@����F���iz��^`����$���%���}�@��B�s\�
p��X.D������N<�)����\2$B�����Z8�J�K~WC�װH��$	wuMCh='`~���}�7�[S	��3���_\7���[�.��"�E��{�����kQ�A�2?<:V�M�9W��I=���`ge���S���JS�N����V�X��g_��q LbO?eT��c
6R�x������*���
�n�M�'{z��t��f5�`�}��liA����MH��U��y��qsL�����Ҋ�W,ރ&;��P�Q�2���04B�Ϣ�6�W�F���ң�S�l]ɀ�G��e���a�ߑ����jtq�	H0�^���آ��;w2�n�z�\�pZ�w����2tI�'����}��籑�f��:�v3������5\<2�G���Q����|�$]��̼̥YsZ
�`10d��� 򄢚�(�^p�Y�3ك����\$NBK�!!�ð\$�v~p4��Wd�x�|O�ǂ������������t��٭��6Y��2�;MG��t_�R����q�W�ryɒ�]�M�`M
^'{N�Ug��إ	�ld�?PϨ�x.�vsA�@���7�1�����,���v|z�\��-C|.Py����1�-�ϛ�CU��rJse[�ܔ��]��(f��0�n�(.W)�S_�o�Q�%��м����[])�lf���38&���=��Y5}r
�j��R�Sm��O�
�H�l�m�Cnk����U.���({7����G��H���������qbm��5�3И�A!�r@p*:�?�m�C��O�\H��#	�/c}e�QA���|[�����=����S�Q�f+b6f���d���G�����T�g1]��k~i�~��"�uUِ�lD=��ZĊ{����]�n��.i����@UNz���V��m`����¬�^B�isǮ�U�f[��(��3)Ce�O���=�u�.Tʪ��_�c�o���0l�AVD����uCC[C2m�Ie�S���ۇ�ʹ��i,�t�;�[�wm�]�]��J�5+�����%p��h�/;y�㮜*Ƶ��Q-Șv�M>��	q�S�xtH)�2������,����wGK��m�������@�Ң�2��]c�EFo�/������+J��k��j�9'�T�J���*yt����"�o�T�����2$XN��*peЋ�ݐtԱr¡t��v�JT&������w��w}7��ҡ@f�A�sN�0J���8�	�������ZY�e�V�؛�&�!����u�����%��,M�)ӽ=��B}\n�?��I-�JͲM�
Nmu+Iz���>���Ǻ~Ū&��xo����]�����dãt�מ�������zHd%eW��T�e	M�;����*I��քz��p�p��.�3[���Qaf�]h�Hvy(���x�����j�Q��+�r�C�l4dD-��e@�k`Λ4�[�w�i���v-u��ͫZ��Q횑�F�I��q��yA�2�a�/��t#������i0HpW@؍_N�^�+2��3��Q�ۃ G�`��á����ֱէo�&=Y��Z���GrvT�@��6�
3`x��$m8z�ʙ��|
Z�aR{pbu	<VR�(��8e�ʞE->4�.����c7b����~F��x/pą2>��`��
����
[ga��d!���鲤�}&&���<�� �&	��k�E��nf�h��,96�;\��
�K;��y�J�=��!����N�*MHD&�?ظ�+�����,�U��s���M�)S�c�]��Վ������ޕ�$ǰ:�WtZRb�/c"��eO���IX�/q�h
�_ʱ�Xq�M-:ŊXb�O��4ZO�_���^���l����;i��N$�X�B&-�@�b�ԏ��a��S�6���
�6� E���Ώ=��|��-c�/�ё����Y�c��!	
�?�����h�Q���Z>Ue ��*�C�2ЎS���uL��b"O�y���Ԓ{pӿ��	{����|����l�τ���jS�x����g��	���!*�����%�Y�|�I�ӗ3m��v�هB��֪���Ư�������H��ѥ(
`�eM�F�y�7��Gٟ'd!.��e�"�NZA��$�  �sh���aT/B�Y�Yz���Y,4�F�̲��I�ҏ���_I��<9Z��Ηv�ߺ�P�g{rx�$wB�Z���(1���'��DrQ�pcW��e(�2I�!��F �S ߦz�yoe3�[#z�slly%�?.2��"I��pڡ��Q�$�x��YV�#��ե���Γ[_�vV��u�8�>q�7�[�bm�"�d�3肕�*Xl�y�����>�@o���%�zU�C�hC�F7�+�a}��� �2��{�)�px�
�p�fm�{���=�`�W�6!�>Ս-*R�0�3n�)�
�����J!�6r�LD���`�V⃈B8��w�D�h�rG!&t[[��]dhx�0�?g��3~A�F����=���8�D_^��M����>������(t�S�����J�*��mP�w���`��N�%(�{�lੰ�^ļ� ,���W��� 	4���q�$	L�FW{鷔�s��vS�_ԧ	��IePҰ��Z�.^��}H��_�$Y���~���ã��C�t����'9Ti\вB�o����Ӟ(a~���JGr�*��ʖH?k��C�����|-�&{W}E�|�~:1��q���	>����/��#�����*H;hQ4�I~:���@�={?V����P��ǜE龈Ӂ��D#�뒻����P�H�W��i�x�o�f��2A`o���O�ػ�~���S>���~�:!;��glfJܩ D�����x�W�AGW�e�Rr������&���0L����9��9�-[?�S]k���K��4;��R}����ڊ*���O��.��H�*qӗG`v����p��qWo��rc{��ɐFS���ldZ[��J�:�=1��\�����қTK�jw�
s�봊������J˫l�P���MIu�L��؞W	�!勒�	
UQ�H�}2��p���v	� ��ȿ ���o��L�'9�i
g��7�!o�>)H\��7*tz�`ǫ�
W�7�n�o��n�4��-��Qk�]A� s&��%�9�x�?;�h:�4��P�!o�c���e'$���4F'�/@B4��Q/P.��	�a��S3]إ�#�d7��͞�z<�u3����*Ӝ1k�"�`���6���շ9:.Y�zq;!��?�3.��� 4|��r���<�N��Ηyu�U�Kz;0�����������aŢ���.$���M.M�n��h��{Q���X�6�S[FQ�"dp�B ��cyt�] #����� ���$��4��#�L����D�Z8�S�م9*+�ډ�z��@+ �>�)x 	��֐�r��"� !�׆�qX���o���ɬ����U��20�n��c�j��{
��FQBb¾p����,v~{�֧��@�-���E��|)E"�m]��!�?^by爚�p��m��sU X'q��x��[t�H�I�X�s+��|��{b���W�B3�{��;��8�R<@Aj�R9l�|����q�,��� �-�J��4�����5Z�x�J���INx��Q���9����y���bci����Vi��_3j����J�,�P(Ct�R�?8�K����oU�x-��UJȎI�պ������'8o<|�����%v�t�*U�9 M*vK���j'� �3L�S�c)P�\'۴(J��p�PsS	v����	>ZH�� �M��)m@|���J����$�W�R��SX㷫��O�d�j���������p�����}���n��xW2Bh���Ȯ@���y76o��fZ�K��U_�:������b[g�_eZ��kyum{s������޺����˗�c*�]��u�H�\��y�a9�˴���y'-	p��Q!���$I�f�ʴ�P^����E��d�<��Ll�l����߽g~/���r};���I���V]{_�\'Wamv�7�#>5=�:y���1���1J���{px��$��bz��d=^���Vl,L�+�w��V��C����[�u��G�6Ie�u�EsS�� W�`0���~��yo��X+�;yK6i�A���
�������8A6�V������gSI4\6�w]x]N-J�M�<��nV�������OE+�$C#p@�S��F�F��L?���c�Q�#��%
�f�ڀV�l�/H���LS����� 7��j#�K�g��8�wP����n*�f0� �����A��X������؀B�r�:��q����i�h�\{M[�Om�6�gt�K��F-�+��om���$�/y��ggǒ�*&��|��A�^��[A~�n�ny3%D':�1b28��=��S��v��6k��P�n��"�k���n(�ܙ'�Nq(�����ϟ
T]�|@;���4E�9�?�-��t6�Eu2 :��RR��J��¤0_����k,�]RxE,�q�V��L*�`��?L��X\D���iQ����nί��	�W�~�����:+�v�+3�V%�i��^�>�^�a8��M����b �M���ȷ�l �ۻ�ή����WQZO�X�4�9�k�y'��V�(Kx�	�P�α���H(����&�
bH��I�EG����>���=%y4ժ�T*�I��m��E�t`�M��!�\�A�G&�h#���$�YȪ`bD=����[A�Ft)�x*}l�p�?�T���6�%-�G�9�����P�Q̧�D�cvÂ�r�mBϢdȉ�`l���{,���\���
���Țk�W�R�PT���4�������0�%|@���H����:,u�
M���$Ʊ����ݑ�����H����<�u�rJ(�θ����[���~�%O(�&d�5�g$�Eq�UĴ9f���e���t��\NN���,��ŗ������]]�wtD�__]N�YY+��1�5(H;���k��x�L�;�mhx&�E���W����������u"b��������5�M~{��M��y�Y#����a{��9㗚O���%R��&%�������㚚�"�J�;e���������1�af6kj:c�M�k����e��Gɗ��%���Ý�;�9�v	���9 ̶��v��.��\���9��M%�0��Җ�YIbV�aº���	#�* )-��p(��p�u,�;�(�;�{W	9��lo	�i(��ޒ���.~h���Y��w�i'v���z��^ `�������m�.p�*>���r��Y��fٿm���Jc��������D�-z�ɾU~�c�J�T��?����X��	2�L���0���1����'���l#�%$Y3n>a�a�0G霍�����Lq ��GK���V�����<Xd�r��;�Wp���H5KB����5�d6�������8�l���_��݆����Z�A,���W���?f�9^_���	}�aT޺髻\S��qZ\��c��M��u�}���a�a��E3����6PvY�0Kv��\k�$s��:�8�\ӟ@��g�H(�%��Di���d��䃊�	bu=4��Y+��ӧ)?;��+e���$�U����|@��<.q^2(�,��$у �9���Nb�}2x�{�
�o���3Z�r�:�"�,}�\Q�&Vm��"3Uĵ������_���Qbv(�W1W�j��y
C��)Kd0i8��;�'^��۞�s"���1L���4�	c�q$�ۄ��c+Z�<�_��._��	��QW����[���N�*��U�o��h�|��I�sl��y���.N؆��[���ӡ�[У<���#���;j�b��%;�#���>�P���x�pKk���O�����[A��Ks�Lo�oQ\��H�z{�I2^ͪuM]��I��ȗeW�<L�^l�[����)���#��S�Ԛ�����M4������$<��(��-�Q�c�^u$����>����Ӎ�e3z�NO�S|�
�����d����*E�2�ժL�C%俤��6 � :n�Z��j,r�� >�Ս�W�)���6Y����;#��>����(�X��U�+�ñ���'&z,ޱC��kf�Z"Zֈ�Rʽ������5�;T�v@��P.������2��ǺD�����.��piy{g�*�(]�Ju`lqM(SԢ�n�Fo�+�$����D��L�?��lWGSڧrG�"KW'mM�N~u��(��(^u�r���hb}E��?�, ����������c�<~�o��o�^�{��|�0o��K��oWv��Ҙ�ic�u����V�Οy�?v�����乺湹���繊�����Q��苸�~��oPgp�Ǐ�rr�?���Z���Y]�+7�3��o�d:`�<Nf���pUb��S+�͠W7����F" ��~&r��&%e	���a��*m]�����e���}J) %�D�9�̀����@^���0dXd�`�}Sk��z�
kGG�Ef{̛�)T�O������E�ݿ_m��A���:���!{����Ss��19y��tGk��h��ˀ��wh�i�ke�fW�Ju�/�����
�����÷�$���v/�����)ޅor=?�g�O}�3ް�ܱO�)��;"r�������E��
7"�����GI#7��Vf=�U�9�iP�J~O�����G؇��0�X�孤#JPw����
��k��X�Y��@X�Ѽ�	�{�I`�me)������1���(@ m M���y�Ο�1�=����*�(�Y�C�&���!����N������;�I(6K݄L�A���H��m�~����N@ԟWQ�m+��н��h����TŞ픣�v��<.|8�Ptv��A��jG�=��=�����ɞ~fQ	��hK��3 8��: �
#�������;8�I�BI�_,3;*��ĵА�H\0���~O�B5����%�������(I�F��.n�q�$v�	>�������e��^�B�|%����l��[��kEwx�O`��Y~M��DRv)���6�	N�Ǜ������$x�@�@��f��[�y�*�*MGl�'^�Zz�r���*�����18Gi���{G�E�P:��D�T��ʄԽ��rb�-�Ң
"7m�'Rw��ޚǌF�˖���p�����Gw��.�*��X�S}Հ:�����e����^�J4O1M�)�p1>ɋ�Mlo,	w�"� P��*>~ދ]���5f%��L�y�|�A�t)p<b�#�.���F�y�6`7��=�����/�:	8������;��jk��׈r�w�)�t_0�K5�H���4������}mHQtSRUgtDMSMMMYƅ)��P�y;�ؤu�Cs�F���~ʬ
�C.��N��E���$�đShS�|�|6���t	0ՁO�"+FXa�(�َ�?ÃZ����O�w�G1�w^��������Y��<i���b���w˿�F
!�?�������bf��׃�xdE��܏0}�}=#ӣ?G��.LM����_�[�ON�{�>><8���������}���`��ԛoH���\�'�V���1ͽ�T��gVG@ YSr���Ʀ�~9>�	Qe�E�?E�"�P��-�ۙ����Ұ3�3�f�Rs����ԧC�Us:M[vz���̪5m����IS�RfkVP�@]ߜY^(ޜ��\ו+\}^-/x�;!a|�ԓ�v�8�S�9Y.'��l2���s1��h��U<GJ��t@��X��o9�������\�l:�Y���$��z���~M��v&�W���� ��F�h���=�q��h��ƴ,2�6�ݧ��"�g����ƽD�AW�2��y�i*X��=�����2)�OHiQ�ZdM�����QWOSG�\ �94�
�\�{�����Wh�TC�Ͻ\�t�`	Zo�E]r���^�7���|�~m��m���t�(w��@dD�"/�1j��9�3���>.�e\ؓF���wȓ�|��1۠!X�؏R_l*<��!ןَN��	��U�q���j�Ji3�i������y�X7�	n���s�*� bg:��Z�2�=�ך���i#��['f�'�V0}�~�jP�os�щ����u!A����CSF��=/�# �8_�ѬiM�>�%������S�,�S����	��h�ʲ5,�D�:��/Y�E�<q��px�=t�-�Cx{����*�䞎֓'����ob�YDJ��iyy��B�=(&�d�ݒ��j!ape��"�����0arJ�r�N���l~�;=5�p����wz0�:U|��X����'�+qm�c9c�hª��q���N����[���/���;rE��V�I��������D��>�e5�/q%�J�PC��5=턆%��0���ZƣPg�ts�z�*>�W���@7*$��2T�M��g/ɧ��+Q�3L�(u��A�?wB|����,�T��'��}���%��Lt���3�ߓs;�<[���q�X.?[�e/ܟ2KԢ��=��viiҋs5RR�;����zt��Q{��Vw���x�ݧ�^���?9������s�k���xq�������������#�ӭ]�빖Wg]���C�rq��	�u�F�u^�t��\�������N}YY����Z1qTdT�ǯ��^�~������-������X*�]
/
JО>^�^^�,z��w���>R]Q��S��=��%u��dԡhk	e	LC�3z�
Qj	��Z�ֹpAr��1S&^��t�ʱ�V_��䔋�a��!H��a�ٓ���<��ɴ�7��u�Oc��~w�V�î��4��}���\�qȐVǛ�K��֚;;8H�3=�$���5�]!y�}�����6��� ��km�5��������tDs�->����ԃ��O�����@80&y�6r ���OTN�V����]1��	�cl#	"j�d���ҬUP���M��.����>\p���q�~zG�2��B�@˺��n�{E�88���F���8�\07�W0n��'D�j�j�du��tyV��Ֆ��� 
ei�9�/���G:�^"�3:�T7�N'~c�Qm�yJ��5c]�Y�O;[�"��V%��@�k=LF�S�]�$�=�4�<�,}@��
�m��Hч���<��"�b��XҦ������!Q-�Ls�aB+�'ʙ�V5��_��X����s��:T�bsjb��w
���cjH ��,X�`g"�z�Õ8nER��QbM�ҥ��d�O�S@`�6�k�v���
,��Kɡ�$���\=�Du��iȁ$��%K����N��t�D!O�S'���+Q5
��0�s��)�������l`0%C�p6ѡ���/:�z}:0@9z:�+t��`
�͹J$.�e'pJ��#J��J��=��l�#���<�P�H�`í>{�i������/�h}ln\Oo7���(t�+��(�|q:G�?g���B ��Ŧd�J�<�cㅋ�����/-D���]*�(�N��'��'I�@��#��.�w���Z��rb�Jk�������TԌm���������wsXc?�ʐ(���̦�:�O>��D�N�]����'����u������/c?hcj?�U񲧵�l������7��;OV��5ܻ.N�
>��W�v�q��q��ΏNiQox��_v�e}kyk�jQ��A����f����1ԩȲ��ę,`y����Q��YCÑ�T�1���7<�Jlp�W,������bF��d�X)��yS>jݶ=��>�}��v�>d�ie�����n��3ܡšfkL������h�s��?�a_��S�R2�rc�@�[��b�\o.��� ������X4M5��a�@�}�c��k�q;�ś���
:j� �J�y<N:}t�������L���s͹`��=���?Ť\�� !!
�m�r�; �
ɣ�W��+1���_�gŌ53�'&}+��O5��[d�:���9�� W�Qz��OCe Ĵ8.���)���`�/2Lr&�Rj���lH��p����Wξ����j��fc�ҋ�G�9H��藯��u��zG��՝-�|ea=�5w_�,�-e�bܖ���C��z/�d���@l���ZS����r(���mՙS� �SvI�S�	D��!������s���ӎ�v,�����A���܆��.ִ�S�����* qx>]��iQ�2MĶp#3�P�Ki�;D=؈?�d�@a}$À�Vl����c��R��&eDGA�ln�����������
��^��0Վs�jg�:z�r�R�	�_�V��'۔N��f��:�*�����q�R%n>^��\Z��Q���&��Y��=,�t���g
�}HT���GJ�R�X�IN�~������������4�/�'��А'İ�m�H�}�c�؇<�EX���7&PL�����#wϟI/M��j4�Pj�5$�P$m���P��b��x��`g�O�����h2���
��$F
RJ�FI�ʨ)%-9@:��S@`��`�%�!�����w<��~x�l_�������uι��C��	��~�����EH��3�����A鮹��h���.y9�����t�6wVQOU����x䴔=�l%K���q\V����w�>��^x���[|^{rl71����ꮒ��tT�F�J$�p3��f;�ʸ`>����HEJf3��J�uoJ]��t-��~�]�����ɨ��:�m������m���q��V����%S�Ө��Ug�۽T��-뻃��9�ݰ��-������wZɿ_+���͗r��^����{w�{y9'�'*߯$��T�]�,<J:����C��FD��0=f��cD(����jX�E?�D����<�Qe3ͯ��e�cSS3-�h���G��L�=I����
4V��8�t�>�3}�����$@��t@�WI|L��i��,�QZ�1Nɻ֟Zg��\WEcHu��	��k�kkEj&�g&�kĴd<sk�G 4X��bP���
.Y��hN��f@v���/��4���>�ן���M�HP4lK��ڐ�ĸ������9�hG脮l �:�2��`0i�<%I	�zH�O���O)qގ/ ���W��
+K������u�r�7A����=�o��M�i�'�J
�T���i=�oٿ�!kf�/L$Vc�f{D������n����T�FJ�!}���Sta���.�zN��.��& k�@ji�5&�qx�x�]L"�b�(e�݀�>��8�S���b0��8�u�?�T��qN�E��uՊߢҡ�3�d�-U��q�/�>�����`ק���XW�a��#���1�Wv
~��?L80�Ռ*������a�_հ��V�!N�v�2M8<Lf/���æ#�nTA�j�SS�Li<�k�i�_�ap�|�i�chkjΎګl�@�xQL�}Ϸ��O,�����~��]a϶!�Jy�ӂ3����EC8�ǡSh��{f�~��D���|J!����R
�Q9�)ͦa���r�'��3ˏ�w�dNK3�"V��uB&&�˥-9fMD�c�sb�~p��䎽uB#���-`fK����npn������ƐUF�evY�Sn���}���A��A����hp[�m��[���֣?�Z}��C�3�Ǌ��Y�{�f*W�2D ���j�uS�w���^�T��o�ov����ѨP��z�T����_��<���y&v�X8�x�:����i}�N�������ᚹk���kt�(�[��^r���j�d~�:3 �������a������4��R����L9:��*�P?Ȓ���,q镉4�7Ƚ�cY�bU�"��
1iJ)D#K�8W^^|[��X��JD�a�("6�0�O$��V`3�Z��{��@�=:�1�k����n�7��L�?�|;��Ӭ������OM��ܮ�MYD��,�_o=z�cYD������8��T���ON��\���5�=�3sF(��k�ĠZ-i7��K-�g`�Ic�x�7����P�6�n�󠝳J6 ���.U��M��kB��LbP/"0�vK.��TZ_W��S0�r��ٮ�r�]�4�~�Z�1�ə��53{ʖP[��!RR�FV��oA3�r�(��j/�d������M���!G�/ќ�dLZm�4f�8;���,�G�J�iHjF���=n��uh��m�ƥ=#�xD"p�d����=�؟�|<�~>��Q`��`����m�/��)ݲ�q�Uj�X	L��N�o?��Ѕ�ٚa�d�Rk�I��;
���%�o�HBo�*���ZO�,��PaKY�C�+Ƨ}؄�Iހ�a���{*���MR �B���7sN�u�(.�5�SG���[��A8i��L���Ȗs���m@��ٿ�����[&�^��O�&I�+*���Ꙃ����d��}����f-�!�� ���3��,p�1��l(�e�6Q�gr{��}�l�lH����n����ϗ�Uz$�l�"���s����D:�P�����$�0�3��� 9$����3E@
�s�@���2٩|aJI�LE�!��åYݕ!�\MF����`U
� �x��Т�=I����*��	�#+��B��9@��`Mr�wO����$Z���@�p^z3i�@��cc����怚�뷒��X:�%�/��#.|����Y�?�����7�z�aV牻��;��-#��,Ʒ�L+�L�
��폑-���E����O���4��s��9o�l?��ۯ�<��n��+����k�ڟ����9,�_Mm�9��߶��>��;���\��:H���lлY
���Hл����󸬡"���o�+�	��O_]$v��o,�~4�A�Ԗ]Ѷ`�E���g�|�8�K��k/Y�lSV����&"�\V�bkV�pK����O��Ә��ĩ>F<c(z�0��V�^�9����K�Nx���Z��c����Ž/t�9�V��w��a�1�G{G�['g�Lgkg~/k.gSru9~S1����������F��R;4��d��������x��^��2�cE:��
Goo��ojf�Y����Դ����29�`_�*�����?�1N?�1.'p�h�^�@ߩV�l�e����)�o��	"�I(_�r�bt;|-\���O�]J�|��H�A#���'�������68b{K�4�*�#3-/���|�S��L�PM����]�pA菝ЬxBQiօ�;f��k#�t���"�]ף�8�R��]�Jʫ�֌X��=������E�X��UV4�Vx��-��l�f�����Y�_�ٵ�"�L���� ���V�wz���-E���W֫�P�c}���܃ԡ?��4	�EڍZdY>���ee� >I4Y�����1�HՀv�k�������<h���%s!*4�"k���鲢���ݲOh-�����* �1N�c���迗(ɥw����Uz;�L{��rߊ��|��V��[b&�s�>,�k9�����G�����qg仑*
�j����~�C�
�������
4<n�X���C��w�5���Bnڥ��
]�x�YU#����=��8����7Dħ@EK�2�P�P S�?j!���I�q�W�������[�Ǆ�ϚůtB�0�a'���M87�/=١�u����0�*�l�)��������]6��C�$��1T�֟��7?�e�	��(�QDCjD]rXZ�[z�����K�����꧋���M�P�?���矆~E֖��MR�u��q��6�N��n���Z�����~M]��<��n�!�n`��P��};��*��.Ho�~���:M��:������n������~Z�vM]��nmu��_�r�Ρ(�в�,�wbpAY�-%�����<ɪ��?��2�N�
�~ c@��W��{�-�3�?2�ȗc�u
)Ȍ6Ƭ���l2�v��WOJ9��j��f煦�A��n�L��������F���6���6���T�4�@Iq����î�����T\#���Z�6L.0p(^�+%��n��=M��C����$^�ˣUt����k4;��h�W>4���i�p>��`nY�G�P}W� ��0��G�,���+���򴡔��Y���u�x�_��� ���ӄJs7P����@[ߠRgĕ�����0���[bK<��E$�6<�UZS�;�W46���I�����=P�OPQ�N�k&��:��άek&�ɳ� ����ൢ��\U+��R�Fٔ��'���X�������R[~i��%����"4ǩ��H6c0�34��/�=�����Ix�*K�p�6Z���8QLv�-��-(���BR0Cץ S�x���S�zq�D�V"[_�r?����C�����YL���[i��ʐ;30�ǖ�4�aE�⩢x)3�8��=��yX�8�u�
Q�t��=0��N�#�g2,�v��'�$d#/^n�v�ZtO�L��ݖ��;e��8���,��WK_Jv�Z�a��d�~n:!/��yԛ�`��_%�f�	���m��p;������1���F[�Z.��4�J�ч�S���>��}�%��ݒ�Ubߜ����=$���W�^qPA�k��C�K̞��$=v�a"�A�%[ʞ�Gv�! ��\C/��w�@��F�mL���HXzV.�
�?��l1���I�Y�1y�%��,p���B.����9���������V�O|�u3����vr�h��G��ʧ�Cx��_N�U���~���d�_� 薠�J�ة]�+p�Ԥ�S*�����K�P<y���#G�3\;g�3;��ám��c�mYyNM��>��U-�1v���9M=���z2��Ω��������������88
�C8�d"E|<0-�����2S����o����=�����C�Ƴ����s���!�������e������4��\���s�z��,��c릻k�y���\��Æ�ۣ���~�Ƌ������7U����|�j񩢮����y��Q�^h鉛88q<�4gێ]R��,�o�Kq)))y�g�~����*�V���!}&פ���?>�<9�#k���,{��̓���8�6hx,��u@��#}=��ɱڟ\��=.')��X��Y\��~���n��q��|\��f���3-��f�ѣߌ���W��/9��#��b�3������۶���i�g��>%��[�����f����E.|^{7ޏu`ff�=>2�H2�~�Ž�CO5\O2\O�������ݺ̃ L�>��J��	ݮ�P�Nˬ4W�ϲ�[f쟍�6�}�^���3�u7�-�\-@Yf�޷�Po�R�a�V*Nu�4FN�����yAs��֙�>�Q~�¸�%'0`�����B��Nfu�zj����f��*��B�g�_����b��)��TT�ľy�$%����4]']K�I���H14Ӛ{�<�U�����Y lF�5O����y�/
m@3hho>q��(D�_3���P����, ����<~w	���o '�>W�T��:t0�=<�=e���V��h�̬��Դ�伖j�ێ���U6�ɁvT��̆�#hkٚںg"Pf���\}�(�X/�>Gp]����8��
��8��.GQ����-hx2��$m,U���9a�==H	&Yh-��8e8[�`y>|Rl��p�J�2F0bMr�V�L� K|`w�(�x�@1��p(�}s0>�ib�+�K�%2�6h�<�zIK��Y�^�g��ض���Q� ������kp*Q#�~�$���,>����T*u"L��4AYE狯�</i��`3�48�c@ j	�lc�Y���y��vO��
%x1����iD�$l
�i�t�]��li���,B��������=�<`���pn��qq�e��Y(��7�z<[��j`�F��m��~u� Dz2����H�j�I]~_�z*�r���r�\r�$jJ���ʢ,b0d�i+����)@N�u����-
�12u��0r��x����w=P��	�jAzNz���l�o�:EP�/��߬�-������.]����)ok?�Z���I ��["P�k\_,���i%�����ߩb�L���������$ڇnw+s���g�u�6�u�'ϛ��<	�t����MͅJ��n�����s��MX^��\^�hA;��W�yȩЧ���b6��̵�J.S���k7� l&��T6S�R�%mqA����!��?�Zod���Op`"P���bh~�Z���31#T7uKoBe_H]�_m�r *��vg+o��cs�d��_�N49��=�3�����?0W_`9�RH;ډ�e�xn��Tˎ����9�|�<��������aş�
'���o��#ޏg`ȡ
�o����FiE��	����
�`���x��Kv�@A�c�c0>��l7�Z���SpV"0R8i�s� �4����u�g��gr�	D
�Ob�ۡ��1���H�˞6+�Ǖ�1b,a[�(�t�o];�s
�ֻ�u5�
�PM���ީ����to��W_����A���H�ǅ�u,���)�Hʢ�Mve�CXQ�5tc®Ѓ7�^j��Fi������i㫿�Obf�C�^8�me4�v?7��0S L�Q@�5Q�A� _����y�M�d�u�� �<)�K׋j!��wv�?~��R �2tHy5~�c��7���u�e�{~��H���9	�8rj�L�a	yMf�waD��򢦀
�CW�ߋ%Bd�[0iwMJ&�T>�(���p�+3
4�ܡ�#�5��N�UI�Q:�'�'��_9���+����F�|�ۯq/ie�A�R���xE�E��F.R}(�o��fkQqo]�	�PF)���[.��5�G()H�Q��=W��ΪB ��ͼ�/��e�PD�
�\^C]��M<���Z�g.�}4�f@SI=��u�1�s���!S�,�.�NC���kwVa��x�C(����q�?���F�o&E�4�OH�3�N�}&'1�O�hCߊ�@��3��m��7:0�48 �%����!)�eh��o�����p��MӋ{��|����ag=�M9k���4�k��������[�yѫ���[~���w^���b���6�Y�{��Uxt��oW��{��sy�u���6z�ά�����������.#<�;��8tT������X��	黯�g��= ���@>e"�1������j����c��?am1� �4�)�PI������K{�x�N%�7{�����=9�w����p^��|���/�q���ݎ�N�@���|$�5j�n�4�;+#!�|l5U�&�"�RI�_&+j\(�D1���A���M�X h�ܭ�@�%���sh?{(E�,�o)� �_t&eƽtp"�f������&��Tef�ts"�}9T]�E ۔����Z�~׿p`�pٷ�hp�9QA,o��6%f�Czy]�2�%@��*��B�燅I���#�W8<�(�������a�=tp�E��c���k�!y,aXS@��P�1�cM?8|Z�:����7'����ik�<�oLEΖ5S?��K�2�G�h䰳�qI��Ô�X�h�eRf���.Ho��<����ݑCe�_�XjlQ!�Hjf���l���T�M	��|;V��:,#�x+����5�20v�����9��M ӓS����ğ�����|�tL�`Vښad�32����h٨�Kgu�5h� $�iBRr�6�	�)9q���xk�`p�C�m+]0�ٰ�3X[��^Jl�N�%٬���U��ϴ�̓�ٶ .���'G!�	��$5�� �jb��P��%H�}E�1e����I+j�,��IV�?Z�%^'=�,︡bD��>{r;L�d\�k�K1`m��Ab3��nf���Q�"�J:IA%��Y*C_�~@��ʘ�'HD�0�7��h6��hM���È\Ǌ�v&V&�����f�rȧ[b���ր6�{��������#LFo1V��+'����*�?E0��Xr�̤����xhK�ՓdJ�g��0ɖ!ٺ�]��1^G�M�x}q���4��x���W�Tz��	���7�<`�۽����k9���(�����7�wA��Ქ|M���k�������J��y�,�~���׶��}Y��}�d�f�f�5��;߫�ӂ�����t4��W�o�U�Y�oH�౟�0YW@2%�2��~������k^iy�oAie)7�f���r9*u��G�:�������mlףc�p;a�˖E~O�;x�땛�����WQ].���y9��,�E�����~S�?y�'�<W`>b���cu�"v<��#=e��)yMz���/�V���������L�"M��, 4H�%;F
��vo�0��X�tqF�������6f/'�L 8���
��*��suC���s�dk�f��GF�~/` ���D����%�!s�F�T�Xa�����<��Z�g@8��3��%L�s����R|ԍ����(r�&�c������Gfߖ�JeP<�X3��pK4fL���C�F޵BcY����X����b�Ƒ%�E�F¿���	*��G;,�Ó}�8��Qڻn�V�����9������2c3�P�r�ξ"���U���}��@��QTzD|����$��P��7|�����Bn������"�b�Ȍ|�,��A��?] f$��FC_a%�R�ٱ�Ɵ��SU�H},8��p��z���ɕS	�g�.�NW���F`9���q0^ez7m/м����nSF��J<!}`�� �����T|�4�A�����k���[n}y�::�\�V1{�(#�X�]�:�3����d��z�����l��>����3�aO�7=g|���8�g����|%�@�
�Ih��bj?��ߜ�7piH�*�
��2��3y�&�6� �:M`�EH����9dD�9�ev-*�2�� �V�I�Q�`'�������N/N��.~IC���]����s��m/����GE��xg!��?I ����N���Ϊ
�
���h�Fa������%�z�����K���봴K��t?K_xHN�VG��6�(���A���U=�J��Ϭ�m�
����S����7�M��v�y^���I"Sk��<���ϛ���J.���6��j��z���f�<֯�����֋gj�ݶ���ե.K[����uk�/è��cHi��<�n�\u�:Pm�����������3j�WmH��V3�� |���a�斻�CRV��޸a[p�kV�u����E�uR0�g��88m�,]$4�D��ax�8�Y��{YOǇa�i7z�v��q��9�D�� A�����
�v��M���%��w�C�ܗ�m@'���[��u�.|R+�XF=�@���D����S���4�j�\���&κ
ޤ�%Qſ�@��&(K��!�b��JA��H[�lx&����G��D�R�jW:�灈ER\ږ�Or\�|��d�R��G�0�H:�Q'd��8,����D�M�ц$���Զ��ՠ���ޔ;s��-z�	&� 9<���L0u�dT��֌�3��~��=z������\{��@d+���aK�Ծ�~>�LD}����f2���̮�M�����mU�y�C��N��+��6�`�A)�D��Ƞ��Z@yO�_���/��8�ve�~@"X���_p���pd�b4����^~HWDۢ��ɘ������Ó�6�he�(�/l6^e/GJ�ժ>S�x�x��з��$/���nب��;��qMo
U����K����$����I� �)�VI�O �k��w�]��Ln!)��&8ʎ*�U����n{��
�vu`+H�H�1,�MKP+q�^/��g��"���sCd(���tC�WŇlh�`�Zz�K���o�B�2�ocQ��!0�%�1lu,f0K�_e(�þA�������$a���I��%�On��#��g�.�x��r=�^���9��-��#�c1�-��b6~;%�e�T�E�$���[:�B��<����d� |��M��E����m��t�b���#��W߱���K7�� ךR�C�}��BD2	�#����X�h���Z8M2��*�(6@�u@4�]=�^c�g�Ĵ��O1l�W����Ϟa�}��w�U97�\:ߏG�=/��置�v3�k��b�	����4���F��oX�ן�9{]�r5�M����D|���<O��{�[Q�������,_�2�1�� d����0<B�D����&#n�m1���ł*�+�R�=��X2���?~`���}�)�B ��ɹ���n��)?�f��}`�alN����Ӣ���s�\���k�mD�\��jDrV�8����P'�H���}Shtp�2!�x>9$Y��>�����lS��"CW'�����b^w�9�4��ߧy/��r����
��J�pd6�?0G��(Cmj:�$	��)}�f������U�dU���2n�zaumԧ�(;�Y��`�s=D;m���;f�>,K|DyY��?~�M%>Y���O��=�=�����L&�ڙ7�v!��-�?���V B1�L1�'A5Ȭ��$�çZyNelO���������Bz�����/g���4�t��ُ��ZK[��i	��ŏ-��-hz�Z���f�E.��3�<>h�*��O��Hi�O��09��64��5������C�j��|:M���H�,	F��:0���pv۽]:�&�ɨH��c�1�ʐ�r�?��S�!_��̊E��ʵ8Q��p�2(Pa@�M����C�>F8���'��:8��]��O��m���,o^�#4B[���p	A!tH�@GV�q���u�q"��@�L$�	���b��h#�G���-��; ^��'>b��A�C�='CJ���)�T���*Mu�.�!o�tQ����(U��7�ސ^��z�����ll�s�%��J�T��bKs�:�ܥ���Kl�FF  WX�"ZI�����ƣ h�҄����C��4:pܴS�������|0�Ԟ���@4�������k̃Bm$<�|��]̦� ��8gҳ]p.@P���<�z�ñ"��llm魞Xekq��tI�U�~}ϻ]���\<a2Z�P���v��LM�������Øi�mX��c��������߯A^)��r��
�K�N=�i��yds`��e����f���z,���V��x����{{.z����?_w�\�B��O��f���p�eu�X����H�i�q�PI��q��0��j�W�ܡ���C``2�L�����N��E#ګ�i���O:�n_閼�'�-L�{e��pC#Z>0A$_+�cnx�=�!�\�$�.�ʻxڧaZ����;ͣ��E���E�����h�P�:��?�6Wmw�6j���P5�_���Q�HejoǾ��LbI�_��<�8H�u3�7����%F�?�c���SS��|k����w��i,_���W��Iͮ�-`8�JYq�yFAF���������P^�/��V�B��m�^�j�H}�k�`��Y��k�g���V�cQ�O*>2�gFpr�YF�P.}j�S �Q�������ɲ��4A3	�nr��#�_��9ut|4X�S�L�7&Z�;m)�t��6��ޱ�P/:ZP�e�`pD�j�L�������}�:Jɞ��8���@��UC">1�>,j����R�؇��Ni��f��i�tR�����9k)ǎ�W��=nz �����Y�a��.�������X��}�XE�j(<8�)@<��#m8/�x#2K����L~�O��e �b�ND>��~�����Ce-\��jM}FE���)�T��<~���h��/��\$S���D�j�7�/%*ҿĝ���~���<6X4&%ч�h^[7�0%���)$��+��s��
<z�x�E�Z��V�Z�Nŗ"�q��J�U�7P��C���8ӆ_K�ͩ�rR��h�o1u��}X�ae��H��e���R7�ez���l6JvRy�6ݐ#�F)0��З$tJ���c�<☕���"a�t��YxV��%(��U�k��&b!꩗��|��S�8��<�8x�0h�S\��1s�~'��~�\�������O�/�q�e&E&=��o�ڲ��x��N�z%I	gK�<c��gXW�Lڊ�e�Yb�����98RR-oof|}�%�4H�	e�P}�22.�ۆ���47W���Q����쫕��a���������^G\�k����t��ֳ�U���9u��5����崘�mݼ�像�	/"p�n�u?[ثo�;v^7u�º�n���)���e��|���� L2q��hUm���LLN��H$�P��pp��[p�Z��ZR�X���u�Y�a���9�1�'h&����WD✉|֚P��u>;W�^���3����#����0���MC�:�\����࠾������l���p�����lz�?����@���$ٛ�ÅV5�ʡ!�hϓ�GÞ��Qfv��_�Q�c��`e�Ξ�nE��D�9&&�W9ڥ[����Í�^�򁗎@'�^X��0L"��EeCK�3��$��{n ��J8�}��Q!��80�W���8�.��ݢ����</�N���_=�~�����EG6�.���@�03]��yo �W���t��tE3��� �=���o~�bM$����S��uN�%�m�4��GȮ�� X�k�F��Ns�+�u�g�����֌[����f�q��'��K���	p{N>c=�^ ���@i�|�n�k�<Ke5%d�_��m��!�Z�rc��l�>5�u�Qa��@�["���8����(�?����R��'4�Sq8���)Jj��kn��(J�3R��}�\��s�gF���kR�V2���B�o=K���1�}778�-�aR��ˊl��~�o�;T�|ʊ�1R*���ފ%�D"�J)�A�pYL�39�ԟ^�	��IMzr��>Q_��Rt!�Y���6�)�$=�0�!֨�B|D|��� ��۟�絁+⳹�	Ii<w
�v`ܵ�6ZQ�9|Mԝ"F�,X:�F�=� ,�%�xIs�-:����uyp���� �0H�Y���p|��bg���"���=��������IA�qhC�"}�GQ�X���v����͔:��������	v�EE.����~2㑽�����x��Wf�V�:�����s��΃	% S;�'��'m%��XV�,�
�f��,����Ms�S��������5t��w	59}8⹋�%�P+٧A�	�[�էHx�����<�[<%2~�;Z'"#�H�%�h+�q=�l�����9�-�N��w��5�B<er���T5�;t���'��Ƴ��=��:�䒶�@��v"M���>�{��ɟ����Y�]��}��e�U��Eҕ���;�[+�;��r��ox�UF
4K -F���%�����}�rTV��T�;�;���22Hyd��?o�K��X*Qw��)U@ۭ��"c��E�g��&���i�����۫���V���֦��D8�|C����\p�JA�T��،�>:�����s9��#�tХ�ٲB���7�^�������^�h��2M��"����ll��/�oC��PB�~sa�7�4��v>\+�_� X\��(�8Л8Z0��aO)� ��(���*O7w����,������}J@������y�c���Ŗgm�nFэ����%����֛��/"����x�b��xS���%T]^Ӹ�w���g�O^W���`�|���5WvX�<��x5��8W���vX|7�l�r���Z��u��Ԥ�Fo���X� g�Xڜ�b*��$r@���դnLp�%B��Y��G2�:W�NZċ��i--�d�t\�\��t9� �,��쪙풜�_%J<�x/���X���U)�O��/������߉G�qv%�;�ăƒ[_����I����З�Cŭ�d���;&��3��uJ��wB|]��3G~a�}�Wr���M\ӬW�TI��V�FƦM $cטCy|��f���\�H�W�%Nb����,5���!�
�΀���,���X�g`���W^RY�mZj37������� �p3S��{Xu�	�_S��fGB�nQ�"
Sc�/2�,�+�wZ���j��%��J���������5�Nݯw-��+�IC�H�VS�CU�7�i�d5<�8��� ��
����'���K��@�_�cB�:��)�Ҷ�Sǵ��Q2]��x����
ˋE�����a��[�P,}������40̌Izj�*]�`��'s��l��:����#�߈�^��?�*�l(�G Ͳg݊k���=3���j03[���F-,g:S<�(�dlca�T��b��$��P�\ø2_�3/��}��uH�'�3��� l��Q��ࡘ]�%*���11T1j�`�y�Ԕv���*���xB�B_�J^��.j))ss�%S��,��Z�݅Xt�d.x��"��K{��.{���6�<c����B�nؑt�p�����5�"�io�`�T�$�j�ɘ��G�<�
�s�&b�p�)��q�̻�.��
�1zQ14g[�';g{o_�I$���i^ ߂��]�>��ܜ�7��U%���ٍ�b����~n��1sX�U����J7�ʚY/�E)�Q8e�<��w���`�e��2�>Ao���c�ǟ����a�V�����J�ɭ�=�r�����4jy���<L�Ӯ�9^+�(����nS��Дf�lm������s��X����f�e1EЩ��`��p����Ti���vԭ����>��� Ao�����jv<�<��n�u7G��}?�K; )8��4�+s����u�����)j%��]~<H�#	^
���"d�@�P�	@>妱 ����Nΰ)c�F��]���v�!\��I�<���R��ٹ@�|\����)�l"ڃjzߏU�/�:��:������8]ȩ���/��S��"��۲��0^�
��-O��Yuϐ��.n��[Z�X�շ���V�4�P��J�[�D�0+%]��+�Z��<&��`�2ӂ�lK�1/��瞚�d�1i���R8�^y���ϗ�B� �� ���_�I+��MCc�a�y7�[J��@�s��P���%�"�_�Q�H��dr���n�|8��pd:��67E��u3 ��Ax�<�����+���"�V���&���^*�G�Ċ$U!)J���3������1�lE�I��_�)��]�Vܧ4+�w�����Ä�t��=ʿ��ݞ��S�Pe�CJ|L?�Z�mƕO*1%�ŝ�34�o��FN;!�|��F��'���gV��`���otXip�P鐕�Kưx����`5�l�B	$Ne�� ( �{�C���hj���	0 �(?u�������[��³N�͝�,/�UV?�ɔ�9
��f����V>��UU���d�ǷħA(�(fQ��}eX!Տ������K?�P�ȍ(oO*Om^M��t��{���w����(-T
��$k�����w:�a���z��J��%�B�`YV ����	��	���1$��M�(g'�2�	-�H�I&OٚY�|�X�Ck�,����R��7�?���Ohs�&�\(]��th����q��|�=���lD��c�:r�c7؎�8Θ�|h�>ʲ�ሔ��*���fޘ����Ð9,/�DD�.Y��G?��/�Q,�`0<�O�eͪq���D(����i�k_�^Jŵ˴�SH���[�[���=��r�T%�Lg�
7X�Ko��4h^U����*��������R^1¤�V���)�	�l���9���L�TY��l����	p��xI�1�/ѭ֧A^������h�7	��"]���������q�#�h<�{7C���7s�A,M��A=]���"����'�?�����X����^_c^~/GPT!K��K�bg:�ܷ }�P��<dFB���4�宐�*
�[��_���w�Jt"h=��<Woշ^��'RU|&�||��9�W���R*�s1@�j�֮qyl�.�o�s��*#�.�ҕսݝ�o�e�[2a�=7���1T/���nG�d9W/�Jd�����R �`�0Uwe�,80�q�,�1�4kUR�R�Gv�2��1���F�6�Z�`+
R�%,>g�Z����iF���'���͖yz����5��C$xy �.+��|t/YV��e�~�m��Z�!��\|l��K��^F���˦@CN�*�$;�ߘ<bmGBfE�ь�H��άc����a�C��/~����<5��:j%.~��m�nPE5)�S��j�������ݚњ�o>�W"Ί�oF
�в��
��|S�F���QcsjA`$[��'���(�_���b/c�z���p�y��>=�@F�l�}H�Gw>�!��Z�q`� �'����u	������6�a��]�ثW���(��!7鋍�a�//���<���[8*�,�K{ʘ.� H���,J��	nj�I	f��w"S���~"t�<q���y�+���Mȴ�'�C	w���~;��{���n�� \�y��b{'D,&�-ʇ�#��g�W�����C��=q��jt@ln�Y��=����*�M2e���͹U)����?�`ކ��!�d}ޖ:�g�4`
����+1��e뱢&��EY�V@���T*�TҦɿT�x�F_!�H�1ԁdyb�q�;N�-
�@��I�0��������Z���8E�P��T�2�y������;Ռ���vOϯ�/�� ���1`���E3Ġ��8��`7�ݣ�\ZQ�+z%������I�y3gǃj�0d���]���jZP�m�� �[���b�ʗp ��(ߘ�b$�/���ǿl�^n?gT�e �zR��fݭ�?K��kz���?d�uX��6�t8Zbt(��l�t���
���(	AB�K�!�ѝҡt�)��x���<����׎c��}��:�󾯘<x�<�}� � �yog�f���]!��p�~��u�8��::e��n�g�����f�j�gb"@�#��I�aP����f����8:����B��KQ�q.pezQY�h����v!��a�?6ϼ�x��bk/��Rzd�6�c<Z��ѵ�L����gv�g��z�JF��ז����r���Qj��?�g���ߔ�U{�|�!����AE=.#�ֆ���:�"e�<a�p��F��WlP��h��z��)��P��f��mL�L�6�a��L%��C���Ô�Yz�y��`�o�ac�����n��L0��B!]��ߌ&΍��#�)�B9ѹ��%��t!�����j`����wΠ���AQ����HP�y������z��VQ��Ϫ�Ї���7��G;�Xrw;)��E��0C��(��`�G��8mKā��L��X��d��}Π"���7$���Տ�q��Ue���0�Q��7��T3rc@���(���D��`:8~ֱ9�U��!�{4���oKF�HX�x��~4a������YT��>����
��%F�mCb>�p	��<h.V�aZ��iG^�g\%�?To��g�,(�C"˻"����+�k����jP�d-�!:<�R�-�~-�V�E�Q������ٸ����<�H=��:������,�����>p���e��LKhF���Pt)e�9o��׽������c���+���`��Z��})��|E�XH�3�_[������x�Ջ��k��v����v)J��I������mv�Hm
J���=�	$o_�G	�V����&d�����ɕ������A
/Z�������TQl�<G����P�ݣ��\���+[�������
ǰSW򣏤'�H>��:���8�܍���"�O������,O�?������]���H�y��՗)�����U���U��)'+���T�2
����BNt㹲��U^�=3�ޤ�6s�O{}̶ַ��hYzP�8$�ACB�-	�Ȇ�����s���6$��z�|����<�(.�%�]�[�y���"7�_#��3?>�^
3�6]�f��x���m��$9��6ok`�hB�x<���R0� ��#n�����c�U�i�?�"���V]}X6͆M�`l�e_�->1�C�oZ�/Yiq_�6��K |y<�e��]���`b�2xl��`4��R�Ⱥ<ݔ[��Cɛ�,C63��C���H�m�B\H�
-��/�.����n������C�H.��b���q/u*�2�ϓ�����Q���$y����gй��M��;`�4�`��7��%�gHÅf�c���b�{yTY~�03����M/���L
�����BW{�sb��|�دj�X[�n9��;���E̔�6=ท�p����k�?�6������`��ym��#HK�s�;:����[�3;�f%y	�	��`���#*
_S�2�u��Z���:,�+�i{k���C��)zG�rC��)�=c�Ig�Ѭ,��)�%˭k]z�2��V�P����e���Dd�藎,�@�cn��:Ll�d�ET�E�f�JX�I��.�ȕB�(�dfAq���ik�I*$4Ǆ�K8���cF�2bݧ�Z1�)鄮�ʘ����ؒ�9����O�K�n��KT��	�����O�i�6y�k�	�z��1G�A��DD
U3� �"���w��� �}��/�wZ����6��*��B!���^�y^ˮ�j���eF1梩, ���!1��qvX�iEd=��b�HbX�]^c^ܡ�\�^�!�.om��� �	�]�q��o��G�I\/��;:`RXeT��3��2�Ӷ�}B�ȗw�/6|w\>�`�Z,4�8����������VZ�5H:�����l�f1`�e��c��R��Ě����C��<F��a]��X]Ԫ�)$2%�%�^�C��͎�?�����02�(k� �DZ�'{�-�D����w&��^���k�Z��m� �7�FHx��G���ѹl}Wb�hy��;����l+,X�R����n(m0�(��&$�D��n���ɡ��2�k�
�;��F���v-�iG> �B�>�����d霫TnX�7gqP+џ5��EQ��g���i,�4�\(@ �����(Y���o 3n�w)�W ��_Om��u%<dSI�;�;�0h���p����c��^D���s/���X9��TR��Q��H�G"E��u���-��o������T�7�ԗ� 0,���:K�IZ��=�}�|ps���0��_��O��b����|�Ր-��b��������l�%>��z�,\��VLi�
�#B�8�(�P!fI�c˟zQ-����1�S3�_Wk������93L�<�j�-��7?�C
�Qgia�{���K1~&Z����ұ�eH��2�_���T�Ҧ�!�8�����S�j���{�N<3��M!D�	-:�J���_���|���eI@�τ������g�Y�)<������?SO����qL�{�QŜ�Ȓ31�?_9�;��\:`[��D[y����Kחg�B�x���:)Q,T��2���GR���������,��1���e&��u�Ne�8F���/����ͣmg[h_o�!��U���#PA]�qc�F��i[-8{�J;XbA��pb�5뀗e�/�$�t#?"�Q���!(Rw��5W�(�7�zG����ğ�HH�\�M~�����'��Ʊ��5�u�����%I!��]V��V�D�:Q�d��A�Rb}<^F�_���/6����<ˑ�Ao���1�x���T���}�y����wg�5�m�Q���YĹ�f��oƱ�
5x^'g�6�l�����](}h��?|7�;�q!�����IE�C�yb�o�Sw�� Xhy ���a�=��v088�p<2�!5�.�f� �q�z��p���f1T�s�	Bn謨��и�x�З�ԗ,i�ǇU��<��b5:̑u�I�h�=�靖�U��?�)�1��{�wi��^�?�f	�zt&T����f7x��`|>$�p#.��\k��u�`_��10��m;T�ț��A�A�j���Vp��~%�F�j�I�_p�o� ��:�����'�^���&1�qV�?�7�={��57>-�zZ�Ù[']S��]�=ȘV����Q,����2���u��P������Zu�h�E輹s5^(�=bU��!:r>Y�p���C(��L�%_����_�����`���7��O�k<U����$y�ޒQ��
;ֺ��7	�u�x���$.0�#&*k=��Nx��Ot����d	UJ&���Y���ejоJ0����U�9�ĝc�=������`�$�)d��_�1: �ғhB=���,W..�]4Jgm���Y���8Hi�M�Y[�-m=��tb:�ޚ��xL��<�Imc೙Uo��A�a}zCq�]	Z�?��[n@���́��F�:{ҙX1mHڎ��j��ސ~��Ǘ�lh���Y]tJ7�U�<-���Ť�U5�h��9d~/Iɠ���-���]!��H��1 �#b��Q�7F(߁��C9�*����ǅ����(�rU���<ND�m�S����p.y�Bt�ã�,��dV?:�JpK����k#N��?���fM�z�Z����ka<�U#��e��g��jB�HJM�i+p������2�Q�#'W��*M��˒	�F[E�ym��um�i;k:������r}�1���'Jz~m��L�_�tw26�N��+;-8�@IѢ�N�f�m�!���%�����D��]�P�j����y%z�5j�A�����\�^����4�M��	�&	3���������%���p}��2�����BEO�m��a��b%�|����vJK�/A�,;���g_��#���G,b��s����1V@�F%��Rsא�����. ��Z7��� ���wMD�&_��Ob���%c���۰�P8��D���R
K�(���T'I@R<�!��?m��:���(�D�e��HPV"��mg����o�"Yj�oM�oa7B��@�_�3l�@i�*���e���<4vHR���5�R���ȣ�j����˳{�-��h@̧�����2F���FV����
�O.Y��}�WGYֆ�z�C�V���!B�����8�ǐ���c�ޒ��0���%�kq���>u�fce��*Ү���cۆY��������x}���B�L�~��%� )^%�*�1FVFr�O��j�������� ���#�:�i��#�eX�\�d'o����l�/OaO�-�կE�S��z ^:�F��G] !��p=:�i�l��ג� �gAr�唀����Mp���fx<��?%Hc:}���:\֍���F3�(7(=�<�U��]��)ϋ}zn�@�BEV*�w�eY�>���	"53�F���)ط f1��,kV�P:-L�+�5��9������<K��@�!�\�*X��h0�:ɠ>?M���|�����5o�����[��1W�� >b.�t<�����.a2����w�C�dχ"�MR�J��AT颕���-��u��~��gJl'2���i�?��2Z%޺��"��>�A�������%u�q<aiM3�nH<��W��b�7N���r�C�X	��<��˷ܱN�
m���~���AoǱ�O�t^��ܵ۫����A���
)�����$m����S" Q��Y���k/��d5�(w�!�	�$m�y�a�u�;�h�a	\��_��#��w� ���,%U���#�G�t�P��	����KA9|O �����TY�ᶺ���ъ����"���]z6�8ʍf�gOE��F6:��7�d� ��"�*����\pۯ��>��vsbۉ�<N�[����5�z�${�ۙ�o>I�k��)�>����;���eXϛ�^�Ml�����fz�Z�gb^F����C�������y�}� ������Iy���{���ދU��?1e��7��j8��.�rgNVu�l�"�������P"p19
����m��7xԆ�:���e� ۑ��2̟Y�A)Yi#C�n߹�k���˷����La�~��A������T��/���(�ߤ��$�	�=~�=46�1;U��$}6��|kb�M}�n25jŏO���@b��B�a��)�3,�+Z�)��) �?i�_1�`�ՙ�q��v��N�1��1��	��D(��&!���pyv��D;T�6e�CrQL�7����{�X� �#��U�|J�R�v�H����/!��ޟS�_��wEZm�*E���j�<����F�����V�p�B|��q�����C����ì�l�|�@�Ov���*�;#/��'-�i�]�~"L{�vP�"�"�%Y��-�k]!��*�|rpwu���A̔��lպ{�p�a�Ɯk�/�_�7~<�}�j���^���R{"�Oj�L��Q�0o�ѿ�Q��뛩)7U������3g�J�d$S
QI͎/�n��֮��<h�]Iz�N�,+$��ez\p̂�V�iP�[�[��9����˒�'�/qOD��Rn�b�Xs:"�&��@���q$��Tk#��v�K��[�$���<P�t���ndN�)�Hs���kT�Tg�ς�W�O��_X+C�è7��z����D�=�M� H�[�y��=D���%�p3�[ܨ�u�"�=JV?EMY�)������Kg_��Uͽ	f>�$�j��L,^� ���2$pC߼WE�ϻ�Y��E7��{��������x|h\2�R�K�Li`p��(Tw��:o2�����M�1_S�}5�Re�J:��ً~��nZTT�<#��o�1�웚�\\R�􏠾��@b�$j�?���xP����*�,@�Ѣy%m�r"0�k������R-K����Y���c��c�aq���͌���Tr4��Ǽ�(B��*(�Trx��9���s���wd?�fR���Qn�(E����Y�c�`pO��;V�w��������E��G#sD#�h6+�R�
�ﺒR���,�_��5�?���g����4�r �6j���ލ��\��A/�V�Jb`}Ƹ]h��Kkt����~?��~���k��Q����/Vٕ���R+V@͵��6�^{ԗ�\��5.z]�/6�j�6�����B�R��P��׊Oj&������VJ\�o<���A_�.�O�V�����&B"e�������2�����N��G����A`��,FB� I�x����KIU/(��v[<����-j:�n��:������O�5�J�?����L)H�O�8�{��X(�����]I�'4�RPQ2'�w�8<��[�Bɯض"o��˹P]�SN 0	b����~R]�W�h+<c^:a�8]~64U�����Ɣ�B�گ��Ni��nIj"�}~���
�qhHd���#�guS{�}�8<�iXO;PAl���:�	'��K�&D�3�8zk�^W�4�#�N���m��j��&�{�����}��i*�98�����%Ӆ�����+Y��a
/�ށjB&n�vĥN�%���SN�� �dH�3��/Mv4p�s�ҏ?���
�T5�Qԡ0���������Ū�p�w&o�H�@�Yt��p��y�;t��L�5��(8�_AG�/J�ĕ4���9M�숯Y���R�&FG�W�ZK*��p�)!��M>������hP��W�F�A� �n��7�T� }[g0�
r��"��: ��?�w�3z#�.-�9�6{�r�T}��D���C��ac�AG`�����E�̈?�����X� ����`r�T�O��jU�*��C��O�W�j]�E�uTk~$���L��gJA�L�uMzh����}xey�y6~�Q�
Ҟ�?��d�w�;}T�U}ywy�zd�l/'l�G��Y /)��҃�"�F�0lƙ����;��C����,����a+8ܵn�c	���j��#��`W�fZ������쐩(�u��:���@�8����5Ӹ���^Y{���+��t��c�P	�q�ܜRɒ�����~��;�RL��I�$S]-V#����N�k|�]YE�������de�K���T`5����O��R��(����&�MJ�o�&�]�?'S?WY��{�j���͎֨K�1�Z��Ղ�녓�y��~�����DdLו�햔0��k��c��Ô^�"����69Ȉ
t�<옐y��e$���=�n���uwkl�n��ejr����a"6u,��2�f�a�ãLTWk��E���P�'l~ ��/{R�7�W+��\ąΆ���n�[���6?���\Dm�ק5|\��l
[�dD��*�(��%���]L���`�D�I�_>mYt	�r ")|M(]����Dԩk|vd|�G��
�3'�h���Ր��1=h���WcZ'����e�u.6L��-;mHj�V�oVt�4��7�1�oj[����#|8P�����G�"g�sE����j�o�.�*�1Y��P��3��aPw:�Yc�/%����'ܸ�'np�Ϫz�h�n*9OE��ߙO����,�z�֐�B��wm�eKj�ь_���|�v<�0�[P�H��؇�#��O��H%�F 7"���9i	�e�Nw��~��
ROd���B���R�<vx�%����[Q��N�,�����@�\����_�媕Ѹl�T1A�KEbF���������#���,�Z7Dz���ސ7���=�����彟�$��9դ�P*,�K��m���]����e:R�T�[ȗ����D*�%��Hn)���0vc�r��
ʵ�B�u0H0I��Y���rD6�x6FMU���(D4���1�8P�D,��P
סв�x��=�4h�}�� �rd����9
bO�;Xh�5s�"�LYs]X�Z~��씾��	�"B? ��~�7���2tn�����O�~.Om�/`0���g��XЫ�_�0�c;�7�R��MA���v�X����o��
��.C��� ��0�����Q�7�����4q֚�>4u=�i��+�-n���Vj�)H	�+b�+J�=oq5cz
�wz�DO� �������Fi@�����hP�5�/��}�(|oin��j���A\�b٭����?���R��?ΎlH`�q���v��~�%����s������ ���hО�r�+>�o�~
���H�ut����'���'���g/�2�x(�������h���������ʤLB�!�0e��B����S��[��{F���E���2��p���3X�U��M���c�l-����Bn���v�G����65��_����t..�t�R|��VSR����x���,���22+���$)��odņ�ᖶv���v�X��R����W��N�*.~��@Z���a��"C�E�����P�!=�RJ/{�Y����QAϝ�~�r� ρ^w��U~��t�h~�Ԗ�Dć>�M�aL)��y�fu0���Y���t�{�ˬ�ǬgL=����w+K��h$�����ѻ���
��/k.Ao+�]�kB�����U���=�R�������.��к���8AV���ٲ�	��п\�������5��&�45�K���!
��<i��W3Ɵ�G��h��L���̀u��-�t�{�" �F�2�k�w�Um��������+&�и��ь��O�;GǍɏK��*9o��'�����QԻ/MJCA
�/��Q&8�����Jn�ͥ���mH'J����,���:)-U��"x�p��C^�\tk b��U:djQ�Q�.�P6�ʊ��V�Z��c��ޫ��`Bq`@�?�(�Ո��p�c$�����3�/��I�F���|��I7p��C
�0jqayd!::�QE�]�籡�mh!VBfk��:+��YԿ�<x0
^��k2����us>,M�b�Y^��=H��mk��8�O� �n���x:�̏>(݃7����Fkٞ9��$�e�L����]�3�3D�'	j�.��13�g��f������*C�b_�^*��H�$=Լ��15���-��%���.��݃�>\�#W��i�]���e���T-u�l��9Ҩ�r�_r�(.w~��}�h<�ډ�<n���=M����d���^���O�ї��@="��'�;����dE��M�>{<)�}�D��H��c~	Аv��q��Dir��{������䗲�#��� ����R4�$�����8�p������g6{v��"[�<X�ОuA������,���kp5_�����Hd�Wn�[zz�ͭ���O'�*dt�i"N#���u�Ӯ�����Q6�k#��R����J�J�k��#,�;�h�V�S�M/�%�ԯ�ߨ���Ғ2P5J��og���
"jm�{�>��O�7K%�����m!�<�����ﶘ�W�iMTu�X����)��}�g0�ì�I�g~�D�~2k��+��I����|6����¶M,�%��}�y/3q��45}�c�� ��u�q���r���e��ƾa:>�!�N�/~��='���ݸ7:yu��4{6�`�j]��/U�X��7*d�x��ח}�5̥SEł}pU�j�S���\���?�i:���x5� ��pD?�����Rm%��!a~l؉znf�� �� 1c�?e��Tl��D�rpC�v��Ҳ#�Q�| HE���=rޮ��*�v�-��϶!p��G�N�%Ԫq���,;���/X)�J���c%��g��o�K���Z7��|��.�	�b����k0�Adz�)$h��=���P���c����@���ZT�E*ß*PDװ0�D��X��c#q�^YIO>C'ItNό԰.}86�5�s����Ł fU��tY�}+�qi�oHl��dxiy��p37:�[�����_��_R)zQ�l�*5����F"7I�B���֛g��m2�Y�̽]�^&��L�/!���|󰶁�D7�)�ʮP�=n�R������:W��DX.���kie����z���[��d��m	I�r�C�F�F>���ی�����m��K
h��3��/�Ȇ���J��Iu�|���H��D��u�����޵z��[3#�������5�Ɠp�?��M�9Br�9��ƛ��'Ӎ.w�[��\'C��[3�Ӡ�}'����ES�,�oW��zAN��i�p"VeEZ��Ɵ��2� OA4��e3sF�D�x��y&���^��/ߌ��q��id����>s��ۺ�gV4��9+�0z6����2P����Ի"��Nwn�Eɠ�M���f(��Yb�����Z7����
�t�����)m�Z�~~"2�f'K��S��,���%6G`A�gm!u$�4�}~��aM�<:�8h�:��@C� ��#ϧ������QG���͡���M&�osl��|x�x&�"W�ر1%�;��e�P�rs�i;��N����*�ۿؗ�9�pd�������"/ў�,�������4M  2r�dʇ�k"��.+81�C��u��!���\5Bmm>�����D����|?m0�}ʸ�P������ �����?��X+���=L\4�(��)D�Y/�ոۣK���v�I�_adZCd�kPq�(���I�Rd��î���#SEv�j�ޚ�3@�\������<�Qf�$ _Ģ 7S8זV�0ߍ!$�\�T+�Ӵ�kx��O�T���NH�ȯ;�Ns0����f5�G�5��g��3���X�rv9��q�?T��I�ƅj�~��cN��炵�aB:x˻x���;������.^Le��X[ �*�}�}j����S
-��XT��3���rT=�B.K�.7_�s�j��1�%u��\��5ֆߩ�].֟���
!RL�x�K�e�ˀB�hPj��v�	��J�v{�"��������+=����(e���$(}��i�D��67M�v�f���/
!n7�Ȭ�d���1cG������;�{�� /��c�6�}),�2�;~��گ�r��>��2�B���1O�T5�L\����2�:��h>\Z1����}1�M=�ȷvNF�ɝ��|{_a��h�޴��{����"�9C�r��Ӣ4_L�B���S����J� ���Dd1yL}��jظٯq����1�*W~��M&�X	�}�F�7L��"|�X��س��{e�~7�y�N�}���|��m��H<x�<wF�P�*Eґ�쫺��c :I��2nPVdC�v+�'��+v����7�y�斦V��f�+�Y��4;����I0Z�bE�,C������7�¾��FG��κA�'j����` ��P�~���eq��W�nv�:'� ��d����40x�	;��״Z�󻔒���tk��7p�$�p�A����V��K[X�O�H��H��N��ѓ/c��ۗ�������L�˻�LkWr�K\Y^��b�����V^�{�l�����NNYj\�g?6.�t��*�Ġ��+��!0'Z�R)M��c�F��8l	��}��*���\�e�"��
��휠z�����<�q�U'�	d'����W�&�F�(��}@K/K�n�$p�H�/�P� �Bk��z���d`�χ�T�o��
�,e�{�=���ΐ��P�$��d���H���;^���]��F�n��`�Vf
{*Gt%Sc���G�A�?��1iKYe�j�`�_��K0�6�G�3�7��Z��wG���A~�yDN��Jܧ#>?d��JC>Ob�l�!2$�8a���P�8�]�	,?����"�)��r=b���cV�n�p�SNZZ4�5�c���y��ߗJ���h9�K���f|�4��|���@��ܭ���ev�}9�W�:�;�c�O�7@.��Z*�oe�vj��O�'I���S�o�(_ց�]A�5��uoc�z�`{~h�^8J3�xj�_Z�(�Р�o`��{XU|�[����A��Q�ڡ}S�z�^1]=\F�����F^+�͗57�i����sͷ�PQN�����y��У�Ac�k&�v��͟ĚT�@*�T�y/������ ILk�7G�bm�H2(51tygeqwsu;/X�RV��e������ȉ�ģ�w�.B�����-�Km~��m��mĎ�ި�����;�:����סf/�g�����GR�`y��w�:�Z�aaa�OOϸ��jS�i�0�lM3Yl�"��P��id�������#i�� s[����"�veƴiG��!�y͟	K��C�[�^�����a�΋O!�/�)X;�Si�&�r�ʶY��T�0�v{Tc?�{�%��k���1�<4���O��!~���}�SZ��� A\OH���pr�'�]��BQ�+��ϟ�~1椣�-�B#�#�j��,ZBB�B	�����U7��JkB'��n�1Σ�Cu���!-?�P��e��i�,�p7�UdZ� �B�v윷���bkG+�ŀ�fj-�8�Ke�J���PX�[�C ��cv��ۗ�j��^e�'����^��5Z:�m)� ���U�z-�>�@���$�R272�G�cM>&n�������JN��,*�bt��*ՠ=���ݗ�!O��㰺�%�q��&��L��$��G��>�CG������
S�����3�����JtЕ���X�L9�nz���'Nt"��Rz!�!A�:�@�V>�w�
�}�b<]���s0�2|�l��tNl�����p�cr��*��}��l�zCl�M�j�C(�J�?%F�T��R�-Eh���@�'����A"e����(Q�k�o��̰���C�����1�}��k���j��Þ�u�R�[��,�`0�D��{��:��i�\'i���y-�K��=�wy)oE	�9͙f��`�`�aˣ+`�G�G�Q �5�s���!�7��_K������ED��o�|̨��|I���<M�!�V��Q�R 4��~Ӻ?Q\��ֈ����o�FY�Os5�!J��M�)(b���t��;��y�^&�vX�K��8�7�����U����`�A��e�01���(��2W�.�����O^�����Jp�%Ü�D�����M�t��Ajˋ�$X��3s?f;����?���v5�)�'�m\|𣖇��
|y]3
����"��<I2n���HF?�&���7��7b��:6Qу8����߶~�'PU.V�Z��TAF�r���F�}�S��c�(�|�wS�EՒ��KO�_��'�ܮRҼ�Κ/���^\_y��.�Z@|��<tm��=O��u�r���uEV�䨑0��l��ԏ^���Bq��I�
 �}��CN����z�g|��bO�9��ACB���g�G�;�:[��[��S*]�03�VdєVUsl��p����I�<�"������m3h��8�L�#/!���k�W�vv?6s�@��!ѿ@���9�I��ʪ���A��SVM�6רX�� ]��'��H�k۵��3��}�$�ӵٯ�-�;��[�:8���x{�;��|��j��6��`ZףZXn�ԟo j9�(�u�mu��%s�7V[��8��I;�8�J{���Ӻ���Hb������������?�A�5� �\M�-Գh�� �"�Z�����I��)(D�������%��L�|7i� yU��X�+5<WH1Z�C)j	�=�?c�_Sg�t������4�r�5:�Yb>%���s�%��*����@޳�5�nܤ���O�8�_G�rt�x�q�s�V�A/y"����E<�!��!-���*�C��\7�#��/����bx�Y��W�i@�q��r䣧׻�������;��(aU��7v>p٘qw�������i�O�
n,,��7��;>&=b�%?�ymĶ]�eq������Κ�T�Mqqk�n�� ٜ����5p�d�wv�m�l���Fkz�c��d��Q�	ZP�W���A`��Q��;�-��=�s,��tF[�u����b�(����wF��K�ʛ�8a�t>h�<�K��rv��Z|Ae�(�o�VbI	��Q�'�H��$MH�^^Om�]yDP,l�y��
z���WD��ܾ��G�r���ð_#Wy�5�i��%��P[&N��7x#?��n�3��Y����?�]�ي���pSt�4T�Y8,A�h��"������~��L�H���R��KdPz	�cL���~�Z�@�E�5�R/"�'�f&�I?�U�h�k�J�g�߶�đ��E��	yNl�3�;�٩U��G�C��%Z��i�p�8�Ik�b2�1P�����j��>�����5[���~����i��=�t�S3�c�N(t[�P�70
`�/��O�Ӄl��e:��:�m��A��H+#_+�J!����B$2�"�	�|�ݍ�æ�Hҭ��X��C�"�ؔ����S+!��S?����R����"��TPs{������7�M�K�dt�&���У��n�A��Wg�C�UD�mߏ�^^�JJ^GNbv�l�4�iLq�,�.���V.�F�+��ͧ=�5ޗ)w끽o�v�o������/z�^�\Sx�P|�M��ܟ0��p����6s�e��2a���K��ⴎ��X�7����Bl&>8s#hj<��}�;u~�7  �������R�ۯ8�8l�lz�j�<zjRzjDzj<�Dj���?b��a��&35�|�r�z}\��"�R����7�vO�{������ք����I@m5�D�6��W����]���賗�3:ƣ�[O�$�6�<��p��z��%'zL7����$oħ�tO2�<X�[Sj>5���O1?��}{����8��<��Xa58n���y�z݁z4�K��u������g_&jš8�Dq*��Bg)�g�s<�L���%(�\��8z��G���s1a���a�
V�0?�0�j�	�x����ӹ;���l�F�arj�~�a��G[���CGk��;�}':zLao-��\�9}1�P�RZs���5���=Ì}֍�D�ax�@6�-d����Ǳ�R�A�,x�Ü�>є@E�KQ/ҭq^���!�Z4�g-�U�A .���z,�|�D%�$��8��A�X�O	�|�8�����)�Њ�K�$������Ʉ�cڸ+�9m�(%��H۽m��I({���B.�}�����c�jv��25��^2ݘ��^OF�O��K���ߙeܰ_e��j��1����/�2����17�@�ϠI�Z����1HG=�j��\�I��e�1Gȇ���&�]+qED��e+{EȒ}�R�VH��?�`�ْ2��p��TNe� qE?�X�:=��	p������@�8ʊ!����Yp�����sr�y�bd��a��ۇE��fZR�p"P�"�T��W*>y8+Q�b��DT�D��T�,�7�#<�������PC�.�?��z[��y�&�.v���a�V2�N�odƓN��6j���¼c[���L��q��F<�~���l��j_F�fi�p"�*��Z]zx�W��^==�gd����#��RR|i���P���(�Ｊy�"�k�_/9y���;~�|ٝ�}ޯ}{*��R��Z.�|���x�����Fn^������� ��DD��v�NY��<�i�g��1�:��Y-������d%���.�ߝd'�5�bm���������q<������%��*��
$�=k�Xd�c�A��c5q�H��F���_�w�eb5UU�c'Xϙ��p�c#�sE�6"�ןd��/�t)�Z�HV�#�
�D��]�g��jJ�K�.�D�_+5�_/i�����z�D�;��ϯ���C��}IP��E���Z)�5���qr1���Ѻ����m\P]��v|N�`Rrճ7�Z�eLw���s�����B1�
����,K��<4�9�)͊a=Rf� �kô������B�l�{]�m�qC��<)pf���C@�*Y��`�v��U��xP%��M�z��Å����kݓ��sTn��>�O�:�q~eAc/Ղ\���\�q�?�|�����x��9�z�"��I�B��z4	�W��M������iۻe1*�,��B���#��[�g}*'�<��q���߉�  @��	�f%�'�3�ф�|$��<-e������/�xq��#LI��E�~�/C�T�C
��z:`% �Y����t8����楜�I���,i+~�١����9�n��
�������5�p��Gů╗Rf���jY��I'�����4�'M7�[p�
����t'��0U������M�a�Ӭ�d�2,�L���/�onr.QD�FL�Z}��L5�Ya:� ��}��ɋ8�%^Vڒ.ƿ|f��q}ȇh�����^��?0x}Qق@��3%=T�܍��:ql+,Iu���0�w)��rJ�$��8��P���ތ�,�� pv��&�ˇ����SH��g������=����$,�0��������!�6ΰ ��N����RR���*��6Z�m�b)n�-��	��ťH(Nq)����Z�š8�������}�?'9����]�{?k�5ߠ*�'����� �n�������Z	J�?�b%��t;R�;��7��^����r�Y�5��G(�w�F�[$�)�eŷDG��L�=cR�խԫ�/lr�.\{������i�U:�)h1��U��VW���� 8UU��7 NO�i73R2���DH�>���G�*�e���|C��[����Õ5��mõ��cp-���$���X�6��8��pn�{,{�������3��Bi����A��q�獪AL ���� ���������JR00�J#�б0ϰ�ί.��]\����<ܝ<�]<��4�-�{��WJ�{*�R��I)X��ْᰞ�����/��[��5��n]�z��a?�(����s{��3Ch�;6�����)kۤ����{`�̽�	i�ߧ��ާ�m���3LL  �0�BA������
�߸P|:�W�c%ө��i��a�>!�8��I������o$�����Y��5�w>�fmX��A�=�0�LY�#s�4�U�_[�HrҔ�LJ*b ��ß_�(���f����?4~V|��y�T
��y���4�zy"2�E{�"W��θ��A��nx��D�N�!Cl:{靻�#r>��]�c��j��}��,�@Uk����#P�g�G�c,5}����1pG,�
��'뱫�}+�D4��;J�@�Ծ����n��٢\��x̨�/G]���#A ��� ��fs�|#�$�YCW�l"՞��܆�_'�o�	�� ��q�W�y_�7)��4�P�l���^�x�[��pX��|��=�'��A�7�h���W�3e�+�\:Y��S
�z��6���a�ȝ�A�2� 'f��X��|(-8��E��h�D��-�T�N��B�Q�a��?m:��.��)�C�n�U���	T!��R##bN���xZ��D*LF�6��m�ޕ�;��N#��%��TL�r%��F�:~����~��5��!:N]9>��UW�ŗ8�CĭH�^�Hl�/���&|@,�h�&wb��S�FH�I�K�,/��˛m_M�ekg{�����$��r)ɦZ��<�l�sߵ��z�v�@Tqa������obm�a�ܱ
EG�}��	��������չ���n�M��\*�SO���,�������V'�`$�tM�̔�_�-�������k�@V�����f�݇�s[T�I-Hτ��I%����lR�L%S�gk���J�)��	ϼ�B�����',�_߷��C�pw�WsEp[U����n�I�������J��3��ʳ�ѷ��kBS�ӓ]h|��Qa%��=�M��2�{_���a�en���g��<���U��[����.u�4}���5��@�Bk���%��*h����EE�O��Ⱦq�Y����91�ܿ�\P^�����/o.ܢ�.��2�e�U�w�Zx�\cSc��j:6�8���`�89IO⤿n6��m�ۺۺ".�p��,�\S�����.O��h�7Z����Ǐ��^��a{ff����Ë��A��5�'|`��ZJW)*
���W�*�?.,�cl�ߡ�o��a��pSu�J��+d^�΂����x�%M�S�A�<�x�H
��GMɢNx�2��J�s�]N����2h$�á�۴�ٷe��6
���Bl�l�Ru5���5��hO|�rײ z�B%�(����}���@]���M<�Z����i��-=	��w��g��ĀF�GY�=��{�m_)���N1eKl�nXx��b�t]eB�����첗�6���Y��d�=?Uv��;5���y�1�j�D�DJA�z���ptq3f�|2�DsD��t3����Y(���l�k\�n��=]�j��n�
]���#��W���LMI����u��h$�`f���tk�}^�����ג�/�#�56���ٍ�8i�o�T��~Ǽ����؊�����_Z��ᢋ���+d!�`��D�@_薚�_[�w��f��J'�c17|)�� ( cv>���m�GO��1�]��^�-��}!� d�x0n-�����? ���U���d���I\�tN�c>�֏�1{4�N�2�f5�$H��*��K<DX�)-uii��Q�/n#��@���z��P|��:ӞDΝ#5l�����2,�qoUOP�m�Y�~7OP�{��v��{� 8�nl��}�ʀ ��t���,��uͨ��S���<�O����5ی��T���-{P%&:��1����L�Iد����%h�~*�C��<q�Ò����������Su��m�c�z���y������������QC������涣��=�ﬂ[�����WWX�լ��:*}}7��#�$F�T��ʜ5�}�ʱR�Q�]�Â�$��֚˷%�"�� =��#�#l�_=ꍦ�U�ۓo������I�>߆�t�]ڷך�گ�lB:���T�̴�$%��O<����4��Blܸ��53��UC������ss���]��H�t�VV��E����xPVz�	}f	6�7o;L�;���'1�,��0%� ��eݶ�Y`NYK�Q+�	��J�Xy�-#F6	�����]mS�F���t6L+q�@�"��귢+K�Fd���`�~/,��;�4'��"������A���wJ���1�j������<���IW'[\�d*�jG�v�A!l�@�Ƀ�%��Q8�^T�5�Zw�C����r�|��|���	����U�S�3?�ݙ��*�'��o#	<�RAj��"���[S���B�ܧ���p{��Ŗ �����^�rPH�"y��J.6���#�����D�X=�D|ĳ�R]�b�N�(1`�W��9� nPHt�/�׬��Z��w�ua?Ά��[�2�I�L�mB�4�t���$C�k�"��C�2�U�W.97�9=E�fKl7�=�2o4#}ܯ��\jR����/�>�9r���|�Nu���\�^ L���
�EF�/z�[#2�n�+v��L��I$Eq<�H�H�>���v���LK�^/�㽧z�D��.$����ʑ�>�~�n,n�n�9��u���\����p`�3Qϊ�c�X^��_��c�N)��.�TK��u�)�E&��o9&�!|zyx]�\�z�We/2 �Al ��)AB�"��)��T� 7��{�'IU{L�\r�$|_z�j��RZ�0�G�(C��l?�Xw��x�ȄDӥ��7�4�jӗ0[<LA$e�i�0<9:��>Qo;ʪ������� �.�O ��؇�r����5ޒ�N��߅�����&Lͱn�Xq�}d����ݩ:��I����zh�Ȁ`/�O��	�?]�\??-�?]eu<<m;>�x;N��M�o��cr�w�W��/��m���Ȅ��H��T��̧�� �s�0�R�xSJ_T�.�bP�����/v�q�jP�r$E�}fV�BY�Df�JFƔ�n�ִph�����7����MHO׹����g����U=�������X�;�V������nۃ���NH���y��	5��Ft�̭~��]�h���x��EY���ɖ	vP7���ùZMI9"�E	& Jfa���'e�&���mJϪ�hB~�Ӎ���	{pf^(���D��o}$���u*^1\�iw!��G�`<��357͢T�&
��5)�7�DX+�Z�Bx�I)[4BmYFm+�kٰ��� .�g���5��O�G�	�=�B�^���B�|d9��	����Վ�w��<RAPY����N��V(~vIk�w���%[3����1�{�yr�z�$pȈ	ąJRŔ`]�������יT#��ǧ�tKNR�`�Z��af#=��L���L)��?J݁*�a@��rV��j;���1���ٴȵ���F�������G��
��'���M��"H�K�(�/��}9喚Y�X�E����᳋;��WB>�r����Whʕ�6�Bo����˅/J���'A���S%$�߶�����J�	C�5�_�1�����r��!��QV��G$ Q_�&`&9.v Lp<T�'��"������� N-�� O���8R�oAfEC�^����Ga��N���j-�t��9�F��y��L"�p��<��5)�&��B�q�@�;��V�V-*�{!�>Zt��R��������ìCO�m�:��Ks������ͧQ�4�����S�T_�{��� j��Ea[��]ʴ��X������x�~���d}��8x�xF�J7�����Q��ݐJU�Я҃�Q������*���A�s��s�M�Py�D\���qqqD쾺�����r	�ǆ±Hy.J
d& wf���D�z��6,��t��!�~ZI��T���͗�Lc��
|���m�Lx�2��Yy:;}X@����V��*�i*�y�j��:��^����������,*z?��K�Xq;�3+�Ģ�#�g��~g���.��U�-E�s�-�&-�V�1���!ŭ���|?&++���ҵR��&5'��5��5��5�b�m�;�C8����!�O�Ea�QZF{P3��P�\Ⲭ�^�Lt9137=MC{���t%�������}48k�S���!,�W�v�]d�ms���0����t�GU����c�F����L��M����o���7k��w'\	�p� 4=��<&,&�Q%:'-��h���k������ w~�R	W�K�X��U&η*p�B��֒u!�>��E��o��}ě�gnù�	���@4\/{ֶ���GNˁ�pC��_f+�w�d�y�K���˗#��!�-� ��G"I!��=��/���;�wV׿f�&�'��.s����\��ȶ����\
Z����ڢ����\+�2#P\Z�j�/	��>��>�M���'��'���L%��S@K���n��E�|�?'�Y�An�Q�Zܒ�|>����1n2�_ˌ���]�a�r��F�TR�TG�!����-8���%�,�OL�S�l���N�Y=�q񶿶��0#�
G<X-�i��[��wN��[6�u�5I�Hy���N��(�p��\*m�� ��`a�I��CaH�`��tP~���"�uJ� S˻�5jB�M�x����A���V$��nԢy�quj�}�<��g�!��f��{s#�Z�d�ߎm7`9���'�j�� Y7���̐9P��n}U�i�᣿ns�w��C���=�T����.fi܊5&h�4w��z���*3�{ζӛj�r�����6HMgހ�\Ң�R+��r���8��Oօ���GJR~o=?ڇ�J7�	�$&׍�,ۚ�F��n$�N�3���9���UZ��pE��a�G2�tM4�[c��5�j����iW��q�&܏��P3�ދ���{!�p��B��\g�S�n��C�c���}�	��������1�����*���iu!�&���bQRU��~�ǫ��>X����{٤]��wy�&�˞=�=8�tjg'c�4AU���me�|A�C���.j�g�z��;�y�����S�w kT
o~0/��;Egj��~�.�������0�3�������.Xy	�؟�MZ�'iYL,
�'�6:�{�œo���5,�I�Y��k�]N4M��\K���<W��T�{��߂ʹ��DD����Mހ�{�G���Z����c�����cU�����X���G��燵�����[.=DG��O�M��ToU+���^��i�0;�z|����2`gqi�Շ9.��h�����VA]e��xc�n�KkrW� �ŧ�j��C�f����,\�ߛ5]ͺJn����|���L#�B�gb:���A�c��H7�7����祧�4=ޗ��_{�?�9��>��/v���[K]pls~F�Ф�c}c�<�W<��UW|/uT��4��aYF�Ɛ�D��oc�.($s�n�E�es��'H��ZcR�c���d�88�oU-DC��-���f�}��K��@��K�tw0z�	�J�<�""�f��p��K�^����D**�)D���5V�}HvA ���)��1�0��!���h�҅rR���ג����xvPn�t�],�b��(V���$Ξ Z"?}-.m?N ½r�eH����@�ּ ��������q�_K��\��~��fƋ$�g�bc�l�=e~�t�z'G��;�j��s�w�VV�����{����8cK�����Lm��4�ޜ���f� 䍉�}�˱�u[�0����!�[Q�yn@�Ҩ{�J���f���i�M��7[��H�Ȥ=�)jة�[�N�0ztD�E	����A���Is]^;#�����	�9�l5�]2���A��g���T~�S,�G������QF2�统�^�5Ю8Ls����yyM�+>���^-4�袑T9��^��^��djZv=D��H�̺�魙�8Sd�E�����h�c�A���Wj��:$��=������p�w���:�$ܪC;b]�3Q���n���4,����,���E87�n�]�j�#��:��Qw�5%���X�Uqfi)_��_d&�t`����i�i��U��i#�S*:C�; U^�do�o���b�l�q�eb��./hrE㙉�C�'��$E
�ڥzk���T��& ��(Qs�q+�qo����,R��i�b��VJ�������j�V裳�9��D�0�<�oЉ)>I,%y��k��4&��kmk��*U0>�6 ��N?��[p��>a�������r��]Y�t�nz��Hc�?YR�և��2�F:�s�;׌���������߫f�9w�����������|q�3]����u���}'8����er�k���R::��O��ģߘ��~��Y�'�a�8Hk�m}�d�=b���x�4y�	x�$:�]��Um���z�b{^�}X���긟xbx��{س^y7y��p�x�{���3�(���,3shg?[���������h$K[�8)+'9I+;OS[��tdr�j��=�q�U$���nr��:4��L����}��g���j��S����
������.�
���w��(��۪y���?D�~�4]������?ߌ��}}7�O�{]��߶�p�սP���6|��#nKq��>C�H_�0#���j8�@2��ߍ
?�Ց���XE��;������M�k�#q���`1�^�����}_A�`J�PD�Y��'�$AA0�oBF6���-�,*�,��X
����-�)����ї�J>�'��Ċ7d��W,]���a!����b��)pn�kty�D�Y4ٯ�$`'75��S�Z�U�#Wo�ۛt���=]���PW��lG��ﰡ����{�����$�m㓓sI��C��\���+�a�R1a<DE�(	��>�d�ZL>k�GJ5^!����e��w�Rs��Uze�h
�e+��P~#A[�]�?�7�`Z"wB�����k���LC�ǵ��̒�}k��t�JZ�[*CK.V
'M����T�P�z�ke5�����g#��_�s�P��3���T��ոHH�}~p���ԗ 8US�Y��(T�YGµ���%� 	=�-�-�i>� �l`!�\��n�48�Ur��D/M��vI������'���eƩa|�#��
��Ċe���p�9��v���>F[#X�[*��~���Υ�3O�k�v�j��w�c��]ᜇ`�@G�f#q�u#�q�J��h��Y_�;hMr��/�r�n�3�*{�Bl��۝I*��)�<�,g��<�'��d�0c!6/!yU�'$�� ��ڒw��J/�ޠ#����p�H�Դ(���3_Q���4H Z��uG]��]Uu��"/���ۧ
a��ߠc���a"��TY�lh��°JIg�Po�����Z���ܿ���ʻ�!8Me���O��o����N��dW�T۟v<V8>.�\o�>�x��!a�2���#��xe�q���������>�p�J;M�s�.	�3)�m�>"��m��s;^U�jO21*F+`���-��,��+.�z��L,�>�RᲲ������c�U���������T������f+*]��|z��aߡ}������i��v?���A���p���C����i�j�Y_0�c��I�`[���]C��r�i��5���`�UL��bq���Q)װ�}oz����UUHxV���[^CSS�����P���dR�M��or񹉄\t����'�Mf�g][��u�΀�!(�kMTQw�ը��"3S�C��\�<���E��������L��n�ڂn���$T������AZ���L-l�m2d�@�>���G���o��yIv�-���ǃ��f��k���iOmt��������a���}��v���uw��?��e�K%�IPٖ��Di���P�x(%}g�)pg3Z�;��9$�'�x��z�S�ɕ�G'k�Y��0,�z��2��2	$Q�md��� #[�u�=� IR�p����`b�Ny�`O{��y�t�H���}�h�j���,褉��=���9��� ����2�G�򱸝�ea'ӣ���n�hk��h�\�)��A�KPq�pq�����>�������u��m�_Ճa6
����gC�Ij;�.J��f��ھ�������YΊ��=�{�r���;o�ը���m|�|��6����Hn�q�QhA%u	6��磚މM�n�Z��h�ܢ^����0ǯ�ZzE�a()�oTT K_�L���QL��nR9�ׁ$�2�b� �f�B�X�\�G���]v��0�j������e�o����������M�������,\e��<���� ���2�dZO�6N��cP�.���Pb���fEI���p�2B9La��[�!s%��^򡤧(��MPy(zMd�i�,��c�wN�J����{� ��g��WX��k�/`_��'�U'�U���H�۳�sPo)k�m�#J�h%=׺gK�[Y)���[�q�w�l���5�s�)�>�~���;i�f�d�wsf�r3am�i`r{�+�|��T��v�a�{��m�pF�����|]��L)�g�s67�{��ʞ������2V#���9W+-�*�����(ie6���C91,�𪬯�״<(·�#4O,�0bs2�Ş;.N ��L��uud_�NC|N�rӦ�8�]�%_�C`R�|���s_�7��dz?���I����a�L����Đ���i]@�l0��zsӊ��Z�J.t�Pt+��`\^^��v���q�&���2�'꟎K���da��I@��(G�wgy0r���s̼�ax�@Gv����S�fw���'Y�e�����gy@I0���H�ׯ�4�R������/+����E��9f�/Ϸ�]؀�q ���}*�r5'�����Rs �{3<yF^�=I�E�Yq̂ֶ��_��>�BV�6��yx�;^�!&�F�U��tm1{)��P�GS��@�A�Hr�VX�[;�70�wx������rK.��JdV�����.az?����M	�p �S�/z�$ު%ε�LF2�̮���^v�!^܀�(�u����1�'��.EI�(#�	D���ژ�rچ�cq�������F���!\µ	;Go3�&��Spw�����
������U:s_��K�F��I���#�=R��{�*�m���>��]���`k3�B�Ut� �����(1c����Њ��@��1y�Ӯ��ˣ'�	<c�oZ��YMBy�-xL|'x����h��?��s���lB��=&��J�8��v�
���6�oz�'_Ӕ�:X�b@�T��!{=�m���.y��ƌH�<f���u�=� �����<���r��
�2	^���P?�z�S	�I	��i$90R���3�F������=a^>%?н��G�H~~�*(IR"(�;XR	�2(h��jr��U#I��!:|DJy5^���xC�&{w�~�ȯ,#lG���������ꁷ�e�m�ױ���|/߸����i�ⲅ��@v���y�F�����*
#
J
�J�r�٢>}Q4�DÙ�[���L�Q���h�Z�ZZ+/*�-)@N9_o2����Z
biB���Z�ޗ�G�x�|!/%��}F��2|��U^�wϟ�����T����ʳ�#a�J[��ᬪ����˽n�V�gͪ��,���}�e_O2�oGi���x$����$��2�DZsH�ŵo�B[���M��c����l
�y1���6���F��S�PJJAIK���L�M���bxG.	ψ��W��Fj:��U6�1El�_��=DOSH+�b��2�β������c��۩>�d<� 3�"��`9p�-	���	 ԝ��K�)���*	N�-�c<�����Ϻ[ 	�G��e/��;�����fU;��[�s��?�5EY���VyC�Ȭ�.2�������3P��E��q�0�b��6�X��;,�PKir������O�h]mG�ۜ�+\;{��jKIUU٣ v�/xa�l�Wi�&��Ǩ0,U�ޕ�Q��s�m�8�8�9���d�<[zq�N�hb���j�/^Rd+E�L���Yk~��7�4�����+�u�\9�0Z�B��/�*��CcJw:����H����	��:�C_#��C,�P�!���T#؉IΤ�{�����Ŕ�a��1���.��-V��u+���(��Kw�}�� ��*��q���p��<#���X[��B�pu���J� ��{�W6�����r�͉mO�Zi<\�C'��Ԥ��Wm��f��'���(�C�[�͜�"��%���M����}A��I��͟�����a�������Mݷwe_H��%�/�4\��v{�?��:��'@&������4���e�<�3Sn6B�!�ō��R���5�}2��h�1jѳ�p8i>p�*��� 	p޾%�#	�|ebg��4��^[��A�hB����X�i�����b�(\�\�i� z5���]Al��"O'\���OY�U��S��9v؎_~y����:���-M���*)٠.���)�肋�)��g��ۜ�4q���@~}𨵠�3��?$�Ik(�X��;�pm�nE���e^y��Ǽ�ޖ��˸7����W�1d���"7�i�o���1��ut�������6{��e\��}z�+O����僁�����sT/&,'B��1#/1��nw{��j�Dd�bMQ2�+�1c����Dභ����҂��1���]]�]TEE���Q�\��2�#1$6*��4�i����9��O�&�(��)_3�Y��#����؁8x5��+�� g"�c�������5n�$�)A�q~�v�V����Fy5�	O/�(u�N-X�F������G ��_h�l��I�,�=�`n��=��A�t�3����)6 4&���A[�F4�u���U�/矁g�r��^N�{;��ah�h ��Gy�-fL/
*$��`T>VAogd��k����P��7P&��/���[^�*�<�Lz���8�*�1FmW�j��9N��ʽ��������=��,Z���Nn�s
P�@�{e��=/��V4��V��!���D`(*�P�ԟ�ҟO��.�����E�<_�z�&q�d/�:W/��{�^k"0富`�������wE����p]ɨX��АR�)"2{���s�����_��]���#����5�9���zr^!_f�_�'���9����\�lU���z���v��Y~	����!�������o�\��/�IEH׷��`��}�A|뿇K�bx��ea�HB��@�H5{�I��H�p�=�2�'!<m��)4(G8�����oHl\)���!�h��A|ǃ�T�a2��cތ���4s�M�sΤN������Gw�f�*�M�z���늣  ��H�`I� IJ� ��`ʠஂ�|599e=1175'C��4Ys__	3+3+�/��iy��Z��Tt��wr�I��6��9�AH ��/��m�G��[�����W��O�l���`���2+Z
+7��r���WA�ەy^]@}�=̌yL6`�0�!%e<�dba��u��Vx/�Ī����iiv]i�Jժ��O/h���V�F&O�'�hrbN�~���R6�q|:R�b����8Y]�>��w;��~�V�s����|�����޸��hx�����¹�n~�<=%���T�Dufݲo�T�Ͱ����m��22".���P�Jv���U##�cXT�i����5�_����
m����HR��T k$�o��S�X�E=�	����_�d��3�a��ϻ����ךF�����%4�Ղ��ruM�5�2�"m����)�7JnND�:����s��o�4Lows���EX��H�# j�e�we��}d5�i�7��CkM�Wc��;0^7O���>�J��8�� St�	��j<q���/��"��\��w#J\~&X�$T�%ڹ24&�q&m��?�"46l'�Y��\����Q��Z%����<с�PupS�$1�@  Vs�"��� lz�I�^Jp�)(�J�H�N���u3A�/?Ol�$ �%�DCUj�
�&��vB�����I>t�R.��w6���60"-�5-r���-3iX�Aş�Jy:cd�V!���#��a��ِQ)�a�ҧ��7\��'
]U�5�&��@z���}Cp��t��:�pp��̪��^�H�Q*����NЉP���p-zG���x�j�"��G͜6-X,�ZYK�c񤿴Xݦ-�A�5���X=�[>�H���CGÂnf�F�L�A��BU
�~�?h3��09�Y���N	�b�ϊ�H��&�uL�+�|GO��ܕ��:�abL��xX��?]]��*C�72*7f/�7<���6�C66,�k�yx���yQh
�{yi"�0�ú��BCeB���CC�Q�CCC��V�zj��NN.�0lu���ےf���3�j*L�k���0�`e��Q�j�����ԕi���ag�LD��޻[�L����V��{
$�V�[�%�J�-�ih��d��PU���|��n�P�uY��3�Ju��6,Ӊ�0��5�7e�fBl�#i�9&"P�^��~o���E����ʰ"#](�?����"��sū~�h%����ddg��`�sY��dʺ�t>�NZ��@@�$ȼ6O�~��ҷ/L�G��/WJH�?!X5�Pom��JZR�;)�����d��
{��Rz��X��J�gp��ߪx�Ǿ�}��oLL�~�H��8�(�>)O���>��d��P��8����n�Maɉ��g�h�4b.M+5qןs����
JPp�$AbT��_� ����4e�؜9�8a�X�&�$(�vo����%����ȃG �蘕��P\��
��� ��qv��2�r�Y���	h�Kk��Aj���k�G��٤�n��+V�ن�����/_�0�h��ɽZh[:W�u_V�}���z?thp� o_��,�zJ�ņ�B��&��e��xXڧv$xɰ"\����uu�����aͲP��3h�'�h�c�lzQT��/0��K]���K�WF|�mj��I��r��r�(C����Q͐�tӽ���]��P����n���(Ug��e����
���,���s?O�NC�T��Ā��-��*�~����I���L��Ok��b���J�r�'�R��+��X��J;�H�P4��1ɸ�=��8��Z�D���k��ăT�Pj���3!*X�bA�q��:m�i^BJ��j*I�d2�:���sq�uKdC�Z{�CP\	p��'ꓑ/�tF�)����5�^7WӐM��c���(�FѶ\�P8"7�}�5���tǭ�e�`�`}�as����[�ѵ�������F��;�Ŝ�s=Ju��J�N�xWTK�{H��m¥��ki��u�u	sv.��2�s���A���Ҽ*DKF.�ZΣ5�$^&-���* �@QN�+��AG��ñp�A�Q�&aX�]Y',�J���y�B�DR=�M/D{�]�|Gv�E�[��"o�V�8��X::>0.E�2�=�j>��`�d�$kjv0t���(m~����^�<�4�s��N./���b���J��(�ü��l�����b�Od���jk^S*u+?h�ˀ1ޞ~�����\���a����e+�Jw�T`�6�V�K39)y-	Ϣ�5(�0"���~}�k���!))� ~�r�XgSe'S����@C� 1=9OC%_s�Gow+qc�Լ��6zVfF6�
��܏��:������ߘ��DXQ�ݥ�d��D���ǟ_��g
�����kk}����q]]�©�%v���S���г.�d��]�e(��#��=���d܄ؠ]�6����P���N��?�3�V�:���ͦB����Ƣ�>��t�˖��zHͱH����g�2s���r�8R��*;
�}�`|IU�˝6P�X�C>����o�a�翹9DÙ�>w��S��9��}su�ں�)�*y<_ƻn�TF�⣸��?����X�ǽ��kՏi�?�z$���n�����x���l��57w�������SBKK㳖��������0�2C������H���0D���9f�� �6��X���Ӭ��U�T�C$�W2N����ld��T��ׯ߀.�	���E�Rw׻����b�}�K�Y��H�6�D0o��*����c#E�l��P�Έ�����"�+��C4�0ՈĪ2�֢�M��v�
���(ɶ�կ%�-pM�ʦG>��7��4�-a���}b<V*��ke�ey7Ge[ɊR��:�B5]�%�*��*"տV��J-Xs�����ʹ�;\���6-Y�8��$��ۆ�PB�n��t~	^R�p��� q�]F;����=*2}X���ai����TV5@���H(7lQ*?�O�D�"�X��u��B"TS��hO�]l�C�<���M
k���%Q���N��x�e\�c)�D�8j��^�*�o��&��؟=M���KX�7�~7w�k)I�Ԙ!����1���OV�ֲ=*tOΪ�+֖_3�P��T+/z}5�:I׃�?�ŕ��lǡ.�����X�R���1$��$�?G�ꤨ���A��Mc�c+]g�q@MD�d�eO�*�_��Ɩ�U�t�JJ�p�׀F1�\�g��dy�����:,x<��}�"Lד�c��_{rp�ۣl?L���NA=*|��ԡ���[�������/��>��h5H1x�6�/�����>�+3����2���K���mS��|(�qm=d�*l�6q{$25�A�aֻA�d�`)��xۛ�	�{�4x����onu9ޜ���3�K�k|4\�]{�/K|��[�:0�r�`�&� 3�8!-)';#"���q�G��;��NWi6���g�x8�8H]�KH����Y�Y�V������7��q�'>�����#i������
���������͑��FFF�Z���-�k���kօ��x���f��;Q���=55%m�@O������-)--Ͳ�
�2	���HB8a��Z�����	�uLlq&�?b���q�����>[j)I��3�ΌsD�iц}��H;1]�@�5���Nߑߣ�gl�����㧩�֗)���DTT)�UJj��Pwp�IN'q���P��p�q|z�K���'���[��<�e���@qg\�?5�P�S�D�U�S�Dtuu�D��x9�A�έn4�X��B�T�`�K$��A��=7��Hc=��Q��E�B
�@�i_5�X�v�� �?6/�������$�u���s��������H��0vY���[�,�|��sM�Y������In&"M~P�k�Q�e�݋�}{lG���)��m��>�@p����ci��ua�^��{�Wۄ��\lV6d�f���u'!w�[�wY\��Z&����E���F7�E������)y\Ҿ.ڞ��(���n���À��'K��wp-g_+�P�R��@	�+H6;	;�d�'c�Yn�-9NF���x��XFyՃԹ �q���yQ��G&��;Q�8�ty����[Ł����� ��7D�oj��%�q<(>d�S���uzYoMæ��ى��e���W���;�"�w��ND#Gx���4�1L���1Ʒ�G>��$h�������X@�"�3M��z�a���	o��L1~x�Hx��6�N�CQ���eO&���T��?_��M�X�ja�Y���"0�Ϣ���!WI�Jzyqr`�Xy�G����=�8D+�P��?1$ֆJ3z�H�t��$�&|Fј�|�i��t���=��y�A��l{u�y �����Y�U�F@|�h\H\Ey=�m:PJc2�6*wtwx_Y�/=��W���_�5[c�OebUf�STQPRVPݧ1�sS�Uw�
]��J��+�'g�����?��3����U�T��Ho���� ��.�D:R�� ���AD�^C���t� �卿�9/�d&3���u�k��/�X��Δ�e����˗�z���z�H��N��OO$�43�����G�n[LLL�����4k6��g�����C��C���!�UC���X��\����[̜{��~�2�!)����Z�+�$�+�I}�$�fl��Y.��Է:���I '�p�6�aHJ�ۅ1I�������O�[��9p��f���88|���,��б�h�8N��OMN�V���PVV���E���FC$�s���xxx�茙:\��O�]I�<�9��JC3�d0`B��I�:�,�C�/�,y(T9���|����mSĖ��֯��|@�Zm���2P�����{���x�m�5�$��jJԥ��M$Oi@�z*/�Τ`1��p&�.F*�ug���P�\iF��\��vı3@G���!�1�(����7���f:������Z��F ����Q����N½��>{Ԣ��ge�ܱhj���}��r�J	;Тj{G��o�a[>X��#5��o��b�e8���[��-�d��w� ����Վ����R#;&}W�3�2�_.�M����au)�7�	��W�Hoy��µ#	rTl�26�L|����L�#�`�IR~���}��,ؽ�{�	�pZ��VS������4yY��F�,�Lo���~)����N1��e�5v�z1�{�LS�k��f��U�{q�?�h\�;�(,��T5�����>��Hz{���XB��%&��J�;⻠'o{�����+G�`K�s��X��'�{��_{�B�[�X��u�jg�{��@ٝ��bh��	a&���B��%���F�)N���������Q\E�C.9Vagfj�ЧI<��[ޅ��[�Z��_p������wf��Ӵ g�ˢ�I���i.!#2�5@_��~dW��b��ԏ`I�#�ڮi���F�ʶB���w?c<̜Ƈ>������<�F1�z'GB�y��8c�s�?ɖ�����*mm'�W>��}@ӣ7U�''�Y���WJ�/���^t��Zoa��!@H�e��� BA����A'����|���9�Y>�n=-�.���nmͽ�r��߿�8pE�hV��Ξd����p�%�SwD&��Ö���扩)y9�!����$��A��r,`U���P��&�<d�vE���:`��a���2���R>�O1d�֦��\�`�ml��E�_��Ԑ���o�������SU��弻y�DEU��EcF��|��R���)-(�G_�����E��L�K�A''g?鐍ѽ?����7���z�L��4H3!;[����H��\��E�j�������!���	�b��t+E��b����^�oS��Z��d}���D��C�kN1�yh�'���ٰ�}�H�ŶnLl佸��Qk*֤$C� ��O�c�=�>�]#�k�῝��|kn�����즵�Ɠ������'^������_��.�T<�z��8����P�wjLw�^���}Y����J�����%�-������]M1� ����QB���9Qq
�K��3&�b �n9Nސ���
5�ۦ�a�v�3t(w�C�x�4�;j1�r󬐶z�wz�OӁ,=[[��#��|68��9�y��j�#����gaIQ�v�v���ܻ�����A�;Ve�/�ښ{��lS���S���X�^ [�D.�����"��L1ULL����hf���6ۊ7G����	BSpLԑ�x-f����B�U˷υe ko��ɥ�����j�[�p��)[2٥�T��.L� '+�vu����([> �jTj��6;��>����ܝ7����
Vd�ua���_'�v�B%���w� �.6>][�H��g�#��WӆS!�,�}C&��?��>�Jzau�)yz�a����w'���̈�������-�xR�A��c>Ahw�z�(H��Y�
H�+�?��З�D��2VSP�r봲�s��U�����������V���ƞxMUh��s�u��������O�<9>:


��P(YII�ˣ�k���:뮑��� 0L�bП���:#p_ɿ�_�Xk�6��(��V��$1]�J�ĘAK�� nFwp|�R=bEt�s��h%�����YȪp{m����K�T���B���lrrz�I�z�g���&�*�ۺU5]��z�:R7�_H�>Ƿv�J�)?�q9�&��Ĥr�lp��������5� ?P�������PG#�%�
7y*��!�O����o8��G��C��@� R�>��x��Z�o>����C4�|Zi���������ȷP_�����?v��YK*[��{�����3��ow����־�H%�x��vj��.l�w��F6�!�)��ԩҘ��+@%��a�,�&@)a�����j�~����C�!�-�A� �Kk>GR=WK�n������Hd�q�f3�+`h��Ć���Yp�? ������6��[ɐz�^Jk]E{ՎcO��m1���,c���䲌T������y��Dz@�z;�c�Ժ����rW	7y�Yt�������:Z�4� 2����[�?dM'/��~cYl�`�����27lP���>�\�^|d(Z}ڱ�IJ�]f<�
S��*	�����r��Ҙ�$��/���{��e �P�0��I_m`0ڿL�+���^��/��e2�J:H�bm����+O�_�'���FGt��x-�d���A���@�mU�,���P6�����J��;�����L���p��]�>3�?��S����i]���	^�oy�&�|݅����e�xo�8�m���e8V���E��S�x>H���_3�V��B����w����｝@џ4R��͜�ڋy/��P��Ie���C�y������)�����C����5�Ԍ�[�yNH��GG%%%G'&&��uEe]�ͽF�|��=��N+9EDHA~iw0�V�Н�N���ܭ�)=磌ܓ$�E�y���,�J�4?.LO�A�þKk���Y�P�_6�k�͹u�;~���b����Q����������&��J�0m�����W��N]L]�捛`��9�k_�H���HP~�ȵq}�<�}���7d�R�H�O��Gr����uX0W�'"w��.ࣱ�k̄xs-�û>��4׎���Dq��,��7�o�x�lki����o4U57�uXP���:�y����i��5�}fs/�)�e�T�4&'��7�|���q3���T6��n�S�|���^v�Z�(Ğ�ϋ�Ȩͱ��c���������餉d�$����/sN�v/��,�hm��ޔ|��*
����◛�#��~�3a-	df�),T]����XdZr4Z����eƱbjwS/k�źv]f4 %�L��n�y���4�A�V�rg^Bk�łs�Y�%�<��5���\��fn�Q��p����J���dŹ��d��ɚ��-�SD-I������B��ّz�ς9�<�E.v|���O��~�ܛ?'�`�#%μ=[NH���PV�\J]�(2�Ñnɐ ��<�`�;��iga�Cm����(��.�z�5qMն�����5�*������?ʟx袩��:"���e���W�G�w�o�4x�d�NPe�Z�uaz&�\}��b��@S�B���r�뛗��/",����z��e��x��I~�_����u��w�d�����H�#>�0L7�>��9A��Y�߱>�#%�	{e��:O��W��W�5r����C��&��+����-Pp')���~��k��ۂ �i���<��
ܨ�sZ��cmϹ*�������r�5 ���ۋdo-Sy��ySZ���.i�����V��<�9�Z�P�@�uQn�����!&BDY���CvY�J�״�Y��pJ�0�fͿ�
���.�l��;��l���� �<7�R�����1̾�<9<�Uckb�F:���a�H���J^~n?�K�&M�Lt�k陌L�<C��V^q]k��9�fX�
Ę��/�Z�<c.�|�OI$X��æ��Ng�(�Gv{�8	��
Ի��rbz� X�P�����Tz����/�b�Ƽ�/��iQ����(�#f�4grG�y7Y��?N�C�Z*�b��ڛ�m��Oƌ��o��c��g�\�w�t��s��I���ݐ��q��BPt!�����1�֝���� �*�������F�67+�[������odH�7WQ�'k<U����2~/�5��e��DX���~1�yN��&�ʝw@�����X$$�P��8��﹊3�tO0�_�Y�A}
��	�`(��	b1T+� �Q���jnx��n�E��*4��q���{���ћ�q)��������Px��g���Ƅ�`�R��p����3	���� �63{E��Q%�*M�GgK�W�y1���A��bT�c0�+�1l�:�G���bDSE�)���ɝ\�n�`�*YM�t�gR�xƝ�e"�lWF��Hn�:O��"�9Ҫ��^���]M���z]�?N~[�Ѳ�� 3]BH�H@o|h��:�aR97J����}Y�Ŕ�32|�g�Ok���lK:*�aޟ��M�BV(Y�m����M7���הa��_���`p���|�+.>�-3XY~��0��H�z�oRR�&p�0d�10�n�;'��Eo8њ�a{9� K	��#( $D��n�81!�6w)q}�����-++����@OOO;;;S�l#tc.ia�< �t��d��A�:��M���J68p#�N�s%b�D�!�������eً�Ⱥ��P֦>�avTr�GdN��OW8^ӽ�4�������?ӟz�:d��;E��I�COwwtt�xI��9�
$[iZzWeb�^��^_���,$��;�A23]��P�  j����z��4mۿyeo�`��O��T݋Pn���:�H��2v��͎X�$�����V�[�_��ÒZy��X�mn�;���*/k�K�����3��cH���W�Kc��"G�Wkc_��7VO/T��k�S��+wÝ:�bN=o�}�߽|IbK���H���!�u������yĵJZ�v~��z��[���t��b���e������㹜\W�K��)�@��g���]�{��֎�ƦB�,�	�ж��I��g�E_��j���Ȕ�,���¿ȝ�f8����냲�����շ��Px����9�������"�5�g��?��M�>K�x��<��Qéڗ���Y�⦽S�����Wx8)��M��Rꎅ��r�������ª�[i���̥`A�7g	�i��#||+��I��7E�)��
L��G�4BC_
�m9j}v����ݚ�}8���w��p\Ģ� cZ�b��x�հ�5�,[�`��X����Nue�u[��2E�[˾dp4bh>����A�oVk˴�����k�AZ��^���S���ِ�`�k`Pg&�LݒV��q�ޟ�oٝ��ۇ#��{�lr�U2��Ge;��p3��8nTÐ� �_�t{��}��J�@D�w�J�Vd�S�"�yE�:В;Uƞ��¸t�m���po�a��a�XO�O���ʗ���4D�'=�5�S�_��ߗzU#���Woۊ;o2�~͠�C^���C+�R�r��MV�א�R^��ۜ��p����Ļ��]|%�RHξ.�:����Z$U�^0��zq��s�v���#�Ov��X����l�®9^��uh�H�K����)++Y`6875xƸ,ޕ����$��吼[%*.�PWw��Db�|=j4�D}�
�'6>OG�qp�R$H����䤥�ɛ�c�;k�򇳝/�}������]YY�Ƞ��p@"��<hn�i���p�x�"��s�-��j���N�L���i��)L4!	L�\oL!3��O�侫ay܄(H�(i��!c9%.lXz�h�Y������33��X�t�  ���&�PD�re� y���ɶ�`�4�<\�����d󣙄n���f��Kl-��B�:��j�C,�O�"��<Nv1���J�W��!:N�~-wQWO�%ty6�l��{�o��oB���,�@ ,�����D>iQ������j�pB��XV��.c`1{�u�Tt�hh2�i���p���c�߫ �����:k���h����&Ҋ���x0�s��J��i�Q}���`���:���1!� P�K���93�Ɔ&��~���;��z�B�J�Z����a=���U^�	\��q��v�{��m�z�]û^;s���y�ba�g��.��m��0���"Q�]��&�5<r��肅���r���,�U����u4z'd��؍.|�Y{k@B�8����ؘ�� �Ҫ�OA�d��Gۑ:}-�TH�xg�'���4s�P[ٺ� �A�pNkFG��r]
lI+�.%�Nڋ9-��0?����b�qA�6O\1W�ǝ6�?�I]\GS^\�=�C���붯�kV�e��~s����9��	��°�>ɵ��z�c|�d�ͨ|�mq�42?^�������y��CQ�AB�3�_��@�%boHN.�s8���K�;�Jv��1�D5 �ϣ���*�#C�K�A�xjf�:p̿\��&q���I}b�N����^F��%�{��7y{rl�1�Ђr�?!3C�>s��C�H~��./��'����W׏�=�D�{U�%'s���_ݠ�G|� h��)%��Wf����R��-�r;�� ��w����h�jl�A�y�{Z��qxy�56z֋׋�ԉ+J*I�Vɶq"M�oZݫޤ�H�[+���q8\AU)�?8@./���.�����r�����Nx��ʹ�m��[����b�]Q�达������� Yy���qiII�Є�[G��q7_��V^Vv$��B�3ŉ&u%�ڵ#J�)�|�T~��|�qϻ�e�q��b�%U�Oi$SQ��Rn��;��q�%.`�9}�����\uf��E��5]8g8��d�:t�F[<���חW�Z���=7�Ge8�S�[(
!���=`�$>Ϣ��ל�ٲ\���)�{n��oӠ���ZgISX9qe��6���	&G-�q\7���J���&���=!����J?b�K�?�����U#>r�>#}��~'�cF��b�)2~����Nϧ�L����ŹYϪ�W#	�'5��!�%��&�Q
��4��n��V��U6�R��j]B�;WZ+�+xK���z蛡��m�=�>���
]M/��]�կQ���rtl��MR�B�7����c��Ҷ�We�rrN}�T��p��bO[����tBθ�r#�h�
���n���
��ۛ[�d��A_�@�ȥ|O��M糈�|G�ߊ�)��lV� SF��mkC|��@�:����(A~1#**T�Z�4ހ�6�j)��%��}� �@�O+0ݾZO~�02	�����z���Ah�Pɢi�)�S\�F�/� ����m����?�P���q�-��*����^T�3���8p�E�л��ZL0�b�<�I�+A�����5��@~q�>N��:(T����@�Mه^�E��Eѭ~&�k��|Ѳ5���� u7�����.0�N���BQ����O��h}\_ �5�4J�oX�G�m���l�C�i߽��X�\*Ұ"��V�TTTI%*|TT�5�3Ӕ��Յtl�t���;<^BJJJNN��"//?.���CFyII�=6�yk�-�7*,���@���6��WS?)�Kk$�k�]R��t�hʉN)r�'�V�UB[ &Y�����~� �pmn�v.�e��*�����2��{��nE㑵��郁��5����)M)uI� �!,�-l���r�i�Dw�55�q?�F��m�&m↪��~�-�J�=A�MS��W���&B(� ��l�4�ꢐ���$a�K@
@��7�I6���}u�^�R<Ć>Y�Ge�M�	>�iw��T����,�&呖��C^>_�䂏�M+A�'��6��s��;B���ۊt�.ILiN!�6zc��t��X�AZ]4�|U���t]�:S�x���i'J��Rτ�@�8;슻�F�8��NV�|;��Ӗ�+�p�c��h�k�P�^�,m��u4��u2R�T�w��4��1q������D�S���BW��[	�$7X���
���D;K�*�#|�a�;'�Ά%絋c��k�m��r�>�ps�4�ݢi�)�����G��0�f��t�|@LT<�ѵ��E"\t]C�b�o0��Ds|{4;a�X��ۥ��/��������Ѧ*�dYL�N6Uz$\z���V2mb�{��^�L�Ĺ���>��'7�w�c�5z+흉�p&�@��[}�Z<�^�X�́�ǚ��(�p�;�$ɐ0�Œ�z�Ƕ���O�=X�����������0Okh��K�p���m���tS!r��N$�?^b+gnH�%��9�ؤ�0�1o .ʻ���j�����K+��9_�[h�\())MJt��1�i,"��T#'Nl\ݢ�NB�A����;%��|y�Ѓ���@��$8�,tV3d!���*5��G%g�$���LI�B.9��`�� S&�u��y�A��We���ބw_D>~��\"լ�(#�ו�f�����\�q`� '3;K!/G)��Lj�8h�T�]{��oy�+��JA+�n(	bC�(6� �m8n�A\�A��f#:+%o�4O�Ǵ^��.�
�,�e�i��,+�� ���O��rs��9;jS��-�<��ܷ�C$e�g��c_Td��YW��o����p�EJ�vA�^��G��A�f+6^\�Ƶ�}����on �8���x�4��TBG��]n�tяg~7 j�j�]i�Y
���7;kn�&+�;�|��Wfٚ���S|���H��)D_���fm�.�I��YM�|+fvnhrM�A�l◜�h{��7����:a��w�n-.�d/���S���'ݹ1�ky!6Ԡ�=��K�ԝ#�e,���T_�1 �U���k&�y�ޭ.�R���"�z5��
��?������ŽhZ̒����7��̫�D�J�V�y�����t@���й�j-��L�Jl�%5�-��)8S��؈^"dwM[���A&&~P_�YS�����z�	_*J>x����X���C�%�)�'�g�]x�n����%+�q|V���v�c$��M���}qi9%��<sL�y%˚P�eS;d)F;�7��o��פO{@֦f���E�\�şh�"�Z��q����p�ٻ����
����ׇc��0�o�ۊ$4����n����e��X���v��_L�|��r�b�2Gl��Ԣ�[Z� [Q��[����%�q���}[�2H*��m��9���[�BC������D�����w�&���5ׅ���W�}K����4/N`�M&Wz��:��GBz)�bb�R%L]CU�����Ғ�+�t�	�����c���C�Yn�č>a���fb#'��I���2�?i��t�T�i�ePO���YP�DKFJ���S3���}�晊X h�&�F"�6�}���?(�:�M��I���c�-/�U��T�����e�5���y���.��}�C	�$�+�=ᐒHX�ȏ֓��,m��� ��F�:]C��$����.0fS�m_�.��n�������v3���Vr��۴~V�����GN$�e���:<P1lq�x�!����їJ�HڿtJ��듽d�Κ�]K�d�^����p��k%��Awt�����0kG|,�(����t4��u���{���Re��ml	�o�,�$,�8�^G�V�뙬�����ϙu�\�k`Y֥L�j����ă_9"�S*�|b�s�p��(�,�#��"%�z�+t	U�'�Wa���(���x%y�!l#�JCO�_���}��O��r��}�9a��;��2e������i��G�ēݓW�pN�6��ƈ_Ri@�wE�"��o�9몍C�K9�p�AG���k�laLLǩ�����%&�͚"���2��p˰TK�i�^bJ��7̈ٺy�I��-Å����:��?��|�*����ӎ^v�r��#�xu���1�ơ�MO���R��G����#��mBv����"�CF赋��&��q?��k��u�J=_ ���_@ڽ^��Y��az%��~_��y�o�����ԇ�w7�x�Y�{���=�ܽ��D������,�::���<�+8
J�Q�,��D���J�������1�D�xOK�:����R��q�$�>�D}ĝz��\���pA��XD������5�ɓ�SJ*�&�ׯ_������)CX���*F<�����X|�Rf/1�Þ��A���O�1�VfS�c��S}�)O��z���WđD�����$A
]���BTS&���W�>T���:�6Y�&֠�l��LCff���$�xW�+*Η�T\ �x��>���� ��!Cx��@V"+�qz� �e���z�'�F�6���o<Z������|�-I2[��Fh|�����>{�L�r/̙颫z����B��C�C��O�((}Ȭ\d&�v���w�\^������8:��w��y�L�R�H���݋���.Վ�D�c���L��oջ[�
�ǝz�=����BG`�oǋ3�RI����1�l�o 1i�тZ9��� �S��Z���(<�4���E�R�F{�Z��`g�^��bGF�e��Ih>u@���%�,�N���vL�V�Um���� �|k?gi���c�ƞX�/��KLyQr|��N�������b�w�B�5+:�:����l�K�������Tv���C���E�M�����m���zC�9�C\���v�l���G&��`��nk"R�/��5
��XYװqڢ���YxE`M�����`]��b;��-�؋�uRZ�O*:�S�@9�Foە{�ћ'O5m������i>v�=r�;��:�,�H>�@���F��*��<��+'��ԑ��.�u��<�P>�d�D><�͓��9���w����o��\����~��B�R��x;����eu��7���k5��_
A� DLHSHU\��>ȯ���6���5H�7մIɍdZ{~�Ą��ɏ���C�ǽ4[��鱯��0�<��E#7��>��u�k8\�3y~?>>VfX�&��kѫad�St��� wqq��T���j�dWvF���uy�[`[��_����K���1�)�Q��K��oͅ��16��L���SR��l�6�đ/"#�X�۷�m���\0|�_�qo�;Oֲ�E��1d��r�J#MLfV�
���hN�Y�H]$(M�"��c��y�n濧�#�	O�7� 9��y;��q&m� n�Y!ȿ��j�l�Vȹ�Ɵ+�%E9�w�渺4v�D��$8r�-H:�T��ly�L����'��blq����Ʒ�Q/M�Z6H�
p�`���߇i�֐��������h����ӟ�o���l�8	��&�9S4����0 {�$�-i�ܛ�߹2y�_(��WGWE�,b���I�3@��Z��7�^����
�����g�P|�(�4��RY��`�g"µ�~	$���U�]�Sa�7��|�'���v|���4_�?�q��T҅*<`���-N����P���ǒ�ʍ7\V]�0J�@�DK1���e.��K˚�{SkJ�����F��L���O��&��ZqhJ�����F�8�����LKy3�Fـ���߮��F��Nl�n��sۊfv����9ܻ�'�3��Ό��D�e��5�[�2F�ih�TrNX��3�+���i^�����b,�Wә�\,_"ui�c^\u�����.��6�T�xQ�Y��/�92��+��5#��_b�p[|1�@(����GHm�9��ة�',�n�����c�,�0%N5�L��%'�c�
0�Y�����I���A���8�D&66VS��tg��p�!@ev�5*"�en�I��+��[V5�j0�rmU��5��o�=���j�n�6Q�[h�����t���Y��4��:!%�Z:!uL�deu�X"�Qyl���l��W�Pno �nХI@�C��:t�3�~��R��K�`�S|v�����^�="#*<�p���YJ��W+�'�G����o�v7A>5��wұ�\W�ur�1�m�Q@#roџ��x�crsUF���G��җ���z�����֗��Za�����#kVa��>���V���)�jD�A�/��)&އ���ZM����N��8����x�����_�T�(�֫�a��|�a�Ac�u\!`���Cg,@fw�a|O����l�3:���U��G~jO� C�w|x�W1��|�-eK�ny8_"&<������S"�?����N��$D,�:v�8K���fF������k�qw�5�6�@�OjE�dk	���	���Xz��&�^�L�t�^�ҳ�+ýki��v7%2[����k'��q�W�=�X�J���>q�X��`n��ď�{5�x�7dM3�0�?z�H%�%w^����;���G��i����,h�b2���(ɸϥ���:y-I��)��m�'�Ā�=�O�w�-����ok`�&���H���TA��"�S�(_�F14��m��r��.�̵�_e 7��1	&��2�\)I(��Q-=A�=�������k,Wخ:ː���Pώ�7��#y����Xn�4��o��e�N6B�苄���l	��+s�}gK���-��|�*��׷�:�7��O���7�A1����1��6�'�c]�bGa��)�s
3D����ۢ�����D!�'�&u�:΂���;~����"�U�������/���G�Z�Jvv�B��Ҟ�삡�]sPGNg�½�X賑B5��CNqׁ�#���z���$�Ջߵ_Q�;�M���zO��Ň3��%���OF�>忏�%NĪ�e����$z�:Х"��=���o��z�Z@y�d��:v���U���,�&s?�q-�{<\���b�{l���k��U��)/�|*2o=�U�wH�(�K����O��y�9R+�zɒ�ѵ0���A-�����,�s���*��Q:�=��?�~j�����sY-խ�8�_�ӓ��ݲƼ��E-����^8C-�C]L�EɈ���yM�^|h�E���9^�Hte-e�ה�G���?O_��BTu�͕+̄�T}�l[�ʾ�'�(zǽ[3\ ��F�R��D�γ�բ�I�I�N)М�!��fb�))�QB��.ս:�(����5W��))L1_s���22F�)���p�,�$Gd'𞰯mzzy�{���ױΉ:o
���}f�)����;鉮��Pؾ͙�@�d[=���6�ν`�Ur0lp���}\RB<7���M���
�[2�;�g,;���d>�[�ɖd�6q����gnc���;X����~�Y�V5���5�ʣ�k�E�G������DMUǼE�D�nu��s����s�5Gб1��m��#sr�挘"��)�,m�$k����C��"��u-y�0�H�-|��f�ck�!����-���T��%��������� �XfK3��|z �P���-��G��{��8�Z��ԗ�,�a��	I����Z�їpĹ�9�����S����)�OJ��eݹe�qY��z
��!ϔ6���G�N�s�$�~)<{��GG�狖�a#�=��_�6�	>��?�b��J(o�V+A�Y,�٤���w�R<���:���p�۷\WOV����֎�oGJn]�`%tӠ�ْK�x�7ƾ���O+����=�n)s���6{<� �����uq�Q���1����е�6�����S�>ܧ�Ɋ�g�|�>�s��i,�;�É�}/}�s��9-!b�{��"0<TN|�i�0YU��C��&�4b�o7�z���4���Nf�S�4�r�{�-���,Ps��e��R$��\�pR��P�בt%	����[a�N7N�Ώ&Q>63AU�'��P��[������PX����,DQM<�@�������L��c��<s=YM��4�ۈ�R;�8;2�.b�	݉��+��@/�몳Er��r�ku!�b�i����Lj�ܸz7?pZҸ�H�y��?.�:�i�N��UD�9�rL�=ᢴ�t~���<�g3&�f��i�?ݭB�؀��R�b��Ԧ2P<TS���f���㸩h�o��bK�Ta���0�6Ad?e>�y�!�ܟ*�l>�1Ͻ�RG��g�W_�C�R�Z[�P���v��6À�'����p�%�'����9Ie��`r�ܧ�ro=qW�ϕo��������&·�\}F\;F3�M�9�)��ng��{a��>�`�7p��rv[�ф��o������?h����Ѽ90�z>��xGN��}�U0W|��!�:u^5��ćnQ/"���}��*Dj�ڰ�X+\�`�����kA��6q�����aki�9GF��Ol=C<��ـ�?����7�?x��<��6���#�̈���*���0���3�P�Nva�vs(�������4�}
���d���(��K���y�x�;��~K^pr3d��J�ѿ]9S��]���%:U���E���H�e�[^���(��S�q�0q�N��<8_ ���P��9b� �`�m�����A��j�C-��B:����R�
�S�i��@�y��!u�UĵF��?QX���jyT%Ns������G�7��M�z�:h���ĭyA9�}2k���ȣ"A`�f����8cU%j���}�]���N}���P������"�r�̩�a��~�+Gy�Ƴ+��b����̷P�=�p�\�g`����p���A�:�;#�����Ʊ�܄&B�m�� � �:q�������6�;�B�Er	�KIW2E���LQ�j��|`hRc%����rf�]]A2��
ӦM��~�ln��&U0+$q����9+����q�$���C%�O^�
6�6��1�E��G���[�3ǻj��>��s��ه�4,ȹ�o��.��8��NL|v����-��sx�s?��Gzg�ɉ��S7d�W�1�J"��q�$)���t�C\��<�NSB��,�t��J~�~��s�������S�:]p@�؀#RPHb=���Ec(�ٳ(�!��ӓ�`�����['�g��)Y�+�Mu��$Ԓ��3`�Y�uw�.���#^K�Z#XR'�bkjm���Z�B6i�kHۨ.�����đ��'��m�:���K~� ��㢒�����Ѽ�����T�8�	�#�*/�s;kZT���u���Eq��I$m�f��p�8��PK�c�h�_͌XR���ʺ ���ޢ��dt���cf�5`�l�v�	�ө���
':}h��_x��K��Y��AQĥ-cbP��U��p�Đˡ�;����I}f�i0gf;�{���F<��ӎI �}���wrA5��wو�(9�A��Ƈ��gn� �g��v���6��<Vś���!������(���������f~���Ԛ�����,�V�	*G�gX�Y�|������3؉�Z�!�� ?��޿�ш6�ά�Hy/���d���������/z}�7��e�`���������WF�O6�(��p�9�t1�cE���
 ��ޛϲ�ưgl1���^��7�q�G����H�Y��!�_	�𘥶;%[�\�Z��$�?5�$YhJ�Z������j�ʿ�b��*"��߿7��%�[L�8�ly_9p��u�I��k����ˊ�� ��7�@����ғD�Ly���5��Ƶ�;�t���!��V��R�c!��,1��$�� �':�{=bf^�<�,�T̞��f*d�"RƘ��i�a�@1�Gѯא���\�L �ʱY9߷�D��x����*��ڬ���c�v�᠐^֯�����)%��8Aq�	�|/nc�������.���Z�����3��iY~Q���(n��֒�MA+)+%��"��!a��y+~����Z#��]]e�;�ȭ{�o�̟��1)i��e�?ҥZ�F���h�}� -����ű$k�$:��k�tdEeb�m�"�	�k�����>��8��ݻh*���CC�$����C��r[Sd?�̡'�lC��h�QV�ny��������W'�N^�ȧ���D�߆'N��Lb�V��3L��hG)wqK����?��O�˷�u���ii~`X��������\�i馛3WS��c=��E��'`*�y�Q��B�`M�x�3�-��g��J���ʋ�❧�_5�D������;Z��o�&���R�}(�\��.v7d1Ep �dD��:�)٭nC��;Sp�+�H������E ��k,eE����C����<Tb��o��g�<WdU�&�*�+��ƂaAeE�X�h�d'	�qH\x��-����E�����j�}��K�Kq�@�����]��ŵP�݃C���Bq��V�/~���u�|de�a&���7ϳ7Y $fď��hk�VP�<���Xc��%��]�B�T��sJr�V7'���}�6{ͫwm(9D�r�xHд�o��٧��',�����j1������(_��c�&<�4j�R
�}(��p�.:;m���Ul�&.¿��f���Y��	��N��+��+�F.8�ԃ����=ѺD�$�ڕJP�hu�z��S� {��;�+X�V���>��B���<f�:V�F����O�Ƴy_�o^װ4CH�w¥D��e�)�֚��֏.��s�꡵�B����QE�LM��ì�t�G���108���,D."&�|}��rN��̳��<�����߽~�:TVJJZ��J=~~~~o�l��o>�-��թ�ד����_����壅���x)3$�b~/�/�|�Ǎ{N6( �.��jb��\��Pu��s[��H�#t)�! ڱ�X�K�cS���i�g>O�\	)<|�QK��)�X���>ڒN�y)\2zER3� RE�7�l�.�5I�`':ye�OJ�(����._���	=��GU�#6Q἖�M�n*z���}6�zo��Z��5w��PE������i�0���G�볜��������sn�K��0'^�6�訪�^F�}��Ժ�Z�dt���Vߙ�[9�,�큪�F�p�kd�lq�� 0�y=BY��*!<]8H����T����yz)�L�7�W8K�� �����0%I� >�&|��� ,o������	�X܎���qW��D�av��Ұ�> �N����0j���2	M�"7�ߙ���5vXf��  �И|NP��|��M�J�?��l�akr
(v�V�p='A�C��>��'�!6�2����[��/�≹�c��_v{���Pt��$�(��1��Z*j��s4c�n�_I)���N;{���� ٝ���2���5ʎko��>$��N�T������}��7��fa'�:������rTI.6��p/������
J��6�98�{��f��-=V�I�"y�h��v�nZ��
`ۢH�u��I�H�91Ӌn��t}�ԀوMAx����} �{�̒��N�J�ݞ7� D])��}�q!B��]���܄�����|a��L0�\M�N�uP��A�Ur5�X8�J�]sb�����jG���0���1���p䠟Q��s�b�kF��8c����<Y�ޥZ|�8��s@D�s>�ϛ�oy[��~���%�����I�Z�`���g�/I��K��l���@�`P9��g;M6OD�}O{���fƏ��Ҿs�����_��oC��K�wR���!���h�!6�\�a����3b�0M?�컍9�|u�\�~��{��,#$$dkk+;�by����=/5� �05����A�U����Z�J��P����~E�P���Zi馐,��͌��n�^���L;o��W����	Լ��{&~����Ppl��w������B����6�dM|u\��u�ſg�mB�X*���F��O�5���I �H�?�.`9s5������X�YC��K���R��s�:�VL�yWWwp�D	��ר��P� �\���(��6��%s��F���ǅ��ƅ�'��/,)��1��(�@E2���UQC�1]@�b��榠�}��f�ϟ}��d����4�����4	%KY0q��6���W��$���Cp=u�t&�{����������ܯ����Gۥp�_N�ICf+�{��>O��E���k����W��]X�ݗ����.�S���J3��AВ�C����?�[2�3�=�?%��fn�޾]�]���h�^��Ծ�:��0�499mW�Z~d�y��h��ũw[tWi(F�E#	��p���?���@z粈Vl��� �c1�M���U~~�u�X��,F��mW놴�d�xv'd�w���/�h��q���+8觎H��sX ф�v�R��a84s�P�;�̠zT*�����b�!��0Biu{[		��U���c%���R����GkK��.�|וS�
ܛV��7N�H��C�� ���K(Ve�os�&�*[��A�X����L̑Z��0��ю��
���[N�B'ciL$�����;�o��σ/)� �W�.��Uɇ*P�z&�IG�@#H�
��W���D�J����'+_�/W����|gku7E���V�w�@Η]/��C d�"3m�\G��k�����"�ރ+\\�ة�%�f���(�Ϫ��a�K�ة_���"���c��\��^v?��_<l���L ���|��w����"�A%�*��D�VRK��n���b}[&
�[�03�TJ�(�7^l\%!	?�YTnN�wh_�3]W��p���b�)�e����φ<��wyG�����=�{:����p�y~V��i'?��iH������S8uGـ�����:V��Q��VFVV�$����e��&K�R��K��,[�����Q�1���n��Q��������iz6��\�/�ב}=+�;�N����E�#4e�/�j��&o��q^Ff>��2J|F���(�:r�L���/���n��34
2D�����s '�̕��Ӫ�R�H�eΊz�0V��/w4���F��}\^Ji����i�
�GdX�U?AO��nb�9���#��.ټ����ܻ��ǭ��Mћdћ�p���x����/�-�&^�Ħ~�^�T�� K���mM����WW����͵&	����ʂ**
���b�Sh,��ݰx�4���s�k��l��R��/�}�唻�/w\U����gI#�K
�T��x���Z�����S���a����v�p�
XV��ف���
9	�.F� �"1�s�z�)1�d;���[���1��9[/�'7/Uwu$Yvu2eg�E�zOF���SO���j�nh"㔏��[�E�zbi����ɶ����8r��^�U�v_oByeS�Xq���ҝ���2nEl-aʅ�S����(��ѿ��b�%��*�^�2�j_����i��ҝ�^p	�]��&[���u�Ր&h�Pg������ıw����v��#�V�f�n�i����o�|3��L.���נ�P-��%��
�����.D�cexx���J��*�5NU���Tv(������Ə�$O)}��W���t��˴�^�~�]�H�i��~dā5�W�9��Hf�	7]1���� �5�/!�d�Z`=��{<�!�kK7����WfxjK���-���a�����ѹ�|��ڜٓ��2;=�E.o�-Y���m�UXnƾ������@v%5����b ����c��2��j�!=��B�¯�����DV��,u8ی�->.ĹWs��9�\ԍ!ӢV��R���o�%�iAj&��쫭�	��������4}mM�ճB��R�*��|�z~g����I��'�3�.�z�2�������%e�)�&�S3<W��hl�p/-' ��1(������/{���l�����;���c9�_�����~���� :���Q��3h�����JYή���׶����er}�����S�f����4M�n����(#{�����ܻ}����:��h\$z�x�vkW�N��1]��Ow���"�i��e�'�r���򣡛�d�7�+�V�vV�ޤ��0t���f��-���](�V�vʎ�.Q*�і5��]�]8_�k=9��*1Axv��)��e��DnRҋ��b�~�]]��'���|�Y��PT���$ȿ�����	1?�R�7��[�����/~m}��.[撹�-6"���_H|��)n�dso����#�H����:�x���g��T��h)�i��~=_�����NE)&�il���Ç��e坖.VU���6��-�4OK�9�R�
�rfh���*�*�r�;/vs@�u���8�
aw �}�l�_{�C$�f��(uj4����/�@q�y���l����&]��
���ۮ\;�k
[���T5�`�9RX��+2�����7�a�M�'6ӗ�1y[|� ՍMM��fX��8��֍��4��e�L)x_��$��M_���jR7����ub*@_@�4��P��Ұ�>|���L�
�C��6�L�i�״�����S����<�(��Ys�:����G�I ����q�r�0��^��^�� :��d��gU0�����X�q�/L?��YPn,Ҽ��c G�n��q'����r�JOz��UP�h:�{����Q%�C �v�4go�h� 8�H���#٦�Ql`������Gʩ��(�tѥ#����'�U�c���hp�֬��e0����}�-�JGJ�¸�_���1��%]�6������σ�1��K9C"���,�z���s���fs�D��V�޵����V<��u�k�s�Y�n��ؾ�U��8����,"S�Ʒ���:j�����%�l͆�~!em���+ު�X��R��uk��t�h����ޤm� �J�B�M���WG�\�|l��r�e�u�u0�4�a�̍��֡����eo���R�nE�a��q�N�a��g�Z��K�8[��W� xK�GF���f��g�a��9ssn�b�g�<��v%f��t���L�Oc����s���˭�մ'���O����������f����+w
8�]��Um�vث�xʡ��ps�t�;�~?��w5����:�[NT�l�~�#�j��J�C@�B�M��Ԧ�vJ�kM����%�UW7HIO���!^}�z��lRNY)��-^�.F�[Mϲd��V#4EQ�LIH�yI8���Б;b^~P����������{�ѽuj,�ۍ�ܻy�\ ��ރr���&OR��A?�AE� Y(G��O,��ps�^$����n|�������������s
)EV�n6P7�T���K�)�St� � ?�[L�pEGis�e���@�����Q�M���U���*�X���\�bFk��1�(��ɭh��x%�񠃽�a�+�e y@�ԛ
���n�!��u>�C��B)�~���p��N3|�1[���`��8�W�u�}֣��� �-i*��f���rX2qX����Ƒ���ծ��3W�M����+��0-��Z��eEz��9���Ҳ�\���	���t���"?_��"u���^)�����k�v$�@p�s�o�_Tu��l��f�\),�IԫC8ш>_���<�!aQ4��:!��fAX�=�/�c���B�O�I|F��!���p�{���H�q�M�$c������a�-վ�$)+�M�#�.�ߜ�1��DL�+�{܏�ĸAj5R��i���1��B�#��7�y[����Z
[T_�"1�Y����Ʒ��Q���QGly3�W�A�G+��=?�Tȍ����I���g�ps%�P��A0��{�P�^+������}�a�R�=��	�٣����X�&\<"�rX�X	=��1<#�GY��$�´���dp��
`^ߘ��q�A�Y�z�m�m���[[;��l-N��c�����پ��O�I@t�x�,F���9�+��ݷ`z�p+x�~=���.1ק��V�����G&=v��B��!��z��'ʐA����T��c��yU9��1�]H�׶-�v]y_por�"��D��OQ�*�p�\{�Y�[����]��*�T=�5!�_��8��Rq��Vs57,�mD/)�:�����5��W���O{�n�H1�>�/����ݢ/�~���m/�(9�y���ƶ�\f{��U�.IUb+ga�S����0���☜/#ۅ��~}^�O��:m��\�a@�.N�9��-�(I}T��W�P���*���0g����f{\񍟋ɞHɴ�e}������s��"���Ju�����v�C���[�U���(v��\����cS~���=�ꀫ͎۱���'���[�����������u��S7\�l��N>���.*`?ig+}����2����x[���E��V
�� ��5������n[: S���$�/X���y�Ķ�0��i��|��Z9��7����*���}QS���R�C��!!r~��������Ѳ�Zz��jՂO��(�6�}b�<~=	w\�O�O��g�O�gy7e�����.����$)n7E7׻��nnN'�'�d�I9C�\�!�a�@aG�\u"u_�[��Pb�G��XR��,$CO�ak@i\QqP^~H)F5:�6	�J]1�"�H��%��a��<��Q&M��P����T|��I��d�C��u����:O�F��{c	R&>�5X�����g}��b�}+�ݟ㥍���]C����R�2	�D�:[NނO�I�pѰ���
è�q���6��jI�q�^ռ)���m�>o:o��oh5=�ǲ}�#�G�<�� h'3V���h� A����G�շ��v�o��"�����i��S��Xs�0�E7�`3�جNB�-G�6N��m+��:��c�s�t@�;9B�7�'�_�B��j�曽����L�n��w�U]Tb�4�w�F�����D`�<��%�giL���؀Ȁ�1s5���W �| ��g��W��h��ƶat�a|C��-$|�2�v5�0�@q�:��.465\b�y�c��-�i�|y�U�-4�ZU	��[EUv��1E|*!���n��zCnR:�� f�fd����B��Ʌ����&E��J�h�w�0aqkh��cJi �!F*��>��Ky��'\�z�\��,�������z܉��E�������oϛ���ϣ��0]HXM�>"�a�����9�H�����t7I�@�65�ia���l'��f��-S�!���J��FI��2(�g�P�m�Scգ��N���i��h��&�q�H��i����}�.n$�R>E���]Hrg�H�tS�V��� D=ZjX����������#ս �J��꒕c�Ĺ���Goȥw=	 m%��1�!�������`�O��F��m"��#�Y&z��B�|Nߨ;��tiA��}�i�v � ��V��d�DWpw���y}}�ٹ湍r�w Q���C��]	�t��v3��K�l����G�e�7��_�LoWy۱���n[;�.�E֫�d�������߶�>�>nT?+`���x���6���M�X	W�է���.�蝑<u��t��L��\�J�ѓ��c2<����p:(?��s>�*QH��_{آ��LH�a�yS�������	���o��O֖ sj�i�oN��	��8۝4�n��2o����{�Բ�l�����~�O6[X���.��'-��<��C��+��ke�>�x���DjS����\��^bSn� ���_*I�8�vmE�R�ū�蔣���6"����a�)�=�?{p[��o�H�g���  �� �Ë19峒?!H	@_�͝}z��?Q
!p�
s V\��sa�qL�­&��+�.�v�> L<��G  �pH�ѐ<����C�rn�!�;ߠ%7{C���,�n.7���*�z��]B%V�8z�v�x�<g��'@����p��3w�ޛ����gR�}�sdD谖�)���a&t�ϴ����>�6�h�%�.s�H *L��`J�?Ǌ	��GT�T6��މ�|y�"��;���y8`ߌ�և'��֛R"�r�P82��u����\��Kh�zٙI#�fr�U#�*=�+���}\�Z��%
�=,P�c�uQ��oM>O�������I��	ŷTcU�WX�LmXJfI��<�ݑF=I�@rw�4bIG|�gn��b�ߓ��&N�B�~5-�<ت
n~��֣ݒN��p;���u�aƅ���ˑ��J�[P�����+hiP��b�jd]�)˜���VL�Pi����uax�U>T�W:��\�5��j}�w��<�}��N���p�{.-��:�Le��h�&^<J�q22:�d^k�Cp�!Y��[؞���{�@-�!�����V�r�x�*?��0��e�̫R}x[X��9ݶ�}8^�!�.<�~��i<�6��{��M��\��ϭ��s�е,;ua��٨J�n���(�Y�"k���K�o�AD4\��tN*�����9�O���2�õ�G����!����xxx$$e"/B����M�bd�.�����}PP�����f����9S��X�@�,�ͥÒ�d>�����I�u�g�j�vi���
���X��*/�*|��,��n�"�d!-�F����6�������N:�Z��KM�D��t<�P�?!�ie���)�49�iƳ�n7�*���r���G5�����ıqc�kf�giwgG}yw�u��=�V���6��0�pz����*����4+�e���0J��j��
�FSb�b��R��|^�EFL68'�B`:������CFL��H���?e��G�\Y"~���ۓ؃�Djl
���Ԓ���wǆ�<����,))�����ok��F�E���;.|�v�z_�����������A-��n�u�]�a�,���w���:=ͅ��-�����a`��<�;&<�-���h�\X����KL�+��y��K{7�sYp�\~��|���
��ip�(����W�W�Ws�w)v�[�� ;�4$��B�y���^Z��x�c�9ce��ʛ���k�V/��jכ�aX1j��
����cS����-vk�;����+�0X�ˆ�-z
�*��A؆<B�&O�{ǩ�BZ�_��F��D3.&�5Z�Cz�,�1$���#Ε�J�����(���X�����ffݩf22�-��I��q	/�)�]؃?6��b6����	�(���/�k���\_`]}���&�er.ƌ��#���]���O7Zj�4 ��-�e�ʮk��P� ;59 ��{���T�XAt��Ĭ���*�,A�>�[|���C�7�sG�O�&��	)I5D�O���avf?$�MUnt�?��ZK:�9)�TY�'ɢ=9x�X���F�%8��]cl���ƞ	��O5Rnd {i�v\����6R$zI��A5x�+�U�Qơ�_0]�`�kit�W7ߔ��:5�$�CQ��\R[��;f�5��ݎ�N��k�ƥx�3�h-�6h�p�c�B��J�`��~��"�a�&�5am;i��y��Nt�DM����˖r�S:�v�����T��`�Q���F�W��=�3�����~����Xzw���,����eI�����������K̷L�[,�Fr����vK�Ή*gr��������}@-9������*KH���7
Ր}'?���� �:���TL^'�v��o_Z��s?\/���n�=T�j��,���;ݟ9�?�w�+x8/x�'��tv�������{�����4p�����t� ������S��7��_5�}Tq��D��֮�ˉ�25�=����������z��,a����(�����}f��}o��Z"w-�Q�-x��*�,&��	�j9��p��ϲ��=L���pJ�<�Ϗ�`�Iݼ ���?��g�͝
 =c����\F��x
�lgLswL_��v{���z$[��O6�k��Ou��;�[[3�N��o�ٛbS�S�3r�m�� p�T���h�x�c���J;�7)�>�vV;��Wb�r�J���/����
`<�
�K��Y�˖�B8;o��A�$���d�.��j��'�;�t�12&�� ��TxDQĕ,��7�ǡ����!��DRE#x�2.�s���z�Uw��[h����/%�Ғh�δ�������[��xE�g?���b�k�J��}��c��������wӖUG3�5_�N�������-�������묜����N��R�PP�[=䂸w$Fզ���2���o�pS���#K��Ai�BДq0L<ɈV퍤o��;��%g���f�	���k�d��*�#!,'��b�7��]�r�i�7�g{Ϥdbo�p���OfZZ8��(���@3�zI����$c0	�x޾� �xI��P�a�#�i�yy"�N%�f����L�L�ń;�Ҿ0z7	���$L˿�W���&�OF�C�8M�ȫ�<����/��������1!�e�JRvǡ��[�ü���AWH|�'��D]%��K]��-@L@mX�y�0���\*/\E>z¯#�a)�l���Sz��,C����l⫷,G��G���

��\d�F��bϡgDNڅ����׸��� ��*�3�}�z��g���0]� aR��h��H��p���O���7Z����D(�K{���?���H�x�I��.�hU>}~��W���r�M�gC�Yd;ό�FJJ�_Q�T%.�J�#2Y�T)���5����6P�y+�xk��є��g!H�@�y���M�"�g��{~k��l�p��֊��v�����c����I��ꎻ������kӟyO��v�D�gq|7��5�"t���(�nt��6��f;����~K��aLW�o�޳�ڤuq����b�=�zf�9Ob��)����J�Zxş�\�93�>�`�_/���B4�mg7�v���H+$>lʫ(�e��J��O�(T���|�	�Cx�=�I� �*��^�Wŧ�3W���F�ީF����Cʍd�~�
|���6n�^Rb�EXo=�E/j5D��tR .r��:.�$��'*S��o~�\R@!r�<��%�?��C^�l����J������/��a��;���������D<�ća�v5�5r ;4~̐_�n��h(ja+B)��f����;���8�0��⫈	��19K�z�j�cn x^��VU�&B�������ۇ��*�*�l_�������\��\�y��槝��<�[r�JV��Nҳ�]@IrCe�0Gc�_�����/v��p8�R�~��,}𝆥^��W�?.�~؋7�Top��H��r��"!�J�\$k�Fn0T���U�
(��icv~��έ.b[��Kl�^J�Ey�S/
%_,:�U��|�X�܄N�^S�'����[��%2)J�|���C&��	�iL[���@��@8��oR���v�V�uzrpQ��&$(���	F�����v�5��UEP�אWje�F8iC ׇl�Cb\���HJq��;;I߽zP������l���@4��{��'��ޤ�-B�"�kM"K��F�1hǺ�-S������I��
�|pX:J�m9��<@Y�2�Z�cb����E滂��@iXj�cu���t�`y@V�[f�x�U�. k�����m#���
y����7�8q���Ok���scv@����L����������%G�0���{�U��d�[����㴚�^�u��!�`�-�dA$�W*�CV;�J����%�XV�r�03�{��ώ2�fC��,�b+A��o��vI�L2��ه��)8�c��.V�H�Cu����#Y���m��'?v~W�����<���_,�>���<m��؈>�U�_����Ą}���vz��~����sg��I	z��
��\�?2�ߔ8���7e��s�s��é�������J���*}�rk�U���X՗���i�4;n���¨;���8�{�T����֚Eǂ�m1[W�9�� ��K�q���Ʋ��-8M	A�i�r�t�lj(������oEǉ��ui�G(�u1-��������C��U��\�����,�����}�b:k�����z��*L��sA�::���%��_���1�	;N�z�+X&�৽�I�7d<]uާ��_��vz҉rq	�@,�a��Q�,C�F�7��8��A� �1���m�anV-k� ���(l��.��P�:��(��F���[��"�sfcD����q����\����h��t~W^��X!	2n�'��9��/��_�/�TNy����s9;\L�������+�,�/��Y�c^�����Dm���|s�b�WV�"�U���ϗ�۠�Vf�֚�a�E ��%�~�I�@�^v���e��x���;C������x:�2s���ef��8}Y�&S'���K\qhX�G�����\����U-^A�
��{��\�ǉЛ�+���#�s���G�k�vrˁQhѾ~v|Tv	����3C��wv���4q!-��I�,A�&��R��9�rq:#;��U���[�ȯ���3��6�gq���
���a��Sq�.��e/����`���Gm����؊����*�yI8��\�� ͒eb3W3�Y+�'��ӗ�&�x�엷��S���Т���%���K��	0>-��Ɩ:��`��H|S"p�"?*B��.��l�Հ�u���7uK��d�~�֚1s&���e�h�x��7t�(������w��[g��%��K
���H�ӵ���z�b�$��u%�RK��fa�6��N��2�H�0��] �J�jG�Z �K��ơc*FFv�5�3Y�M�-d�ԏa��6)l���1Gd�+M�#�+�6�&��ס�~�����O;��WM����g�k�g�*�k$�?P�nF)��.�:�Z)��ݙ���\�6��$³����K��m�G>��h����0ȏ�pY��S�X�+���ϓ� ��*$��Y�>�#��BO�� n׷�_m5G�RR!=>���]Ga`��y(��1����M߱rg�µ�����f�F����|j��nn���w�r��^D���8�
9�����-//OLL ~G±�]_����#����.� ��bQ=RV�����n+h��vg�\�j��i2�{�$�/䟕 �3[f3+4R�؆�1VU"�3=�`u*�g*X J�-f������~L�=�V�7�f��8��M��7�Ȑ*�����W�`���4���|�~��sx�f�*k������4 �xA;Q���I��K>�26�UW�"�;�q9�0�"�;2c��%�������T��,[���L�p���,�.J�t$N����r�2���&�4�<ڴ�9%fg=�ʳ'+��ڥF��oT�����
'd R�Č#1�ͨ�zޣ0Q�=��q;_��,J���V�Ɂ�/��+��&)�)�_Ӄ��#�Ps�h_rD[^ ���R�aT��s'x3d��1R�S}e9"GE�^r/�ꜵ����^�낗��'��G�n�Y�▩�R���H��K<h����S��=,������H;p4�R�Z��g>4���]���X�aY�%xjD*�)u�j�]%vQ�k(���/?��c�+ o[��xe�p��ߨj�B.�y�Õ�T�~����
�^�f��
o�/u�䙩�.�#t�c���XO�����M.e����d$a�sWc����x���
؂:#4,�/�NIC�:�[R�5r�1M���od�=@�J۪��d�5�6Qϸ�N��{Jaxia7��!D+"���������h�\�m�I�j���J���7�-{���r�7|�|�>�f\y�a�p�n���q����:�.�W��<U��):�o��nÛ����=�_<^��ߝ��O��=�>�A��u�����u
x���1��f���,�:���T�3E+?]5��v����/c��j���O��t�uMz���D*zI�67�ΛC�� J}�����N9��ε�ͲE��Hq���{K ���l��w+���a�h�P(����t��L��O�j�ƥ��Z�w��N�������ʻ��K�&�^
a�=?��,��٥�>3QmˇnI�����f�ҝ^b�DH�	P��<������DMTJ������ʈ����qi��~6�[��&�qSz%::��[G%6�l�U���$i�hݯ�FUR0!�D�K��I��],��lJ1V��a���Q+jt���f��D�]4o�3���n	��c��}I�7!�Eidi%��Ce�����t�W�e�<G��q��4;'��c�e3�y�m�}{6���)���=����c	u�Y�� �@����K,�4��j"6�f�`�rv�wwqa��^ ;J'j�'�8)5��mj麝���#7�-x ب(���s͞�Q3���
�}k�AvP}3.i������Je�d$G���p
\�=���@��AZ��x�c��W9L1T�o���!H�1ZU6�b_�k��
���z�&)7�P�qO'�Xa��?��QW�f|����:���4�RԠ�U�Z�o��B��D�8�.�P��Y�6z���&��m���{vI��!�U��<�[l�$H�����
R����m�:�\�"�H7���^��ܜ�^J3���]oώc���gR�~E�ʦ�TpS�I�OҞwc��s�0�o=1�DgS?J�J��p�d<�.e�$w�e��N�(y��c���T�'Tӣ�ue�K�nО��2"S�cy����6�|�XF����5�-��M��CO�B�s�}�衰�hM�s�d�Բ��o����+`"�[�:�Ly?��G,8���>�������T�{d󬓜�|���_�a,�aS� 3jYΎ��>�;J��/��X�mg��jt!��M�s;F�;��^ξ����)�x�#�V�?]q�T%e�*ې|�w�
G"�f	�Mu��;���*��v΃Q�7��u%��%Ļ�.
.���g��u�I���xEE�1 99�}�*�I�z���m��	�ថ昔���
<���5ZM�]&�Z����r�w�^g�f��st�.x��뫟.�:�xE�ݎ?����:y�}�@���Ӄ`�c�P��ӛ���[Yћ�j��r�/���_v�EN�����P����x�P���)��py.�[똓��VPUU�ST���WP�S�c(�ɐ���m�;�x����C����/��~���M	�$ 'p�Y>?o���+�	�+�����賲\��n
���ϟI���x
uDc��}n�!7�WG�a�'��������ث~�}ݭ9G;�ؾ�dNnM&`�����2]V�*㖊�2JaZ��a�zw8���Z���r��b�+�qlR�����7��X��a 2Ώ��m���X ��Xըq���9�-���=�#=C�F.�C?Y%e���ɐ�^8A3#��{À��	F�_ֶ����^�CZ��&T�T���%�+O���mZj,�z�7���&w�����K%�z�_d�2�mzO 95�*�ރw;�bA�F
uv^r ��2��!4�)!�(�Ru�>(�o3�S������>������~$�
pN��
���ت���ש@��CGc0�j܏�l��c��M|�<vRE�Z$�-=��P%h��8M��Ǳ�x}:����q����>{��u%ڳ��.���[ffVWf�*++K닚��<}=umd]e�f��+Y�I˵4\�K1����%��L�}�]c6��E`���JE��qv�r���
���ҕ-����&&����jMД��d��B�z 0�iF"s1*P��f���BMt8����j/�}�Kx�a�p������'��Bw�8~I��lP����$��HH�"т7�?jG0$K@Z#4�os���	Z��V-��W���(eX��& �b������H�YƩ%k��r#��&��߾���;{�
��zn)��_-L r/�+:�Sj�E��v��r
D	�,0����C}`xĬ��le	m�	\��������@@@B��1<5�4�tA���75�(�-�<)	��uCt�4�~'B�"*Y��8�`�/���ţ-j�Z�L-��x%s_㨵��V�1��|]�t߰����wVl#�,i�R�g������ ���&!�����r-�����%���Xx啟S�K�R���&h@��i�F���m.��[�� ����P:V����J%���i���E���;�O������4HvV������a#���vLT!���آv��֣C,�Uwc�G����۹��?�׻�w�N��NO�7Y��>� �%�����WK�w�w�O���{�ٲ��3��ܺ_��r2e�/���\��´�4��y�L�x:�XGTT�`�R`<��ĉ��ԋ��4"x�>==���-t�yv��w.�>i�$�?q�s�d��n����!t�z��L�ϫ_eۆF�Ȋb��`���~�w�=��������pk�܉Um�u-:�?�gYa!>�h�p)�v�\)q//�N۶*���#��.�x�����5�B�C�������<1� =�m^�[E�d �y-	�砃E��YO���~2��=�n��+8W�� p�i!$�2ƟW~t5t0��KM-N�?sm��K@+��lAp���I���<�������ڞ�ɥ�1�Pm@�)�Y]m�WN��Ǐ;�J���W*�Z[״5���f+���~Z�̆�4�����NvP��u�I%��*IjP�����5�L$��,��SRB6>�"?�3��+)Q_H�� �X���JzK�XO�f�)rk�>3���"5�T9�������l=�6�Z1j�F�N�R�F�F�=#�ޣV�P�F�����޵G�U�֦j�_��������7����<�}���z���UTo=+Qʻ�j�AR;ݚ�
�k �D��_2s��B�*�����i:]��	F�I���Yc�����0V�ķ-�o,E S�ݥ��6�a�d������G�������Y����:f_�����n�����Eq�猉�˨ď��ԯf����18��� �.�{��W1�d�s� ?�i�����%�(��_�{�3������?�~2��[������"`���*���4�Ї�����EGo]���Cyl�]w���'|���H��/��k_�J	I�罬�G`j-I�@"�_(��	�=͑8N9���!]�����CQ�YRh�Sv�17I*TL��#��.Ȓ�����G+��]�\��#��γ!�R��������"�&�6��ܞņ�����r�fwk�I�i-(�y�+�Je)'p��4p'V�bD7���f�^��n��H�D�������B"2��;yGc_�љ�t��b˽TUgz�ܸ�c����n8�7���&��O�����[��/�P�M�)�f�$��sd��]�5H�c��GB���fmʭ�2As�'I�FJ+�:��iS�OF��7uoif��67ꖱQ4ι���};�)���٣���t��9�5���ԑ��p!F��W�H.��.;��_bK�
��W�R#ɪ��Opo]�V�n)��+�q���jw����]KNG��A!��<��U�6�����K���ڶ�dU��<��GM�7rj՞e�0�0�ϵ]l�Og��xS����PF�S}zL�@��̽� �s �o�N2�8��%��yKr�˥��;�F�O�2�'��gb`[��íϼZJBF�7l��?�]�?�yv{�����gMt粄VԲ�A��AK^��c��vu�����=^}��kOE���332f���^��e.���|���r�����D��i�=W)?�Tj����t��� �c$Z{1���z��i^ԙ���]YX^���\�0�)JC~I����!}�|���(��(���p��G�r� ���S����3���c��y�O@`<���I�o�)/8.S[q���R�LFZj @,�N>�h��R"7�UL#��O�H� �#�+�EV��K����,��V;�����a�%0�i;;PZ:�+�k�H��X���Bs���v�C�ٿiJ8�5K"{ �#�w8"Q?�����Kr&ؓZ���d\�@M>��M6W�z��+�k۹>��i~1hZX�}�L�Q�Nl�=�+�<�e|�f��Hy*z�g��g��;���[�zx'xh��%c5_S��I���J �]��L����V{t�"$(&�����է����.P[����H��)���
�����A~#�W�R�� )=��7������y��S������yꅿW�X���(���t�k�H�����H5��a4	"i̥)�L����^硹�[�=�Q����E�/���q	*(5��G��vޟ��L���,{����ꙢA��� x��n)�+���q2�hr�O�D�$�[�&�:���rb���9��	���n\$�2u�nC�z#�vA#��T�?�0�/AK��w~�c�� �V'���T:�}��S�Ӧ�i�³���R<�u���l㼶��=�̢�A��C8����>���9�V������:�~��E=�֕:���aR�8|t/�eoj�n$�����
��Kx���m�7:�la�|�s��z�1����m�sk�:�i��$1�&!o�'�u����J	���O5�����T�݂^��,f��c�<�'����%G�?�Nz��J��0��9h�~T�	�L:�>f�S���^��	F0A�^�J���D���F�6?��a:�r��s� ����l�+��]�$��R|�lz��@`���yh��.Kܿ��i��m�346;)b�_$�U�JO7c
����"�6ۯ�r'Jt",����[S�b2�I�{%�խ�ő�jC���I]�ҫ�'����ǧ��:���扥������j -Ϯ��7���)#��"?��z��mHrPK�h���Ե�g�VG���D��qE�w! 0�0�
��o��]m�����%1��Z��wQA���q�P�eA�^�A����(���A�ՠ5@FAX!��7�L�u;l�|����r!�����t����M!h3I6�ɵ�}n
�YK����7����Mi�y��,VPJ=�r�e@�+7)�/��H'8��,$,X\�1%R2��y�IR}��c�٘zES��B�����1짉"�D�:��g�1NU>B��N�ݏ�bt���s���pN��|Z!'Y@\�d��6��n�W��D�B6�qݗ������Mʏ}��]ſP��P.�|�}\>��}n���_��_�ۀj*��!�r��$�Oy�����:����P~F2X緓ԞX��p9�6��õ� Ŷ�W%vX5zP%N�P����%�%'%'�Cq���mهr��6M͡�,ⴘ&`�,TN���d"�Q����z)��T�o[*�v9�����D�.W��[/�o.5�VxLO�z�Z]������(kD����Y��'�u|��, ���d���g`Tq�����K01�ҏA+Ej��a�_�$��23`@���o��L}w�F���ҖK�?3�<\Xn��;��l�X�=�����^|�g���r{`Ҳ����t�$hz��r�|*�G�J�kTk��U�_?��fW�E3
XtV4��9�R�d��l)�
}�]�����3�~�Y�'C�(�7?J��<�R�0d?1�_�'��t���H���}\QA�ĵ���cE������o�������'�����}��]&���` ����V���;!�؎0#���o��luR6`U�p��*N�TG�B��[��^w���2z(Գ���Fdo2�J8�����Z͟b��[��m�q|Dn:�5(��TB�0�	D���uj��p���)1L�mp�Ve3zs���)-!�:J��&������A��$i[�,��v�R3�ҏ�u�Q�%�޺;B%���-r?���]�\}�!�W�q��"�⿁ve�C갥J���v�]9���m�M$�re��0�s4�*|���D�'�C�Q�^]$x2�Z�
\V��db����E�X�~ٿ?	{�y�����H�A��ً@�G4�tV~��4���d#��kN���5�=o�I$[�����&M�k���?���rԕZ�E�(�gG���_��E��@=c��Bgs��*��
�/��O�R�
I~��������F2�� �jAv���A��N�������zu�	r��m3���]Uo�Vy��Xc�l��⩲�)u�QiU���^���z��y,�u�TNInj섙3�XZE���HC~�%tٝ�(۞K8)��9x��=�-�|�a�0MX�in�#��t��I4����q8�C�ԭU᫴��D
<���	��K�T����A�q���v>Ϲ��n���;\��(;�l�.O��y^����W��5�MpZV�9H�$r ��]%�ob���I�@���4+�RC=\=�m"Ի`�e=}y��C�����#�70ݶ$�/l+�n]B̻vf�v5ߴvR=�w|�^Sv�6�q�K�z�ŗ�3�/2�<�r>[޲�;p�ڜ:;X�=p�������9�G=*:S�v�йU
�*�]�7�w�v�n��3�|���#Z:zF �>�]`��m@Z���m�`+H]�o���e�!22����^LJ��BO(��b�ꈨ�t5����q��.��Kf�x���$'1��c�¸�D(t���P���$�!4,���Im���/ɵ��z���F�i�����G���K6�Q�7@x~��d�`\����'��f2P�z������4���>��M�m�..� ��8��?�8H�*��i�Ӊ+Ǟ3��}��Ӽ{��Y[^�wCj�_P]�x������}�)���&[���:��z}Kӏ��Qn�
�[S9:/4/X&�FmF���E,X��<k�f�z4���#����үd�`52��LTdU$Jq��KSY�Zƽ�^�e�qsm�J��}FsZSqL�RV�IdD����e���4�|~Nz`v$��ĒU-<vh`:C/1�O���m����:��UQA��U�.��uD��"8�iΎ�a�1C�W3�����Wv�'���x,Ѫػ:d��}�8�����g�c�~��j�)����j��P�`�!�ǘ<����;�<^�m�D���G��ԇC�|J�a�?oay�2�?��0���̝28��C��R��Ӥ�,3Ľ�. �\cyv��c&3𖡉���i��֩ rc��{{D��Z�U�� v'7��{u���-?�4��B��.Ο,x��*h.��*w�?�G�U�t�}���jQ���4а����� N7�խ��c�Nع�d��[Vp��6���/G)�²���ޘ$���N"A{7��7|7�	�G�mWզwW�AǏ��W�n.4����ދ���z�[Cy�)C�Qz��A=��;:&�dJ��#��5Tc�c��q_��	�]=��K�M8"��������X�Rq�����枣��� U�"Ӥ�2��w�RB��JK} �Mq��f6�id��&��fUD�n��s]E��sSp�^����;K��3��v�'=�E�|&��XVw�_�a2,����Ro����G��ؽ�����ۍ�����$���oʶ�Ǐ.��Lk�(_�1l�0�k{�'�`.]�u=��'���x�3N9�m.㨘}X?�^|'�2O����d�&ʨ�'f�҅S �jI�@���k�me�ʽWq&�kK�?��+�xb�a��B�I}m>���G���KաO:S6I3z0F��E�d,�}u׷����ӕ�4�w�F"�y����wfS�O*hW��{Gy�RҫA|����9�1FB9{X��`�"���DE��{����D��`��THl|�����EUbY�Vɢ9��(X[���ܑ�D�1�}~�C�.�m���Lp�ҁ!�����v��/pk���`�-8���Z�$��Z%���}l2Kqa��ά=��ԡfE��v�w�)�?U/t���|.?�0�g��-�t*��3"�"������E���=[��lu��;�Dz<�׀�7��v��\)�e��>`\�)G�-5&�u�¤��q��_���#*��4h����{�<G�%��{���?��py{�U<Q"��"�^�{�֐φP9�Ԕh^�C�~('���u�q(~zn����"�M��}�z�|Q�Rl<Ԉ��h�Ma1K���u�НO4��%t�
��)`WZ'�	�Ǝ��u�Ѿ�}�%�,I�?�G�'�@���\��M������>ay����\غ��dt�}�+�����L��cC��8=?	_Ԯw�{�4I͚�Y�l��18���ˣ������G���ZE5�mޡ$\(�d��e)�W$�(�lj�ئ�1�:;;�E,C:�׷8���%CZ���Y���.���˻N�v�4�N�4� K�E�Bx�i���Wv�C�n��wepvä�b�T�PS;�R�8�z�d�|���V�j��H��>�!Ar�7� �PV��� �ȏb�2�ʙ�A�Y�z�N~�7�p 8��=��n[��J�hl�H� �_{ﱵ�,��ח���c�Ё��+��Wr�&�PL#��Ɇb�yd��H���8;�Tm��`Q�j�X��^�|:}��u��|�ϝ����Xqrj԰��Pwl)�^2�\1�1�A�8�$i��
r�I���O�ߩ�}��w��m�3�٣{�x��nqb�÷�O���E�ʐ�q�wg�-c����L�����%%�a"`�#���Ra.X}*=(:T���ԞԴɌn:i�򦑮�".�!�چ�CxlT����Ǜ-�]�z��U"�ʬ�9푆��(�D�'X��"�����w|ǌ���	vj����0�7�����N%FN,0{�D�x�0V%�
/@����V)��%�>��Hj-t0��\�^j24�;1Cw�
��1��v��������DZ�ώ�\�| �CXm}�~�h�֌�gxyL:�ӟ���v�j��K��{Dr!����h{T$[5��M�����}�Wc�-!KbH�P?B6���-�=�zTyy���Qy��4�Ja-e��ޟ�o��m�Hv���9��k�.�n�H��Q!,ќ��F��ύ v��f��`)��w�v��`��@@ߘ���:�Þ:v��x�џے43��1� �k+������7L�Z�oI��gi���X�Z�����='ec�7fv�Lփfj�"�+EZ\M	Mv�U&���ú���ﱄЈ��D5���SLA��W��r �\l#���%���w�v�(�,��o��_�[���&o٤��&���%l����b??��K;��web}��������L��k=�����Ф��q|L�pp�Ԍ���4��K��m���^�]�;��ܝwݝ_�t;�
18�ɹ�k���|�Fq�{���2� x���`�m~��k������KÙ�����z�IUN���
xK�U�u�X Q�k�"%�S�B�`,���A�
 M�ųh�Cԫ�J",ꘗ������w�Y<$�����#&$��+�̦��ӯ�	ߒ���#�ۿ��R��K��Wu���W7u�G�?�f�v�g���,��6��g�TԺy)�X���mAM�oNRM��6RM�N�t߷\"%o��	�lJd�;�3X��R�WM~����f��c>�>��^s�ܵEh��\`�^**�|0�(���w��=�nS-`g��&��K�B�P �2���c���9����)�a��*2�.��Zr�?v��FP6�u¡�'
��{vi��F�D�K�Zb�����T:+k^T}��$���mc��q@�a��~�K�紐��!��u"�yJ�R�;��aJ8&b�q��Qb�����&
���q���߇��L��]�sxtpW�����(e�n�E�㓥$�/���/#��H���qI�D	���&��Z�'��)�;�✵��i�=CO���.&8_����;���7��Z�t�����M�6}.�լ�KDj��P� !Ǩ���d�$���y����;�Y���;	>� ��naL�o�˅+�o�����6�<���x�l���������,aC)�&UE)#�]�H���-��	�q5��LK�xO��I�B%z?����T�1�l��ǅ��hT��iw?�O���sa~�RH�?�[�\��Ѭ��X�`慺���`�A�Ė�0wz��mCA�xrL	# 5^/B�|�����"/��8�P�QD�%�W������4�����R����ٚJ!�vxI��Kw��9u �=���B+ɦ~��V�VC���?���NTaN ��GE�D����-u�^���eD�m]��վ�{�#�ү���ʰ��|~� ,�V⥨�.�`���7��!�<��Ia��o1}`)�V�^����HZ�Μ,��!p:ٙ�{1�d�>��a�k	6���	j�vG�$ َhC��]׻1j�=z_)Ґ���C���-�?�)|�M�=�u��:���[�'�M��H�,�_�g����V9��8��/��AG�a�U+x��)SX���JGc���>`�˘�c!�d��˂ {xa=��\�a��j�yh�,9�r�K��5.��j:C�P�<��h����Y
���"[��[��?�����/:�l�4�5�4��d�\�H8@��h2��nG=؂��)إ�,�Po?�����X���(��#c��97��ja!c��K�
��R�gC��-]�޲�ۿc�
�����\�z�c+P>O
!YEMa��XN�2��a��o! ��������|Э��Ϣ�;��>�ZB��= G'(4׎��E	�Nĉ����?+kφܼ�p�]�;�FY���	�#T'kh�H�a���$�k�9�\��L���ѮT֗;��t�Jf�<��?}K@��CR��{]Ϫ<�L���e�%��-� �g!JA2,{Q!$е4Q���O�<����e���)�1/hB ����Q2-��h��W��o	�
e�2|�
���C�(q�c��Qas��U%���o�� ��ǭ� ��!!�۩�?�x#b��GlÞ�fi��t�V�x�+�us�8J��5���7�@��7����]��rw�l�Y7,_~{�1Nޡ�Oz��h�`�Ǆ�]�l���>��ou�DG�\*��I���d���q?}�8�x��n��ǩ*���u��߲z�� �!_4��Z<��L�V>�n�U�]�obJ��+��tb����-]A?&�R���,4�Y�����v�O`��߇^^\����~b����yӠ�2�XA�s��% �TR��`�F�>���6���qul��^�!��C��=�?{��X����+�����=��ĘY/O�Lx��N|_�b��z������<�����ܿ�=���c�<�E���(əA,0N��Y�ϣ���$T��m/��x�'-G�製������ێ�ѥ�?�K������t�Z����+��.�ϜL�
��2>!�~�X^b���;Isnvm��xYA���S d��"��d�	Wʄ��+��#��H�rY<�b��^{���p�����g���;gl�d�&{iu/�"���3�O�e9���*71c=z��`��0�8'�pOeZ�^\M0���̪NtCϊT�]}3��É��Κ/|���LS*��r�vF���;7o祱6z1R�F��=Ø�2A-%Ϸ��_Bw�Ձ��}�o�z�i��A]�c�0$!��X#�7�A�j8�f���������c@r��'";3Kp=i�d����A�����*x�'�����xMS���$�����)�٥�Z�|�k�"u"��3�P���N��(��~¶�x=_!�ap�,zq�r��	��n�ʗ���Yc��E���A��a!����O#��![NL+���O�k�h 	�O61����A��!�X�C��[��]V�0yE�o��L���1�'�ۿ��R5B�����r��,Q��bM��^�y�>��W�8�EO8��0wB+�xe5o��çZ�q���h���{�X��Z�_�"�G8x�%2��.ڨ2��]��L:R�Ldqm�e*\|a�p�:z'W�b��0��"{U��&(">�.Z�xS����V�Y�*�p2_���1��|�tXм3��e_<��M�~et��r���?:��� 0w��Nz����FK��9H��R��QG�H���eƣێ�뛄�㶻�<�W0�̕�*7��N��^a�NZ����I�yL�m�n�9l`䲋���f�6�����-�߰��6���*�`1?ƅ�VI�sX������=���1��B�-��iq/�_y�ox��C��3����3���-����3?����u��H���#,���FR<�mj�jʹ�5����Z��/Ew�4�^������'(k��&��ƑD'�`���G#Z��"7����ai��7�wL7�Hh�l�{��ùč&����U�0��&���� ���o���/�<91�!~
d�i�P�W�	�|v"ڜ��!'��������V6�T����hq�:[��(G�I~#,AmN���O(c��#���##Q�H¨��1��^�$�����"]:�M���rQOf����a��PK���+�Wvxc�h�h��,��W}6pG�51�%���{��Y'$�9?^�p̃�GA��)O�˫�.��Ta.�lq�xcA\n90x����4���846]UVd�Ђ�NЇV(��([��l���%lz�I{̓�|>Fb5��L ��$��ށ�k�u�Ag��$��A��wi@��1=*p��;ɓL`��5pM2���C�S�]�}�8"*C�vC~<N���VI�l���.�!�����ʇ�j�V���v�#���l��� Xn��S�ڬ���`B��#U����W�4쮩�S�f{�C�-@�����k�]��a�7_)��f
؎0�c�2����84R�K�5�L:7:�]���6у��yX�-��KӐة�0D��#��c�#��}�]�.}v|����z����v�&�������	�h�D�/��}�͒xc�lig�g��d�Űi��I��Ma!{71Xk����=��_�L9��H���\���1��50����KO�h,..�#�U#�����.�ְ���5d��Kx�I{����;n,�����k<�s�?͇5ԕuhRj�#�w|{�$��s̻"�1u����?�Tj9�(�ê�,쮱"�Q���s��}�oM��-���ԡ:���z9�"�L�� ���C�Zր@D:�@�����&�WI̪ٝ7�YeN�S�rK�w[x��'QR8p��$�k��O� R4�Lِ���Ih;Q;�`8�T�z������*֗]��c��Ջa�I~3���m@&u�ȵ:	�G��5�@8r���) v�nߖ��y�*�A����G��J��$D��w�j�\RE�k�,����-r�vy�2l}?3d	��h�~�9�!��i�����?�� �=v�B��I�a�3@"اǦo�Lgr���ЧȠ���__k�q��Lȹ߯�����+~�0�b�]k��K�7;"�`�sI$&x����ԑ�B����W׺��)�l�}ɝ�u�#�L�P�|��H���I�f�g���-�I5����8���K��xfc}b<0'�����'����M7J"�'*�nl��w�6��r���vRX�� 8fj���iy�4) ǲ�l���ѳgaz2d������L��%e�#6�8�[kR�^~a���c"��I�V��n;#m��
��s8��������}�;9�P�K��5�%]׺����Ig�n�̘������7�-�5�<d}! ����w���6�X�'�������O��ә/������,��;�Dq��,�r]��@��<ZV��ŤU�v`��:������䬛R�����z�E8�MRr>%eg")-�b��1d4�i_iRE���T�#�tڅ�����ȏ_�K;P�߿w[�7���>~���#�{�~�}�gh꼾t��_ʻ��C׺�������F����c�����9/W��:�8X�ե��T�6	<��ǆ���4�
�E#ӓ�efi'��6�E&�� �2�%�������>�*�Q�f�@Wp�ذ���a��B: ����;F���&\��F�2���a���`�wj"�+C�ē��"�m���TYȈS��H�ά�Q2d.�p�F�������%2ɞ*�	�����V��Ly�פN`� ���nLu.c���� �������q�c��)ﴖ���rՍ�`j%��a&�{���@���9��<�h.ь�-�	儕�����瑮�p��ƅ��l׺���'s�y��Ǭh?�������A��f�?���b��8���3b�����]A4�uB|�q�n�yT��<8 _iul��Ƙ!��⻎���c=��z��0���J�o#��	[Vx>~�x��k��tv�)�l0�u����ą��|ȼ*��������nD��Y���V�v-L�f#�[�}�įֵ%
&����@�$�����A��l�@���j�p�X�� "��fw�h�����V�0�j��őm�����3>{�7/�#K�7:�h*L׫|�������\�*��.�BRS특�5r�L�e��^�5�@�4+C{:�~�'Z�ƥ���L�e,�S9���w�ߟ������oLz���vp�(˞�ƹɿ���{ӛ���[9([])�����g��b�lq����9���Az�/&��� >!��bϤ�՝�u��WX�F�7����EYQ���B�~[��w�*b2U�[+�u�\��(��7q�4����Ǣ�R�D@]�z��?l���F�p�l����tjg��`�-ZW <�����R�|�p��4�Ha}�x5��wk����]�-$&�����Df�|��W���%�~��`��>�(��a�K
p��;�������xn��l�Q�%s���>{���RlJ����af��W�����W.Zy��9x�O�>�$��i̅mi��w�|6\7ڇ \?#��2F�My�����9���ye��I��a&c������az?ҿ�]�D 26�@e�/�F
��bB�S�=L۬~���$��qr�GD�l�(�U�퍜't`(��`�}c�� أ��C����]�X�4L��oQ)Z2q���q"a1Ƒ��b�b��}/���ן������k�-Q�Gb�b,'&�u7���ʣx-v*���^H�W�1T#�4��멖�
��{A�B�i��gɤh�Sj��ã�Շ��AE^�v�!D����+y}��3��h�V��^	��>��`?&S�-����{v�%�����7/�w�^��'�_N%28��U$�M�%��בl�`־O� �6;� O��3����-4����3R6�j�l$[^��Zb��G�;y�2:�q�� �j���1�D�3����������nNMї���W�Ђ#有r1�{���7�R]��k�D�j�1#/�1�a��|�'����z��o��Y1���$��S�~��>���t�_��5��='
�ݜ��J�S��;	�bx�V�v�Ӆ�����v�Y03��FN99��Q�Z��Mϩ��Z���T�F��R,�\`�u^�����eu��h������T����d2��yL�e�uyZ�w�J��U���Z���@�2�ҀjjB`�'X�M�I���e�;ٻеyG�偬-�<��^�k:��V���n?����T��N�ߞ��g�f|�Yn����5#�-~�kY�q���j��>0jZ^�\na�����*T� E�^����]����}�1a���k�ܝ�1aٟ ���KH{�DS�F�88�PO{�"8#ߥ}xE	r&�@�4M��>�߽E�Å��Վ?쾛�[6
���t�����ʨd�`��S�N'5ĩ��*���A 0�ך�P�G���@�z!i��Ld��d��p)Zf�OW ���,f�����,`܂����3o�����NLM/.-�_��NX�>�bby&2se�ڎ�_t�jj��5R��tں`|�����һ����<`Lߥ�Q	�꽍�����5��j �����7m���6�b��^�PyN�~�;��0F��W�w_�W`�Y�l��$���/� KmH��vԶ�S��r��b���Kr����x����eW��a*⧮�aR
L+u8�>�?�y�#�FXgQ�b3q�g篼(g�aof��NNoMs�mbW����%��6���.���9Kv���@�^��^�*��հ��o.��H��
"c�/x�&��";�$+`X�]���їܙ�?�4V���m9YL����SCU�9�j���U���·�a��,��5��a��!~�E_D	1t
����i���^��r|B>���?mD���O�l<{]���6��{}���a��q��`I�!�<����5L:Y~���zL�n��3��ܳEYޔAl��ˢ�[�R(��6��,�8��o��1wV*#�,<��J-J��V������t�M�� �.��J�LB�
�İ��B��fJ�+n�'j�Zp�������2�;��k�RU+t������3�w�U��D��\g1�����p����)��u����^�MO�v'[�q�Ds0b����gO�*�Wx��C� [�S�PO� ����V>��GGec;�1����(l��.��[��������=���  m���O[��:)se�x�]#/�c'Y�?�V��M���� �?T��6�h���d�c����E����9?yA�ԛn���NuY����J=��=�켗�dA��ߨ�bu0���~���Y�۾Ҹ�﷡K�(��.Z2V����N�ZϜ��&�޼��-��ߜ!i�8�o���	�w��a��j���q��ѣ�GAL��W����}[��N�N.
�(h*L�␞ӒVO�5��U}�L�70:���������#K�""�%� P�����O)z�%���d�FS����ru�����՟u���1���d��g�d�F!�&WT/?����Z�_�eI���j���j�-|���F=H"�-��g�Z�޴���׬-�g��[�=��p��}]>���d�.����u��Y[Z���Z����B0�L��W�܀��%��ٮ\%dS�k��O��lR�"(���"������(R@,Q99�	x�s�sΟu����jGƩ�MO��@_���F���B�,*��Hԏ	'��]����Ui!c�#'�����ɿ��][�8��u3�0��O3�vV�-���%A�c����H�^�ـ��Ǔ��@"xUiF1�r�5b}��=0��g/C	c��H� u�����w����q?�/�.��0�~�}�_�Ðb��g��7�V�'�㯅�Z����a�F食��@U�v��鯩�_����,�U�j�>4�0���t�3�@�^�l��M�$��z���$�,C�5|Y�=? ]����I8��lZ~�_]�a���m��#�a ����Bw�,!��5�r�-�U��w���}�� rS�6:Y'q
Cm*�N��`	��KG��m])�R-���Ӏ]�Y�be;�� ��K�I0T.�ʅDTV� �ј�aLn�4��lQ:��n��aa�τ ������{So9e85[��'`�}�1Y�e��ڗG6���47�4�K��\�n��[��#=t�/�"��j��Ԅ-���������r;��J���߂O��C��c��C��M��.���Șp�ez�XZB��q	&���L��İ�8}�Cs��\J?���^|2�	�!t0���|�����}zkL)��������.1�P5Q��ʹ�B��G�j�{DN<p騃f��wV�%GUp��נ~c��X��RT3.3s���������"��(�l��mq(G�O�`��!t�����^Ok��&�`�M�0�+L��{�H`#)Ep?�cg�W�%� �џ{�4]���&��5m����� ���m��T3,��=bp#ͥ���C�����(�t�� R5REHJ�B�}.ݧ�֊5�A֦����RQ
�
��J6݊�R`��H����\h��=x%\a\m�LL����:�o�T�i4B�"�[�z_A�SUM��R���I��b^oL��4�B���������� ����]TcԆE�}{���[�ՠI~�K
��`��|� ��!�v�J[�h3M�w0Lu�w��;�����i��Cm_d�h�T�w,��)Dt5-Cݱ��q^q�=s�6�L��n{����Ի��g�W�����Rv�&ח�p@����Q6k��(ttLB\<9@�(!�EFON�BkU��5I{T���İU�����_�X"S����6a�P���0up���ܬ������9?�����!�y�Ք��U��9-JO7�LbX�4[�����3��֛a�(��'1(U�t4D�V����:΀k��y8,%-ls�~�aҕ6�)k�t@"#�61�|�Y��:$��By/4��^�p]�^�'�9�F�P�#b���*��f��Hc�`+h�~Y,3�X�Y$.ą��#�CIk3#�
��(۹AP9*�{$��,�����X�)B��b�׋��(��K|N�(���8�%G:飈"D���B'}E�ͨ�*qtf�������~C�:[��q,��]i�~��W)l���ZGLVw��?�d.M�Tr��~�iQfF����Z��v�w�q��R�}��\���Z�?#��m^���	n��ˮu��v�	�Gz��O��.\�`>�:�kS&5�:c�%-�`�Q4�g�?���+h�F
���}��vl�x1���B'�+��#�AL�} ��7��Z�G4����a�g��G��V	K����XxdIF�4��}�4&�.g�6�����[)�8^lEZ�>���&��Kn��Z��gU��ocL%]Ao��{+���Cܝ2!r��b�X� ��ą&�ԍ���1�ܱ�払}�e����%���ՆS��~v/�+R���N�
�U����Sʜ[/Ppxe��T�y#�v8}륳��gyY��P�t�i^�o��{�^e���3s����FN���ୃ�����cQ�q,E�	E$�b4gs�ݻ��U��b%<Hg]nl���'c�g�bc��Rӧ��G����U��<>������eP"V�p.���փ���pNw���J�Ce4<�k�:�,ؐ��}�T"�WT��<���r�̻����0��������V��Զ���CY�Qo����
J��
(һt��
K�tw,��4" �t-,���"]K7Hw�oy��<3�0�ss����<��	���םRB��%F]ϓ�%F������c�,&p�?ch��Z磫�Mf.&�B� 1뿑4v�ª����Xʧ���`��W	!H��
 x\�
 �G嚫Ba2�w���a��1���,y�\���d �{ƪ�3d�ڗ�P�e ��
��ŋ_-N;�(�ւ�����W������4���+���JCˣ�~�\>e=߃�_u�9;'2��Aݝ��=��񱑹��
(o��/&�i���h��|����Wp��N�^�N�\�
d� ����4��^BU�j���殅I�'����F�h+@���DP�F;�zc<Sa��P����w_����s��1ľ�nSleb#��V�!�p�;��B�Gぬ��$�C���D�+kH�IpI��,�����X3Ա郹;J��:y��\��Z�9���l�1�$T�����8�@E����+�Dե�4O�C����|�@�lo)�k��(m3i_4�Q��_12���R��cO�i��)�f�ZH�D0�xrD�3��iȄ�,A���Iv��U&�w�\?|-���Xz���&���ań��_*�H�g�!a��,�m���*�Ǐ��A\��*��B�H��a�-Y�5���?���ה�a����	��pؖ���o�'3� ��/4o�(����ŭ]W=��|3qT�����}ois�Mb�.]����C�r2	/��/ˍ1 h�EDe�xG�L��,�\l��s� ,2eK�}#Ϳ��K��D#8���P����a���P]�e&�TN�5 Ǟ�7�&��x�4�k6�&��`rQ(��ņ_�n�8z����^=���һ�P��߻;�n��uH�-��C����̀����u���Lq��1������`�!}Fj��_����n���)U���l���`�����j|#/�%��z�|�v4^4��Ĵ8jJNO�/E�2�{���#��Ս�s�:{���s.\��b�Fǫë3[�g��7�.Vs%Ľ �@7��סc��^{��>�ӗ7�,�`�����(�|�y%�m�G�9����2� �_��H[������ sH����IV�}�;��xd�um	��W� �b��J���`���͙��˂�A@ФT�Q�"�(W�+#�Xz�\���Y��ʱ&*���t�ܬ,�BW����~�o�Ղ��*t���eoaq]ibu�ӏ4�Т
�g�Oj�) jp��4/�& ��ac�Y��\�`�K���k�������c�E۽և��!�D��<�i��c�IY_����@�+qBO&�{�WdPs�HZ��c��)Ef"`�gu{@fૠhChw�8��m�o�w��W��� h�t�I%C���(:}�f&�V�R������tmؚ�oK���v{c�������@���3g��?���^D�?�{�"��c@����P�.�l��@-5?^)2Lt	�kU���g������n*,��]n"E	�,�z�%�V rc�ۡ�'���j�r�3�^��l>,��B�R!YE>*j' �l%|ng���Z�rQx�	�d�� \B����'�h����Y[����K	�����	��uQ:2�r������{������K`D��t�7$��k����;�(S��)6q7���
����L�h�:Τ1�@ ����dx�A�H]�n�j�� �7R[�d��?q�A&
:����ל��g�6-�O�4��]�ގ2y����kʁ�]���r��M���b!Ų#�R*#���W�{��ϽV�|�����}�f�'�������������y�4��*:B��`}�I�>�8�Բ��q�z���-��t�7Y�qm ekiI��#I[��q��f��V�"?�<I�-���_��v�\��D�%l���\�mO㻢����\��y���E�j(��ę��Z8?���Zh�7��:]i}�p>*�K��Gщ.��JD�'��xgg�D�P��P݄��NŃ��P��*��BV6/�0Oߡq.�p	P��a�YBQaL��YHq��ga�c�,64����Ц�܂Z�� ��;��?�Cf�%@�@ �U���oR�c�����ط�*�޸�����XK7:Y���R���^���gU3>�P[xa��v���gZPgu
��Ջ}�F�V\�\���c����)�*-�8���]:��� 9�ҧ:y����X�^H>1px�d�f���#�ƨ��Z��$(��알1�A��3��h��j�\�����D�\��c�9SF)(렢�����4����� :M�pt�㦗��S�6�`O�0�:v���掍`
�$�{�n.�u�ػ*X����p��`̪9i�l�Kev��^�������K�_b;��wAZU��Tk\���6B�yWCT���n>R���@b�/ [v�e��D_���uQ�P��[\��3^�.�{������OVq�����\����4UIq�2�Z���18B��jH��2�P�3�VH�p���l�dP"y��� b��:�����XG҉�V�_w��֫����T�o��m�H�ם+c
@�zu`�ܳG����=R�zB�X���ÏQ�-���w�_#d�\jS?�ǵw��T�����J��T��d��rF���
��{O���I��e�t"������JF�p~��d�����v	��rn��Qo�V����	�����nC;dv�7�ޞ���7ߌޝW������7���/Ӕ!G�b��b�k��q��p���IL���H�!>M�GȊe~�;">��Cgooo{���l�c_ی�V�S����@2Ȓ�2�,�]S��������ާ���m`;����
��h��$�A'�Nô���F�g�W"$�s��N[u����U]�	�3��f�U��1�x{��}�z;��:� ����G��g]��Y�`	��s�0�[L.�Pa>��s2��d	ee�c�(J�#�M-����ae��z
�`Cm�`P]�'p����l�_�2ZB�}�^MĠ1�q�Gb����C�l6��;���x,�F��{'�S�v���G���O���8�4�`l�2P��tKJ�^u{�,���؂��kB�k� �$�)��������Fv��#"�o���R���f�'�hR~����ŧ�8a�X3?
2�@���C�,	�q�Bb/�>ףU�ihq����Ch,�u}z{B����%��U��'n��d[kS/x��%ɝ��E������DV(.�$%n^���`���V&]��������B�.��(:Ā�و���s��F$�u�B`��f����?�o���`���FR8������ڗ���|�&���K_�gQ�d��=�H*�򗂶���N��P��e��dJHA4����i����+F���$�k����X�=��piГw�����l��%�y´߁�r�8�յ>�F�a�ʹIG�X%�7��W�ʜlA?������Dge�Vp�a^�{�l�s���ZǛ�!��tY[��頠�l_����{���LL��Ӷ���G�6��b)o��_æ+׏��b-g�|��,���TaL�ɒ�=�i����q 2�꺯R��>����,������R��n�#G���3'�o����̗����Ȝ��SkG�d G�7���zb��w�g��)G^t7_����]����e"/v�|���SC�a;�.1�\�_P(B���07�MMu\�Y���5nK"��b��+�/>�����}ަ�aw���v��ζ�L���݅�y�������[�3B���\Q�m�-�axn���t&e�S���oa���.���e�>�V�IW��wU�.Y�Q��+`�3d�}��,��F�K� ,`�h	��à:��m��Bd<�9TY#k�Ơ�"���'����V
r�2�)N�K�����n= ��>s���<�x�wd���}x�Jn#X��!jt%A� %B�}�h���-d܎�ju�Ό�)l�>0jOKŹ�$kI=�"v�պr�N�ȥB�3�r���a|��ơ��6�n&��6b��%*�~
�	���yb�_8]��Jrt���n��R�~�J���礆�l>�� [_��ԝ�|�Y�GsMK��H���s��7.��`<��9l@z�	�Ap8i��b1�+�jv��_��R�;���� �7�q<?:�Ǉ��i�=��5���v~��(Ȑ&m�~=ً�r@����@l��m��~~�N���ʘ�Ҟ�a�8��xv,c蒶��d0�l�,{������MQ�o}���P�ֽ�Y��4Y,_������5����������ONˤ%�ps�9�5[CV~3��$+��GD��l={��p�Ӱ��vT���2o�s��%k����7����f�.=�z��=x,���B�{�`F��U������s��Qײ_��h�ΠKR���4y&�5�$���<��FI�?� D�۠�� CR&�|���R�D�&�C�>nÎ'�-������laI�>�u����7���Қ/�i'ش���}�Q�ޞp���Cm˝>Os�ϭ�����MyW"��b���)�h��6�����w��wg��Mޗ�6�Q��\'KjF|����`6c���ׁ��K-$����W�UG�)jϽl3�ǁ ~"?+���kײԛw�J��㋜�sӇ�s�{�;���g7I��Ŵ TV���|����xe���މ;ۣ^��.�D����!�W��c��o{y����w/N.t2\D�(���3�zbE˦�& �AVw ��`��x
<h�Li�JarP�m��K/sl��~q=΁Si���c	�� Aֹj�H{�/g������\��r����qF>�x�9��UD�zov�}㰒Cy�j׼��՞�N����lF�y�}����
�xb#�,!sa4��D6����7-UX�F1�J�U����'$A����� *j�.�X�;�7�[�sl��.�~�u�φ��+G�+��V]�e�p��>Y+O�[���X��|��׵jT����!|h�UQ?�<P�e��C�?.E4��2#�tą_"]��17��_��Vq�hƯ����V��ۄ���z��]����"^�|�r����Y�2�p�?-�g�4�fu�P+x_rSܲ���ڴ2�Z��D�S2q�J0
����y��������VH�jg!^���-�Γ�3ݥ�͓+PѺm�?�3?E}:^5���TF+�P��{�<��(C�B��)M�� Y^#y��9+�X\^#���#�-�*��o9z�_�Y�QښV�P��s=���W1�ء.5��ϻr��߷ ޛ����I=�����m�妟v�Ís�(u�8�������C�~85>��wim�@�59J�!oo�l�>���z-���h�Ӳ��e���l��~�&ü�_�]`�Fh=J�m�[Q�x�Iz��_4�Y���.�ޓd�&f�Cu�:ކ4)?m����c�V����5Z��:�S�Ҟ�����q�e �*?�U�55b\GjS�̪�������"b�b��J��ul�֊�,��N��|-��d�-)�-��PS[N��/mB{p�g�/u ~?� ����{�M�sn`��TK����}%%%��]�2��9tK89,�uO/Uz��Z�9V4Ԯ-W!N����FŮZ�|.c�'��\���,�^���n-\�ǵ�z�6_�i���.�ݞ0��M,���^>�9:һY�k�GѪ���&��]N'oW	�c2&�u+��w7)Z�"*���fO���w���:$�$�xO𜏶s��K�)ۋ�-Z�3b3�?d�}���yzzzx����0H�<F��0+�
[���4S�8W�q���t%�<��I�2�w�0z��(��`_і�/�.�%(H	�̒m�|8ܒ��?�Ȑ����Yr���dȏ��뾿d�e�S�����F����w\/5�N�皧N]��\�uW�ZB��M�tb�]k'[�lQ�ON�A��K��������]��D����)�k�/hxn	a��GE~�!	� �':#��'�������H"̈́��޸9���n*�撬�p��-�
�@`x���5��hN�l��_K8,���Y̝�AD���@�w#�޲�=}ZO�����09�2���c`[��	�����7iO��e�TSV�@22��?	8�3iJ��%3{������H=߀pӗ{���	M\#ݞP���m�
 ]�����Qi�q^.
���}���dp��(���f����6�-�����b��:�J+_d#�8�)O��v�qɳ�[�������Iel=L�&��ʛ�gQT7=5�0���+�̕���h�u`�m��/���R<aB��b^�[Bm@ �*s�4�Od�J���	{B:~���fd����(��]�ջ����:������%i�o�\ֻgSy.����LffH��b���Χ��5 ����d�R�i!����i�A�~1ȥ�ɲ��:������yu[���м�8V��Xμ�~G�� -�
ѫ�d�~f�?����wh��4��9���i2\ZT�m<��komc`No��"�2Ō��=䭢��0qK��ԅ=�lBW�.3�2 x�Cz�@�{ʐ�UD���d4{Õi
4����s�G� /l�P΁�n�pHKc&駱\�L�Q�Ezfdxw�����{W�ߠ�1�3Q����<f[ӧ��<�
!_�	��5�N^��9y��0g��2�]��Z�I$�mL (����]Ȁ1ՇxYt�N(3}�� ���Sh��x��-O��B�e�D4���p���#�Irȅ�Cz>G~	Q#�#LX�H�ӌ2+ )�T!��۴������p����������xm}��')--����lN�y�-�y�(�I�7_/U�b��ۖ��W�nB��|��v���VvI�ר0�ý�z}tw>�v�m볿"v�:k:��Zݩ���.�F'��b�߄������Z��x\8�"�s'S'�Yr��qD<�d^8�{P �RE�&?3�<������iD<�3�8����}a!�\J�a�IZ�g�L�p-���E�vw%Pzy7��� ��x�������|)��^M��4u�X�:S-x�_�����UAg{^�'+���35.;=&x\�G"���g�����Gd��&^1z>�cTz>��j�l��n��b:D�
m��F���lQ���esm+�%��S��Apz�w~��Ebԏ�p�#�W7����GP^��`p�6���ʅ�A����A �.�p$�	�*�Ȍ�27i�"����,��s;	���{0Ή7��X�;��~,߿Z�¦��� ��u��q�{���Թ��=U�Bk�:B�|�!���Ƒe�bC�F��?�� n�wV�1�/�����@���3z{rK�W��Fy� ����^{"��
w�&A�<�k|Hl�&��fԵCkH2�?L��xN���?=�$��?�#ũq�s,��PvA�'���h�R�q�J
M�����|p�������/���`1�A\�m 0���p�tۄ�����7�?��c)ۉn�M����kKA��-"��Ǡ����Z"�Ǐ��`!K�'1�EVK��Ed&�4�H�@O���t��4y�[�="+�ø���:�����]��S`�Ky�OV|xh��k�x��܏��@���cs�@~�J���c��c~V�ÁQ<ЈH�0����¯����|&8&.��}E�K ~\:xQc�s��x��=+�#�:7ڍ�@�~A�EA��S��=�"n��ŵ1
��\��Pbk����>g���e�x�#ty�<,���c��f'�}��������7�����h
�D��iA�3{ �������|(�D���	1AAA�7 V>F>��-�Em��s�Qt�P��$��nSf�"7�v��v��u������%sW2\��!���"�����V�z��~���cѻ�˛$�����"�5V'?g+��M��"d�u�|�G:	�,��F�D�Q�� (`lX���	��@���cYA���1��H�����\\�M�M�����+����;��e��W7'�?��� ץ���������
���s��FnU��W{�7z^�h�`��Vǲif!�����A�����0�:���gIqe!��-���u89�Ϊ�k�yiq�a�������)�7���7n���D���!�r`�t=�[c?���Q�a��9��8\G�܄TFC�ou�q ��B��<Nb����@�,橿��ԽaL��3��SA�_>E.Σ��~�!jA�}���8@��iL�w P��@�)6]n����T(����-{(�z��PȨ�
�_ ���:��JD������Q��Aj+(��߮�D]�ܗ�u���l���9��f�|s��X�j?�a�d�CbW�-k�h��nΒK�,a���5���)��`p@$?�<|:�F���[¸�X�XM�#7���� A 3�1j�2ZtN5>C.#1�)ML��Ejo�� �l�Ul��n��Y����S>�������ʒ��$)����:��|����)��*~g��Ey"sν�<�<^;����GJ2��lثW�Eu�a(�n���&�Qa�Qy�i�`��|7e�b=���i�JE���a�H��L�%�7�!��{�@.��,y���Q���-�\:�-�w(SI�Y
���`F���%m���:Z]��,s������tCo� �IЬ{��hs�T�kh�?�r�m��P3\���=' �(>�*�{��k�I�Ȏ`�,��8���-�@kOS`����� Y��4[a'���fo��S�J�Ԍ/~�7���9\� �+S�$Z�P���Y�����)?7_���e��agz�J����w@`˄�nA"$W�n�.6�շ��"ݦ��UJ�׶�ǒ��x�DM:��3@54�����oGv�"9�"�rg�n�N�;��K��؅Wo#�j:~�f,����*����M���m��Ϳ�?���X�
~no ����=p�=i�?��݇�q�=Nk��3U����)���*��G�����4^<Y�2�3p�f�s��R�P.����d yڷ��<�{�WT�`Ū,0p�Ŕ�_B�=
�d{�4�@\/"�U�$`�'Naʅ�.�������
�m!��	*'gH���p+gp4cFI":��ˊ�6gC�s#g��/��v�F|������kG�NwW�7�T.\��p׸W�5z��艺��F�����z|��c��/^��"�J�m�=���P��6��jN�n[&U��`�P��\dw(�n2y7��&ˮ."�oz4t���F#ߋi���vV�ˢi٘R�#�*偠X�E�+ꍥ���
��<�0�ڏ����N�<#1L���&��p܍a�u��T�b��L$�mPm�ݛ�F����AO��������9P`!b9+_s�W���0��<Ƭʓ�v��Z��;�lX k�u]����D���o\Q�=^��=�3?���A��n�x���Ј���:�����'�2���E�bY��ӛ@|�Ңl� |0��!#����7�T�'M�#@��rj%r�w�լ�v��G�$s'n��8L����U�;'��0�IWbn�dH��������;IC��PzmI�4T����H�n>�������髬��P��ݵz�ZS�H�J�{��hJ�lQ����Uo9'&�7��.�O��������^�ħ~��/�DY�c�6�T	s	/	�W��f�>���f"[����X���9/����=�B�i\��{�SPzj"����x�{Y�C|V��6'Xa�.�y'��*8Uڿ��#z�����'鐪*:�@	��v�x����ϻ�G_�B|��[K�;ы�QbB(�& �L�V�Y�ܳ�tQyX!�N�Y9�����Bcb��_h@8Il���K�����r�j��aP䢻t�>�`�%�K���2����MD�G^��1��/���R��\gEx8�oq4s/���y��Fs�O����B�B�����+��w�H�(��v�/vׂ�S��<��O��o�n��|��ߝB�"ۚ��NG����GmoWr�G�.ҼV��n՚��n����R���Q��̃tl3Z%�c���#��H�H�Q_�ȁt���^�v�d΄�b���.q;O���z���$XJh���r���q�Z�\W��C�Ob���)�&�S�α����x-��	Bf�_���?Z�Yn�ٶy�̑*��1���&|o��r��2ͷ~���������jJ����_�\��r�3��Z'%'���٩T��FN��Q����4�� C����Xaύ74��z�����P՜���'�iK뱐r�EݶL��r��b1-���*pa!HXOwո3�­�̙F�\y�r�h��d'���'&u�|a��s|z'���ֆ�(T}����,��\�Q�/�acV�Hՙ���
��o0vL��TV]vL�v���4d�y�{��"x�\y�O*t���=��Oɤ��c��&+�mf�c G.M�z7�r��c@ 7�sg��Ki<�p�2�B�^��Y��-G���gY��S��mM�B#zы��X_�07�!g��:��a�ƯH�}�D���:#�|%��ģOF���?0M�E�Κ��}�X��սE�攈�JZ�*>�T|��V�<j0>��d�/	<��ӊߥ�"�BZ���p
�VF�g��l�Mh�M4�ղQ[׷Q�	�������t���'�p�O~�9j����8�R��K���c��~�o��ާ��n�s/�RrufX��Urm&�F�T[�f� ^I��d@�v�p�9�?%Ӧ�/_s�XD���HN���
^T���PŖ��I?��g���(5w�^�C&���*>���y��E�.q��u��¡f�����.� �m�v,��.C�ښ��e`�F�׉�i�0��A��6C�q�"�1���m`��0�*����j`��{�*�_�l��=��#W��~u��DӴ_���$�w~������Q����ŝ���?��uYϞ�H�I��G�Q��Yh�N��cy��z+$bԙ)5�k�2U{��yx*+x�u`ag�X�_��0 �������	83�w��9mͷ�凃�'���ŷfb׽�}V��|�X�������~YΝ��r0.�W�<��y�Zka��u���1�A�\Ԩ�K��_�[FS�/B#�z[g$*����`���w�?�/C����A�!�5`R�����.��n+��ό^񐭴4�뀨�S�����>���Z��Yo��qu���o�t�l:���u]�M�?i�:�]�Y�����z�:�"K��D�a@#�T�Ac�h��;��r�� ��݄:�����p���b;�MwD�s�� �%>E�z"8��G�:#�?�4%��3�5v�똆辿����4b��$�R PƔ���>�}�ܠ*���Q��g�) lE�V]_�|c���/+g.c��Aj��8�<��Z�,�k�)�wК�)����J�c�V���n��M���5/ϛ���ϼ���5͛�F�p�t��S
�X\��~�q흍G�pqCm4;.���d�9B;�ǉg����t��0#��N@�THI��[�$ �0�'(������Z���c��IB�E�_¹jz��'��FdƣV�䲬�>�Vx��CX���O�<�MM�^����?��i`�#2��:.��jdᓳjfW8�Y:���&6֩����1��NaS�.Q� 8�p(�咵|^	7�/Ed@_�#��)M�Z9#x���E��i�n�Mѹ9��2�dT=�����X˂dqZ���7�
�i��`Vx��BZգ��;�+�"Z�@���'�ZBk������� �go7ّ��<�Yq �+^b��@]��T"�hǠ�n���-��~;T
e.p������C=����-�P��dLK�N(�<������� ��=�W�{��E��5�q�Ḿ���"���b��3�b��,��}N!&�^Z�L*��؈$�j����R����L8sf-���DC�s�'�`��A�O#��^I�����wЮÄBٕ	�#y������������]HsT�Ĭ;C���)8������Ƽ@���<�i�~��%���w���(�뚷d(���t�\x����	��y󆣯[����ט���lE��`"�c����˻���u���=�+Y߃����uߋ3߳��1\������.ߛ榻���+̾�W��W�j{���c�7���:MvA�}��2���B=x|�r��ԧ�I�%�OwY���k	g$L�.�fD�6�A����>$=rؘ_K�Z1A�TL�m��)a�ϝjzpx?��MZ����m;�d����3e&0E�u{?eK���]�r~�w5I�b��o.����ki���Ʃv|��+]m�'|/pUK1�0[�~�?[�1ɒ�;M�cu���x��&ў�Q�,G-������d]_:Q�-F�?E�cw�,��.�W{=x%�z@"p��d��X����P��⨿xɤl��7�A�x����f�9�Y�h�"B��|��>����nH#�,xwq`����P�!��/�S�Ea๸A֪
��'����2����dݑ�X2��o��9��/�c�Ե��S�k�o�S����v�`��CR0��1��U,g��aۛ��_TmG%��^ZN��4�6J�?A�, �T�/��&���K/FRڤP����;�����m�)Y�%�@�7�tI�G��CяsX2XI�G�`"��H#{��uF?đqы&�8Z�^�}����5�e^���ku�kDPި"�h���P�����A��K���	�W�֤� P~�A�rVh��FM�>�dg����vO5�M��xQ�Q=�5u����~�߻4�CF`��E��Qjo��A�ϒ:�Ӯ���\�<|)�%�G�k^k-d#^����_�]��������.���n�k���*Ƶ����^����G��A�?����UT#_�F�ӭ�	��}�#����~E�������:��������}%���BF+3cQTؑ�t��̈L�d��X�����*b�P5��f�HL�P}�)������f��=K��}�@�fm�g������}��%�MME���hmUr�F �C6�
������P�����ߕ���}k6d��>����Q�e�1"�ܝ�/g#n��fHm~�`,M'��3Nz'e�@v��m��F�dEK�,\�ˬT�T Lg~�]�����l���N��t���G��)8%�Y�8���E�����gZ1E��/g[@r����Q١�L
�����ku���?��l�R�-V�0�9\�e�`�/�F^�ŋ�n	�y���-��7��?�:Z�\N�^�]|��pg�r���G�|����E�=�z��MWo5Gٝڀ!��©&���N�P%�%���í�o�� uT���\���`��G����X�ы��q��v�J�l���qvXB�����J���iʂ�p������v���k��������D�}S���C̈́M��8�gC��G�A�����ef��|��(+��)�z�=,Q]|z�u�WH�jDm��n7�k�������ނ�]J�w��͙N�󍃖�Nƍɖ*�`��,���a���,u50�t�|p�*��a�M6�۾/ox�PV���W[2��۟��
h������>�/��p8���y�]mE�'� >��q��o$��\d��9mRguc48u6�~�2@u.���э��w�s����[J�ӑ�tU���b����f$mk����FM�X��ƱB�ns9Di]�XR\x��:Z�����s���Eg�
��2�V֛����!�YY�͍5͕�f�Y�T��>�
C�6|��Hl�$��Y�,{ƚ���_�մ|�h�q[, ��|��ܤ���oT�=�Wpg�Y��R]E�]J�t�E	�P�c���	�@�@�@�"mC��W���nQ,�T�YJ��ꃭ�F�S���C�̍��;k�$#�+S�;�[�}�i��e�r��Y���؀Y7'y?�t$�PV�U{���va�<�	@�>Q���B(�����d�ӵH=���¯QZ��je�?T双z�	��j�Zt9�ĝ�B>TA��S���O�y�!����@�,�:Όz���xz��]zb2[��L�I�Z�]d�:�3�u���W��#w�['����7���==�=4j�h&3��c����_3-R�S���U�]��fI� ��t�h3����F��ℍt�tKCW�stH�:�o����ޮW����j�[�SQy���S~�G��'�l�r4dd@�+�F�I�]^`2��������6}�/2+���n��q\�`9��\�ZA��[úH����.]M�0>���̌�`�R�Gb@~b��\7��0%����B�0n�-E�i�.*��T}R6�J�u�ˣ��i��SN%$b��Sk��tLq�`�j�����?7Y
ң��?��{i�o�.�Y>�;n�>��%2j�L���5�c!���ތ�3�%)lذ>X�m���O�*B�:?�E,��_�k�R��zN/��]�-�eэ���:�����0&��,�{9�g�a�D[�C��k��J��X?$X�u\7��h"����fc�L>��a��?�p�V?��X]���l��F���X�q�<㦰R�F��SՉ���Ak���o��v[﫭�O.P{D�q��î͗q���66��-�����p̨T�寺[�����"���t�i�Hk��h�`�Z_5c���b��9�K�	���ǐ��S߀���--�?��f%��I�)�<������"��,��ꭍp�,G�A�����a�T�*��������p�$�e��50̴PW<��y�������*�`�?���r�k�J���~ا���^��|WG�4,���]�&�j����7�Hv�O�0���R��t�����w?笥������pk£�:���Vokws���jY�����#ど=���(kq�W:u�?g���M=���M��ד�\���Jáå��J\�K>���3D�J_ކ.�$�_���H�g?��D2�diw� #)���ޟ��Up���uNr�Y�1� P���gE��B݌�Y�*��v_S	~k��S�H'e���ѡ F�J}ߴĊ�6��'��ۂ���j�qs�Is���i"����\*	��y�D龯�{��D���[��a?ds��LT�-�_Nf Yz�f�TR�\�>�P�W����8�uV��̰VU&/hzB��J+�d&�f����W���6ȺYM�����L/����V��R�T�� ��h�'Q}�)Nx�Wp��qɁ����=�U��.ú�_�����M�)�z��9m%ퟓM�tL�
��������6�x0��X��2��d�+9���h�$��҆G��A���F�	�n:��H2y��dh ݃R�@V��䍯�&M֏��&�FS�2`8��ĉa�Q�~y�p�o-I�;4	 K�k	�?��s��v�M�y�c*���\�s�m��fg����hĂͲJL}�3ʱ���j�:��ed��Q0����Q�TO� 9�ć����1������]eФ�0B��)HH��z�dgzE�mIڄ��R�i%����D�Nٷ�&��t�3݈KC���TK�?�:���O�_���|'�e�pӞa��/f!�^=y(����u�V�����klsc?�N���,`�@/7y-���a7}�W3㘕)�%8��������o�4P0̵�'�鋮Կ(��Y��̓Y0I���0eղ����L�?b�������~��P
��ҒxޝuSh��!=5!Ƙ�� Fױ�+�8I��������f��xA�Su�.4��k�Jޙ+'@��L1p\Ba������v>f���o� �[��
�?��>pHOH����<��'x���^�������Ƹ�۶��͈���mk�u��\��� ''��M���MNN���WLL9��x��\�|ڶ�Ͷ�u�ȼ��t\����I8�n G�����M���B\��u?h,~�N�ᬥ��mNk�@��el�!�IP�5&s%S��PC_EG �C|�:�ںI-�`��q4L2�ek�^���i��~,O
"R@�S�r����Y�Q_�Q_KdG�C�YY2�+�+��`Xn�٬@m��[�RO+�Y����)_�mk�����͚Z����ҍ��B����=G��Jˉ˫+݆���ojj�����^�������{����A$�#�I�/C��P�(�X���"�7�����(�+��I�>��Fv6s#��_NzG�
�Z#�~�����d4k���H;>�nfMPl?�a������a4<i�	��Cu:�h��-��ሴ�k��|H���Z��J��ޭ��,7���\sԂ*�Ps���fu=w�Y��f���S�f[��Z{'�iժ�1k����UJ�PԊM��{���Fk�ޣ��O|>����=��8��q��|�_���u���݃S�F;e���;�Hr
j���=0 @�C�W����Z&;���Wε?��B����1����*7t6%�� @&	���}(��bg��$i��d����~�B�i� ��-24��k �7�RC��r�^x�/nn�P ��Y�������S��Q�*�3~,;�ӡ2������`�]�v��op:J�3&n?|�=}��N��L䐼t:��Cs���"�j)����U�#B���`R/�<�*?T�!9���\j����^�@^��>_-_���W�E����{#�3e��juF�E�����x}���c��_h8G��@��kX,C�c�8�� 3���䚤�.��|7�1�������h�K�&�ҏ�3�dXa}�w�7bi�
!j<ń���@�Y%�<�=��B ;u�[P97�Ii��"��<�'��ԝe�H�����F24�l]���O�RE|?�={��t��1E�q��ͺ�;{���	'�v{D�K{s��B����0����x��^ڕEU� 8����0��'���t���X4�c�*Rv�gG�p~2�	"���zpٕ;!���h|�;�S���B�7�����y��e�����m�땆�Y@�;@{�B���|�Gم���ȋ�/_6�Abuuu�uB��i!��r�_������?���L��:�5um5�3%=�NU]�O�NlcL�\��'U(����.��)��^Cr��'��yD/n�]�4�4� H��'��O����_���*xkP}?�w�T'�c��5��d���bM߂�O�������$�%�g�S+ŭ'�a!��Gr��'�)��a

�Y�<�EJmC�r�M�Oܑtu}]Ľ�s�,���L��
���㖃o����������?�_NxuY}�ooe��=��1��f�t||�[�������ej�Qi�{�El7Q��g�vF9�?��V�A�}qH�4��%�k�*-���*NQN~v^�.�£�'gQ��jgS��8�g'vMB#��qP��1�������0P�&M��M���@KJ}�Z�I< ۳�{ʮn=L��M9�:0=��A��|�o���z�Q��#��X睵�IĔc��8��L�,��oX���|66�b
��K���4�h�(��l��&�Y�Z�@�*�� Η2�WvJC�?��ߨ�$.������nS��dr�ԇ쳍��� 0����o���)�Xt�8^+"Н�r���e�7�c��_�ICO��ߨS��l��D������쬥��i�:2:�]~V_�{�-��������s�Gz���l2�?!�h;�O`ޛ��R�BV��Oj��Od@I��3V�f0���;Ģ�j�����vJ�[�[�|�I*H���Dz򤌩�/_���	�V��Y�<]�j|?��Mh����?��P����O��׵��J�k�����/}�-����5m�2��r�m8F�2��X�51"ز�}��.(���d���1��c�茅�O����i���@�N�ǹ�)rt������	֚4�]�F�X���D(�O��Kj��^�\����W8�'����
`"�ծ�̲��`h�B)�?"���z�nM!-�L��4���n%�a�y|������IEMA-�\�r����  �����IpDVF���&���8�\J΋�g�l2G��U�������6xn�x&9գ~��ފdqYi����'f�O���T���}�J���`��I��0����Mv��%;��9 rIݢ=;<�\�8�����7kv���d���vh��p��=x3M�<�!]=����^�Q�Al1�&��`R%�a��hn��V<έ��2�!�����A��[�,	J���� �a{��h�M+���b��\����8�/��Y-��t_�����-���I�Fq�(��`�3��5L��h��;��~��mhhHNN����p$ȧ}�pf������P�w�s6$�r4�����5��;w�c)ȣ����_x�8�P�@��d����:��['uh|�`&Mm���6#�l�J��?Z�����L�7M�g;�Ӭvا>����2&��ZF��O���]��*Χ9h��R7]��m�����Qǡ��YM��-=v0���buY��K����u��Ec��3�ԑ��ݽB�w_+W^�'�]�9�|�*��2����6�B����!h�B�iW����ֺ\�~̤E=7S;Nʕv$B���g�������h�j��;H��!�%�~Q}Z�;�K��Ӊ�d��(;B�sK�{K��_���K?��R"�K�����޶�6܄r��Zv�kșB�2�5�C-��ڎ��W�uM:?W����屨�ziq�0U�%��z�J /��D��.e'�a"x�Z���.qg	(�m�vIx`�j���e�$���n�O2c��xs��"�X��#`��Q�LQ[��t}=���w^�%��"��*�"�cy]?��t�	�n^!>�nC�\h}�lc� �:j�P|�z�S�p�U��;_{�n��7�^���D�0���4��^=�1B_�5�J��ĸ]��l�p�*���Z:�s�$��Q�y�3�R}��c+�HA��NV>@���~�,����UzM�j*z;L��d�a.�ֱ�^��&'^���6�˥G�a�(�Q瓮��k!'_E5w_�6?��SG�.�|2�v��[ݫ$Z��.#!��⿧��!40Z�;N�s�+Y�U7T`Ûq�Ia�9�0��,��S�����	U]+�++UEDx\]%��6F�PY߸Ž�==��La0'_��կ_�&$ �iq��IN���x��"������Զ���K��E6�"e�1+���"Ϊ�Վ������Vhs�.�Ѹ��c�R����?��6�[�D��7��Y�1�s��t̋͟�iΩpU��_�L���c�3yN|QM�r8i��ͺ���>t�@A��"]u3k��z�~�IM�nY ���gY}c�>1�$�>L�Jh��S�f$�P����e�֞�8����I{B<|�BBϬ�����+)+�� sА�0�������ud�q�J,N�k�2�W=M<6#��0;7���Hr��xT-��/�23�N��6����W�e�e>*�׋�}.h��]��7�2;�|�S��R��vp�1E�V�65HS���h��WG���5s��ړ �7Xoo�����.��vAR��g�lu��nϴ{ڛgG�j��Wa�������s~G�uש٥�AB���_l	+��oZ�r��F����##��%}�����nWP�0x�E���~ZouPG���CA���fL��̛�4�E ¼����p��R @�� ʤ	���Q"��c x��/7@�/қ��v�a�b�O�9v��c�u�"4a�j"����3�S�C��1g�����*�$S`�S��Y��N�*c�k�Z�b���L��{�3w>
��	�w���(�{5�3Y�;��qkd�M�ic���0�w_�kc�M�|�-�7x��W7坫�߭ғ_���I4I����[�h��,9�ˊ��q����lf,>0��, *&E��ʵ�!l�������z�n��FZVj����>���`�BM��n7�����r߸���u�[�ki-KEz��6�%[�UDY��Ih?v��sl �f+/Д�v�)�|��
6�Nz>Jq��7�s�@2SsA;���󩵧"���e̠
:x��Р�*ɦ4!��X�ўr��G^��5��%���'kwLv��F«\�3-5�y0�������+͑��Я����lQ�3݂j���C��ck�����ك;;:;�ќ��ٔ|2�#��ڃ�^p�F!��e�$i��e>��=.�@[d��Y�U��0���5=�ӧ*1>>3%�uGT"b|�\[�(.Ε��ry9��;��"�9�S���F��L���C�,L��%��]Q��ƕ�4bv�Ѣڳ;��c�^(����QR�i��g��۷�r��+��e4�yGt{j�d;y�\���pT��U�لT�U8���"ړ��-\@J�U�&���!6�� WlG�I�Ҳ`+����D���Z�0G��Yl?�B�O$�D�E�`[$�uK-�O���L��ސi�䫉9ΆWYt�57��#�v�Ҏ�A��	��zJ�c{�}�O��(4(M+�:��hȯ��;�g�gw�(�(N��R7z�Q��|��O&د�b����ű5t���,�����!# �|�@nd+'��s���j���WBMcBa��EP��<�a�D*`�ч��)ceJpF�&ݣ�Ug=ɹUw��R�ھ��>�..?�V���M�u39��ۊդ/��;�un!#1sn��#��*�(A���Kc3sK3��P"���֣�g�xj|�ɹr  ����{K�'tXN�}yo�$��r�z�>�B�[.iT�K�S�?��Q%qش�d�n;���xYR.&�s�f����x��w߿0I�8�}x��@j�*4M��A�r��Z`�Y
:,&���� �>�𹯃�5��DA��g�����^2�q�.$�Ys�����mPX�iEA[ >�N=�le�F�Y"c�P��6?+͗�n��kž�|V/�х�=����d Ef+w�j�B�b�����@�t�K��t�n��mE��N7�*�|R���#��rp)*��<NI=�� ��-���4�}iN��p؄]m�B=R�p5t�/OR�7��I����(�IOX%g��_P	�����gQ���:�Vx�m`�`O��Ov|��wz����� �ڤ���L��D��Hʙ>&�aλ�7�H2p],�s	�}��f&_����.���;a�oL��H�J����m��:|;	�(T�gd`�w��7��>0�p]h���æ�f�*��:���aq4�߿7xbUM"�w�qg�h��b>���H�`�hҝwt��-h�p��������0bbҋ�ѳ���i?t�{(U�=h�<<���}Φ�b7v���m�=���z��)����"�1�`>��*��~�̠�
���K����no�������ݯ�Ho*L�^S:(]6=-��ѶA��]1�J �iK�k4���T}��Wv��e`<e���O���4���BvФ?��5������ɩ���޴z������*ݶ��Ւ,�M�����h���ztt��������*�'�X�D~a^p��D�U�ϼv���J�u::�DF�y�������3��C'D��q�'+!�`h� �K��T���h���*+��;ֈs��z�BtX�h&n'�I)}�#&?]��fu�CnpLx3\.��%�;�՝j���O�r �E��'1�7��ay|��r;�ʺ�����''�����R��w�*��
���)��L�ҜGˆ�t�H.&���g���tI? ��H�Ja
Ԇ@Df�i � @a2�t*�#
���d�$6�ō�_�@�Ô7Kő޴:T����3����9,<�D@}�@�^�m�!����e(��-�A�1w��!'�u��1{Y�Аw��,.4w�Eb[Y���~L�.[��%��ͣ�����,�/���<�KЄ���j����Dw�J1Cc���9�����'.s!��la���V�V>l�󇭼�ޖ�-I���a��䰬EV�JZ��@�0ep�ฏMPw-d���{�Q���+�GLv�c�9��=~60���/�g�v9\�����)%wX�w�� �����&>`�+�����త-7���r�칡�����~@V���Ox*#p޲5�ʻP��,���1����y���p�1/��v�m6Ľ��<q��4r>���T�~"W���.�����J���$XW�p�{����et�.��l�ce;�
�'�i�1|�$xs^Y�b�RQ��҆xQh��
bWd����4m�Sa|kMrĽ���8�e��G�Zp~��0�*��!K��rFg���.�����?�8L�ؗͤ������F`�U�U�\5	�s0��8@B� ]�Ze��o�9�՚������ڏ�ap��u�j<��%h7��'k�8�����wdN�B���!Խ�%������YB�#y4����2�7�����_HT���1e����r��w�J��,�"�g�XEC�f͗5lח���~蚕�Q���t=ʽ��Kt�YO��d.dޗ�:�\X	aBB���y�R�$|V�a�é;;�lk��}(����Vo�_gQ�'u(T���<0����0	4_EUg}�0x\	)������pG擑:�9{��Ps	y�NI�Pk2H3
c1�"��Yo�k�%��IZ|�Jxl�W]r�Ĕ=�k:�6�,�Q��g��ꐳ�ҍ�]D�wM��D�y�=�ڄ�Z��Qv�T_������9�Ӂ����? �L~�X*�k]2���q���C�z�(	 �P�rGƆ��k��iB���o!P��Y�_ԙ8B�e��Ξ��hH��0=�7�S3�ş�MA|�����	�2}~���$���*�	�Dd��#7tSNkY���R�z���"���p~/��G��	'3!�'��^�@�<��Vޮm�f�̀ ��58"d�G�]��$�鱗�R�cqӽˇ�ט�J���>iUz��#I$؄
��#�;b������Ĝ�t]*����$� *�ex ����BڴA��

MqT�Ő��ۯ^�ᬽ5"2��N�đO���^'�������x�nYx!�@���x�-]ٓ�2��fEF��R�ğ�Nx�|g�c�{�=�N��MŐ>68�]�����kM�$�ux��M�	�N'D��D�>�"����`<�G���e	�[��F�rUQ��6co��t��J% �g�.�S]��I&,nq���-��#�~�	���"�B ��5c�W�K:�~G�duh���S��-ΐ_�RK�������d�
n�b;�m[�eO>#\�^^�0�h�ru���%����+���������G0�%*.	����n�/�p��/$�7�~;�C �xr��T�@�خ��BQ�F�
����j�҈��l4�$��+�����'�c1A)N)v���+��.w�]���h�)*
�!K��᎘� �� o8��j���H��`���i4C�������������ԍg�����v�a+S~���-ǔYȈ��߬��m�춘�y0��䍌!���NENy�����v0�A���Z$K0��@~&�8I��R[��t��,č����P���X3��NYRfǊԅ.�$�i��#R�	���2�j(ʹ9�9e���S�?���M�N� �����P���[�Mn�3�*2i5�P.����0��.9��F�2U�%ƥG#\K�Q"^:H�����#<�/�u��B��E/1*�%�hh�Q�3n^a��HP
.�8��4<�l��B���q�x>n]M�Zv�ܾN�g »�_"=�������������`n}��ِ��Y���7P��!G^9�H(6ʵ�p��TZ�~��5[(c0���x���Q���|�}ʂ��2�N�Y����&�˚4��+3���Њ;�f����i?��R�t"�l�	F��~�-��tT���RP���;Qy`�7|���X�u��k����q	W�Eq�&'������w���V2�0�y.���{n�L|��Ծ&;{�ra��֞��Fj��N ���͘F�o��U���D�ǻqV[���V�j��F��n��7�IX��2� X�*l�`�B��
B];Hۖ�w>�����
�{�bWo������Q � ��pL;l�}M�f#f��
ۇ�[~4�U��BM?͆v;��C�E��q�{�b���]�\Y���f*z�R�_��_��;�V}J�!��G����,#sY��gz+i�~�Yq"hz������@�g�6M_��VPQ+��'�?u$i�S3�@�1	l:�l��n�9���1>Ϻ��8�y�*��"za0�yO��W������| ��0mBJ�z��2G��j��7���-nz.� ����6��7V}��A�IM}���V�a���
U��Xl�(V�B��b�{ú~�#W�Ҽם��eϘ�7��\e
�B:�}��K�!Ab�ඇ#����o^�����&_P�*r��^'�MQpԤ�I�e�*�vO&+y��b�^�,���ob'��p��> v�do��^�h2a@�����q�j�z���%�κ�f�6|~��Hgn��~���~Ph�6��Y�}'�yR�v���ׂ�Ւ�j�蕓�[�߀��3����}}ꪪ�~��}2��
���思�jA�Ii�+� +�(���c���9���@���T|@-H�(��%'�{���"[M�p�k{�$�dcl~r�Ȭs�9o9���r���jS��E�*�霗�b�p���{��7�����$��:FVGK>�aDp���r�˷� 62��/Z?JR~��?.�xQ���0H=����s�p����	6�9�5��Z��D�����-mu2����4�鄨^�j����¿��T/'F���
��O����ܞ1��+��7rI�lTT�Z��c�N��u�����8H�W��4
c��b��b˦w���~>�g���/i7��,�9�H��;�;�Oi^S��!}��qb���=TE�RN8��u�$8�,b�uģ�Jgs����X))�~��e�art},!D����su� h�a��D�YkRwz�t����^蕚,�ܰ1nBf΋LA�\�S��'�u�����C^z����*1ّ��{�I�#�3�MЊ��[�X�M�e,��ѭ�����k��z����U�/%>���=�5�DMr��g���_tw���L>C��	�ZA� ;�Z' ���Z��׍���a�1�&�!�=XK/�I��KbN**�����v��޽&ۋ��1<���|(#��yx��5��o���9���X����54}��������O0TA������U�%�U���XY)�=q��h_SI0����۫ʟ�����2��6H!�*����	�\�ۯ��5(�TTX ���
ua����+�|v��]�	ğI��?���{�XLPLT��A�[��Ϛ���Ҫ$�R+K��ډN�bK��6i�-�N;1h��F�X���"o��S��v��͉+��߿C�I>�����%$�km5]2 �u�FJ�y�~x��6�cdi�2;B���6lll
ƱO��6��s���4�
�f�Ԡ�JDiu��ԡR�b��B�V�/��st���yr�U��+	m�\�PK�hr���L����Ǔ�����X��ik�ut��GR��p��'� ib�۟���<;�4�o�\���
X_m>�8h����j����fh�J�|��昇�2γ�R���,P�hg��L�����R�E��kN�}�����ȅ8�J�1�	�d���r|���~GD���IAA�,	yQ客`Eb�M�	�r�W�o������F�~4�j_��� ʑ,'�ϻ�Q�
����E-ה�����'ht��� ��:�IO�����k�s�J����ۼ_ǵsS �� �ɚ݆�&�>�*%��;��
���:e\j����~3�g����pa�rڅ5��ײ����BџW)Wu7����A��W��,��A�~�Fr�0n �DT��Pkz,%�#�ӄV�Z�V��ylI�9�/�x�L��*<�j�i -2��$��i�6�[� C�25݉c���PY��sP0��s7+m@��+{nUG~�0x���Q�t��Ax����ʎ�l]m�S����S�5p��BwU�Cy}�J���S.҈���B�z������%0mS�\�f��L	x��K�O��V���6����k�l���w9�^(|�$�X��R��-��"*pQ��2Fs�uթU�����o�9�����h�tb�6�O*ȿP���s5��v��R�>-Q \�)��P������$�ރy�v/�{�#����*�)M�g���޽~�}��f3(cA�Kj�Mz�4��4m}�]��-� ��%j{�!�����r4����I�s!��!st�w{?q��Uޠ��"d>S&k��C�}� �ΔR��&Kahң�(%��v��i���>�X�tv�|�z�m��O�c���Ltk�F{{�1��X!��¡T�D��oG�0 ����0m���zzjH��� H��7�Er�8�����ۼL�ݟ@0��\C*M�L�ϕ���̎�a)I����NG��>{/!T�'7��~�[oϴo[��r4+�ߨrn��)�l�G�588Wח�����ђz�}������� la�sxeX��o�T|����|-�d��8\�V�؏�BɎv��{t��BPZ�*�� �'��u<�����͌�8i��t7������"�{��7�� �!��j��ПJ��_�9�:��9� ��4	jCbh��\lXP��OhWU�,%�R�䵝�Y��G���O	���i4e,Uuّs���d��su��l�1���iڨ9��_��yGa����W��Ѵ��A�g���k��o�:�����wY������h�ܬ�����M���޼>+��)ҳVcVK���{x��hS ���ֈMגp�J�����e���;>�����c����_x�"�]#�Ȏ`�'���&߅��[f�Z��R�~s9&b��QK��G�+/h�u~n ��[����
"`;\ bBh/�Y���a���_#Q\�jJ�b;�P�x�4����f�"�Uߕ�����k�b���*�G7n�*qY�p��""$�	3K���,��)f��fm�=��=���vb����8y�}c���t�穸��G�}zO���$W*Y#�;Yz��l�C7�.!� �&�MP[���s�s�[��C��Ɠ���K!k�gɁgѮ 8S+�X�<2�9�{��"@ d�I�&�;��Js!1��|�\JyMmc"�~�ܖ��y��ʈ�Ҥ�%��nh�e����F7I|Ewy+���҂ƛ�{�=�A��8�?3QN�?�����>�vue(e~"6�Rw0�ae����z��� �{�jN�s��96�E��[n@���gNU��h�g6�)y*ȇ@ߎ��@��ɯ�TdT�T����s�>���s�#�:)8a/I�J�ߞ
F�WjA�F���C8B�R��U��O~ �{�Շ±bT���#!vV���谮ZT�y2Yi���Q�LxH�3�dCv��RE�J��M���!�C#W|Y�^dY
�,j�9%+0���*>���n�7�*��l8�5�"�z����
�/=��M[�K�	�vn��r{�U�ِ��Q�1@<I{���B1��}� ט�Ӑ�% ��w��
eB�[�A*����;�F�ݭ�x?�G��������E��=��7�
��9(�$�1H�F=����&hi%�;@�/1��ĉOa #��2������l$hrPxp���i��K���@T�5�4��45)&V��]δ!�^���jb���=$t���IT+�?���3���ҝb���U0�5n���O��ϥ$�+���^q2[	C��
�YS [Ю���8Ώ?��Ց��;�1�"&;%�t�5+V
<�A�����Zm?Ǜ��!���|�k����ww6�J˯r��CK	��o�X;���u�zV��?$	,aTSA�B	PVoG�"'�P-v�^��?h�Cqg4�H��ޭ��|��2����a	��Qr-��W1����S�"��[�=Lw�"��1W�ʯɎi5����-�^�p-�W�G�zC9��6��" ���3����0g�F�=���_^P�� bGY~�O�!�����p�u����a��M
�$���x�Z	 �w�g@�M�(ʙ��e��q�����+���p<��� 2�4��/�o/�6�ӓ�pi�� ��3�l�w�[�Zy���]�I�g^tI�s�ݢ�8"���������#Ʈ�3�7n��B�TI0�H�r�{y��ܒ��,L���!�����S�i$�
����S(H�X�Wt�� |�����N������)��ڸ���c��CZޜ��)��*�;�0T�7_�o��������5�S��l�K.(��(��؇��W����d��|��v�$c,B�`%��M3��o����/�(��TH�D��<�;�]fFޕ�_��)4�:���A2 ��4Q�ӮJ�Z3` �8HY�.�U��+�ɞ)�쓎!?<'?<<��	�y�)ԏц ��F�'�lia
*�2Nv��GсZ��;�Fh����q�>^��Z�f�̓L �-YAn�FP�.��f�_�3�sA'�l��j�ǥ)�K���Kq�Su�֑0�R��ӥF�u��z����W^��_��~~FGE�n��P�A}��UFZF~$�(�Loj7�^�T �@����M9=������vL�����,Q�[�:z��ˌOH�_r��}�P |r��,i�����1\�F<(��B�cEyK2�	�%�P����*��k���5��y��1��T�#gz��+���|Q�puk+�-P�r+�N��B�g��/|���q4'zu_�I����t��bxUm6��ٛ9O��ktz$��"��f��c�]�~�+�1s���Is�bQ��\Q7��ہ�+���`X㣲.�@����S��J�*4O@�)�>���Ejr��~{ْ�e�����`1xLZ�Ww�'a��ħ �y�K[f���{ U�� � 2�������]u�������ܭxA+������γ���p�[�*��˙C�1-�@�F��j>��3��Yp�����ʀ߻����N��2k���A��9�=?����8�Wڿ�����R��`d�BM���U�"OF�a_Շ�>�ъ	��%�U���%�s��<�"��9�	��ɵf���.h%}'!��n��c����>}����H�(5,$��e��������R��h��V%V�ry����)Ǫ�f�el��n�����::Jِ�tO��"�Ȱ�=O��b�����2���lg�nkˇY��pvO`������i��wz<Y���r�3���Ę�ݮ%�.dɄ�a]h�IQ�� mQ�B;-ci�И0��`yn~-�p�I�0
�Ck�����=]V{�/0O�FRdb`�_�ͷ?�%�BRE�� ���G)��L�L��ၯ=����ܿs�����KMO�6|/���	d�����9�DE:��y�T��1s�;M�Ev����s�m�Q�x�)�g:�����$Х���f�p[���T3T��;��6e}�?*��z!�"��B+W�  6����2�/�v��?�%�S�,����[��y~�8Y ����-��~&�Tux<���S��� ��7o[7}ڧ��^x`�,�k^{�\"fL���[Fn�C�E�!�E|�z��N����+'Ļ��h��/���m���+Y�+��I[�=X����8p�(җ*��W�/r=@O��;M"nFK֖2S��LR��a���jŢ9��?�LaRQg�x�����Nqn.>w�~���6�^c�~����)��y����uJY�4�l;��G��҇V&G�E�ڿ�_�,h�^��������H�A"R�ݏ��
3����!�xb#&q�;q�n�?{��45������센����v<j�
�i��R��/MDZ���>[f����%J
�$�#���ˣP�o)���T�{Ē�kw��J�Z����OE�����sU��ݥ`�����P�J�ݐ
΋ġC7Ϗ%�o���J�DQ�Ex��D̴�H�G�����AMΎ���ԝ��̼���U7�X�
�]?�zN���A���<f�*#2�����y&-q�(Z<� ��o	vP�e�7�<�e;߶��l7�^��6(V�Ļ��\=��W�yp�U���(������h����3Ͻ}Q�ϵ�R��%�)���U�2J�1�l����,!�҉�Mƨ�C�9��U�uRQ�תKs��y�v��:!�l��ĩ�*�+�'�_�@���b�|�����	�()�R�z������������˗/��%�/-��x�sTێf��G�R�4�$�G�@э����L�"ŉXq� d��rZ.�L���]2
�����᳴���$�y4E`.I�J�ETjj*U��j�(%2���/Q��ϙ�7��J�N����o�A'���� �:�;t1���ɣ��l~rJLL)ș��)���7r��¹�']Ro���ұ�1�8�������v�()�ޗo|/ߚc�^'�+!-}ۯ���-���$k|���ݶ��1��0'p�kSL�k��w�C�����H�&"{X;�͸�p�m�Mj��!�^��	&�0�k��p2unu�CS�Y���J̬�z�OiMDw����55
s��,Q�(�S 'U��V��=�b�H̜�M�����;��zr1��C/��d*��\�r䣥gb�,Mn�c��6���!GDMU�9#Ǒ���,��⩆g���	��P;�8"��[^�3jz*�Y�PS"�
�ʵS0�w�{fx+F��FFM���y�+�_��,������ԇ���s�����H%�!^���P��O�h��tQ8�J���"��{�H�XRFNKY�L��K��q�ӄ��=~�^�{�n�@HWʡ��l���m-���#�Q�u�98��hӑ�f�٠
�2A�y�}f`S���_19�H��\A������ gO��<�~��/l�7r��I�>e3�f#���m��EP[�D����9���q&�"�5�2��0a�O�P0�c�QI��)O$���՗�VJ��F���2*����<$$��+��jI��ͳ'I�=y3�	6.�_�CN���C�34�劰B��F\PL�_bݱ�{+��򈑗'М�\��3�~�?�EL�Κ~�,����g���9�:������v�kN1�J�,��Z�T_*|�
��d-Sw�����u��+�e���Mc�iO��K�w�I���1���Z2� ��lRf�\��cHل�n��,�o��~����ò����D���J"�tycf�!�)���%Qt=q�`��p�L��n�Ό�Z��b����̟�tVH�H��o�J��Ic�V@���i�t��`�c������oSI��֪R�~�!ģ���9��*�w_�.�j�S�f��&0rų9r?�9Bd{&߬�x���_*i��~]�w�8�`*�ti��o
Ǐ���3T���of]gU,m�\�?����B,4<f{3��`�M����bR�&.r�]e�^-��<,q���KJ^u���;�H��d���T�NQ�:?��rww��)[HI����]__��P���ШQ1�, W|��ۓ�r/HD�"3�����Q�A�$�z��N[��Q�ѷ~�A�(i2�����z�41�bU�	O-��w�����+��x�r&��_R�����5"�l\�[���������c�������`�+��[D!��D��8��;�,�M+�M��Q�P�է��R��T���L��5W�܄Ն[���$�N>.��N�|�:�}	G<�����7�m��'/��_4o�6G(q)W�!{L�Ŕ���H�.�Hn#��u={tj"t
5~}r�|K��C,�y���ÿ8?t��D�!M೾����i풍큹}}�X]���y]�F�iL�{���e>4N�We_��Q�+F��I���Pe`�����}Kj�/�L�V^%��w�N�[F������I�(Oq}����>�n�4Yy����Y��R$�SuD��%v���|:�8�_Y�	��Py�`�o��R�����>��Q����t�B���O�޾���������r �W�1����l\��49=35���%/��4�㳸K]E�Hy}eEqeEu�������eo���Z=X�x�Y8���r������ۃ�`��m
���;w����$O:;^�+Sv?
 ��w���֊NAE��W��h���|�+�:KEE,�e^[��r�E��w�m�z'Kq�B����c݋c������8�E�.��E+ǁ)A���T�VV�+���K��A,�ڂ��]�����UF2G��J 4$,�ި%S�����e����MkM�D"���E��l�HK��^�w���X6]�ˣ.%��xA��FD� "�ذ,R�F�ݰ;�xM��7@�h��hx��}m �v�s��,_#��uw����YV-��|��@��6�&�gֻM���k�}�:Rvz���`�����':cDrl%�_ks��t!U�<��?���^���w��o~n�m�G�Y�6��DF� A�ف�w}k{~���0��^,�������wWd�H��%��LTk���+�K�cgC�8u<�T?B���/�m����`�\����wu���L�[:���*	��+�����@���8��<C+�7�^���躬j�X��{|{B��6�*7�u筄�VD!�D
W!�WW�--��&����`�<iy�� %3����0��QM���Jǔ�)�

Hmt�R5��1R���R�k0��A�ctHHKI��<�����y��_��ٽ�����($"yS%xJ�*+�j�k�R��d��+�nmN+_�b�='&�Ge�j��mF�68�Zl<Z��Z\���P�Iߩ�桰�Jüe��Tz3��O�&���NN������%�����A��-J�D,.����f:�\�g�{=XY�8���nI����0��U7ּ��A�e;������2��
�fx�F��a��wH�/�>H�8�nA��9�*� %臖��%p���=3�ӣ߾
��t�!ܜBO�D%��%q]������u���� ~�5�m�*�5��+S��$�0b)OQ@�W���1���{eb�F��T�`���`!���q;`�ǯ��0�zjPG�L�_tpaAM�[3����ˎJ[R�����܌�G���\���6��0�"!p�2I?v��1՛�7��'v  ����������d���Յ5?�W�����b=�ț�c��x~���X�84�������φo<S����K�@���Q��xb��[����j���M���,V����5��y�����z�fg�*��9~�lF�T����P�Q709�ǂ�0���`��7��]�E�Lz�$�S{�����p*�ͺ�;5�Z�W��z�R-�Y�ڍY���m�V"MoQu(�JqsZvc��{Z�����I+c�#�H+��FC67# :��o6-�ߊDQ���l-��}L߃[�X��+�����$pX(�a���k�dw�W�``�㻽��6R2���(N�^�!%�9s^��#�b�ƤA�w�/*��b����R(I	�F�ˊ�}'�+���H�b�MN�!�p�PB������g�����Gʷ�F��=됞�<ˊ�{���[E���8K��6�NG���8y��(u����e\�>�O�2���O�k-;���iS�K��tBz�<UUUQ}^�ףA7q��#��j*1�6J�>�i��>���<;�D�f��L��N���N���bs�5���HR�ɒ�wyzU� ���K��6�Z( 6��w����l-Y�ɯ:�[��S<�	�
�U��S��0��7_�ʪ��7N �2-�4N�7vwg�I%*���*q�ضW���U�z7� ������fh�r�?X[�!�t��xO�Puz'��1��<6��5�}��� ��r	�
e���ᲅ��Ei�"�@�B��.%ܗ�ƈ�����H�����f���߆�#<���lz�|����������|sWG�Ѧ����Qג��Ǎ�Sa0,�}�)<7����AT���s���0!��\`&�ū��\����'a;���S�&s�ƳP=d�	�T�솫�u���Ѵ�@B�щ/h'���
�Pp����5ي�sF�K��S�p�t��Ls�:6�n�1bG0�f(OjEq��4��ς�ʵO�|�'�C���GY��h˿n�X}��c�5��R��[E��5&ٲ�9�^A9�t��Z拁�P�:O����bEÑ��<�ZI{�ZF�=�AL���+B��$艒��Ȁ+���}iJ�1���`_���Ci
w���Ӣ0������+�b`��_g������Q������s�~pZY��)go������k�;m5Y�fٚ�ꮒ�궒����j(��\'�^�Wz[��w��Y^��C>��s�5a�.�u�ӧ�_�^�v��Ҙ�&9��%㗶�>���6vv/�Ԇ���%�W�bccb&�B�9�G���"�I�����v�&Ȳ����`�{��`)�P -h,����������R�s��;���~��
X��0�t3o�v+¡l@IK����N���m�A�>Efb���>�I�D�۞s?;�ŅVN�z S�5� ĳ��_7�A��`�9g��*�=Pk'���E�G6JL�B&�дR���&�+��B�	��NiJ�?i�����(�`���qr�{=�m����nK�r6�{�BC��p��R�����w���H�/���;倉���sZ���xӣ�V7���?HN�^J�1��^�k=�k�m}�&Qz^�%>_k���+]��a*%�Ԧu������Jo�F}D_oͥ����U���hT�Aȷ��+�=���u-1���@>!��$O7K
��A��#OQ��?ۡ��6�U�l��2�>�`�Sa�t~Q4�32�dϹӣ�@��N�d��(Z�l��uM:̭X0
� g�\|%�I�|�W__#���
E�'�xEv�1p�` �`O��������Ar��G���p�	{�w��{�|�]z�yd��n��PV�|��b�?��^�z�I���\��l�JO���Z�?I�h��u�A*w�}��j����G/_�����)����60��uhV�>��ό��=3}A��P��$ŵ���^Շ\�n�)r�]r�*�^�&���������&.~PW�<9�$G���\y��{��99L�zo�_�[�
����s���Ͱ���{�/�Χ�@�T�Ig�M�IX�pt���Y_)���B���P����ޭ��Å��e���ĞH��dc�e��b��ZL�[4���kkU��;kqM��^��s�#�������hCZ]Zg+8�N�ф��r��v���3n:;.��˦��e�g4�o��6s�g�-��d607E[��/h}�ڟ͘�� -��[t~��K(n�t�;W�;� ���g���"�̴�O��<WV�5���W�1�8�#��9�q�R��#V�w����.�ޱE,hT�3��=($k��8�\���:Ҳ�J�g���Q�QOy�o�+����/�n��б����ֱ�;��{�|�r�9m/���;�9	4�������v	�@�,����3>�i�ȶ���E}����_y|���������;��a�Ιu�@�$�]��h�"�����v9"�i"� h�9�e����[�TZ�xY�.5iB�e�/�]�G*��+��������������0X4������=�DW�ʅ��U�����RHn�J��b)���S���{4v_���[�=M>�v�Ƙ(>�_rQ��Wor�J�P跘7A�AFl`�U��V}����X��+� 1p�f�O>�fd��qC�s4S��� �R�σw���Q���˴���Pvd�GV=V�����T�!ğ����HWĪe�x�K�\��`F`y��6�(��Y�� ��7� ����ϏN�����JT�VX��W���p� ��81��p����A�V��DX2�#�f���|��x���뜵U�[[�<?� �c,�.�T��Ȣ�Z�9d������H�^������*���R��4�>��������$֝�\vd��,� >H�N@����a=��q6�
������6|
���%a��]�t{�XX^���@ۀ �dw��Q�C�d%�HPPY�L6���+��evJ��sI:s�L�����+���v(���p��F�����!..�����·\Iu�����s?���L��=E�Z�<V�~Fk�646�|�mט�˻�Q����M�l�l�lE��h��-9\hf��
飂*֜�zҌ��$�D/jk7'08n�'
��N0���<�u[�(?�v�Ar}[t�F�޵��U�T.,<�7�:��H&�&=:�2�./�������ͻ��7��Q:07��|�(�>�z��՝��ak�S%��;h��A ('���\R�,��YW�Ӥ�崴Ug$�7�Z�OY"���nI����C
������D����6F�{�w["�"�&�λ�o坏V�8u�T��#�f@��~�2�?�31a`�3��u� �a���T$0���vL�6���u�T��莇'�n)"F#�^�.�wO��&�Z�DX��8�Y��4)��Q�I@	��qGzy�������.���M��z�W	�)�V_^���,T&�|�4~m����J�� ZQ
~̉��WN���|�B��d�qO�pi��="5�i��`ڜ�EN��~`�Vt�������rz�y�Sk���v�΁�o 	`���\�[�*�f�[Smar��㮸&Կ��",u�7�ʯ���i��=���{א��{K�K��Y�Y?��e����r�����ޙ�A7��L�R_�N���m���0t��L��,x����["�:�}�xY,R[V�{�o�z�Ն��&�U��e���(�a'J�/����%ر��3�]nUxIy4�����/U@/6I�%�M���IQ����r��ȥ��#�R�G���
">���g	)x�w���L�B�|������]���֔f~t���+������I�r�0}���Ybeȷ1=S3����h�ǒ�%�K�*�!;p&_�6-'еf~wN�{�@��ô�Qd���kh�������hl����Ypa�b����
��p�,g�����+P�Ȃ�H�4a��*ώ���؈��cB�ȡ�~��Z[��U�3ư���"u'6jPGC��3D����o�������vZ��繿��)&`���MZ�R�W=�EFP,*, *� 6�A|L9f��'#��x>�
�`-o>g	�B���qhƛ�+�ǲ�Lq{�Q��};�S��yƜ� ��^c%�5h�:)�jL�yC�c6��,�o�V�/g�$����mk�b_5���	�R���
)^�3$k�bߨ�Fy��b�O�Mş0�]��T����v#���O���@3 ���C+�e.���9����f�Qk��m��'��-l������&�+���g�ZS_b�@��.25@��L*1��A�����M,�.9.���,�t�����X^�0)&���v���B�؁MX�1㉔O�66�y�.��&S��M�O����MV|Sleg��pF̀F�5�NҦч=���\��\F�t ]DJ�������������Аٕ`$��1��5�}�"1�F���G�7��L�n�����:��]`�jZ��G��݅�O�:��p���{�����ZĦk�W�q�N8�>�|Al��A}}\F<����s�Y�֤&Eߨǵ%%mL
%����
�-�!�-\��j�)�/-A�	�=�M����g'�ݛFFRhSp���g5�|B�	��Е��0�GM�-g��Mc=L�I/�{� ��=�>�	��,����%�VP��e�+�5��<g�t�P!�#D+T�Ǭцe;V�3Uv<��H�Z�GSj��n�D�;l���/�i>����g�C��J�$�1`CevP����F:B������,b�-��ߡ�<��[.��7dG�=~/�=	��B�]�Ix�ؽ�����*�[Bʗ3W�B�g�N�ߜ����l�75L$\�ְB<U��OoQ	�G�Kuf��b=�j�����#��Me��Ӂe��0fb��wY�Ļ��A�M������R�0<�{ν1�G�TБ��N��=_�(���hQ�v4�?v>���)�VehFR��[2�G��Z;@�����K��!6¤~
�OҊ�t/�U�eӌ�r��'\9����~y
n�;�����Ny�����	�6��Tw '�d��س�f�U��i�Y�Ij(�N��Zt�uj���B�8��,d^�5��;��LS�#��n�[���Z�.�������jZ��p��[>A�,�bL�":�]}1`]z��{iz�1Q��M�c��v�޷��E��Z[�C?�3Bł)w|������M�/{3�Iٿ��tV�lx�J@bg�L��-$�����4�iü��B0xP��̎�;cjK⥜�����$�B�uu�l� ^��Y��$�;+��xV�$X�Ld�~#�I���c���E�MaM�0���>i�5�n$���!�qo�?�����d<\��՞�:�颎ҟ�mv��i��4���=��s��v������1pR�O/�3ȕ�J$�xH!� v,��fxU+�U�+^&yg�5��>�,GmG��.Ӣ!�1�6�ԫsT�Q_��T�7˲�̊�Рēa�gX�n��Yι�L(�q����>��چ�`�����@�uڅ�|���I�N'ST�2*�?�]��ܢ��i:\j��-��q���9��Qe�����$6hq��J��(�kw�C�'Ӣ��*�/׹����v��ߎo��3�f��އ����k��g��r�X��hݷ �1k�y⡨vA��#,&>�.z���s���bx�2>{	����cw�$�1��R��TI�	ᡬ�{88�h\�mSI�#�G!L>ȋ��3�Hݳ2���Q jj��;��+eyܣS�~S�n��ZhRT,)푖���в��uO^^J㎯�#�3��P��?j�
:Z�ݨT>��Q{f�'�p��X����vA�.RBI$Tx���2�uxJ���V�wgk�Ώ#Gǐ,�%��G��-���Ճ_��狹�&Y�����.KU쵞�V�$�u�`��\�l�#U������tjX��e���d�ϒZy5j�[%Y/޻�}�IL|ߜO��4LfL~`+gE\�r";�=��G���B�K���Z�BSHn�X�O�h��؁F � (jΝ27�Ry�|;�A6�ʓ��1^&���#�N50}<�>����f�~�;�Q��hʜ�8f��կlUkL��p�@;���_f\{�����r���I;u����pa4n�G��믞/�g��zN�4�F~d��N�v�lY�A#����`��=����`B3�Eg��j\`B(����-����� ���x�ؼH8��胋ᾯ�#-�8��>=��={/�+\����mxܻ�D��:*�Ԉ'��a)��v��!��P@�j�N����="���o������n��G��i�$�?�C	t����u�i�$C4�A(8pT*���*f�A���1F�a�G�4$�|4�@:8�^�)�Ԙ$�Y�a8B�,�������_0�|�ЄC��X<�Ր���0HDY?CQ�����x	�t5��j�Dp��t!����$Y~��=��{��|�QNA*�G��ݳ��QF%�p�8�����Y�-�o�eV�4���vU��^y�
 �O�	�y���7r}_���˾:t��J"xsO3�6�]�뤹ʪ�߫�ec4�\�|c���V�hw���2i~��ѯmЯ�F��#*���:_�3�`{������Ҩ��y�{��bࡴ��N���M��K�=3�_�N_����$���
��:Zju��r4�����r���,��&�p�+�$�BWX���I�i�I�֨�2��%��s�)u�lw�ܶ�j?j㩻8"R!d��0�D��u��R�ZA�������|�^�Ge�%�i�g�ɘ�r_���,��ƺ�(���H_�FZ�`	|Ke�4���&ҁOl��(C0�O��|����b��diB���=�ar�8KAa�!K2����K�϶�~���z�r�C ��c��A�q���B9@9cԧ��`#�&����ǽ�V��:��q�e�J���&��[���Ab�T�`,_������EJ�(-�}��e�q���O<C/"9�i����ް^QBe��L~vDx�đ;���9''{�E���n���( �	�M|�T����+�wp(\���rT6	���H����(���bv�����v�d�qF���{�k���}�����$��_T���>:�);�m����_�y>t�y��u쿞�+�Q�O�j��j�����8�DQ)�a~�b���t�G�`�T[�8W�a�[��\� @JI��2��K�	Pɟ*��oݝ�͋��v�?k��)�&�DT�}N�D;"�A�,���T���(�q]���QQ�v;���Oϕ��Q@y�BԖ�ɏ���L����� 5֜Ql�(
�-��<b���a�'�(��!t�x;g#��m�p�5,�҈u�T������>#O
�"�[x<�J�{%g�1�&0���z��C+M�H*d�,{�=�''9�-��-xb�YD0qY�_ƒ�����c"Xװ�v~xt�3�(�ޚ7"��E=���!z����P�Rر�vW�}�N�1��1t'8����{d�;W�<�q�����Z2}���`P�,��.D����(�b쪢��b�=��
��k��Z8�6h�Jw��0so��\��.���S���'GA��Q79s�j}2&Mzd��E����P������c�{������KK�YY���x$��ՃD*f�R����S��?�_�A�R���&7�6�� �L���ڗ:�~H�����`��
I?�f��8�u~E|���Ѐ����9x�H�t���[]=)�'T����Đ��֥yz�����,�U+	� 8��/v��b��\y��3ˇn�M��TE�;"Ma�wd/��CdpW�Gy9�3匶<�`�|�qn�h�Ǿ���=����"����É㝟vY:;�����5}��g�(.�����x���?��1���:�Ǡ�a^P��L�a�xǩ�i[�l��1�yHC5x���4ޭj-!Do���$�{�A�T=�ص2~�$~���������4H\�̲�ٗ�i�.{ЄP����=�Cy�+߫$�{P����B߿����8,�9�H$k��	�����4t�А�3�7��l`z�g"Wp ��N����F\9�5�Ґ9�)�%ls.���u�����N�o%pp���hH�$u��p��(u�s<@�1s��� XT���,���x+��1&�괱��R�F�2��`:o�;�����A�b��&z���\^�ȓFjg��&�
����g#y9�?���T��3���N���N.HD���^jb/��s��./�s�@�ؐ��,���-E�N�����e�؄�}08 �z��:�T�֧\x�	rmn՛}),�Wp�e\�	�A˹��|D�q���F�?#�٥"'#�!vg�����$~,�f����C�quB*�k(x�T#FaV��N\A�8��
����� ����C�|�D�:��Y)V����S���� �����Fl����~dAn}�^��౏�,9�'��Y��UF�F�����6I�Y�\����������(�T_�'jd"AH gL)Wt_F���:�~��U�h_3o;�㜢�?�r����̻��ܪ��j�ɴ_}����3��cjW�3�������4o܁����N����ZǶ�Ǫ6Oo���ɒ�p�xos�Y磚�wʔ�	���nk�}�kס�u�؎�fZ>ؖ0����3�w��{���7fƇ��W�"����L;v���X��Β����ތ���W�uS�ɖ�8_�2y�i���u�ayo���8��/Хdsk����Z�"Us̒�j�#�L<��'#�$$Љ?$� �q#��Ehlρ�! K�m�r?] Lc# [�J�dk&�+�h:c���o�����C34�`�(��A�L��%^�]��� �ٱ�4|eHf3�Y�qz�������=��\[,�434�=Y�j��$J�ڿ�2�4�4�¬Ŀ�ujeP����%��A�㽯�-�$e�$#� 򁓻N��n�I�`D��"k؝h�\9G��Ro���p8��h� �h�}�t�@��
�F#�q�@G�>�ƴp��<�7T�Bt�����/��U�|@=��d�f�Ȱ-l��"w�V��;:�������{��`^�v��۹�URum��'�&iO��-�OGֆZMA
�*`츠�#S<=�J)L֋_�]�$�>O1��Oz��*��1�w�7o8��{��-�Iގ�`J�0�g�!0�d�%-��}�aO,N0z�B���`�"~�̯��o�n�����D���� Z)J��փբ��쁔�Ը���B�,�B��Ē?%υh�~�_�&A*.8Z�[�,u��jt��Ub��)#Z�� e�/�T Y�G�dG>�`�Oń,䶹8t����'-G+%���RI�ME��u˻!��ɞr@X��2,�5�Z��`��Knz;�#M�����y�������ʧ�q���}.�����ҙxZ@�Sע+�0�j7�3_៸����ᮈL
8m��H����0��p����h;�)�n�ys��[p
��=Q�=��
w�\�����z���OH�py�}��sٍ]�7:�q��䵙�X���n]�J�婯L</F==;�FY�MҔk�l�]�_��X��W�wu瘶��l�A<�K-�̢oO������T�]����|��f@��ѷN�γ�W�����K���_�7��G��DfW�]��2�{�W�>~�󼆿T7�G+ظ:X��d�5���)|��{si����Z����c���n���W�ZW����Y� �q��k��0W�ķ�_4�"�DƴP*�ɈJ�d{�庰f%��[s�jr'��& _��l7���� %�,T;������.�R%o�r�+~)왮4n���g��s.�i��	i"���쎆�D��Bؠ�U��Zm�U�Ÿ���vS�F�������EV^5[ī���d)n�%�d�����$��)�I�"�"ۈg@��4���e�����Sv{>�'UÏ/NiD��*�fw��������~K�p��^�/h�)�P��AK_��݂.&���!�'wh� '���Q%_0v��,G��%��*�o�O��d~��NK��M��Y��adԏ�����f�V�͏���O?3��-?|�i�X��B]���T=�����k�&vݾ�QN����ӂ��[+�A�ٲ��Y�@����j���q�k�]��MGD��	���JS�B��B�<~���YM�,<�{qN\�Y�������k�ͮ	2��$~'A�*XR�����*E{+�������3�Xr�,��ҙ
)m�~�F6,���.a	��g1\�[�ि,Ew���ƙoC���<�k��9�T���X�e�e�������w�[��ߔ��m�$�r��5�3���4OR��D
�G��6�#L�N�	�k[;A�1���=H"tN���~������8J��7��L#�K��J��?vO��~1�i�U�����φi_�pu����?���ˍ&j磻����~���_е����u��֬h�G�Ɩ�U��{-Qߓ�6}֮`!nV�	0jf�Mz�����k��?��t�. >���|�P��F���Б/F�8�
��9me�S0WG��*�{�����x<&���L�������� '�e���,�p5WN��{��-�w'���Ļ��o�N�so/Ӥ�*�o6�n�d�7�r�K��Yn7������;}��]����C����yů����1'���'�r�����q�[�`^�EE�'QhB��픆�}q��g����e,�矤Q{�H�M���B�޲Qkq���u�W��g�q�=���X~�3e9-h?��s�:�V�\�0=%�66Uo.�g����C�%H'O��.!Xw!�_�/.��+ϳ���o�&ћ���0_���~��U�۫w�G]�����k���>�Wi��c�S��x��V���e<f�?���z��F1��QO���IyI,{]+c�8cG?���8��Yj�1���e��a��cȱ�ǰ��֐��j�`AQb��bR���l`$5���������i��0���nlM���.�����{ѭ��7mM�%M� @�r�/�¬�WҨ�������+}h��@W�V7_1�*<��	Z��)(
�U?�p�[1�	��x��L�p)���W����R.�1��5Y���q�!6���yO�{t!P����˅W%f��f�=���;�ႝ���N�"���oG�0(ÃU��v�y��̟�'�c�Ǟ7:��	�	�mR���M�]�]���y���q���m�I�!��qý��_�z�T�&�(�T.l�`J������E���
%�8�t��y�i��!m��#�z$c�1���/@%['Z35���9x�����,XW���S�4��)��½�Zv�8��i,t�����:�/������~��Y��V��k'C�N+YO��#����S�%��G��_��d;���>��~0�0>��C�������gꅸ~��H{L��D������/�-�5�+�]��x���!�!���9}X�����U�d�c��RLvB���{�}�����Il�T�u���B��BBQd��3�X�3�6�k�q�]9LU���e��t��r�y��"���o���2��zG�;Oc߱���q<	������':#�]gr٤�̖ ��Gm���]ߘ�jn�m_>�HNM�`�b�MJ|�&�.�+�L��pL��R�=�����q:"a�Jy~��M?ck�8�D5 mKҠ�yg��Sn,
(��	/�$��f�G*)�,}��dV}��ĕ��-[ˈ�pm��BQ���I@a���l�d��<���]ɓ�w�n������w����� �{�:R,���{=�*�1�G�|H�ڰյrs(��X�+�R�lc��õ��`,����j�uƞW��� �fQI��b�l�1�4�8�cm�a6"3�P+6��m��bT�H��<���!��Z�>��I��Nȯ��]�;ӊ]x��8Bҏ����Ҧ�+kƤ���E����W@������7���?�5�j:��}\Nm�@I�$\�����a
SNK��i%��`��ƭ���~9ڦ�6a��m�zGm��b��=&k|ҀV�aֱX�E#�����;<����E��j�! ���o'q:0�|?5��-�`$�M�
���j�܃�8��~f!�<��|��Hy�Ӭ��f
<�A��p��*�.���e�2�F}��H0B�а�Pܟ����*��	�	T&�OڶE�(*�3���(�#�t�1Ao�ox��q� �׎���w%�}��	�au����Ψ�»sE�����KO���r�������yS�̒10D1�޿�+~�Н�������<��p�!q�H(6{-�t|��]VA�(��ހ�D�ƩR5<�8��)H�HH��X��Ԥ'<�"W�m=����
��1
vb|="�{�~��ͥ^��*�����$�d*qJ�(Xa�h_������dM�G;fw
Ho���e�0�&"�b�ʟ��������$z%������A�ь/G�\G�����W�*T����Ʋ���L�ɽ!��������� �j0$��dg�j�i�]��ja>$Z��b3�+D��<��[���j3�tC��{ǵ=26ɺ�\���,��\/8��]����AÊ���z�����S�ˤ���č�O'��e.�8�D����-<��ݖ�^<~]v�������0���o,��_]�WV�_���|{�}�/��P|j���2D���-�g�e����	��w�:*���[����>ͥ��䭲tu�ɽ�Ι��K�����=���/�uGoUdeeel,�f���� �P�l:p!3��n��jd������Z��j��`B�+�"��U\I������m��0���a�����~�w�&�P���p���^a
9��y��3ӱη�<�r��a=���
w�WY�ܧS%�>����9).��s�5ͭ�Ͻy�m3_�2����:c��Sv<>�X��R'�R206�|�O<��e�y��A��b����XK��z���f���$�ö@r�|��4�&�Cr'������4��z����N��T�N��U�Yu������Q�	��@ＲG����(�����t0qR�tKt�ח�U�ix�����o*mI���3i%�2�yU\�o^L�����C���������	� �����^����ϏL*s:���7wb
�$��y�,���.u��lv���[�#�nBЗ��w���G������������1�:�
��5���u����z���+��������ڼI����)x���/yA�p������# ���I:��\��9R��&�Ő>�F��C��V��]�9,�����$�k`��(��'�Ƀя�����-Ǐ˺Ӎ_ӧQ�F�ы�#�j��H+:�IU荧JO����ߙ�{0 �˧�^�b��D����gf�+`n��$q����9w!�Y�T��u�2j9��𵝋O_���zfC����<u�k��%��DYeu8��F���CF嬈�>�Q��>�:�tן�]ːi2ka�� ��[���-��oh��?S'@?�%�� ��9�'"��D�+L�������6_z���nΚ��3�!�U
�/P\��4ZX���"k�a�L���NT�RcF���]_o5t�3�*�j�ᷴ�j|�"�*�����W�p
Q^�n�ִ��K����r�$�$�Y0��dy�>u7��k���Ǧ^����n�M9�0ί�*����V>q�ߛs��
D߆{�a�߲�Z��Y_�+^�0�58Pr�����SW%ǎ�������������¯��β� T��^�aT����Ѳ���{���F ˹�iLɏ��2~��R��>8:X;8\_[�9l
�ZnD���&�Ӷx�g2��wk��G$��j>6�?ㆾ�\*�����K.�LQ����ꓢNݧ��������A�i�,����+׾�x����]g��d���ρg����yp����ͺ��q���!Q�U�3e�ͦH���o�nN�]M�u�]_l�ܨ�]�~��4��w�Xǟ�����&�͚�K.��'
���ԛ��o���<�`�s�$;�a٧~%d!!�%!���W>��N�TǇ7�e��շeRk��j��h#��#j��H�>_u�$��}��'d R�`��W @#�qګ��d�m���n�r�3Ӫ����f!D���666���΃؁����7�:�F:#?=i��Z=�MI��F��+oN��^�?X~Tde���2n�4ٝ��"��sh���ks����Bڰ?���b�g��]`��γ����?N��\N��+u�����b��-?���U�&M�A��t�b?�ZG���C�MWZ�K>��z$�;�J0�3�^��)�\���,�z��Y���I�IY��s*���͏�:37��n,�I�H+F��^�sX���g�oZ�Yu%�(����Phak\u�1�.y?;��&F�R��������X/*�N�����-H���1)����ܒ��l@����OW���o��˼=1�.^��ݬE���fi�@j*��Ū����!�Uk.%�6} ��6e@�s�݁�?u��Ց��q!���c��U0R�$�=m��ɫ=��ݟ��Еh�`_����1o�=�f�Ї)�Z�n^X�ޘޝ�+`��_y��*"YPPa ̬��:��(�@W6�����~Ȟ�t)J|"����vZ6�^�F c1-^�j#�G+��%���?HWD�^��' ����B5���8T]"�����Y��88eq�i<7��`!l�oν`}~�$�v����}V�ρN�g�O�s�yD�p��]0��u���i[�<ۿ������i
K��ɭ�jwF�#De�58zЄ�:�P�&.�툨Q&s''<�R�5%7unqvn�?Q�gm�j��B���JjW!X�A\����M�߱'����`}�������1^�����H}&�Q�Z�e4yV�½D�"~$�٬�Yy��Nǿ¥w�g�����!�'�Z{���v��@2�\��Y)���I���=9�O��3���<I��:d§ؙ�&�(���(T��Y:j(�����W����W��l��VDeT�:��f���&~�}H-�r��Gi��[u$�uX�u�t����ꡨ�
w�U.6�;��Y־�B��ؠ�E*L���l$��m�P�n�2S~`��@��Ȑ����P_�l��t��b���Iݜ�@ʭ�s����ѣ�~�o�gN���ƿY�[i�~oj���=+��9l{����N���S��?́7�뿺.��/ϻ��ﺞл=�f�J{w�����߾���<�J�Ɉ��x��2.�X��豈x���z>nn�'��A\�q��o���ݟ���O\�]�.�=
��5���^d *�f�v6 �(*_caI�Է��)e%��P��
����
�C:T>lc՘�%u>��Jx��}Ct�����v�8�&Z`"����3vbmS�[�a-bDt��u�͏:N�-W$�	MM�u��7N�_�FW����LK�1���'��Z��ˬ��(�u
;�>D����ce��-:<�*7=�*%y-4/΅�,�o+��{.Űm���Or��j,�#�����d��=��A��(��B���m��v���-����v鄳ޘ8�A#��*AZO��%��Y�P�t�6k�h�nk��=���?����0-��4?��M��y�a�iXQ��d��^^�]�=�健�ô������]x�4���������Ʒ�vN�Qh-h�!�^�z=:�qh"�����0�2?Dee�SN��Z`L>g_���#,b{_)Z����r��ځ���:��6��$
�0�$$G��(�� �5�K@�K@`t�tJKHIF�Hw7���y���������|�O\�u}n�⎑�IdEۈ�����|Ĳ;x��{��5�U�ދ2$�����B�|E��ċ	>r�p��S�H*iI�����v�+z�O=�	��!��X@r$�0�����4��Q�&�f�ե=7K
�8�f�sE?�VTë�;Q��s��X�_Ĵ�M��+J�L�Z]�@A ����g=cE�^���]�,yI����'i�<���zpບ����Z���k����p?�����!�� 8k�����Ԏ��:�'�@���?XB�����arMB�>j��Nx
V�[*�}�I�z��ƓS�SY�T[�Q)g�8y��V)��)�]7(
m�i1O���P�L��ic�r"������c��.���7�P?*�T�HO*G���i|�g��s=�a=犳����^���]�M�I%�J���0%opwp�x���vZ�u{y��=,�{[H���z�$��n����ھ�t=�vS`�zO������ں�۾Il���LW��[��v�s��y�j��	&��׭��,��dE��
�5E"D�2T�:���6j&��UTL��qn�5��vݞP�8�w+�|H�ǬeEn�bv3]��?�𙭳�'`��Q���Wk��)�cKK9 �RY.�4�ݵtl�g�~���7W�w�l��{OL�:�!���mh"�aD}�a�o��L������X�ι��l.^��=ɭ��%�G��<��#4��1(n&�t�=�|F�g,��G�	o_���ꬑ̔�l�uSRumFS��B)�/� ������[Q_Ȩ�z��b_5e� �J�;1���O�ԟԢ_ )�,5gx��;D*��Sc�P�
���qL����-Q�:�1�j;'�B�@�"t<����fb�l�������~%r��k�_�z������c�1��8�I����ᬹ�q]��r������r��(]����4�]h~���'�6ͪ(EU�U��!�c��E�O�O�m?2St�v_��x\ٶ�4mI��"����b�><�-�{r�-��5�K�!�t=c��E<Q�y���*p�;k��{���#�)t�5T�0�@P�e��]���Z�<��� 7��\��H�9��>P-����:T&�S�����@,���K_�|&ϐp��8C_���7��!�I�-�o�;,R��]��¿����s��Va�T�\���)?�:�5��5�[��]*)���$���yh��|�r:�����M��N>1,�~��5v�	-�Lm�b���M尞��h�i�RZ����r)��5���K1�+�1�_�u�e��KU���a;��<��1v�O�Ø
D������l�x���Y?���tuw;<>"&!�ʇ)��3ȓ�hu�R+�����.s���9�5Ƴ��t��]�jnoj���\PK�����g�b�"˯�s���������+��er�����6����}�}F����Ov�9����r/���n��,��!z���c��������1�ĄG$�����'�N�l2��MՁC���B�O�S�9zK�K���%] �˔JE���j�PTC�MD���GO��݊8���3�[���7�H����5{�r=��7�n'�b�5�'Kw�GU�3������zs�f{�ǜgCCS�)��<�zRY}RWؽu��&�j^7��n������<���Pq�>Xg[n�U��R҉��XW��XH4�_�mf�f��l��sƱ0]ݡ��5�'tuy�K�ӪZ<,Y����@D��?�x��[X�Jy�n_+�Ϟ�`��u�|k�2�Jo9U=B[#�\��sZ���q�� «������Ӟ����,G0��T��i>��|�<��;�^S}lj���a���>�Z+� �ު��>j�>��ۆNͪjNi�"X��A=g'���m��LK�$��%NIͰUE�8Z�������I,+\�W����nH�����|�����[.����laد~$�f3��7�6��g��g��i�yfh% xl�%B�����!G��UϘ�<�eM��lПgPhW�I�a��KC��w=i�<�x`
l�Z!t"�Jd�F��E�%��֛��!¨��
<z\��p
�?�y(�k(%�28=���^���
�k0A�F.X��j�bp������b�k��T3�`	F4�,�׻�K���h���u���C�:�~I�b�sg-�%��t�v!#䍎;���uԨ������3gs_�r?l5A��xm��U��7�Ґ���\��.�f�����f T=��_X'��FG�U[�VF� T����
�6Г�(������c�!ж�/L��v�(�5�4K�.������^YZ���K�����^~�������H5rx]�wAM��;�͆F�dNk1g{��1:���r�?"�g�7W:{
ܠ8iq��������A����b�帲�]��5rS�����f-za�?��v]�]�X9��/,VE��tF3����;��!����	oR��[Zۺhv���!���NLMM��4�Nu�IE|w�����>�Id�T�h���ZU��[/��;X���.�5-�U��(�t��
2���U�i�N,�"���4_���u�ۑ2��#���&K� ���C��2Z&$j����G%���%8���1�Y
�����6�j�i�q�q͟R��[��6�*�Ɍ}�ޫq��r��t���>pR<q�{��O���m����_E��C�r2-3D7�����2i��iG�E�8i�0ʉ7���~��Xk1���?���@�߱�ԭf��lе��C3�I�уk�"�+P���(�O�ZmSrx�1�{��`��W��p�u��?��R��>n�Rvc�C!hJ�	�Y��X��O��Hx����Q�t�ז�Cxń�X�����ݕ'��*R;y�
�+,0��V~x�����**�6�6n�׶�\��:AT�,D%������9��r��Hc�H�>nO5,��+O0�́-�{/Foc��+F�1�zbO|���(�Q���sp4�����P7���z.��lT����y��Gہ|&V�X&�Z�x�VCf��t�x��0;�b��i2�e�:�Jİ6�Y�c�dl�Q�-���!�����0�/{�rЌ��"�"!�!�s�������	�KdL~H���u���Ԣ0ś�p�71hbS���oa�V"~��|_�#�(|��¬|1���řҴ��0$NF� �&�X'\e\��M���E�6���!Z����Q���/���an���<C���kR�������]M��y�]3*�{4�ܜ��OB-}֡�dO�oz�3���G�n�n�����:+q9K��ǍYF2�'���n���g�W�}�$���Vز�{��_Y�����mX[o��QZJd�S%�`��2�U��3[�k;}Vt��pxk�M7
�i���?�HH{�U�湎�ށq��mƱ:�pc�1���d�u�!��U����GL�T�хZ[U����� r ��J��ov����j�y���QH��o�?F�7�~��/̵x��&NE�H��6��Z�W�z���W�+��h�l��H�U�y�]]���Di "g떅lb�nj��EYbZ[���+<�5��ᇒJ��;?y�|�
�k%�hd�h'��'U-�[f̈!&,w.1�_�Y�(>�ﱊ����z���;!^ Q
�`"��[.p5(�D7ڗ�����K	b|e�_�����MHR/y\/ylLed2�%�qF�5'Ͱ�"�l�,RJ��.����/<�^��g(i!XE)��n༑������`@Kء8C������*.y��|�փ_3}y�TNx~�q�I� ֏�ݨ��Z�`	�GG1D��piC�Yj�C�;Q*M#��V\ ���4�I6�D*MSYVW���V�o��j� /�j�hs������;j"S�3v�>o���\�&C�MP�I�W �ծ*�*^�h��tQoWZ�������*?�\GKR�(���1��5�> �*eѸL�Z��K��T�?�`��d��˔`����)߰�J�"���H����Ъ!�+D���@�~��x��=��&�xC��H�`<��Ϥ&iLe���A�^��m��PSq����--���y�dT��۝߂�`��J=(.��~��=��HCk\/��C�HL�t��dcc�m��C��Ψ�1�2$�D!����q��Ґ8m&Ã;��L��d{j'��	A�����,1ߢM��_�ήr�xMw�#m>�d��k���$�~���0�{J8n�Z8�r[y�jE���n��t���������U��]4��S9�z��zb����g��_\��q;S:JP�8B��_�g��2�Du�8�q?u�bY:��ݺ(�ʼ'�9�Lw��J��!վ�O�@h�*�۲]�֩��n���ʭl���F��e6/�`Y��'�C#)�1222A�E��_uI�MO���� [�ξE
���� Zh���z:�<3�SPo�w/cvҞh���f�ὤ��g,�z�4�1ye	o3���$K���|w�b��6Ň��1N��$�"`�k[�W����ظ���#��������Éu�tEw��-Ie�2Gu��9<��p��I�Ba�a*�aE�Є��Ø\�R�X�	;^_��1Ԁl�,��� �Ȣ ����)� -K%@T�K̠v���`��؞��=x�b
V6ѷ71��ӗ�3҄ �	Y��m�:۟�,�xrw�א]S+}�-�)�����OR`��N)������@E��nLW��q+2�iƉi�i�4�'2&{�Z�Y*����<�0
�`s��|�M�EO�}����%vt�6ѣIN{D���ŖU3'�ܵP���7w]�WŁެ�MlX�jE���r;X�t潏�g=����^� �R����r���������kl�E0���X��:��TYΛ+A�aG�tH>��E��n�S���q��Z�������=�/?X�B��p!��a�T8B':/䭨O�7(-�aaEV�,�*7�v���#L3Erb3$׏٭�|p���&�X�A�x��T,)��⮵��+lէ��:�&-���&�h]#����B0���4;o� 5��d�{鳦���FJ)��i'_L(��0"7��%����D��@�uܝ��1Ǿ��l�k�����������0��7���������o�%�n;�o�0=�1{%ߣӾ���N��2W�{��cc�
e'u�w��;l�P�*��vh�Y��*�9���	L̦-�xz@In
���T#;*Y���SV$%YP�*#�m`C;J	�����m�_�� ��OW����mU�\Ҋ�d�m�Q��$���2�[����c�Xk����������u�و��?����`���%,p\XHDj*�����iԧ}"��Tҍ
�&�J��L�V���s�O�z��>��D-�v�FP�5�in4�H��S���3?.��,�}�@�W��& ���q*�y�:cB~�R��e/�e�⿲wa4c�W������a
l�wS�6�˚��.z��9�G|�L�i�`�/�@x�
�Y�#�CMVX��N�X
���|p�|��/��W��4�x��$��YK(�	��M�na�ޥ�m\�]�b��|as���*b���;���Ag�s��3�Nu��I�<A���@S㯿@���L���e��.�w&s�ف�&5h�FɑK��:t����G�0��?�K���;�ZZ�Lj�S��g���&Fhkd�Z��W��9K�_.YB�]�*_4<U���%�1��Ņ"�w|TO%HE,���[�;Vy�U�ruBF�% ���	��q6�+����A*X,C�����E�EH|�x�	�[�/FXTX{#�3��(򝹟,d�Z@���8�F/�^�j�Z
ED��WR�?,F6���R������0��O*!���� c�j�R�]4��8F�դ���̠��0�g�|;����U�tL�`K�w�6�9l�c8@]u/D��0�S✔�������vMӗ\ �"6�I�h���\�Ȝ���ړFٛ�^� |��p�����-Q����	���;~���F�%���a��6�+GQ}�v��r��{0'C�����!���ևl�JeO� ��\���Q��L��	�Csf�K
����Do�FYK �s�������{�O~6?\�z4�kx^ĵx�x1�m�?t�*�P��O�:l�~j U��i�odL�my-m��m�������j�p+�J?h�KD��g�eB�>���y�����3��
C&�,���b��V	���^��|��Lb��F$^�ߝ�Щ�*�]����L��\�ޟ����H\�s�]��^e��^�K�����2��7��C��Ƈ"]A���
����N��#����2��H��"3N6�Ԭ���a�������xy)�Y`���F��hWڿ�	����'�~[�:����0������Ԑ��v���N�v,|��EM��qy�(H���&2c9 ӭgۈ���D��"��.���VV���ݦm��ԤO*�}'���ܣu�u�IM������b����dbA0��(��ʆw��WB�w���x7~'���~[G���ei�h+���χ���	�U������M, ���BA��쩗͒i׾R-}��"8������u�ۖ�YV8���9�̣���D7| ����3v+�L��.��%�m��?�Z6�*>���3z�]���2[�F�#���n�PBP�JomT#�� �a�x���	�O����[���C-ܥ�*y5� �֘�˃��oh�- c���NP�_9E���#;��!�Q~Y���J$խ�a��wN��u�L�+t+&?C�����j_NZ��y�~����XB��YXHF43��6Z�5G���6���m��IP%l9�	�|�ִu mʪ��liCxG��~V���^���0�z�����@�ڐ@1�O��K��#mȡ��*��yt#T*�^���0 �l�j��UP ��yD�!�\ț�����s��h ����_?-��q���q��E[B?M4�C)|�R�do�����q��7H��CU�4�mv���vq�EM���T��2�|�l{um�m4�A`4�-���ՄO/��qi�"�����~fV��~�w< ��N�b>0���,��6ϯ���v�|<d�����إ���Ce����A�|��F���ན���IL{k!�Y?)W}�bߑ�s��m�`t7\�W�J��0?�f��kI��.���2��~[�iѰ8���pY��ɍN�C�����,�|pY�
_��Z�]���^w�9V�r)�M��=¾�cA�J�X�KBܬ�a�/
�C��
K�(�̫���$�]g��\^�^\��^v_3�б(�-��ji|�F�ZX�?G���M;A�j�{��n��o/�.��|vI��}}w<�uw��{г�>�v��xw!���b6��w}�v�,�v���q�����O�2X�cR�.�1>�"��)�\N��������+12�.�5��>�5����lJip�B����px^�L`�4 �)�x+թ����Q�OJ�B"��q���L~;ݞ��:��N�1��b@(B�S'"ה��������:Z�፸�h�]U-slFQُ�Y��:�^$���G�NQH�~f99Y<�b!���AHO�E~~��̵�����y#���!�ʦY�����}�4njg�άͶ0!�44���'�Q
r�M<&�$��0u%-�9�φ��v����j�������"	�j�",��Q���
�^Z��LUЗv�!r(Y(�,��Zҿ��EWQ�'��b_L�>�X��oWN�!c��TD��-}hC0�s��?�`��0�+h�����)?���T�>���6�eFC�AZ�gQ�!��� O��m	���>�MFV9@Le�R�AP�hch��1.����2��7��l~��4�w&�<�\�c����5�qј�p~��r�="J~�#.�CԋH
*�ǝ/:㨌 �}@���8�tj���!&"�Ұ�H��
i���R4y2�l޿PR�Җ�૘P'I����4/{A �։�_��b_^	l���uM?�+F��s�-�;#����hwiX�dn � k`�u:���0����T���S�|�O��w��H��H ݠ�����i2h�*�4�RHy�*�M�^�Yֆ��`#տW�J}��1´����Ԓ�ct�rH�J� Ȍ�A���~qo�Ȅt���f܌��H����w�P����SN)�M�p�̎��5p�o�!��Oz�JK�+ć8{��t3T-�SJw��!gZ�-�n�ז��ܤd$8%4;;�7� ~U3h�j~̑�o�,�Vѣ��`����j1��I��%et397e���V�_"d`��i�S�����iOF-l~^A�rޏYK\�I��(�]]��Q��]v��;4�[�������bf�<�Ǟ�oa<#�<�lnǺa�5��Qg ��핮��<�����1��ܴ�m��L��Ǉ��A3_v#U��#��J�IÇ8�����`C�@��t�7 ��7 �\t��K5)K���q��*���D$$�������&#���oW@����//�=Ɇ��:T������E}��]B���:7�?Q�G�/�sf�de���ŝ��z9���/JN�F#��f��a )8z�x�-��~M�6�%j���b?Sň��ٔ26��tdT��8�K����>I��J[qe+}3��ݿ�N�G�۳��k����(��D�Up������h��<,s�$�6]���^����_�Q8UDa�9������vJI{%���(x;�����L���c���l�KW�v�QMK�rE��茆�����&Xě�1��q5���KG]Kњ�r�=	��UW��*��u�Jwv����� G/�����|����{ԛ��6}_�Bk��%F�F]���z�I�U����������P"�:��ß���~�\��A/y��K�B�BQ�s�_�uB��ݱ~�"��O�`���Y���O�Z��]Ϊ�5	�W�A9���C��_nɃ�4 }d,U>�,����S�(���!�_���y�E�E���{��*d���XK����z�遄`I{��B�AY����H��<��� �Y��y��g��<�,}�<��_�@�}Ƌv�����h�$4Su��3���5Je'xd>o��
����B= �PK�6;(!$P�K#h�]BOC�����v�G��=�+�T��*��!,R&�5���We��}7�s��d8I:��H���
�i�	6�1�)1�^^��iOC��T�D�E���T���U:��
�Hk*��:��X�E߼x!������͜��(3�����n����-W���0���r+Q��Ë�R7$�fO�����ͦ��8�Z�8��߽�$��ug���5��V�A(�r@����ߙһ��:�ٱ��&m��H�pb��	^1&���2bS�0��ҬQp�A�}���WVJ���3���995�L����ݚ����fژ20���K��e�"�!A��.���'�~�?8���m~.��0:�K�655�x�ca�s������o�A�@o����e�R��# L�4/�}�$.��r�t��k������d������љ��j��J���R���$�nO��T ���Ҁx�:׶"�u{SF��&OWͪE���3T�.�X�T�S��S-�l�߷�u�6�cә�ՙ�u��&g����d�؉���j��YG��v����C��I��b9��v=T|�Tl'U�Ɗ���*��ꄇ����"+Y��zi�}��b��]R	|�di�e!�4��̆_A��j�Z B>ї>`�t�-;uE��4�`���߶����+����cy�L�@?W����'( ��A�*�s7��:����E ��z[f�S��Xz�WA%�Ic�x��敥x?�D=���	�ʆ|�|ǵo�h�f<�7*t<*��ɡ\�͚��_j����k�R+����_�L�'/2�%����w��I�e7�����b���YL�ǻ�,��|N����Az�L�&K��Z�r7���/�z��H��2XՂj)��O��]rV��e�ĩv|�����o���d��]�u��®�j���x+p������������_���f��Z���shZJq�����Ee���v�f[Y2?�IkI�P�q�@��P���B /�I+Я��g�uU#uGSա�J���/�N����H�c9�;���;���;��9,�m[Z����!��!�^�7��"*��p�Gs�E�V٪���E��A؏�ޑ�����,&N���Ą��!g������tt�Z�6�uv{w�K �+�>�k����m���~7���V�z�v�Z���_ζ�v���m��ß�y�}����H�h�<����W���� �!M��N09[˧�1s����
��y��1�c�f��]q�N�u��8DJƕ�}eu��StR����_����ϥ"��s�wRK9̬.�}�8����- W��H�h�����FE ;�u}S��Ir}u�Sl��[�z5qخ3j��}��vt}j�y
��h~"�=������{�'wLK-�;Z~�i1x�2^5۞H)�*(yeS,n*{?���J=��	��ڹ0���&N�ݩ�u��y�l[-2��y��k!ڹ�Q[E9h��Hsb�S�Z�xl���ȃB��H�q�Wa��"��zqA�`��/�R�,�p�?!6d���h)}F�p���9�dL'.0�ٟ+�LɘQo�P�i�IW�q�0ԃG���`k�OJ��3� ��<�?�O8f��{	Wsl��J�'�' 3���}�~:����.Ԅ<Q�l���i�N9�q,Sb�'a%���6Z�q��^l�"]j:�s�ug(9xL��K�_׿����C@��nl����,C(�u~��g����u,j4ўc�-����I�. (�B�jC��`{�Y���:��ڗ��_�����שF2aP��7S��>Q0,�@��5k*��3T��X��~�C�A�] `��l��R��uT|��B|:����#�͸�a,E�u|��'��i�B�j��1�KW�k�,q����wL�W~dǮ��3 �v�6��G���;ϣY���Q64������Զ��TFY%4�pK=q��|<���?�w���x����
���F ����W:�A��Kd�]�;�;Z�ϯĩ���'7J�r�4�l�*9b.a�H�'o�r���J��F}A�bK��-k]�p~<��Z��Q�o Vl���1�ߞy�6�/8�'z��H��T��|)�cF	�h�W-�9�k8G�R��٫�I��1�].+��|IW�Ss~[7w�p"@$1 ��	1�A��R���M@� #���r���Z���u�+�-9;��'�M�G��7��e��5��R�����sy<|w3�$gp;1)~�i&$�Ƕ������rH�k`{���������ٚy�ˮ6�P�K)���ٯ
F��jY*EW�c-�p��*F+�?��ʀ==����ĵ6��:ԯ�dr�ȥQا�2��\�&�`#�K�G/"G�lw���l&�r9z��89)޾�YC��W���Nw�tJ*Zj����W!;Q�h�j������3#,6�����QV��Ĵ�?x�`�rtŜ\E2�Q��ޝ����B�X�o&ގ��f��������f�Q]�|!G�AE��k�W��djk(�#�ǯ�-�/�X��%����[���1� S�{����[�:=U�2��!�G~��s�e#�ߔJY���+ꤘ��8��=�V�X��>��FuZ�e�]c�oh��)�2��C�'SD0W��d��]�=w�L3��fƼ��������X�P4"�҄�P�	�C����P�hc�@y����L^��PsR(9�w*ӹP��[%][�������~K#+QoW#f��"�?���*+I`2�F�B����=P�AB�ʆ۔�I	3��
1�����;��r�˩��ݟ��ձ+���Q(�p�?��v�Y� �$�GݺQp#�E�?}>��Od��a�3�eshΑ�����AIT���4zR�H�`��I�PY�gE2[�<�V��0�Xk63T�����0�7^Zb��1��K�n>,�qiģ���eQ�B0�/�SL^����B@%W�n�!>�A�v�[����P�?��P�>=Ҷ�ElM!���`��Q��+,<��6xA7b�q7�	�a:�.��O��t������4���~�L�M�6���S���{#�d�Je�@�c�AO�&��z��j,����C�a�U����+�T�7�n�ug���6�UV�� ��wg�3��c.�P�4�4�&!�P�P\� �� <i\�W2x����鴴�,��
��m������":J��7�!�g�7'x7�����mWL�^03�����Ҷ�?�m����\�,۝S��r����Eᑜ���i�ϟΛ�����]�6.	ow5]��qY�Ȉ�N���1�����9���)r歎�7�����o�0�����!H�P��ԗ�k��U)A�J]�����C�أB���~��;����NNP#?����]c>�>�����T����)
Z�\LM��ZO���,֥������9y}�т����?��|N�s��%�J�����9��͎	�В��1���������S�AC=�4���[պa36ɼ�v_�!�E�i5		�Q�e#-�����~:��Xv�~~�w*|)x�&�{�����
(9ԱTl쇵�YMmづ�i@K�Y���V2�e���2.���ё�W;v�d�����	LC`8�l��+O��ĜV���o;��,鎘O����u[���3��w��P��@g���<�.۝i�4XE����K���&g����]�O�����9Q��)��J �P��/��t�	X^r;!U�ȯ���9<�6��A�u�S,)��_�D�-?H��K�Rj(#I��(��FQ&ht���D��Ã����pI�ڑ�3�95x�M���{p� I�P���T"�U������w�Ɖܻ0`b"�z������.<��>�FO���r�19�Dg�w��b'49�0�@�M�{<7��P�
��
hp{��(�Zm��� ��t����F�EWȋ�� �� Ǟ9Lh���S��#���8y���k :�=�����#��@�H�^�'�����}21�
u���W|�4�M78#u�:�w�B+�M�P�|;G�$=�j64�^fԗ^7Rnq�;����������W�퍕g�sW�fW�V�XO�XhC�DF�z�
�
/��	�0�BU�L��p��z >�`w�1��ں鹈M�}�ԏ>��Kh�n����Z�V���gHbaa����e�ja��5W�yl�|�;�0��<��k�k���\����Ӟ�0螮�]WZ���j��N���)g�]���v��	c	$��ǩ���H��{Yhp���x�U�z��w�cM��zS���mT���r~��Aqr�H���d���S.��_��$��Y� +f&���yğA��"��EET��j6nE8U��9y� ��+}��w�,�d䴴�����Ʌk[Jiwll6Ǡ=C��t��j&����/�[���r���ډ��o
(�!��m�>^���m���L�Kȃ��,��{�t0��}<��*,�����:�EhUڬ
��Z�'J��\v��j�k��i<�o��6C K��U����X8�v
;('s=&���{x[��2b
���s;��
��^Gx�������&�*�1�7�|��
KO�M!e'���{�9�S�E�g@�#�2u5�rE���e��/�=@������@�eA�ð��=�ph 51.�&:�[��7���2$|�B�i�����	��9�I�줪�G[��pl��脰�lqǊ��gy1�׷�gҩq����ܰ2���;y�x�b����
"��}?s���M��!�@nC��#��Hb�i(�Y��3"�)������ߍ�.RcK��)0<l��s���y�L�4q�ZT�Z��P���-z��c��7�0������j�$
��P}<v�Kc�~G��C*9��% y&cƊw�-�����Kg)n��SQ�Bb��Լ�3p~TC��>V@��yJ����_���	�1����A��$�#M��~o�-E�T��V_�.PMbUC�
��E�� <i��N,��k����X2\��H�l�˗�<�_/g����М��ϑ�X32���;�L39��"�B@���^�C�֟y���'�����)�K�O^\=m�H���_+%l�G�׭��+���"�y��KE����ɺ����\��|&�R5�� η���%�i��'�Rcȡ�`��۸SI�J�q}ܘ�'�ˢ�+��a�8o���(�8�V��<�	���k���"O�6`+��xw�"�4����D��2��oM���ꕯ��.�A���D7����hWn��/N��\X�d`�
�*zBa��jy�����پ��w��cmCF]�rV?w*��g��S�U<�CK�\.�ר�]���AWn��:�E~%�%w��?��H^�F��W�?_��N~�2�6_埘��߭PY�mU8�� ��K4OJD	x�m����c���}���M��4�-��H��%�����#����p��?ݧ*Ӏ�f��ɐ���紇B.[�fy9��ܟĶ��\�a68�M'G�\��D�nNk�9���|O[�ofۮ��}/v9��,��R�ey�l��N6�j�7�m�ܷ޾�zos��v3~���ه_oԜ[�V����'�\�ɧ|Yn��ٛ2bB�m�R�!��i�8�<.A��2��f�KBhE�8&�tec��{G��MO�~�ڟ��hM�[+ڔڪ��1��>�[�!�_ڰ<Q[�y8K��	-'#)]�=��;�Np/�C�[�0�*E+G�����\�HO�|���k�j�B��������<���`���݆��|�GkE�I�J���j�� b\�)[�)U��Z7���E�Ͳ�햒��TI�G�%f�ր_�|8�_s<uit�m�6�V=e����
�B�A�o
��k�\P�Su5U��5���P�<Ve �{��`g^Y��ޭ�$#�R9��_�e�VF�b��w��OIK������V�t�Wb�˜_��{Q.�A3x�o�{�����@��m�z�e@�F����G��?�O�:�*��i�ûo����W-�����ôM,jV�Z�|���}ɯ=�;�����#G+���@�e�|�OF�,ˢ�T�꺳���1��Z�`S,Zk��yv��ixwӆݦ�w�kyOi�]�d�vȻ�� �1��������-r���r��T���@�!���8������N01T� �"̢&��I��%�5N��|�V[Z���[�����E�������H���.;��If{���3�����������R�ؘ�IV���9�U �%4�f9pY(���\�t�H��\�B��Nx���~UK�M�1¦=2�� l�k��ɠ:(���4��=jE<xL���(`�����C�$# �F};��@��I�7�{O��e#�5'Be�T ζg��DĪ�| wkW���N�̆�B��.pܤ�T�X"��ҕ�1��q�Q�U�?�<{+y�.o�͂�8��/+9������)��Ԏpf��'Ij_�n�82uX?~ P�QcˉL��0.C���Q��0`Vd ���!xp��-ε�e@���Y��
�gpnChQJJJ�Z$��f�q��������;,"*H�J����]U����w�NnN�-Ϭ��P+�
B��<�!�1>�:���n���K�n��"�/WK���u�'n�$Z�Ӳ����n�[�O������P=i���7N��j6�����PP~�[)��w�W^!*����P�u�ٰ���L%|�LLf��G.���G,��7J1��հ��;������F-`B`g��v�\����6HG���� �"����v�,���Ny�E�+0���D6L����38�϶�� �����壌*����\��|"�wY����g��gǾ���Ju����uNI�}�T�o��i�T{��?��T��*�� �l��
L�/nmfP,�>^�b*�-}
��#��Z��ڳM����V�mU��CVJ��D�V]�	��7#���|�^h���}Є,zO!,��W����_�h�S�a��cNY5J>�m�B;q�3�zB.C�ث��H�'OlͶ
+��XB-N`�o �4���m�n}��_aDޛ���&n�&�:>he�aq�W��Ã���U��;S������Emx�&s�~����}����/�b��c2������=�p !v�l�9��ۗp(/G���R�d�8#|�g����5B�o��0*�͉�Ow�>�bV[¸�^���Ǣ��y6��x��E��
s/�*���˟��(Q��������,���u݁�NR�y��¬�$O��^.������]�'�r�½���+���������&��o:��FI)٤[Ba�L�)��!�R�AS)�n��"�����;������ݻ?u]�u�O����p�HC�)	q��8}(.)\%�X�(��s�s1�*��DF}�L��*ذU�Dب�I��"�����~-��e�(�����كP�K�j�\��J2������=m!��⭢�+p�!�ϵ�C�����/|�2��Z�$�[y���i�$@��& �ek�hq�m�'�};U��rWGS�p��^�n!����k4 ��El�b:�@ ���WL�μ��_�ɷ)(�Q1m�KZ@��`�V�$^��r4M��Ս�6�s��d�i���Px�E��YhUȹ7�j� ��x.�y���}3|�W;��1�
�:��[.�Z��������]�P-\i���ܴ�_|i��L؆J��0��gp��t��p�n����R��,Q�}�"s�`�����[s���z�����<tlEAX+����G!G��r>>��5Ε�H���������3X��|y�`���ۨjӷ3y�´F��i@�����UT<�9�o5Q=��iC��͑�L4귯1,�g�XC�9ї�$#����|x{��B��	:y��Ƨ��;���>4F6��^OIyf�趐J�y�v5�)����rה��Ъ�����$5�����ڔ'W�
�3?����I_�����1P�ߡ؋��P��J����X�ʨR	���s��i
S߬�
�Z�
Vdo�[�Wa�#��+n�^nQ����:M�(;������� 9IN��� �ֺ�B{M%���T- �5H�x2�(�RHC��c��J���o�yV�2��WT:hS���.����䏴��DN�$�����������ޫ@��p�D���篷��u���ۀ��*ej�WEK6�Ҁ�m��oV���rq�*l�ӹ��2�G��� �	x��;C� ��+�,Z�>�L��¼�����T��:��FH<�B	��m��@н1k�|[_��/���
�<��-�t1�K��'���D����#4�mc��򤝱:`#F_�t�����S��aV��t��Rq�	����FU�~8.��uu�)�}s�I�Ϻ�$��b{X��ү5 ���l�,�vژ}����� �i��`P�_P�s��Z_���#"x>���d\��L2��{Z0N��5�=��'ܒ������:�|]�}c|]͂�>qp$�@J��3B�w[ͳM����m�R�`�)E�7^�b`��W ����m����*�l�!�.���{6y(��藕��5�u�,�w��sngk#Y��x&���#���2wg)�7���'��w��WH6��+�p��N���hY���'%�~sJ*s90�r��t�/�ru)x���@AH��3Y�?ō>�l7�ծ��̿"����f���e������m�q���T�wk&� �^dmE���W���{q�`W�C���������?c���3�aI��ә�\4��E���NE7:F&��� ��-�;V&���{{�01K>��O��4���D���'Y�66�@��w�Ku+췿��k�44z//Øl`����&UB������e�rY���_�i<���(��/�ɗ����z�zV[;T8T��S�đNA�Y׌���i֕��na��� 8"(dy��L.<'s?q��.��n�;�0����1d�k�sk����꒡�o��2���+���A>@?p���N�H�f܇���
)g��/�ic�h�D�lKx틦�5��8;���(���h�[�ŉ���)2z����C��\���08Kz}�]iSq �@ �?˄�� g�
: J�#GsG�Y��C6�4���WdP��X�P�-�8�����}�QTk��S��ڏ)�N�HV��9�\0���`�;�������� �񂝂!b�f ���).�7y��f�D!l��{4��3���4�Z KU��@b�b	䇓�F{lDg�6r����y{��+Α�Tb`�2.1p�OSE��u2�����y�4��	!�ZM9�>�o?-	d�Q!��7D��X���ٺ�kњ�j?F������	Bx�4n��heA�|�{i���"g�.Wi�-�Zf��]l��i@q��A�:��[[>>�fg����N�ɛ�����J��-��ߦ����w�h�6�� �(+�m�jՄ����ŗ0Ѩ�2��:���T��BUf�J@�M�9���K��R#s�ػ7+s�A�xՕp�䵣!�Sl�r�br�~.�qw�M��r�)����f�)�r��j<��r<�j����x�"�P�\�)~��~�_I�6j���n�|��tP����?~�(|�p�$22�
�қ=����3�}���8D���H}2R�<>��������b�C��`=n!ꧾ�	L^�Rje<���,��-ߣ��/8�ޒ���Ǔx�3��_�>�����o�F��\��{�N���O.ѯk���z�c��5��H=�D�|ʾdu!6���-R�����qv��y�Ή���|I���i���_�;�R��f-s�f��t�>�`Vd��V""�U�rk�����^Q��]�}&k����D��Ð�,J� r $��Ԓ<��|�=��1^�T�����@�VW��8H��Ɯ��C�1���ynŋ���B[O�6Z��;.v��o�G#���ӥb��^+��$�	3`<m��.+�G�f�h��GE�ۓ~����ߦ�h|�W�$%�Á$!]
�8Y�O�mu�u^l|TJ�(��"z�/���X����)�Iĉ���&p���y��C�*d�@��#�\�2��:�xQ�Oq�iR��Y̢j���k�'�����8"h�kt�z8;nG�� K���s̶Ȇw9��9D�C+�2������0СU���Q\chq8	�ku��ᣗ���|)uT�����J�w����_�&�6��iWذ&q �b�p���K�@;�?�! �Q��ژ:_�o��B�E�W��0�@�J��s:�{gޮI�,߿�η�����~�zU�t�(�2;i���O��)@"�Դ�w����7�)�R1�1P�����W����ᣬOs����������.��3�{��Hܫ���_�/�_9�.��[*2n�ED�ܮZ__���2��N�ܟޝ��v-���^�j�����#Mn�Zn�*�y���usrmr��x�-s^��%���Z�s�4x�1R������7�����������FJ"��������@���ͬ�ƹ�y#I���lS��0h����!�������B�#�'�o݊k���G)	1��C�����K(3A�(�=���˺�.:Y�f(ib�����vi]�^���rC+�M��<��t"�z|ԯJ�eܮ:�`X�RC�Rbq%�)Ψ�@"�z�B陪���(кϋ�jËk�c���8��݇,d=
'��i�f�;Z9Rg����]~�'݅
�6���a�B����#Khęz��=��U	�@� ��9����>��l^B\�d�ο����←u���ۺog��{W�i�֮>���"�5"k�Y���-'P_���B��U49�#�_��%�W�e�W�}��à��_V���cO.XY�"ZG��#��K��Ҁ�?_⹺���ɱ�|$��ES��j%f,0���Κ5���h���}q��t$؍��K5f�T�4�3 "��I>�U!"j=x�ꥳj����?!�^�����1ݘ uJX��i3Sz�%��Dy�h���n�D�:�4��W���0�s�~��2�H�6����~(�n����e�*�ɐQ�kp�F,.z��ϴ�u�u,��@��[�>g��¤sk��� ���'���B������U,�� N�������[d��N�,x�'�	*�Ǌ�9F/��϶�#�s�&ɍ�&�S��zZ
����\$6�$���h�}���U�r@������ni��a�K��9��@T~���r6��Hd��ClW��	�f����?_�,x7��onZ>a��cn??���y���c�[k�����ޖ{�=.�{��r�x��y�K�xw%plw_�w�cr�O&�
w"5��eo+f�{���K�e������+��*q��[���'������,C�;�".fR�"o�5��h��8�VF$�����U��u�n�o�K3Mabk �۫2���!/�v��ew��𻽻�;�.::���;�|�*��?a�_T褼�4���AjV�Ö���|T6���d�qſ�滥��gޖ���}�A��u��uމg&�>ۼ�� l�nq
T���ѡ:�(S'���s�uT2x ���+>���P�O�5�PUHV}��@!�W��6����7�/�w��z\�J�����\��:֫o���1La<TC��9"Ů�8�fB�5�@6:@�x�7c���'�����DɜT"8.̣��M-t�螃5R�c~���nZN��/�����m֌[�g,�z{$���w����V��"?��4�x�i����I���y&Pp�Xp��X���t��-���������'��ۉ�{X���׺�V�{�7_s=�	Q@ň�������W�ͨ���\ �sݬ��T�"�$[jC�+Q�|��F�F_���`T�cb��(HG�&1��dҬ�P6V6��Y�: #Vtd�_6�f���b�c?���1-=���*߈�L�������C��/LP���b�1Z�	UP���Hg���}�:�v�m��n{3o�ƽ���R6.S��p��Ɏ�3<��V���|b$R�������!!3�'�)$�[��]��mY�`V�|�8n��Aĩ��?z��W�6���d_���@�7_��ɿ��	�5���B4�nP��ǧ�W3�[h��L�,���p�o3_^k4�M'HqH�� ��\�|�|M��+���1�4V����р!�x��G���C��o�:���$������F獂
|i�5�˰*mJ��^�8�0NPe�NǖH��0�#�ӡЯ)�6N����5�n-��G��2[��	��+�E���&%_&�`��)������=���ye�1�����&�S��/�H��BU��T�Ƭ����iM�SW�Ǯ��qs��q������,�ϓ�}]�VdFP=���>�p�J�:^��/�@���B�I�������$���t���&q�Ixp;B�q𐌜��K�칶���Ϧh��iN�����mK��o͗�ݰ���!nb���|��'���f��]!w��������#�5U���ۜN�LM3ށ[g;_����扟�?�+��ֶ�~�6f�_6l�%���[h�*��/�i���!�?c|�}ˉGB>��4lU�KI�GI�GwdW������k��#�����_m�y�俳l��[2 *w�7�.Q�ZD���[�[��A/ȣ�H&B6|R�A��eO�ִ���Ee�A��r��cz4ڬ���t�4L�]�q��ͻ�aO�������ح��$���������H|����-j��?�d��!��,&�����Ey'9@l^�/�x�>3�P�#��,VͭI���K�zmt�1��yZBx�\~.���kZH<�g�e����0�UZ%Vq�J嫯���S�O���kѫifz����yY��Ξ����)�{ѫ��|�#{�ʬ��}Hf��,C!`�BE
��N�D��wk������$	b2�l(]}QB�J�3����3��U�aE�Q��7N����ٶz��P�8T�nQ�)Oc���Kn�	�ք��)�.�yф�z�|����Z�P�/�@`�
��k��u�!kQg�M�/z�}f����m�]Zn��:w���W���
v��[��{%��4�����s}F�^�F��a��ɫ�ro�����/o���>��h[��e��TR��6d'YL<Mt<��9}%�!�~^;�V�_8h2ħ��Y���$�W��^�����d>�:�.�Æ	�1�
>�Ǚ��W�����8�ʑ�/w^	,|q����_�h�'ξ�ڔ9��ڪ`��I���^��4����HVw�Ϲ��������,q�k��J0c��J��>~je5��ڱŏ'�����ۭ/�n����gT%��N�Otv���R��X�S_��<%`�U��hg���y�iK��d:vЛ��ml^�V�ռd�1`c���M��7 %?S
R��M�V6g��a�'�ULl���V}i��Zy�N��C������?�2�W�C����ޟ\�07��:��?�ًn�)�p���y��%s"er��Z�����yuО�'�~j�F�b��L�9H��mO�;�L�Ս��x\{����������eC����ާ�7Y�Nlz��h�jx�^Z�{A��t���Ğg�=�H����{I����}���ϻ���}�2Vs���h���n���BxWr��#8��p�+���V�x�a.��?L��O{��\W��!Z|CQ*���>TZJ+h��j�O��Y�����G=R�$�Qؕ�0�a|��Φ����:�#d-��7#曬���!��sg3��U��CkYicn�;������W��O});W߄�~XY^{҆�2��3�w�s�w��3K�� ;��&�j�x�!�/�3O���� ��o��1��3ʹ���ݾǵ� �n�+���ƥD{��Pc�6=d�!��	g��Eg�����g���^e)*+y:��{���8���vT@��v�zz�c�Cn�Z�P�`�����ȥ��R�͢4I����u`@.��I��ɈM". �\�m�4�~�UN�X��K!��mT�*��̦Oӏ�5E��&�`1�l-���i[��C�M��R!)qK�q��E�5��~���7�Њ"�`�����EJ�+����*�#Av�O�:���olT���[���L��(Ԋc)��V��**���"!��|�B�2��O�c�_V���c���[ſ�G[u�À7s�Q7?�Zs�.��NB��g�{���@��)�������O0��q8!}�c9k�8tu{c��he����Lȍ�|C�W݊zfT�[.�g?e?y<P��:���Y]��W��k%��zl� D�'�t`�ݟ���޶��5N�~���	$#߮�/~��/?�)u�t�1�oq����:@,/�n�½�]+\�>W@)�V��b7fx�M�O;̚[��v����D�T(E�(��ŧ���7*cw��*���
���uG�Jf釲���-:���Fx����Q9�S��lh!������B��q�r�|�C@���ׯ� w���tL`E���x��������fyfo���R雭�k��l�ۅ'B.�WI�g��ꌿ��	���s�y��TU��o���y�p�B+\��B��K��Gn勌+~������#�@ �ErX�O>9��Or�(A�9� �>�J���6g�*ad�c@��F�yB(�w��t40,�D�ϒ:��E�]�4�*��0H����Y���7d��G�x�	=E�=A5Y��o��=�,�W���/����8���$�3��aed*���������s�h������s�y����	C�?m�5�j��P����LA�-�1:$���ū	*�ؘ�ǉ��B��c�a�XUQCRѿ��ݞ�����Q����d#���P�D.�ʕFmţت�u��� �)q��Α9i�UQ1�3k
�������'���E�M�|k�����g�{{�]!�V*�y�x.��v���}[� �k����g%��m<=y���o{��O��YK�E�2ed^�DwVH�!s�|i����"�F�_��%��̂�B��8Q���f�*k��l��-�����Bk����z��� ��H!}�O� ��?u&��
������t-x��A����C��;L�GWm-x����D���D�G�����H����C�j��	���l�K03:��em��	�/��ߔ����9F���L��`�f
�����:%�ޗߟ�'���j�̋���N��gY�`Q1=����E�g�,��=%��k���;�8S< ����Y��<�@�;#�P����<L'��g���Vp�Tn!��|�Hbyn��r�3֗E�5�I��;|$5�N�0��������n����
u��L3C#���*��b^[�/r��LVMK]�+bS%��,S`hF$:{�(��{����'񓻾cȐ�X��';/�˚��3Jx:�W[�m8��46V��������l8�Z��0_�WB�0�ԭ:��TG�vc�����$ժ�ӉԨ嵲����[w�WVZ!��MR��?u�6��~풷-�v��ԴT�V�OC3tJ�<{��V�d�8��~��W��R6��qh߲���+\�:{jϿ<�usNwiTsiB�Ƞ�F��8Oe�����s�����7 �o��Pμ��V=A+�Aӄ�+R�,.��N:h��[������I����T 	�U8͟T�cӡc�_#3��3���v~�^S�h���e6��#�'9��I10F �D�R%���I۽�c_��~�xY�cB�t� �?�],�¶�x���wI��4�t�W»���1�{�՜Ϝ��Ӂo&���A�֕;��	6��#�O��tTXLI���\��)�`{4ݝ��f��J�T?qw���so�I/I���,cK��N���Y=�u�h,F�	u52��")�U����_�\S@k�䡴�d=�X������@q�LZx����Ѥ���g�H��gDO>(6���u�*~*�Eck�2R!�:����b
���";x2P�@��v����0����b�*L3Gc��jL����ϑ��j���ܟ$ʻ���6�g]���l���������=���&ʐ��<�.��Np'�*��m��T9�0<��U�;;Vܭ���xI��nd�C#������Cr�zj��m�p�aܬ���2����C�o�>�:�C�
�n�-̀���4��J�%�~U�j��:�7}�����h��:���S�W�6O2��ss�L &�Τ3���Zk���%������^i�	����v��2�b�9�=5�Uf�4$��yu��y��˯��AԨ}fR����AqM*Կ������<h��{4�G�=%*��|L�=��5��Lw"%��'v��!~�7�9M�����bJ$ ���ּ$��G`���(��y�c�|���;g9����Œ�v�#U%�R���_<G��A�]�d��V�Ȭq×څ1�_y�$��Q��3���m��~ݐ����:�i���V ��S�D�O���0�:y�F����? h�yG趚}�
���.K��*�~�M���-|��}^�y�ب�p����
<�Q����0 >1E�����+�EҌ�s:hq��b��9�Ҟ��ͱcR���n�=:��3���c�����<|�Mc���xh�1����D�$�M����e�.)V�!M����_�#.���,.����KT����fa�������A�{�����b�U�Ȟz�4�����yi2����/�W?�R_�F��	82H�T/
Eiұ�G�U�(X��<���\�N�8�ȹ)d��⑓��بD�����䔏�����M��E�:a���1����l%�M�EY�-
�E%�yţI݃Q7C�`g.�o���-0=UN'@8��4㌡�6������?{��ﴗ���(�զpL�g�.Z�{�8����1K�)c)�]O#�����U�����$!$����'޽o���$�`�䇏ǅ��o��;���FB��V���ܹ^���]���ױ'��X��`��i�=��=�-��_��
��͜�g�Fߕ���]�eF\��W0��`�<jz]���e���G=}>5��> ���^���pY�^��h�Nk�e~�ْ����2����������F���Լ���U�]G?RZ~9��&��v���*�%�Bm���䉹��r�*���T����!���2��椊V�+|x�f�&���49&�+���t7�\�*���2�[�ӝ��H{/f�Ij-�k��H(ե��c�[�3��qWQ���/���ߌ�$��k���1���RT�����%����y�G�gҍ-Ey�c�P��A���Q~wj����nE'���erV��w���l�h(TK���	9�h:OS��
{�x��߄O@�S�wn1}��S�;b��R���}]Z�o?�G}7��u}5V��Fo\j̻�r����9
��ee5��i��b׻pEw�S1��ă6�2����̓��۫�M�pgW�4���~�ݢoiS3��Zt���.��fq��*ɮ�.��f��m}��u ۻ{�C��㙉�v�&)��Ȱ_��\�mt� v�#0E���pĈQ�y�`/�a��[�a�� A���ӟ���Y��<�!�	����E�#�ڃi-IY_d�Z!�/8�^�❐���h��X꨾�����[aW�t����8)�a���n:�|ݩe:�`?�v���\3��Cȡ��!c0�ݛ	AK��w�Ӵ�Ŀq��e������As�j�>MO���=�'�0Ȣ�\zئ��4��A�A�8x9�C.;.U�n����~Ô$�6A�ԧ�Ze��l��n��KMp�d A���a��0���O��}��#`C�iv�)�2b�����;U �LA�p#p��oom���N��Fz�K�=KK�p
};����n�����*v��&P��ԕ��Ip�R�$J��e���g�u+9Kb��d�Sp�Xz����'��}��)C��a
��f��59)�!�j��
υ�+2�pne���?����]Ƨ	��6�e������Uݳ �M�F��E3$0��u.��_��I�/u:
��tD7H��,�� 6N����&J�I-bK�S�)&��"͇G�-G)�>�͗�&އ��{'�/V�Vd�j�g2nt�'͡N��n'��"������x�C�0����CG��m�oPO@�u�ȴ�F��/�/��;_D�bv�E�>��ё�S��D�;:��C�@������P���	q�p��������^;�sZ_�'�o�ȩ)��Sb�=b摲��/z�T�o���T�VI����ibu������zު�#��hg�ҡD�3F�M��P������L�P�gZ��N���5��U5Ɓ��"�d�A4����Ϙ��..���0ۚ��z"/I��xHb�~�����?c�����(��C�]�\����}��`}H��|��D�/V&�s6
�MG�aO�GWTn�Q�2/l,&��=��L�횆K�hP�"�yf�K'R�Ҟ(�[տ ���y�w�IM���t��Ȟ9��͗tH��S����N���,pۜ�<������Y�ٷ?nNСj�GЀߌa��c�O��F��!e����z�2�9]����\~� �֥��@�W~�O}�Z�)�0]�ùr��Vog���r@h--�@]�h��}2���hC�.vH5n=�2�CKP�詋s�z�GQO!��G�t:��4E�,��SYn�ѧ�h��x}�*�1�u��9?ێ�>D�!��M}�{��u(�D��
�7t�9��t����x���fn�Uxl�[�hx8�u�_^*���"�+��S5!��������T9neq:t�N�d��]�CC��3��r�w�������v�9�x��������K�)�Sv@@��O�圄-~�I~���P�TD6��l*0��q�s@�gh�1�B�k_�q����U$��}Bﶷ�������!>S��ȐzM����2q��	���LS����Y�o���S����d�e��@�A��@��
������d˙��M�����-�}�Ai�ь���s Z���/6f{�0f�Z�����K�|��S�RFV���^')�ۺ۸V暵���4_NH�6^m�
��^�G�71�A�\P��G���l(@���+A>bäJV@m2eeoowhڕ�l3��2ق4_ع���[�VUwM�ba�JP�#���a��q�s�| �L�<ONc����̲";&tEÊ�p�����u�������0у��$ͧ�w5��'�?ML�ׄ�Hr�@�
{���ci(ZG�D�ɤHn^2H{m�A{ �*�־I�/(Q�Ak鱽�7��O�4�Ɔ#��U7תVSJ�e�$3lS��D>����d8�U�]��	FC51��r]t��ՙ�K����ݨ%c�_|(�˾��c��8�vw�ӹ���߾�B˨�O��wNW�_~f�^߄�6,\纒�X�26�Lϧ3/�G 6Vjd��UM�\�wT�N2�\���0�`8|���&��V�D�pe�C�{Q��$���C�G������18���׵����.;0��h�D,[ ���+L��&Pe8��ְAzJ�T.\�4P�ҁ^в.z.�z_0�����6+�'�]��p⫔y�� �	�i� ����4�#bpH�a7�X4��vŔ�W�-�o��T*�h�aYPtC�����1t���tf ι3+�nkr;��D�y5��f�ć_�F�ڼs��6�D���A�c�eXv�4��~+�kY��P�3������v��	�:\H���B������,S���e��U�@OR0���1�)ΚޒN��A�m����O����R6��ۋr$��n/f�)i��T��k��7��r/�������R�^Dd�}s�rƾ;�:�~����h[7cW�t���@�A��]~�Y��]G����q�z��E~i�����eB�]����xi`�n���)���F�3����$���g(oBq��Ո���{m����it��������$�Ϝշ�~�<��l�<����4�Jڼ]0 .}�Ș�m��'>�H'2�)����R�)).����7}R9���Vn�'�^73>�����-��~'�G�����K�V�O��kb�)'��]2�?���Z�w�E�caw`a}ee�*֮����|^����C�@ ���� �S�G�&׫:�~��N���e~���;<?�s�`�=�ߨi��M�T��{[|_�Y�z��� ²RV��gmC���o�aڝe�+�E�܄$�q,cm0� ��V1!�y��Yf�`�(e�#*�;���.�Lm��綐0��f(�
�L�I���jC���ΰ����V?q���F�+���~�H�_(%1��99��Ξo�q0˄+�����Z��-C�h�F��0܏'�{�I��-JL���������G�[�cH\/�$���I�	��tq-~�]��y��?0m��ܚ��\�j�$>�T��=�����g$��E�򕘍��|��a�=�ņ�G*p��4��{٘�����o���n��A8W$�(��j����-�7!�D�5:�E[�~+��Y�(�F��~l��n��k�eb]�쾏��Mc�"��,40�u�5-��K�HW� JV�t��3��M��e��L��SR����k��r��� �H��+�m	�>q���4+�z��$��J�`�ӟ���6=�m�Q$���W#�L7�U���r4���򢒤������	���8C�S����<1�F�xq���Q4����~��T�X)B��
�'׺�5n��=��Q:n�)t2��D�b��H[�5O��ru��(�L<
>/�����w���䲍�rʑ2����%�&ʟX?��^��Z��h����ss��2����:w�6���(���}���P�\+�%s&�h<��%�XU"J
��e�6wߡW>���!�LމS=�ӿ5��� bᑏ����j�v/_���žw�݄1:���X��#�L�Պ�0�F ��@�>,�G��vAbd_h���G�����Y�
D��턁���R�E?���v#����2�����;��q�ݪI���$c����C4)y-kt�hZ�ǒ��U<�5��B�a#K�����c�m�6��[er���Qq���/���@�n0E�������h��&��]�����ؾ�~	�={KC�%�P���Ӥ��)���y���7����2��̓��T��=�'�u�;;7`1���G ,Yl�,�:g:G
�H!�T�ܐ��S�oi(~Ra�}���A�<U>����L�����yZ���k:z-�z�ܕ�ע�u��$SDO�s�0@K�ء.�QZ�	|�|n
X�
7�^^uϩ�-�Le�i�FX<��j���Q"X$>�ų=�N����fa�������������b�	��7VN�d<�� �{�����L"��A�c���Y��T3'Gv*Q!2|s���ka�|#݉@հ�([j��r�Q�q�_X�I��^���_�Yr�2�%���M�P"�b���c�Ǩ}��d���à����|�Ʋ��s�m���V#�[�"��WB+?7��.�_B72B�N4$h��t�ǲK}7vP��uS��Z7I� �cv�P�.}X������y���J��s6�֔c:ܥ6�2/�lY-�̐�/�:ݭk��˱�Y���L���Ɂ�$n�>�����U��gO+�q��<NV"��#����7p5�����I��m����[��ȗȞk�]�}\�wY�;��^K:�|4K���UM.�X��.�Yz�WZΝ|�	��M���.R|���[	��L�������br�i�ڿ��� ���?�u���.H�x��H�D!�s�%�]�k��;�2%�0�x�����W1ۍ��d�2�YJ��r��֒�4K������l`�RZ�}:�ZI����Y�VB`%�ӆ@I��ivل�LΦ��a��/�S��ƪ�,��ֶ�Tkx��s�ڨSW�����SP�S���]`<nbFpk�D�h�}=�NG�"0�0�+z����XX�:��_;���)��Z̧�\�hGŚ�Z�S�Gk������T���p��%����W㋳�h`.A��ϋ��D(��1k��/Ņ��`i��� ����cJZ��b)��T1��<��^���T��7�rtn�.�*/z��;⾫xj7<�Jk�&�U2��*o��Վ�kb#}��L��h�֭V�,m��1�L�5����؇~�Ozis���ȂϮ�M�mwz@��3���)J�<6���i��x�$6���2��.g�k��W��%.ˆ�s�9@*�4�����j�d^�S���I�?�AK|_y�@0� �|\gO�P�|-�$X����(�&%�J ���Y���2MK�T]-J"�*N�o�o���<�"sih8h�EzE�q����4��@ίC��q��L=��/W�e�8N���9 N����S�|�I"�z�%)�p�W��� �X���;R�$��#eH��0���2�@�O�Yj��{>2I�,�]���I�XÆx���I�ല����u�דt�Ƣl�6'w��{Ȥ;>aI�:���3���o�f�cJG��%D\1����Pa����2����2`Z�GT��UϧW���&�`���2]hhu�8�}+���z����.����bd��KH�,-e�I�0xC��P�����mrf���ÌF����박��B+����`�O\-A�D���]��OC�/���C���hs���6x�>O�+ה�4z} "��˚����S�pk+Xm0����"�	���<r�@[(�ug�mNs�92�4܈��?��?,�P��4D�tbBͰ;T�5��3_T�>� O!�yjܜ~{�1bY�&����ge����8O�C�k��k_~t�8�R�b�|� ��@^�)*���A��~8�64@yp��u����m���(K��I=/�,/_���\���4dX�S	w&T	n򢤴���!��	<�qMi�i��/	�xë�4��w�vL ���VYse��y�ؠ�X #����o?��}
�X�PK��-D�)������*��B������8#y.v��Y�܅{P�׳)��%a�FP�c�p�)϶�l-�O�>c��K�����ğg�Bж+PL%x���p�`��U��Ul?C��<n/�cȧ�� �
M�}����5��޼(��	�Q�����x1��vH�����c4��
T�8��{��z�9�	6��{鈮�`���-���}:>�@��\�u�x�8�:^d����tqǩ�z�9h�٣�)������o��et|x�o~���jNy��F�h�-
�Z�K'�ɔ��C0u
�+3�Va�# `�*{*`�Ft�3t~�zI���vE��4�f�b�O
  �����^j��]W��
��K�Wƺ���. �!��۔~.�e[���u"�M��t�܏�è���a�(�1OҝK�h�=$�s�-�K�kV�'�!<6d[�N�$�i�>���������g�Y�,c�����~�/,�7��Y�����n�i�m���(��;����=*��sL��W��M�^��~k9ߛ�$e�����D�>���V&Kv(�C�4P琶�%ٯ��'
�?�>�m`��Y��,�v0�~�P:Y4����}�5���Ye�}\d�Q�T0J�v�ax)�H�旯6&����$2`����c���x�p6���;V��3�����F��A�R�Rb��j���.-b�
���nb�R�G�Z�J��T���w?�q?�����\�u}��������
7��K����Z���8��s"�}��I��T�S�
[-��.��h����ܴ��|�T�����x�.V3�N�4Dg��o��S��M�_D5�';���a��I�ۉӓ��3j&A^������Cd�T�L���/V���c�?7c5�%<�	Ւ���I�\����_��9��u�h�w�(�r���������ޛ���$m	��jѸg���i�'��H��rG�?B>L��p��4a��ކd
;&�ra��w��Z���6lJ\[bX��9t�5����������{f��be�X�������������/?�7��Z��y��˴��O����Y^�q��7��M���Vdj�;g�-V��#^�h�RɄ;�yM�j��-\���u�}�j�<��4h���'��9�2�������~�6�xRQ��z�����>��o����xь�L���9Ϗ��'�s�S���"\?2�,�f*���8���'��O�E����Șp|��躜�i�ʲxvν�#]�������V)ܧȳ�(ks>n��`��̵�y�PxҦ�
����6���-�`���M�X����x�A�:X�w�4���~�[ J�q+��C!4����E��_!F�b���b�D�E�%���R�a�_��x]'�H�"]b)������I�����Z0��P�֎������ ���+�/g�5�i���*Qc��O�Ju<2�w�H�1���>>��7C�����ψ�I <m�[d�I��� |�,�@S51
��ԩ��P�>��"��Q��&<F������~y�������ʯ�۾�s��㔉��~R���� ���16��$\_�s}��[O�)�e�.Ë�k�*Oo����Q�*��^,'�_m�!P�f5��5c �H0��ɵ���8�iv��FL���:�M_�OnNz������l����J�E�8�����ʁ�@~���|=y+���=I�û��}�o�������� ��?}LL8�\s��/���#ױN�9�&Ng��	"OS���	�jv�c�ͬ��q��Q�����Ji�*�]+1���
%>n�<��9����
������D�j2��=W�����6���*yß2��S�z8	o5�^
�h����S�$~:JmGD���o6��=��:4�{�S���w���������Gj)�G���!ڧV�������=T�vJ�l�e��6z!be:��Ʊ`9GIw����� \���k�� ��"�T����V��q�
t���R����5����̎�)�~�2�rk ��E�/z)��ǁ �:G���ܧz7����_8������ʹ�U�NnN�+j���ЩiW]��_�)j'��M���R���`�`�H�bwW� �Xa�i��ZO���Kz{��_2lL�Z�m����9�޺o��okn�N���w�&���+���)��M3���J R��d�Psz׬>VO��u����w��ݯ꿰�5��kWj2|�4$���\I�* l,sx%@T�� j^YJ���������f⚐QS�>���tV�|8�r��祺�[�{1EupY&bw�x��7� צ�n)_��<�D��b��+f�#+a�������L�;��8��O"ر>�}��޸�\���2{�+!VV�8��gi���I��u��`���������"gl��3�6ӡ���e�c�h퍦��
�m}Z��R���ֵ���y�;zϙ���	`�[T�bp��a��º}Tp��ky��������*{��u����Dtl�+���ل���+n[��Z�Y�?�67ך$��:\����x�"$�6�:'��k�L%<>�O'mϙ�>��<���n�ǏU�06_�n���@"��%�z=|�#����'It}�J$�Ap��[a���s�3�+%a�ˉ5���>{�KL�4^O�KJ�)EWt��� m5���	;�&F
��
�"�X��\_�_5)S.�f�7�>�$�{Ku����u�O�kBt���Up| $m����U�ꭢ�+�k�'l�Y�&��9���?ӉI{yW���C��=4��b$����l�B��ϐ������l�ک�|���5iܳ�9^^����Q5�?��LX���G��.�d[`,Q���6�04�/����EpRm\ְ�XE��E��w�}�7��h]�t7r�Ix8:׳����u�N$����>�~6J�~Eٗ��г�D��o~J�BBy��ҟK�b�K-|��<�7���|Z��������QsC��
����
�e��9[��ab9���v�a��k��"p9�󨆳��u��-�,���o��Tx�~F`��NK���s۟�	�b�y�P>�ʛ��۫�)X-a�)�}�4�K�V�z{0���&�T��	KnRW��Q��+�*�fz��������������Ks:[��f~�^��K�6�z��З2c�`��4A��������NX�L�&�t����h�������B]�e��rɉZ��4��Kj��?I���&��T��
�	�l��O�%��\���b�2��U�[ň\CG�N���Z��M��/���l<T�����*{c�ւ$(���#v1���V�O��>���!�֫@,����R���}i�挑
����hpSU_^�m���}"�}�K��������s��u��.��+�����M9A@�>(�L���ӂ��Qi|��@�j��=�k8$r��޾������U��M����m�{շ�ţ��d�Pr�2S�8�ھ�Z�Do7�HQ+��*P���n7�p
I�+��C���3$r��s�!+:���0=�0�>�B�V�S�t]��)�v�bu���_Tc��k!�m�E��Hp�Cŕ�߲ڭ��&�����!��	2�C��34�O㘈�h͠Xgr���4f�s�����R���^k��!�Z���d	ֈd�F���HM2dn�	�28~�?N@���}=~��P�����{�M�Ҽq�_�����i����yb��bXsX�c�	�?�Pbv��ܩk���[�-`E&�u-3u�ff	U��
IȔ�����i�ћ�CۛM���B<-���8q����F�ʣnl�y*�<#M�ȝ�JE�MY���/ ((@��9�x,׮�֏��L@�!�	� _7���lc�o+��9b�t�:*-r&�h�7�|��0��Z�R�]&���>]���8V���i�ݫH��ԏ�-��Z�N�Z��>1������Wm�]b� ��#@#�����tzd��ö	v�K��p��ޣs������������_2]z��wZ�W��A�=k�~_#�>-��34�YT�g/�=�%0�|i_U��	���w��d��I�q��������o�*�c��nd�Ekn�׉�\{�����8U���O ��n�Ą�^Ngu�a�Q3f��1��%��r��׵y��~�ٓ	o�O��l�X�6|K��*��	���+I�(�(�&���U/[�����`�_�������E�c[�Ѷ��;u���h�5��VEo"���� � g�hi^0���<TS���� \U�+�W9��~�}���7���Tx�fM�`"�:��o+G�_^��\��T!EV*�
��f���<�����GZAG(�;�^�$ک��w��k��������V6�~��_\����E�/�8����IS_{�1�M��޳�������b�h�*s�d�<U��G�@{@�g��U����o�k��Jy(�$h��{��Г=b����ɡ7���}�}̿�}���P��L.d^r�I���z�d����#b��ţo�B�mF(D_m��=�ٷ�����g��z!ۻ��"j1e���E&bqV�eUIg=�"�{�J��r��\�$���E��I5�UT�������M��c�t_���R MF���������+����RLqX0Ci` a�(%��/�g&F�+�բ2\Ogs�_4Ot�
����?�U�����Im��e�����AS����RҢBK�,�`K	�~��z��V��:�W$�*����S�a�X%�����Ƶ�r���i����* �R�>�l���7�u���Oo*@��g����bg�%\"	DY�C@B.7���3�z�}�p�~�w�i�#!Ĕ�xA39�� |6�n;�?,���/�u�(X���(vv�@�Z��d�e�mT�G_V���6�O��L*@力��:���0��-\�R��u��9B)((������KР�>� �9E���{Ǯ��8}'�{o�ϝ'���"^�]?����]h}�� ��iU6�yS�nG��=�o��c� �$����L���:�����{-B�=	�(�V&��h��!����*��<�_��W�.���d�*�<��@�(��奺1����V�A��d��&NWx֝ۚy�u�O�P�C���h��
]�| |h9H��n�V�iyd����3�!��PV*��ݞ�Q�3ydK�Ie�s���7|έ����Wi�䯖 �Lc���� ��Ny�6u�ʧJ*�Y5��4٣���� ւ�{�2u\����5i�_Xi��)OiB���I��'��H�Y�bv� Š�+~��Ξ����NpM68�,T�������C�y<�5-ܴ��D�����~б�Ci*��X��&γ_̐	��g������=w�c�6���q#dQҺ8"�L��Ș�@H�:sU��|!s��C���O�`�������rQF����
{���#��-�r4�������t������V	3!h���J��ߥ��$�8��;���g=H$��u�wT��x՞n��|kg!sU���[��٫w�x���!D�Ʋ;@yc�JynB;q�5��]�SiN�ǿ�^Q���6�WJ0�vd<�	F�!��q>fr��#�j�
T��T�c���ۘ���Hu:�W�8�fy�M��a���7/U�T���vb�:b�$zM�������4�(3,s�a�{����H�o�H��C�H��G����k!S��D[X˚����4F8=��J�(����|��?��_v�Wx��N�:8�O 6��'mX{�.��NQhն�#��SX,�NU���:ΩwdoIQ��8�襡�3z�����MT!��^�T��9%���^7��Wðf)\�e��O�L�xI)��֌RZ��y>���:�d�:�zW���f�A[�/t���F	 ]��)��z$���8��J��iG�tt!��:�n�:n���+@o��ՏW
�����>�)��e�x��U{�3/���<4�m��g2���\�ź�#4��Iӫ���y�V�xϾ��A�
SL���������1굂3ψl��Y���f�-��cQ��!�d��;f�޺��~읅��ǔ��Tȩe�ʛ:��:GDľNK�u���,A^���/�ĺ��G~ʶ�J���:cHO��R&�?vÑ� 5I�y��LiouU&d�K��_��f3����Ga�7�<k� ��OW�B��16��}ja�Rוu�j��-����>֩ryN�H$I�U?�M�^��p�$�����k��k"��č�I_۬oq�\g�tp��r��"!�����,o)=�v~gp�)��)���u˔�6�ET���۴,�~��[�S܊"m�5�ї2��{3�A�LK澰�]2j��E��Y��"~l�w.4��m�u����[�Z5�������ť�WV��l���p�#���'u'���h�<�^��<�o��J�D��$Z�m�~�U�J���r��7��
՚�e*,)�G��w.+�Ѿ�Ƣҝre�04�����GG����P�+*�sy̾����^5�K��G��.Y���&�Z$�-'vmM�E�'�I�[�1�=�v/]�P��:� �up�sc^�����sU�)r4�r��n����G/����^s����&�2��LՐ~��f�\�bj$z7�_Q�{��wQ�p�|�"ʤ�A�?�	�%U�cMS7P9�!��Ҹ�����->0J��1��E�d�j���q��-O"������:����5O"��U�g�e�u�p$Һ_$�#�(|�m�|�W;�bBԨ�''L�}�}�w5�[	���<�ߩ�q�
K<y�c�L�xv6[�6�3�"�����(���O��@�W��u�l7Qv�����e��ᦶ�]m"4�8�Ie���ԏR�@n �@�j�s��_,�ͩ3T�X�
S4�XʒR�28�hR��Ѡ�D�}a�̷����,g�u՘�� �g��Wz2z���)���&��������6��
���uL?��p�a"�6Z���f9�2wŶ@�I|�����E��I�?�y����>�/#u;3�
>F�.�6
cy�Ǿ�������e�~�&|��a�:4*��4��V΢�{r]VE&t'㼗$*ݰ6��4.=v��ʓ���hf��W�ȭ3�M�e��5m���m���~�N9pQ��a:���)���ҹQ��<t&�C�f��h�,h1A���y�C�?��Ϝܤ�݊z/$eǲ9�w��^�4<K�܀�������z�{M��)�����r�g��WУ�jJrr�b��\}O��:�:bm�2N�m s�H��3�t�}/�Rf����wu�{�Zg>3J�%7aL:@����3�U�����/�_dW�l��a���Yz���S�l�U�/ŕz���ݝ����o�k���7���y�"鐦ʪ�A��G��|	��%tXzK6d���o����#!c#s�W1
Gm��F���9u�����ΌM�z%��~Q�U�1�q�����PC��C2�HTSA�������jǞˇސ4��2�h�2��/|ے�xU��Dߟ�b��\���#��%	,��M���17V�T�Ѿ&�(�v�;FyE�v�:��֑�h�ӵ���"���4���g3��#op%c��Ǉ�t*����%z�K�7j�g�$p0�x �����8
TD~�*��Wz�fl#e��f�}���!�_�G�ۆ�$�R�������D9��4�۔��HE>r3����M��sT �AE�x�yAE��g2��_��N���sM�d&����	���T������L��h]Q����?�!uQO�	y�v�=^�]�/�i�i4� ��<,`�o[;w*{�.�\#[�ۈ2	�28,\�Ї{}kn����NW8&�9�}��*W���l&4��<�6��N��}�؅Z{��87����g7t�d��?I�#(�����{1��=�����-E�=:�X����st7py;���[kbF��Mx�
���}��^��O�A�F��
5����s�f2�$�ѭW��<
��ԵV�ӄ'��Y����R����� ~Nt/_�M���$�	��U�E
yX"HbDh;�T����❴h���o��=:S�r�+h�MnP/��(%%�3��S�'?i� ���]���#;�T�F�Z�d֩�4;4^�*���V�8-ՙ|@�SA�Ht	*��ckGMXJ����Tde˝'��L��u�tY�f����X�2I;����5��gTSxTMn�t��<JC	����@�X1���
�1�_� P��ђ9N6�8#z��[):�V���X�P�o��H6��Dv7��m<9x�����{V�I2Euy��ڔ낡d�E�g=^�$+1q_c��{��n'T1�[�ѱi�����U�Q��{�W� ��Rr�I+�ΊSv�h� �=%�l@���s���3�jr.��y���-OW�Avލ�K4��T"��X�����#�����].5c��{E�w�&ٵ�ȭ6�3OaM��*�*Z�5I*<����Cc��҃Iu�q	nðW���r��`��~�+�8���_h6  H}K�H���o�.6����zV�2rKѳ�y�_M>�J�2�C+�j�|q���ذ�L�"�����ͬ�w�k��^9=.lzjaC�w��D���׉֞3����樤���k"�+z�(=u"O�e��dK����l8�;�Z��`�-aX��\陓�g�܈�^��߂�%���u��͆D������낛���vVS���Z7U �Ȇ��ƛ�Mz���.#�q��:�th@��#.L.
a�zWˇ�e�k����j]�oF(�o��9�q`ڏG��5`ݍg��5G/ o�gX�t�<�Q�zG��t�F�����k���]⒈7�I�\+���H�L2���9(�\��iMU�6B�6�	VT�R/�	��f�WN�=���U���R���.~
w�\R�]_?8 �\���6�D"o���:ޡ��gGpz�mj?J΂6���6��4	��=#��4�ܧ&�{�Ech�zG��x:�
w�2(���i0�6���߉����7�B��z�׎_(��I��'��������b�u���%�������E�h	���y���s��]�S?�qx|����\�-�.v�+їbH�J#�/��qW8E���^|QT�q{h�3i��j���Gz����$���w*@�[���$Z���U:�����R�A;y_fN�gs���;�]�JZ�2ߵ�%��|��i	��DJڐe�Ŏy��d�f	iE��/�i��kO%u~�?��p� �$%���}?��ԺK��	�ݰ�* ��n|�mb�x�i�'#&��T!�:�����P���ű��9cμl^�
Aw�(��_��doW�)г��~$�S\�w���>�x �I�>? y���e+7z���05�����io�Z��Ut��ί�r%E6��l�T�ҋ�F>�����?�n!���-�J�M�r�UpCrL	�8i�(-�Up�hm�eg�I�E�+�-G���jZ�R��h�w?ץΠ�t�»�����x���t�wы�T����UޖĜo3�����晞���I֦�/��.��Z��S��?0G>]0I*�%��B�FӬ?�M�NB=*��ݐf��3uAȯi�����#����/#���G ����cq�#xr>��sc�&�%����>�iA���';9m���a�r�d�`	Ս�5�������Q=�1��3s��=I�E���ǡ��o=�N�U�{�������F�����[Ƨx�國�9�_�[�V�?�+Q�~9]`��(HA+龍�#k�{ܻ=����s
�Udǯ�J
�h����u���$_C!,,��
�G��wb&�@=T��a�T��]j�q0� IP�=6s��&X@�Z7K�q�t�z�D�&W�!��厦]f2R��2�򣄁UXD���߂����81hs�ME��
�����4�ɖ���UI7����D6�;��#]�P��d�8~�Cl�j���2"�Æ-���i��CS��"�޲������?� >FB	k��Y��sS�ޘ��L��p� 2-�}~�N�H�*�A�l4��=�>!�v�?6O����<JMXp��(HѸ��̩��侕#Zq��Ǘ�Ue-}�D[i�B���f�\7M��o��7ش��m;��k֨�e��1��z�H#P�	�!��v9�����)t��+�B/����8�:��tӻ��*M,�=�i���}\l�-6���.
9��L��y����ZzvmUҳ6o�F�4�j�<�.�z�W�r_�qP�R�����w���4M�ɖ�"��Eu�Ko~X�r�P�F�x�d����sF�FFE�{�Ͷl{8�
J�˨������rl�P4F�z�L
q����e⺔��^L�&�?�.?I��9�6�8ir�F���5�s�|�G{�B�*�i��	T��7�����oË��Vr�k�˫a��e���b**�:r޲R9x0�	�,Q�կw��Zqoη9��x��^0Q	ݳԩ5|���?�5<�٠��N�r�S�ܛ�f����ݏ�@,VcnG~�TGuH��Ē^j�]�۰�V���r�!�=�����vS�ć����n��"ү�)�}e�~N}?�Ru��oR�n���zX��0��I��5)�����W2o�!."�Йyu�{��t��3�
�/��:iu�^���T�{�Y�=�qyu:�'Y�a��dW�!��ܰ�y�a��,T���L�2�	L�c��
5���I`�1E�wn�kh��AԷ4P�8�0�+�^���O? ���+f��_Ӄ�Ȑ�޺y���Co`���;�p�d�8cb�o�&V-���H����B��1���p�C���i�ٌw��`�����1�[��>�{����δq,�	�d%��{�&�$�7៎\�.v]���D|G�I�9�)HY�󀌟�0�|@+�~��ܰ+�_�-+g`����4I�n*�DT�HY	�g�U��pߦ�p�Pxn��_�=bү��Up?�1�)Ѓ���M���s��=5��b����d�J��s�t�ЊN0�[�}*�h"��8E���a�?�-���_\�����rט{�~�Qu���{U͌�麬��B��H��Z�x!�/6�fUtO(�.������,���ުi�ј[U�k��+]1,��O���⹗0�IG�z��{��'�4�O��i�ip�A��������q,����\��Ö�ᵏ9ţ,��Ǯ�����
V�Ηꏊ�vE�q�mI�N�܌So�~�p&��� �7�r�QHh;f`Z�̝v'�C�����f�@B�Y�S���mbh��ni���bC�_G4!{��	��r�����t�d���r�ϑޣ�U�j��r��}�ޖk{�%�FeN>�Fڹ꾩�گfUy�M��>��@�"�w����Σ�L|w��b����5	��\���o޴J���	/�W��B$$�B�蘚�����t/h����ertt��NEKS��#T�}�4��j���	�s�J��&m�����,��B<.�Xt�	����wVP��2��~��@[�3����Yh��^6a\�Z��Q�,x��f�T0g�����&p���������0��\���5]��1r�;=��{���ӑ4�yV��k��	�Jlm����ȳ�R[��$ry?��d��G�&���&�OM�cb�CL���+b��av!����n<��9
N�H �
S��'�N>�bt'�Tt�� rW�l	��t��BKI*N+">�7F������FL	�Љl'��ތ��vc�D�0I��C8?b�)X���_Cx	&����bܠ5Y1��\��W��2��,bd���H��]qD��:w���e̡h����x�8MiOF�;1�*V(��օ�a��iE�JehfTC�����YT�5$�Q�՘u���>u+�)��͘�@��s��
Q ��:�3���f5"�k������vKJ��Įj���ލ)�F������n\oc=�}������뎭y@O����_�7t'k�I�;�9S�x�:��wA`�EOlI�
;���k�<Q�����[6�4�͛FE��Rm�4}s(G��f!_��d������E�	-|������N�cߏ��@E�l�c:��zX�t0]�Sl�0�EW��~;�(a�E�?�щ�)����=׀���R7h�S\����j�����K��oͶ���x
	�KZog�S ���e)�Ƒ��/���Z$7H���Pl��K�B6pޣ���~�G���"��e�據O�����x�z_�,LSպ�[l����y��j>�R���I;H�x�-GUkߨ������êN9�nd�ݥS!I��펿*_�s�����L�_�{�d�����q��/�M����j۾�>��1c��Hf����+���榟Z��^qO���T�C��Q@(�w�5f�Ο����d���&S�4
�/�nO!�|eX���;�H]����n�Ϥ��?5���*x�����_�ָHz��,�����}��>�ۜ8���y��7e�B���k����pm�A�����ܮ/���|�Vi��$�%z�i��;l��}/�+�q�ߦl4N˖�{]���/�R������y���#`����ߓ�z������H��p1:
��B��G}k�h$؜�锐^aᇵoV��Gt��@lx*��0�{�q�nе�ӊ��xfl��4�0U��&Ql&��LG�KSvs1&S�?��X��J�)q(�P%�F(��@�/�B��G���1�f������l]���N���<Rr5i�+٪-����jT*>�.����>B�+PX-�x�kI�9_����o.�xK��#
y(,�Mq>����[��|ɏ�xa�
�MKA.�O:�H������@��(ٿ�l��u�I5��:��\��`3��o��18���)#��({;�_�y��~+]�G�[�����Gja�yװ���w�ߟ�}�*�"��^��W��d��O�Y�ro����%���F?�Y�]W��ָ+zh���uB�"��F���y�L�ce�7X�"�c)a�M1�Do��Y���v���25�ߔ��B=Q�!�W����ZG�5�l�̶��=R����jţ/��C��x�>������?Œ�͆�k��>R���w���~$�%�N�8��m�ٹ��+Ղ��P��gŊ4E��I�Ɔ|��F�Vu�#�Ų �Ԭ��K�����O��U`�	8��T��/<��j�)$)��S+Y�4���y(��#��[��Zu2�ۗ�b�dq��N��%Go����k�,MΌC�˖�R��-��ĄP����i� ە�!�&=ɶ�'+�ᒒ�>��,g'G����y'��4׷�N�'O�,ɔ���i		аYB��u�z2���j��xmǞ�6r��S6LM��o��S���.)�9�M��=�Ci���ҽ1+���D����M�vzU3oNqhJv�3����}t��!}JL$����L��B*��ŏ����C#�}QC��Κ�▪�h*��.�l�'�6y��Ѳ'�Ztߝ^�]�R���X���KC����| ��hN~���PAĂQM�FO�������QO�0�"G�ผ�r�ަ�O0����θ��M]�T>бj��?[����,�9���zqD�I��m�v�i_2w��3��h���.�Ua�Y�=���S�ݹw�ۯ�/l���t���?�|�����g��g�"�׻?�PB�&��O�<�����Q�Q��	���; (��ܚ���t��Ś�}̊�(��D6@!f@�07����&�X��1yARC�0����q�J����cu���7A~�Z���E�l�P9�|'��tR��\'�.���5�#��e�i~L2�}��H��b�3$���vHg+gJ�a�s�6S���x����s�@C��u
�O��ÒX�gǱ�)�sD���X�/� *.6�:7�,�f/��W����~`�x�[-+,��h�e��b�}���Q���H��*&�����c�a��)��)f�GE��Ɵ����\NɅ]Z����=���V�+���L���Ӝ倻jP�&~�����|�x~<Zm�������G�2i��M4�\���.�f���i�-o��mlv(��_��wx�ʼUbc��o��},.n��.kR��Pj�zR� �=��&��㙋S��{:O2)���ȕ��W��؟v�2F�{Դt8ݢ�*Ђd��.6��֞-����-KpJ��M�C/��%p>�!ܴM�8I���>�F��6�]_a����Z(�
���?|��9~�;���0@u��~��P.�ŃNВ�~�4��}���O�3�w�������l2��]�w�?�f�� mҤ$ �IAĄ[1�Wf%)J�Z����I�s��9"o�� ~m�������΢k�hƽI�i�����������C�l�I�&t��G �2�)~vߩ.�� Q�6UP�)���-����]/Ev��dd���<4��t��<e_0n�>4�KI{p-}naoYҢ�ᘏ��r.�I5�Q�$��7�bk_�+�,�y����s������JG���˰{��et��FR��nl-��5��'�*�������X�?�VY�h��p���~DY�Z>Q���dc�Ag$��N񫳱׼A`���f�f�t��z��SC��+����O\S~reL��vU�l�Ngɴ<h����+�<�0X6mwC��+�x۲�Z�p����Y�g������ѰS��a��-�}��W�ٵ�d+�` �C*��cR�Q�f�t�i%�s��E���@޽[�ae
&��o�FT{��usI��2\��+cb"-�2�Y�l��Y�
��|��u�W0βա��hY��z�Z�<�R���)l�3��%e��ܢ��.S9m�؟���CQq���d���Z���8�%��>�I�ؘr22��YYIɁ@2�X�c�">fffv�Yl���lkq�7KT��h��N7����q8�u���JB��=����$�������_�����}�nE����̟��΋I��_D5-���|�~�w@Ĵ�Q��\8y}�Q-���f��LRɄޖ��Q(5��)����!(C�J4�I @T�߅��ա6 ��T��,ċ�&���5�XAV`���ӌ'�����~��79�du����t����̒S�8�}���ޮ�{9�7�*�]RakL�48�R������(��M����vW���g�?_��I�^A�~n >z��gC�s��ݹ8Z��{v�;�������|���09!��M�0��]͛��z�3hI���?G��ph4���e��w��:;*���wm�kk�x�	��!�^N�P�2O��X%0�\o�zT���r<����u�2ҩh�/lM�k�o��M�O!�=�P1�bV� �q�鏊9Ӧ��Oգu͵��P�*��d��da��^ &+u9�{~5��������7�UH�����ۄ>��>�<����b1������:�;K������%�l�%s�s+����)�y<�ڒ�kny!�Yխ��"��۞�5�-�������E���d�����3��_ӳkD���>�����g����;J��A%����.F	��vS\���l�bj�]���`�)���|`K$�Wd�_;Fc9���d���S㨂I^��K@��7� �஗�0��c����s&g_�[��%8�0�Jv�
�����~�\���p8`���`}�Z����fy�&�F]�����i��2��kk�K�P�d����V7�X�2҇ճי�)��e��Y���6ӑ��ɢ�rT61.SehߓNd�r�ȯ!�>��p����9�@-aH�gOBns��!�X�),{g�f4���n����z�^B��y	v�_�m�U(��#x�mm;s���@ްzU�I`�$�j ���\�"�"Q��U}�\gH��<��n�F�V�r��
�×ĸm���a�����TIKn��'y��*j�ש�^�A�M( }E�^�UAr� �Ca=k�-1S��I4sMa�u����]G:]6z7�]�o��tԎGْI����c������.X�\D��y]�����5���`ŕPu�������Df^!�	F �����s<'Y��V�i.�Ж�٬;\�$eW]j�`s$VB�1�+�aǕ.�'�X�������팰�,�<"���h��;�JPխ4m��:�o�h�8������#�jZ*�cZ��%�[N��浨Vo�8M�4�L=��W��Д@�1@[X�H)��  lЮ�.fq����Y ON�L@��f��x��c�^����Ʀ��S>=���>�~��c)h�#���$�]z^�ԯkJ��C���n�6Z��� H�5�0_&ݲE}tqA������_��^�L�?�ј�V_�.`H�k)������\�3�Sx�y�w�x#��<I4�KQ��N {b�0>9$��=j��4�U�bw}��[1z=k�a����es�۷�PP.�;�!���kG��w7�x�18�,4�l���J���n<-vq�ر�bӆ��8������n�'z����B	�]B�����d��%� n�����;c��:�� 0'�O�bUQjy<�^�|Źt(���G��5Y(w��ԥ���7>�ݬe~ˀο�`�`m�}C��Km����b�}��<�����^q��˿	�'>�8��{2x�h��7)+�"���Ԗ	�ղi��*�xˁR���s�<���k�M��"ÎM�?rɼ�b="�������s���A�%*��gf���GT`���������0�s���";��9�!���
/o���fw��L~�]i/�Щ�q�����l�ĪI�=�s�h�����hi��`g;�W��eL&�6�`Ԙ�3{�^�aW�����9��K��z�W��g��]�5͛�����Eߨ�/�=�(��L,J���ݿA��&,�^�dL�xD�����E ���,�jϩ;��t�/l��o�#���F'�)͉��7�T�H���[.(Kw^�YS��Lf:����M������j=��0PL����~!+$�{��!���~���X��Q#����J�Y�"�آ�Ebը��ZU�b��F�Q��Z�bծ���ʉ�������+���{\��z��}�p�h�
4��A�Ǧ���`=��e�(��dW�u��(,�,�c�0�>L�&�HNz�1|�}K�Ҳ�_�3���k�x'�~y.���o�i�?�tl�JdZ���"/앫��NxEƢ���W�B���(>� ��+2�G�V�o��5�)f�Y�it�aAJkX%:VL�ċ��n��״\�b���#F<��$��*��%�.�����XZE�bʸ��_���$�a	��f�?e�@���q��2զ�@L�`0��C��C�۾#~��[a[N���eȟ\D�.+=�p�i@����c�\���c�ȉ���i)��ݥ����6.�����Q�p�y���� M�?'7u/L��w�7�2��x�g�]'�(�Z���=���	g�8N�����u�+͵v�������H�֭�%�N�҅?�W!_�\��e콢����$͘���P]L͝��ޱ����X<%#0��3�v�#�|����8��g�Sjt穒PS�5�E���"�!�&!��,*���O��n�S���K�� �D)����Z��&zO1�$�f���}'�7?%Ô3�v-�U
�e���#]W�2�[5���od�l�Ka�y�]
s��!3�As��g,}9��;�w�Dv\��lc�^�Ɲ(x�ܰ]���� ��}>��&e�V������R�D\4Gʹ5�:&�·4�Y
5�x���F엻���~�R�c�Z�/��\y�}�*�x�0�^�;B��=�=��d��x'85�[ +�ʍ�)�G΅ⲱ�dM����u/V�1ӪK��q.����1��`f{��G�@�gͅ?�nh�6�h�Z���y��V�_�y�^���འZ��������ɣ��ㄉ%XYh�ſ�b6���	�Skښ�T�Q�<,��2K�E�z�?��ls>߹\㌿�37����$U��ܪ�M��WR����=�T�u6�����f��m��In�Ԣ�	Խ������?���[��ș�*�1��K����Ʃ��4�s�a�x�t�5�y77�����Zs��$��I�<i���F�8�Ak]�$�7�f��"U�k�Ȭ7|�*O�ˏ�/lM{P�d&��X��[�B��`�&Zh��8�#6(��B�/<娩DW�M�=g#����� �{U�l2~��l�s�
�bқЮ� 0��R��@ys���_�f����j�V���� ����Q��Ž�ϐ�T�k�	^�MOMs�>����$�h�ݎ$9�S��.��tF~�s�c�<{�f����7��{�O_,9f��+�#�x����L���P�.���c�S�7�S�Rp@yef�^矞��m?ӗ��"���^�p� 1��I����|?�w��wӤ��_�?,��c�%e�5���J$5��B*�^blk~>6}Nf��7��ڴ�U6�f�����o��������$���Z��b�ځJ$L?,�|�m��i%o��_��w�4�am:���r�:_�$���;�|��L������2��	�s��Y�]��b�Ȣ��Q��R�@x�2�&�j$UI��;�3���2�8�J���!�3>���Z)@f}r�V(�H��ʻ���%�[�]�ד�>���S���U�<�& �%L���yUsw�\��@)zN>`!��b��@���ZÛ���KC�ːʔ��sk�rwT��s����z$VK�*#l>����1�����ށ����ARQ�3�9����(��t��U��0hd'�(u�#�e�oMwu#6$���_3�X�L�RY,�]�i��=cťU:�BdUN��p֪�AKoP�FT��u��d�3ݸgC� (Ӆ!3�aZ���(�T͚5�Z��?k��N:_����<y���3�����8�#��ҕJ�^�������C�w1�~~'L*]�9�懓���[����`Sf���d���i4��v�����U< I����O�\T�r]�����_�9
�h�+~/WCjdn)����%�������Z۰y�
���"��֢�f�ܨC�ROsh�x�w�%nj$��������v�O�AK���,�^q<bx����͎�4�S���j���tFFЧ�w�����)#4��t�7h6�3��h��뎴�އ�:�<+�Q�T�aK�Y���v/a-�:2>�"2���jR-����
�$0�M^����b[�[ٱ�nw���Z@��	���׏�_���BRM� +�������wDA�y�T7�2�mοD7��e�S���;x�����T�V�J� 6��5����^����O�9��R�u.�L&ù�d�p�Lu
=ATF��<�.�$��䎣}�����Vn��V0gO}�3�
oWyTؖ�s�P��]/_��wBIl��r�m�)�����5�b|�s
��.�KG&��ڛ�$G:�M�eA��c3��B��[���Uv���$<�u<�h2��P�1�ڲ�г'n��)X�baY+$<5^�`��b�$�fe������^�a�k�=W�vSw�l��������J�Cn����8����"le��@Ո�����*��m#�Xf^��IV<�� ɰ����~W̉5��j��z��� "S�
�t���Q4g����h�,k��J�F1���[�P���Ļ�NՄ�;��'�,j���j �e� ^d��� ���z�+;�uw[c�vR�i��*H^�}��9BЭ���5��O�>an���9r��C�j���v&\��⨮������[L��G��R"6BW�ל�`կye�K��N�)�<%�C��I`ޑ(v��zD�TX�D����b��T�jh�)�z�j���?S{��YK��r��q{m���B�	��S�Ă<%B���w���~�o[;\�~���מ�E#FH��H�D<�]"a��W����y�3r���la��/�T^T����l�B�H�خ>�� MA�A�e'���!~���e���z��
�U�B�q����������/�g���kF�~W��|�������z��y�^̳}�-3U�s��A#]��^��]��}\1T�Y���-`��xy�Z"�4�#�!� �����* 5/���VS�A#^�Db����_��{����z+���m즃�i��=��o��{��p�&��� ���74�\��a�2[&��i�6�A.Y���
�%C�"�ԝ0hW�&^�0f���2��$���+��x�:Z,�-��=o+��]���4k�עd�'�$�V���w��:nY:@�5sAK����萐��b��v��^��Р�-�4�GȚ�|��j+Q)�d�<� �~4|�a������j�������QK�\��o���
ּAl8�?D����Xݐh�!8����M90����F��WY�5�-�s�,�NFBb)���H96|7�&J\̖S�4��I�uBx�S<��y#1qF-���`c�|Ia;�.y3��(^Vq\'E�E��,5H�D�&�O�<��e�˓=�Fw�"�M~�!F�R�R�F� )�A���tq˅s�-	xdW؛{g&���c���:��AJ���S�Z���,�p��ޏD!��*�ڛ7���u�ѣq��~��I�2$jU�r�d]&�.v7�V�j���" ��H����g�kQ_5l	VI������q� L�'>;iZ�T�1e��b�3^^�VK(��j}]��q�����ǩ��d,)�2(a*j���[�~�U�{�94o�r�FŲ�Н��R�R��\Õ�d��gyv�?���^
��3z�̧�ԦrxR��^>�c�yi�erנI�#V<^��*�!�?B�'�4Έ?��d̦d����S�C�&8򼗻�q�yg�����-˚���b��0�@�|ow}�����@�&�jʅ�������q�4�ũs|M����A��QW~�̏��c&Ib��5W
<1f}M3��?}��������3�Jwy� Q�g(���O���W���/��߱J�N!{�H˲��J�B�q�C^�Tc	S�,#W*�W�;�=�P��z�c��:�� ��a9?�M7�
��1�	�ŷR�ŷ�,�_�/�]���-H�q�c�I�r��6��1܂':� �M���z�h�b#o^�����b��?d@;� &�2�+?�e�`�^�mJ��u�俖��1^:ޅR!��'�.iw��8!�"�������1�$�jE��+Y_��S�cC�hט ԩ�*D-�AS-�`����
	��r�G�^��O�Pw�]73��C�z_P����Lyy������#c��1���x���yچ�T7�XGV����8����c�
���G�|�n�A 5U�_�� ��:�鯐�mJ�Ww9�y��:d�묆�?3���������LsJ^]�\�V~�C����d���ĒG�w�6�K>��Cm=�YC2���[�ٴ��ٞ�Qw���]-k�����fx���=X�W�=+��H��,��{�x�K��Bb��
~]K�t}iI��<�y.�T\�����k���σ�W>/����%	ʸ�"s�Rs��s%�����_��s���*��YT�%��@.|ț�%sg�,7��F��mQ�~^�;(��o8�_!{K=]j�������^Tʟ�LU��ċE�c��x%CP�mS}���$��4o���:ʘ�ww1���gل[�#a��H�T{�k6<��j��������$T��mv	2����F(�%���Xek�o7�g�}]Y����+�Z3Ž���?u�cTࢲ�h����9��CB��t���S.C�y^X����u+��YLOȍ�@�MF��0e}hh�����j�jY敉�}�J�l��n�Y�+�6O�3�K�r�����N�4,"uq�<N�s�D��WW���ܹ����,��U�]'�u.y>�U���wh��SkZPvMS�V��^�We2<�e���ޛ&�9Mm=tUq(��L����Eb������L�M�<m���W)x��\v�9���X���6���D�4_鈞+v��2�dFj{;D]yr��뮤�C�H�p��$�[e �2tădS�h�<�=6�Mvߡ:U�����U�dg�y^r��nx����.a��*��E�y^������J�R�S��u�^�j���n?�[d�'IB�J����}%ߟB�{
��T���,A]�V�,	Rď7�fA�ѿ?�.�*-X��)��S�D�<�D���kn�4�m�����W#^71�Zu�<�%>3�H@є%���_�!�	7\4�p�В�뀌��]���0��~���D�;�_���*�K���P�H#k�>��N�H��:���\���e�����찏��P_���<���m+��r�KZmFY椒Cjf��$��}Mk��U����͔~>�=��X��H؝�<]T4��ݣ�Em��"�S��e�k-BO����NƷ� ��A��� �k�#���۰�@!�~<�x:U���bU������,�`xKA���/�'{Kn�b�V/�B"X��2;Rˀ��ELr����\s��� 	~A�Q��F��N;ž<�ݔ)�m�k�4Jef��o��+>u	�G��[�b�%�d-\v��3�e�Q�e�+�]]���SJ���vb���f� ��C>�l�\� /��[!��ꈌ��P�ߜЋ�9��:�)S����@3�t���~�n������,	W_XB#7.��OqY��CL���lEi��9L�;^/b�*��k�6�����i1x���KP�N�B<\�8;
��q��T�i�-�^���<�:~�$/�ײ�g���f�t����vsGE���P}SmA�:��e��m���D	��3�Ta&s9q�B#C����߭r ��Y'aL��a4n��"㉨�GȌ��e$[5�Á��]��c<������L=B������ ̠�h|�4�ۗ�8��$4E�0T�"��g�3���|bz��[�"2��N���	�^��h�T�&A��EŰ����8-���������{C�>���ã,`���d���먢�A��e�c�m�W�2�f��v���^���\���^��ܩ��*���do�B}2��}�Nrmڂ���l|<�a��+\�7��╦6^����,�;sw���g��<��L�{{˚��:��X��yݭ�*Y��y��{E}�� ��9���-��y�:&�}�<[G�_!�ם�,�[A�6�=t/aZS��7�c~◮~C���^4���(����J��t�z�ʥ�����q{u�^S��c������O�����,���锿��̒�#U'I�o ^G��a�|�l��r��×�O��9/�2F+L�D��ܟꢯ�#O}�����:�W{��	Ih�h�$��Fճ��t�ɋ#Z�����5x���_�3����A?{�:6���ЯsZ��'����)�Ip��Qot�B��&���Х�X�*Ɓ.�? �*�v���ю���
���S��fs(^����E�Pyo��K�Q��Ty�!8aw�j�*K_9h��[0�Kg�i�w �8j7��!�W�@LO?�޴��r��}�V�91,�zuJ�#g��K,KWs,�WLUl��G��J�t��ԇ�>uP���m�L�ʽa_�3��`��+�r�5�8���$���Cs�{4zE�p
(0m�>��A��{�wJ�����k��T�ΐ�,3�09�� ��@F���*Rv�+���݀�T�EL�A�l(��"��/*���X>%�)(?�RN�EQ���B�N�q�rK?J�&?��#�� �Z��Ɇ9xy�yZL�>���Ҏ���~��Ѻbt����~O�4�ӳ�і����#S�ȱ+^^l���LC�m
��$���O��؀a�	�&���_{4�.���>��Ѩ8�W�:� %�o��7ݝC� �e�����?c����(�_(p>��S��]�l�Z����q'�e6��������޶($8H�����(��anY���{��������ʪ����ۥ���Gu)Qb�a-��y��Tr��L�/�)Z�-Ki��L�z�� �p���ӗ�]3����O�0��G�]l�d ��W�L���<"��3G!�I��M��`L"w��C�Fϲ�h�6��k-�S�>�"�D���b���[�t4g4��H�ܞ�s/��@W����X'�B��}
<�uZU}y"�ʺ��u#ʔ��Q�r,f�~�Y ����ڦ�^^�"���B�#w��.�PlwY�6dO�[�u�z�@�",�@��Ȓ����|�b2+�	o��A~�{nig��V;�nCb��d�~�M��x�I��nԒ�pC��)�J댉��e������>�K��՜}_���a���R1M�P��yo���R��Ȫ�V�	�
6`v����Ɵ�<ge7��,d�ȰʻS�K0q&8��6׾!q������/�Z�y�*�P[��*���ibe�e�����l����[+�1.�<���rULg��.̟��������D�3;�ŉ��u��K>0�O�f�戥�x,�L���Ӧ>��n�ND�"���xs���Fw�0���Sq.I0��L�'Ϊ�"W��$Qq�>��;��3L��ԒJ�eͣ����_���~k�"�e�����RW\Ʀn2z9���1����F�א[�����%��m��y�u~K���Z����%��K�R���x��pj�w����'��^2��es�J�[yoF�y��5\�vo�����8���\Ix�M�N��H����0�ƽ�~�Aʱ�a9�ߣ5?Þ�-,��{������?�ȩ@'��8�72�#z��]�E��϶U5±Ԥ�ذ�⽯$�-	�5��� ���d�1��3b�i&��Y��ԃ�s��ڍGOʱL��Uҟ�Q5N^�1��>��@t�j4Z�b(�o���S�t� �s����d2���ǾP%V��؝iܤ�ѹopR~�^]l
x63�Ĭ��n~�������݀�oq�-8I@��}d�������²A�JG���M�q�8;_�"�V%�v�T���A��Ϸ��az�J��-1���h[�~[n�j[�+?㏛�l8�[�u�9��B�5Գi��t�w�f�/7����Ӟ��Ay�33�<H=t�^�QlZ�EMJ7�ܩ�g9N҈,��|I�%�x����n/��R��J���t�I��2���9 �|%� �\�����'�A���[J�U#A�{F:��\CJ�Y�Ƨ�B��p� w� wտ��^?zՕq�>����{�K��lj}�%�xEh�g��.M�ֆ�£��o2��\���	��b��P"��zԲ�ɢ��x���A��s��[���k0�F�9S��ћ )��ME/+fE��R#��ލW�-�(���i�%��G�i?���e(�n�Y�;x|`�m�7�B�ٯ(��)�d�2���P�H��P0k,<�)t߼��It���R��NZ;�(
���YT��p�o�(%����e��Rt{��|���qN�'3RC�U��a��Dw��#/*XU�e ՝39��K�@Wx��i(����/c��i����x�0+�fJᛛ�-�p�pb��:7:>�7,�m_J��Y#F��5��t��z�Ĩ��r5���<��%�֔;���4�x%S|N�J�u�4n#�Wx��"�x3�����֕�*~�H'>��g➖w�Wïoo�4>(.��JP��#�?j�כ.�du�{n�;H�"�J���͍��b̀?�;���.�:�m���ܜ�$&r����Wd��t��%�bT�����A��Wf���ՙ[����u�x`@L~ w�n��((�WR����`M�]�1bRE�Rq���R�#��ޟI�?����MG�x��oe���]�?5Kj?�+ChI�]m��Ռq�D�6�A%�	��H�f��ܔ���p�8���d���ޮuL�L�R�I�; �6�J�[G�G8^�DOS��`��S頙_���Hw�CBx� ��\c�܃z�y����� <3�XV��t����M]jU_n��>5�����B��oixz��؜.O�3<����eڹ1�&$�M��
�&�#�M|�noWVT��MG�A�AQ��D�`�<F�p���N����OTy��`�^�I��������V`�iB?R1��V����m
��-m̱�ϝ�~(�阧Β}����)�K��]𡊕��1�4�!F��o����e��Mx�4�5��@��w, 4���ր�E��fa�����V�]�B!�y��ש��_�p;�Go���:DS�F��V��i���k��[؁Y�E�ڡ*�\?��ϭPd��dn�ή���rDGI��6��-��5�F�Yj�6���P��&��D�^�^4��^���$�F�H
��`?Cay��u3�$��LG��s�h����� ��o���}nn���rc��@�hd�f?�b#���%��[�U�D%���r�(�:z��c��	V�'�%QIxn�";��i�j�Qǣ8�r0��&����_�'%�zYn�rf2��G��Hu������\?N�,ɓ:sՌǔ�"vDk;_��x~�U4p���]ޚ��#;g��}��Q���
U�m!Ɖ�6���ʟ��?B�L�p�:y3 ̃8��n4�6,b.X�{m,�������Ncd[�����f�H
^RO�Y�E��X�DF��3��Z�R�2�>��_���"ʓ�&
땏�k�ұ4j�<W1���q9J���bR���M�u8inL�c��DDD�I2�^�	�'�7Io;��{x��\
rg��-ӵ�d�-�.U�D���m��̹�;d�AB��׊� r��-,�� q@���n�*K�k����$�ַz)36�����T!'����	p�V2Kon�3R������xz�����M�ؠ:�|Xr偊�����kys�1C	�in�5co��['c�5K�Mf\M�'T�A�9���Kw�����ߠ!p�8��QBu�7�T}n���q8V3�@�.ޤ���q�慓�ᴐ�]w����V���dt\�@��Ϙ;$#d&�9�IX��(QU'!�����R��B�� �B�kHzs�T��):����N�p�H��Lη�P/���Ȑmҡ��ӈ��]�Y�ɨ)y<�bN�Yʤ�o��s,�0J4H�X���E���ҒzR ?���e�n"+��e�v�ޢ�o�АY�ۓ�������<���հ5^LJ}�L�_��.�T�:��D}�u���A6������$�M܎����Ψ���)LT
��YB�B�-7z;�]����g�T>��$Up��P@��O4k�4e�r=�ABS�|�EH����f����N�	�H��	5���	�^���G�O�����гl�/�YO=h<���`q_��B0��/R��vCn��zy�'�����$�
�s㞭��QR쵵\�כ9�8Mh��������:��sX*(�ܒ��țژ7@�F\^���A5(���Or`>��K��r5����E늯��]�`�lo���3ϻ�1�ƣ��,�;YW�F�"@�q�>g�LZ�S�� 	�S�#�FpkyK�QhL�*��	���HTԢm�YQ���]}ð�	[�Lz���ޏf��6���w��Np���Ru��S�V$����-�A7�F��/�ͼ^�uGe�=�!���0L�j���-�w�~DA��[�T���~]>��j��qz�_V�n�4U4�̘���}Z-���,*��Ma�+'K�Klͳ�����~�U	��+\K�h�y���F��yC��jf��$�LQm�9�5>��,�~�NIM��b�4qk*^�XV���1d"�|N�����c�y���⫢Y�<?Py^���Jf��k�g��Z8)n�]�'.��W;��K|"ׅA����C@bӃ�vvnB���hឥ�9��'"��x��*�_g,ne���z37�ǰG~ѳ��B�
�;����8"H=����6_�o'U󢔰> �B8To�G�n_�i	���R��B��� S�*��d��w�!
�����`M�u�&�v �;,_3��$��Kdʣ�s��Vg�.�$�Z�����ޡU��I��I[�#e���i�`<z?70��Cj�C1��3}=�F*����ªgQ��P]��ҋ��˦1�e�ו�����&|g�:\�!���DL�p_�V/F�
��]�����	ۿ�.+�S��v��u��*��lݏ6X���܆\��m�<�O�_�#"��Eu��Y��FH9}�8��kr���]�*�l�*ǭ��/��vD٣�!���qie냩�F�L����g[.u��}r�le�hL�.�t�����>Vn������0�7d��q�Z�੶M�}�~?	�-*-AdX���i�!�fa��sY���s�XHR\H���3������� ��>cm�afYo[2 e�u):�ގ�Lz��O�����[�D�d��B	�{�-���p�[��H��!��[7A����`��v2Cv�v��N�nj}>� �Zw��en�?�q�D��;r&��=��P68��t~c#��]f������2�i�7o�O��)��p�dg�u�W}����y�V�������g�D)�<W@}�Y bs�`�A�H�H���}f�1ƱrHw`m֓Q�;j��=���(!�P~K�s�Ա~\��i)f.�.�ڡUγ�l�l����b"*�3����6�S��['�����h�+���I�@]{%9g���d`�b �2>��ޔW�K띶٬�Iũ�)�s�gR/��%G3IcʢYy��,@ͽ�(�����)Vr�ׁ�s��^3s%3[\yX��a�%y�\�����o��uP��Ц��3=b�C�N3�s�L��t��u,��Ł��wM|�FJ�#��Y]#��{��um�A,#ջ�֍y�'���J�1(�oՒ~f?Y8�*�)xGDB�����[��%�Fż��a��=����9�n;��Pޡ��e�5F玡c_�-�D��&��y��TR�E�?TDzO�j;����[���N�e]�S�#s�,HH���eJ��7!�tS|Jq2�a;ެ��I���#]s���0�j�hWb�s����D<�DZ}H֛
˰��-Z���7�\C�Xz�m5��ԛ�ͻ�z܊F7��L]�c���z���[�F���r�M�`8��&J��ܾtig���M�J����D���XT=�[
T�?�f��Eԓ|-�.��� �a)Q&��H�5�C~v�~U�6�HhR�G��(=c�`��o�rl�V�s�r�_%X+⪨�ae��GdW��c7̶����h��Wiu��S���f(%>�l�o��Vur��|���W9��7��z���x���s���s\-�`L�C}Z�ۇȯcǲe,r9D� L[��c�S�i�t�\3eC�-�a���P�iN��_}��ߣgxc�D��D��i�
~0���s��@�p��N�H,L<ox���pjYZ��fX�TnW���Rt�o<��GL�_Mk�\s^N�&��]���꿩6���b������b셰{�}[��;��nx�q{�8��WB�F���i�?�8����*��8���&M�v0�z�I��1�g�̆�Ȯ�|���2���q���Hf��*o�?+?�I�� ���e.�$wǯ$2�;uA�܅2$��@��G�ݽU�혨ȣ;�@��*7�w����@Am��1۾ٸ�?Xh�z���Y������`�ZF�a��[�,�Am&���оX�%x ���l�qm3���;J'+�ȃ��i<�ǧy�V'X�����S��,A�sf%�-=�k ~�����F2Ǯ$���e���ɝ���c��LU���|�f��H3U����������W鐨���	Fh���1&I��叐��0@��.�~�LJ&���n)N�KϿ�)ɍw�s4�d=���p�� ���.P�"`����E`kƥ���v��P�
]g�0�/�x�aOQ!�h�1��I{T������� �~�%~��W���D�9R;���W�eb}�d��v���hF꜃r7ϳ��&c���j���zx��MꝘnH�]�v'x����yDa�/��Y�ԯ�@96?���ԉ=�x�畒Z$7�Y��'�d	<�O�ۼ3!���N�����}A�1/��*�5��m���A1����/N�&B=��$:�S|�������6E��/����|����k�	�����ʙ2Ψ}8w���t�H���D��~P�
�A}����:�eq6W���J��\��-1g7K�Y��S,B���
�����o̐V�ǻ'�aV��HY?RkЪ��A�L�m�����	�;�[�
�>�������E4FT���|G�x�*��Hg��3���c�3f�K��	�h^��9���n =�����VoV[(�Y��J�.�C��]���\�șM��~�-����?��	x�<Z닎����}�R��f���D����}�����?���r�Pw�w���}�i�c7�
��N7I����'{+�e�9�^b���ҥο\]ڨPĻ�8g��_E��G��|�������땝�O?>�|b� I�}�R~��C�?X=
�2{�V���j�|g��j�u�B2�Dw���+��s޷�7:�o
1�	��jy2*4��\����3כ�m�1<��@H��NBݙ
�~=x_��ݕ2�9�lN~��a(�~����,����-�:��J/E�! �rp�~��
{ �Q��������{�I �~��	B}%��ܠ�SU�Y@?,���:��Ao�<�ur�e$T{���gT��~H*�Ԙ�*LK������ i��`X�q�$4������󤺜�����u_0����ۍ��.�W6�+�@��J�]������E�稶��6;b'&,�}�*���eF�ީ�<a� �6���O�C���S�C�;e�dL��f��P��d��p �3���'@��U3)�?�j~"����w�M��j	�\	4h�;������J%�'�ևL������O��un�B�1U�K�v�	��-,9n�"�a7�=\���>��ھ�+�Bs�g�Zb�Λ��wU�'�pd�H'O%��(7h��W$p���#(�����n�M�����_�P�e��K�Y<�c�e��A;F�4�g� W������~��b�5����?�W����B�wV�C�?%����Kp��������,j`��{��$Nz_�u�r�G)��Q��/��{�7�0��>=�� Q1�x[T�1B@5ws^-�ְ�;�?*k'�Z�3��E�G<h��C��#k������3�A�`�����Y����]��R�B����.��vH��^��wǺ:7o�L��qI[0�a�{m��қ�����Ҡ�(��X���6�,��H��܋w��N*�_b�e�tc�>~-ԋ��_�`�7�����P�ĉ��s|���)_�铆��8T�Ϧr���n�3b]C��\��P�����T�r�i#�<�˖9cf_���ܒRM:�Sma��tG�bc[�nY����ٵ{hȆf��A���OG�,�P���0�c�`4�HJ�޵`��|z�#Mj�S�}Z��U)��CSf�����ҵ����������e90��_՘�V���ґ�Z���@�s����J���>;�^����~�P�n����n>�W��� �+.d�����^��	��C���Sm�{��D�n"ē��ӿ^?�V!"}l�]�k��D�������5�'L>X#b��Ѯ�8h_ e�Vu���]�HWi=��o���i:M�f���_~������������G� $E�)i	Oȶ#�-�����ɘ���4�@��$�)�<(JnQS/�yY�Mb~.U!E��.��#���$��(�Sxc炤�*V��C"�!V����Ы����y�Ӈ�1}#�#��k?��[+n�݃��t̫#�Sd�qR̿З�Wσ��>_u�(�]���zO��LI����BEo��ua�zJ�fP0��%F�{f���83cj�܇h���K'��Ǧ0t��i����1~�J��^���K���y]-�|�M�bW>�8u�����f^�"^�"^"����,"�JJ�g�[�ʭ℗gM�Cd��!�r`���M��R��c��w��T)�\lPv���X9yށR� cDd��E�Br�>G��^x�b݉IG�t�$�c��@~��O~��37�Q��`}��#�w3zUa�i��yÎ�f���,��	�ꦀ��ko3MR4�R֝�!^E�S�ݺ�!�Z����L��(������{���"�;��07O�E��L[��N�<�靸*zl@�.ؼ4�/5�a�w�3��z4�:�Ȁ#�u��k4�˳�P_n��
�|�DD���#r	f�eo�ӬH��,�!� ?(��f�i�mk[l�=�|�_TfGp�����B#�������"��m�o\��Ա������v�w�r7˹�e�۩�j.�<p�G�K!��<<p��w���cʜ�p��i��HE����gMuFĹ��>�7)ԗ����l���DV([�g̿�4r�:A�^E�s*�#%�:����,�pje�gb�8^�*%�x��1�e8E�TF�<0��<�PfMz���0ՙ�D��B�!��--�����n��:�:3�����)"����u�@�&ta�.zñ��Jv�� 3�A!����6���K�y���\�Ѯ�٬W����Oc~�^�}�#z�lM�@s����ž&�ea�����e��������Wj�rX,ٵ\�F&�b��k<L|�EK˘1!���e3��3�k�1�ڻ�������ˠ����׿_�֣����n=�A���
2�s���=*�k�Ҏ۵�a�J�1;��lj�1c�2+��Nf���uv��bl�z	/�{���Ε��Ӕۂ�~}��Hpӻ\(H�|zpq}t}�yr���v�cLMOXk	Q����z�����rܦh�C�G��n��u�m���q�ߧ
"|��GF[�w.:s&����5Hx7�����X�Vg�[yL�u3��`��=B0Ե@��f����ߣ<�W�'}0�ust�#����(�A� ;c{�;��Օ�U?]H&m��{�RU������è�̭���'y`[)�*��v��Q������Nޙ����U��NncO�zӓr��I�:�X�P>��<�q� ��<�A�,6�Dޅ'�Qh,1"Eɰ���"M�KA��5���U�(�x`r��2�����F����#�dnDA�<[��yXx��)��j7Ybb1� y�2��{Ē~��g%�����2�����g[H�;i3T�|�e��n	��Ƃ�<���a��1�C�m�ElZ�ܰ�K��K�i����sD��4)9�6�G��wIH��gձ�'�P�wp�R�v(�8��R������0U���W���؆9�ʶ(�8��tG�g�i������j�y�Q���J���"HEJ�KS$R"B�^C��
��@��t!ҥ��{�CH��{���w�d2��LΜ�^{}v�s������Vː���!�*1�LA��Jy��w��]cD�Go�ׂ>ʦ?�3��5�����yN�gґ�W_�lYxs��=��G�j`l��~'�Fi���X����qʾ1��u�s �W��Xv�^��vY�飝^yy��s#&Y}[����C��1�2>x:���!pJ������M�N*X��)�!�!}H��@N�uڜ*fi�ͻ3�q�e2Y��Y-N�w�濍ȣmo��oj�(%��W��T�t���'F�}n
�L,A2u�5wŌ�H�z �W����d�dn�= :eX܇��K���{�FI��:�P���t��Tdwz 7R &��	9,�k����0 B	d��}��.�|o�Y���(�9G�?���=g�+v����s{��}Ιi/�*Ȓ�g���j����`\V����[��O]\����r�a�M$�¤���N��g'��8.E�׭̯[Ι���3��3&u�E��&��>�3����D��8��yO{���>��ϡ���A�ϱv@��0�l/�֏D��ns�,v�+�]�K�-4O"�YF�%�<�B�\�@ŵ��T2q�r�z���J�s_A ��a�P=J~���"ds��u��At[�=���-#�@�7d���ˀ��]ǾP��⧊!<m2.%{��Dz�_�c-e~�s_e�:��X�s���o�W6+���
���^�n������z.��#,��Áph�r��l���]����7��Pu*6$��5�� p<��C �Pu=U�c�����W�p\����qF��[�u?lsw���°[��)�ףH'Ѧ���m\�u�{�[st��=|��o�5)��䓢N��/���}t��%?��N��*�M�KN�a�9�|72e�Q�������vM��Lp�sh1�4�qK%��8��p|�i\���+��o������(&���<���Z֙�wh?2J�}�ⴧ��O���,�DrB]Kd�tT?P�~�����T�F�$�8���DS��V|. �H��43�gݚM�bI#�U�ا�G&��:�?�\� �'͌�'%��<#]����u���,����~'?���9���r�)n�.�k1!��|a^ķ��&M}ӵ�z�cd������@�����m��M�ܓf[#�ix����m�����?Q�����r�c͡�B�x�P�^�,������0�U�[��ә/��c�;`a���:���H�ʱz�y#�)��pZҐn[t�mZ,�t�Q���\~5�$:l�f�~�m���R����[�?�+�ꝸ�b;v�Z�@qz�˫f�N}��_�t���1/�/��W��{?D8���m��m,A1Dd����'b���
yۢZ)]Nc>n����)�<���{�)xf�{����-����ڨ��h����<;�f���q�~+xB���2�]��i�kt�c��FwY#|s1te-��~�ʡ�7)x����4��=����G=$�Jk� ie�zD�-KW���@7�4C�+�[$���]4��؄]�Uh�ܖ`Z��}(�Q�[e�|��Ϋ�m(�6��$�R`>�_J�:#��+���sR�Ƚ+B�����V��Vd��}��-Qs�Su�����p?dO���1���\9&hH&*��5u�C�%�N"d��.��Տ�j&W��g`��R$A~.Yr4<i<���g�3;������y���?��u��C��r�M�Qu���S��m;�n`�m[0Bֺ�/fF���-��:�$�,q�N��(~K'���
��3�z�U��j�%�6W�y�-:���\[瀙�V�}�J�"�I����|���l��9W*�-0)*Κ�ª�֭_��B �Hj��H��J�Y���l��EgF���o���5)���UNJ�i�t2/,*ހ���<�8YȀ˝^��׎�7�����a���2�/���q��_�g�I*�������C9yg���V�?�c&���.O+����4�Ĭ��8Id~'����2�,���wٖƠD�@ڞx�5��Bw��f��i�!�Ƣ�XF67s�Pxi��e��x�!�]�ۆ_�±`8�׮���_M�R��k������.�+�M��x�/R�=��M�Mt�>�}x��������K�������\$�E/�}V��W-wP/\���^���c�S�l�3�$��Ӡ�M<�����zg�����������O�%�­�@	"	%�9C�����@���E߄�M�˱/��9+���ۃ�ބ��ZIo<g��$�-����9#��V1^�"����>�������_�}{�#&����Z)�o��>���o�t�OUOY�ߩB�Fb|�m<^M��Jlh����#�C�Yd�������k��`����Qd':`Q���%�	Z9�]��߬HگX�f(y,N����ż0�
�,�i[��j�]"R0�VM�)-כ{�E���a+���U��L�>'��Q���8<��ݻt�ZΉb������-j�/��8�!�j�(��-��]�����[;)ZV(�z`1�v���_4��W�S8�7W�:�]���3�l��R@�/yu�g�ڻ��#��߱�^/�Te��1�ן���J)4J�;��hv�+b�'V���4M�~���6lmUF��̽'�Ϟ��t���.
z�N�.�yO����N媠ǒ�I�����4k#���l�{o�J��.�;۰aH�$&x�#�&
&���1t]�;���g�|	6vgLݜ�7�r��My�7�� [l&�#;"���3F�2��_ĺ)��/�GveEd60$(?��J����|;�������s��f��u��ܜ��Mu4��|<���7�8��W4v0���+J��_�5
��$D���[Ä�ֱ���#��s��K���M
��a2u_�I�E�B�����Z9!�R�?$%D��vB�=�T��>�[�؇��x=3��U�'Be���^'9(�%P�_�J�>[���8�����n�v�-|��r�8��ڑ�T6P��^ �l���Ѹi��$��fK��Х�g�7��7�&&8�1�b��'�ʾu��@��aoH�U�qbk�X�kŏ�����?��k����%0~��WQڻj�@�h󳒁��]��/�U��0�M7_�:n�(�7��E��,�tc/��T�#�<L�M/R�͓�;�bؓ�6�yp��<ᗗ��5�O`�k�Ǟ����I�����~U*���_f�g�+�ZI��#��P"oPc�Q����+Sy��
?�ɾ,٩Q�6��=|��G׉�0�H �_�z�qM���EU���&��]���P��yI����4 _~M��TI8G��]���x�
���~Z�
vō�t�׭
��
U�<�c�����S���]�d�y�^D�-��w'�d$�ؤ0��~`c�����*��jpFB������R����>]P���M�Kˢ4�Ϟ��x����b�k!��\*	����qQ�t��RO85Ȣ&�ܳ- ��������@�/1d�G�3�!)C*�m}F �P��5�C����:�^@��ڞ[M�tQPfm�Q��j�)k޶�ҩ�laTF1�H�J�EP�=��
bzO}[��8��L��ܪ�i��V_=��2���w���>�����D"<����\�<��0*N����q�*U|��B;?�l�������X:/��ӏ\/����>�����pzx�^�����nk�5��''�ݷ��b�	c�������>H��	h�� ��ޘkl�Հ�&�����b~�W��QR򬮚��:�X�:�������d>_���}[��=Wr=��=�+U�v�R�r��Q�K�_��{N�8�jǋ�"�R�pC��.��s�p��in�ޤ�m�}�0x��n�=P" S����<K���E5sF)�V�b�4�f�<B�K'!�hN$r�ꆥ�� �T�;�;�J���&��ݛ"� dX�d��\Vыg��`��鈼lVHC���D�a� ӳ,+1�:�Xɭf�0����7�{��z��3�D���]~���ۻ�#m&eo=�Ƚ|�$l�l��Ae��*x�ke4k�Q�|�CZu9�0^Do6k��橥*0��)u� �R��[���1��� �-EL�.�A���N��-�����n��_�u�L�>����/Yt�����?Us��3�	+��R��-���Tɣ���F�(�Vn@�2- ��I�E{�'	Pu��˘T���!n�JV	�'23ʥ������-��!_�ukY���)��t��N�9|������.�iM��{�����_�z�50�7�C���D��oOè�i�O���I����k!t\�	ߥg��\��۽��rz�J=�����no���M�/�-Bl-��՚ū6x'�DS�c1�/�s�G Lc�W�cMq�����F��Iz~
k�>�1�B�t�Wp^U@H���K��S �ew%P�z:]W���[�\a�[��dٺ�r�Ⰵ��oey�	�U�ej�X��;����*�r�'�_�?�!"�Q���I�RB�S��Ѧ�K��ξ�o�nm�|�a����M���}D�c�o��
�'�����t�k����,~�-�By�}�=b.DW%q��SjVD�#��:F�u�M)*��U����z#	��m���Vy�[�[�J�5TOP����ْ�6ȩ���V$(�VtG-S0R�Ig"���f�2L����A^���W2�_AV��J�^�$1*a�֙��s�{he�drD��Zjn��KLۭ���q��kh�\���ޜ��������n0�ű�^���8"��r�U�l%����͂ߞ�m�#ᕮ}���m<0l�n�orٿ��OS6�-H���PR՘�����R�m��_ʄbِ��6��I�������<�.��8�^^�TT����Æ��zy�-�>.�:�r�h
cuZ��l�C�����1,���D�bu��|IM؞�j�]x^��5���1]�Ϋ���-�5��/����E�:� ��W�z�&#�3���Kj#�Tl-�yK��)W3',��<�e�l���1��I�WZ�mut115(�����
z(]=��e�+�f�vBb�i�j�
|�Ƹ���W:�
ع�;j�a4���jc���A���Q�.7Q!�v��P:S�ݛ'�<�e(��nh��fud��h�s�Q!�:��xU���l�Lg��U�N��u2����53��8"�����w��w[js��]�Ǉ>�"�����X��<�%����|�4��Yה��(O�����H��SA�X�14챏N��ʡ�J$�K�yU��.6���Dk%���\���T)-@��MF;B7ҟ���]QyR���.�1ǺW,�`0g(��-|�&=�f����t}| Xx�?�<����٫6_]�x���R{�\m��P ��ɗ��Y�Y���W]h���a��v�Ը뙴'�qZ�&���t\Ji�剞Ӧ�:�ZI�ԯ���3_���5V���f�}�<]qd|Ek�X�8R@�~i�d��H��o|�№�ט$�Ý������~Ǟ装��ٛm0nk�����ۿ����=�HQ���X��
b���k����r�۹J�vZ
�!���rl��u�\(�-Ɔ�#r�̴,��q��n���+�;����?S ��6�9�2��Uk��q�V[�Jxɹg�����I�w�ȖH�)�oK�Rgk�Dw8�,|�B-�v,�RI  �m����Iϛ�D����uX�y�0��;�UӨ5M������7w�*U��N�	����7l$�-j�����m�NN�q%yt(�>��a6m�Qy��P{/A��#A�^�s�D��2e������-�UKJ`�+�z\����"*P���9�P�dm������A��3a5T�Q_92%�7G�
�H�٧�c���ů���q��oq��B���k<�7�����]���7|�o�i#�����K\�wO�>�����/a��ʏw�۝���WE�6��F0ƛ��d��?f�����ܭM��?��@]a���Qw���g@�,�9����a���l�O!tBx�����k��׳T���� �؎GTlY��_��Tq�1�qM�ߞ��a���A��m45eW8����n"��B{�LgWų�����8���N�2$�B�E0
uO?H��UD��.)��a�"�t�Z&�t$g^,�G���y6-=Fٶ�d��]�/l��	_'L,�����r�|a�^R�����#̝CI�0\�Ys�B�Q��^1�� �������M�1hu.�Ph�皰���w�0\mXJ��L���=���t���6iʻ#�*zG���?gF�+Y1nօt��8��c�!�}��Ia�w��W��d����d��qu$��$]/�cf6NpQB�͉��4i�����2�A���)<�y/ɻ�\��@!��^��ى����N,�v|���u��'KI�^=�/ �A����~RS|-�S�X��n�˯�a9���#gуK�����b�|�}'��8%�QeH��I{X}l����^����g��~cs%]��7h�jG*�Z�߾=�?ZE���W����k7��/�p10~� (��>{\jrsŒ�Fj{�)���<��x}o~��u{�|���(g�ȫ _�i݈�-�n�����%L:��T2��{���s��\�57�%3�YGƗ�A;	[��2�&;��7~Ai�����x\�1��p�zv�o����G�5n6�8�
����s)Bv��p?K?���ޫ��kM�,������i�3�>��Z�*6��A1��m�mD'�E�hh��}Z�r��Z��&*)�����@$�Ň,�?��mE�)���I.P�(�}6�k[e{n���S�fѹF�oF�����������4���~���g�Vu˯7��|~w���"��_�Q%���EnPSй�(�\�4�:�9e �ǷÛ����̇�*jti��?x	�];~��Hh��m��������a�����O�.4�hq<h���b'�m�E���f0�!=�/�bVK�!I��+(ۊ��#��ܗ�$�VF�I�6Qyێ~��I�{[�����ϼo��C��������L�`��]7��G����
>�,j����'7�o0Ȍ��-�|�0m�єu���p��$�1]��MC^fA�AMR����InZ]�T67�U�Ñ��zvy  16�-���]	�L�U�M3����<�J|*����i���<"�a��te����3�?�8c�?+�[�Ν0A�n��ӡ�мE��O?p�G?3���d�X��e5w���p�leI���(nI`�G�t,�8�N������5m�ͮ�{{|�l�FH2��Q��$whlq��9��x���r�t�s�*��Np�^��|\5i#��{O�N!!��j�3iS�v�O��S 2�|�&�S"¿F �s�H΍��t�c��}d*����(����^���&Dƶ�4�j�կ�լ��ss�vem�������j�򔲇���V���D���3P?�q�l�[��l =T|��O� ��u_ș@�'����	ˊ]dR����Cu��@*F$)g	E�?�!I�U�^꼽x4��P;��A!�cW��Xh�L ��P�@'c'�8z�2E��G����44�vl��oɈ�T=��K���Z��X���K��&1D��gP2���~ց5i��wF�{7�:�y,�o���%�ܡ��Pl�f�D�{�g��{���t�ԿUl��_���r&�5�J�����Sc�#h�W���bdZ����T��#���Z��b^�Q�����u�VM�u�~��~X\�>��� �|lzk^�աI�@j�va3Z����ض��߸�"mRTt�o��`;0�a�kՋ�h�_�H�,��rH�~��Ab�+#
���נP�!8�cX�nuT���I�x׍�n�$���^��Ƌ�rUޒ���<�$��g�4�@w,�W9��'�9������	:��~�6I��J3��*�Y-Iܬ� e��҄���J��b���%I�v��俙D W1IB���)�aªH��b��4��?�����;��1�:���y���Z�*��Q\��G-��a}������A)�:m�q�P��&IG0sΛ�6�N~�����)f������X��.�B�4����	v�d��xٺ�n��<�ݭ���p�:z�'K���n��{�����x�ǝ��/���S3��O:i�����ekv�b��n�p�C���F��1u�z��I�o�ŗU��b�������F�@ �Y�w!��e���}T{�v���Ӗ�uS��~ϐ4�\8��o�_�i�+�Z�^�7�}/M���|�&�D��u�?�I[
�n&���[�������E��Mo�=lF��ϊ���c 4�ћ����b�.>�^�CM[�12��SS(�a0u��h+��+�A1��CRw|a���/��ү���1揳E@}���Էrp'��������b��D$�wk�U���%Ue���K��vQ4���Zd��V|%�6ҵ�l*3���=z>j�/�>�<�%n���E���wK�$�����	��:���Q�k�@K���;��<�FѾ]�y���u��1i�9T���JA$����a���_�1�R��g��OVl�4�Q�)ګ]�!���In7>3m��f��1d�!԰��C�%��B��ϒ�^T�a�$OĢC_?y~�{�X�n�ϒ���oͱ	�Ve\���Vٶ0%]>�:�Ş6���my	5�k+Nz��P-�i�K�B�j�Nݱl�@���ySC�s{����M���m��y�>)Q�IN��%���)9�*�l�q��?�����G��8��9���m���B!^� ���p9���<���$�j���ʩY�j�j��W�V7��;h�k�W5�=��n�`�sph�,@��+��,���X�X?��*��~Fe�������ڷ�a����ӓ����\��3��<M���YK�M���������>�9\������7���SU�Rm:m����m7��		�Mk�M#}��M�kP����޿�$���DD�C�M��8JV�U�Н�IΪ.DJ#���#�� o�:?��2�;�'��%�i��ɗ��V�n�n�)�,/9��zj����M�ڪ���>W[_o�4a�>�88)���CK��}_zoA?��L��5�9 ��|#�X.~B��;xC7������c��Ud������{O4k�|�UL�TĒ����F���&�Bt�F%or�?0��'��$�������;D���SKjˣN�o��a��b&�b�M_>����n�%����y���28	�؇�{����l{�ϝ����D���,_�.�g��߿<�P��:|�*�^.�:��%�p��F�W+�$&�%=�}Y��Gm�����9��r����?d+�	�^+�~ܤ�i,�/a�?�[���V²�g��7�v�u��ͣ�]��X@��S�����Lf��8�`;�����:���)����$�r�b�N��o�|� 5-?�P�	í�ě�����m_F�]}�ҧ��7� �g�BOj�ߵ%gѮ1���� �k��E
������(�k���-[i����	g��n��'�����_o�����HOk�٩���ޅ��\7A� ؾY[I'?N�Q�;�w��m8�d����.��~���P/m����ُ�G7A�8+��y:|O#�Ӊ����wsbt~9�Td�34��%�>�^_�5�iX�B�m�NbA�Y9� �g)�P�_O��q;*g��ԑ�SB�h�}��_��^J|:��#pu�/?������3�
��҄&�&�L�l�V�(��$:�,�ܹfHRO;�{�)��b�C.�}��M5朿������BPY��/���I�J#I���b�q���	I�y:���b������ӥ��Tۃ�y�p����:K@F�US��YMt=?BZ7�����-�+`�� n
wHZ>�E�$ǆ��X�� �a��)�G� &{ǧS�|�@��1���O�&��W�Y"it�P��	�m����|H +�ٽ��v��]yGm�(#��~ft4	_��ھS���=_�A*&VPEE�k���{e�*�Bv�������w�PZ��b���B-�)@� �A��h��О��@��q��",�y2p�RC�z��HR�9H1���C�ˣn>���D����_x�D�\��0�ѧ�D����W�Gj"�c�r �t�;O�����ξ�:��)�My�41�t�/�����SF�7=2�o�Ѿ9��a0�E�r�"�s��,;c���T;���Y���F��IL���Ú�E�~��&��1!�|U�6���Pg�Ӭ����.��}�L�����;ϳ֞�s�'��*��U'���O�N��L�����,/��>��1����*���2���=�H�����.�h�ֈ>���CCM|���p}�]�-g����/r�褦��$w���[8N��l��S�`�  r��
QL������	��u��0&:1?V/���4�MT�.��3u=5V).:6lS�A\RDwB�O���O͋x��p[�����(ⰛD$ݳ�[m�?�[{�~�<@F��c3���d���"�҂2�� ��v��������U�8�����Qf{m�Z��E;�u�`�5 ��?��
�?���Z
y�TE�xZErP�tktM�1�������:���i3R�)5���.'���ݾǢ�^|�wF��uy��{�땘������n�X���wgױg�������o<y���ƩkB������/qQ�9(��v�c�z���v�F"q-[�J��7M��V���Ⱥ�c+���Q1BM�\��.�%-Y5fklۃ������M�����ָe�E]���m����)S����Vr����׳d2�(%߳x�	�j���Hˤ�+�[�ޢl�@LE�z��ܛٚ�,��)��O��r� �џW	��SfR�x1Oo�`�� ��l��"��_2̧%��!���/����Ǌ@�DG�x�P�Pg���x�Nאi:q�`��B��4'W��_��sKN)��Y�J$���0�n��0q(�<��yHe[W�/	��|�S��[�ݟ����	�&���^|�|�X����C�b�:=Y`�!*� �辏Ɉx��k��vO�v_�\�{q��%�]c����.�S-�����y�+¦aD��9$�̆{�t��j��f �Z0������_q�V�9�	"Ufȕ;
|�L�|�Ο��˼̐tg��-/��6����Sez����-�����z�}5��Д?#��&ʧO�9�'�r��	����YE�;�8�}ؑe�Ӭ������[c��4`D�Ϲ��M�ks@/�l�M.���i�:$��:|��LǞ��#rJ�H�V��-p3QA&zh�a*F��4fR�]f�k�9&�H�NJ������X�9��fk�&�\�8;N�GF)���Q0+kT/�rr���_����#Q�.V���mu���4��{�.�ٍE�Q@��] MxkP����2�Hz6�+}B�4_c��~�v�C�\b�-���]��rڃɫ3�*%�-i_�f��Cs��,�6L�4,�S�C��A��C�{�K�Ȃ�ɣ�VD3RŔ�8�(�Z��`��f����h� �O�(�(�
!��oT�=��f�^d7���
�v�o��*���c��>Wh����a�B�P^T֖��y�%l`W�cAA3��H���դKb�\�gȃ��B�x�:�V��]�akc�a��o>��흤���|�[n�Q}3�/)��/]�����__��`[��bP�h�So/~�i8�[�I����ő���HY�ެ���5#�0�Iec����6��b\E�<	�=����0��w)a��L�����r�$�;3��O�9�_?���]ç����miS�{g���L��=~;�zm}�3}/qq� ���O�Ob'|Z�FS���b�[&����^Ϣ��E��.{(<��ߞrü�T���$\wf��wYE�L3.�Z�@4��6���ޖj�{@`�p�C)�\��SW��EO��n%�W�?y*Ҙ�S:f�G�}��m���;�9Hm�N1QA�Yl�b�-bl����oDչ {�ٶ�/���}�#ט�0����t�A+��6�o�nBEm�k4�{%Wn�
ҭ])Eg�C�/�m��JX ���m�|��'F�����.�9�6U葌D>�4Q�o^���a��ޟO�];m��!8̫%yރ1��m���^,�b�i3��(��Mޢ������?��w�){n����bT�����",��a�8(�g�M��`�8��Ԏ<�?�d�� �^/'�_��E3=~èZ�U�!�.)���Q�u
����W*���4Z;��MN����3�ɒS�PD�ڧ�f��l�FcsF�UY�i���mdD�����;�9L���d�&)�E����k�;Z#�I��/�\Gk�յ�a���
���n+��݄�Vv [1!��S.�@�s�7<�*�y��W������K��`�@8B�u͹�.K	Xn��>{U_���\dZ��u'm4h�5Q��t�����2�Ok�i`���Иro�8��3�E�?r|��9V�9��kp��G:��&U9�a���w�fr�zWF?Κ�{�We��`
�X��"����>A b�_�{�4/�Ŵ/!�Bz�C�z�Gs>"z�j�iࣣEg頯K�;no��]6�eG"%\
��cxuxӑ��P�k�H��������6����k? q�`��(���_��}��h��d�@>G3 �D7?�G�%!�� ;<5 �����]�_�!�g�wIE�[&Ƃ'6�;㓝�Wg6��>�:�Ug�\���������2���~���%�{��$#	�, �i���F{�o���M"�s4�Ǳ�� ��x�tZ�{���_�:/(�;�B��$��S�O�ҽ�ĤtK��V:$(��}������!U�N5M����R%�M9��~c�m��t<p?�%�b��M�@��]�o_;l��������ӑ>�f:������^��d��6$�Z�c�%���1fݾ����ϴOm1�#�(KL�1I�������Y�~^���7|��c#֔��ԡ��n����$���m>��?��t�mZ����¨{����ڭ���~ʹ������T�etz��Yd����*�����{?���֘a=�!	��	�),t��\'�?2�("5R�� M��G;�8�гNI�0ҹ�����4	7	���W�g*����fr���ք?���Xv�C��lJ��\��ZoזzT�ZC�����aO|�ԯ=�U�^�<JA�qZ���a�P�U�z��O,K�Z��ݯ؈O�t�YT=��엑��R��*9�(⏑3GfQV���	A�G1Q����Ƿ?�Z��!������d!y��f#������o�#X�zIe-i�|�byK��-Kǜ���ѡ-�HGQG�΋��v�_+�P�$�ŐS"�gE�e�O<�{�\���>�����}s�sU�&�ƕ�Θ}y{�k�P�a�o%���얬<���d=���QV��.f�t�,����^�o��ěu� t���"�n���#�ǧߑg?�|���y������N���O7={*F'��W4�Hw�<�?��후Դ�ќz���R�	�g^�R�>m!�,_��������Ёn�g7�;K�m�i�i$�4�������n�	�!Ӟ	3�������_�BI����F�?�q��g���&aÀ�u���1�V�V�K�Y��SwG*_r��sV�(ݶzE�!Ft��>�,_d�:	�B��ݧC��R��-^!�2m�r>t/�P��Zj��DD����ǖD��#���[����j ʌ�������s��^П!��E �TtW�%��U�q8��{1[!g"�KW[�;�*�ဍ�B�c�ߺZ^
�?3	�v�	s܌���2�����ĥ�zkx�쾿���C)O�ZXᬼ[\����1oI���*�c�7��Q-���-v����3�f	��I�\M�Q�ϵ�mCc��T&��[F�g����p���4~��������K쬉�v�@ ���2޹7��-n��9�-ٙ�M�x]l��q8���ܮ��q(�׀7��5&�u�I���s6s��s?�/�������o���߷�D��Ǖ�����ת�b�N2V���\���J���f���ݴ'���M����]G>{�@����i��qW�d�k/s�g�)�Z�W��fE�İ�c�-�ho���j�L�i��ƿ50�Gڏ���0|͜�Ya!�-�! ��7���j\o^e^ߊ�+�"��n��ݡ�@�W2�F��L8D�y����}�Dm���oEAAŻ�����(4ٷ�jiX�s�x3kz	y��l�Ü�*���.o嫣�A����#�3_@_�������,x��\�X2�;�)B�b�����EA6���'�R�C�i۩���#���PY?3��N��Ѭ��:�~�ظd�������Fηo���O9�?�I�|ׁ����[���,L���B��b�^�0e(Ңs(A�N10��x���e���q���q���K��q)�o����w��qM��k6������̎�{�%^ga�t.^�M���`Ծ3�5��d�ۯ�%LIvn?�+�"&�����v�����%`CP}C���S[���O�H��D�yJ�ٻ�%Y��V��7{A6y˔Ү晘Lnp]��˦|�*>Ku�^��S�6���.j:i�|Q���4+�T|%����O��\35b;������3t$)!GY���*7:�O�i��<	�n�=��\��[@i��t���`���sK7e�ӑ2SX���'�����������=e��4��r�V�'eH G�$�Af�C�z�����s���v������@p�ȃ�[�����Q����[�lGC:.�\s{B*��y��F�b��L���P��F#�m�{�{P����ax<G��Ξ)�p��m��M�^hu~�h�;K��|����-���u��|*~Y�@�Va�X�4`�����
8�h��<�y9�B��Y
����WӞ��'��\y<�q�Q��}�$)�R�y4(aң��aL�<m	�6�a]Or�'��o)��X��&��y�G�\�9d����3n�ow�w��G5�~��7,��MrC7����f,�o] ���j@�V|�mZ#z��jg�=KwN��{�L�N���TbE8](����;5\�_\(�Xq�*������E���d8i�S�	S���0�8�y� �L�oHyD"ݻn5U���؆���)�>k��N�T�:W�+"	� ��[�اji�9�����ؾ�Dr�WX�1�m���
_~�2'�la�ժ�뫷O�3�~��!"�������D$%ӤF|A�n�%2c��΢=���+OOE�� :@��#��H��Hc3��Lo�ͱ�7i� +�w����q.�5���N0@Ɂ`���o��� ��h�V �?�E$�G���� �/�2I��mr��niu#�v9���M`���r������pE�i���������� �ȴ\��b���:�m�V����;6��4S8�<G6+��?�,zɸ�ɲ��˜?�9�"O䮟᜾f�������o/�y�~��IC��hlQsiC�#�ZBl��V\�K�hs_�/U�ryUc}��n�~_&��}��`!�)���Y���N������֠q�Lrƃ#�"ہ����|�=��n*�w���"&��K�l3�bN~�%��"O���~��^=��d�'9�;��↛[��6y5�:6��ۚhH�=,����
@�40g��r��!��>t��oV��=L���L�7��\��9�?Q%2��z�$�%�!��W��:4��?$j��ad�e���k����Øϊ/�����~����<�w$閔�-Z��؂{c�a���tLcd�V��ġ�Mg�Z�����k%z�����L�w�r�6�8�q�y�pGP���ҙ	o<6�tN�R��U����h]��٩�#6��B�pʭ�azάH�7W��}y�+V���Q`o�V�T�~
}f2�'{7�t�����'����o�&�7w�Jr�|4��{�í���s�����������,-�M���E�g"��5#�la��@1Mԃ�wYS��^>`B�}'6&i�Ϯ#aQ�j���������\;ƭΡ�]|+�4��{U#��2.t���tq\r����7���b'��]O#��y�h|Z)n�}uz��?r�t�W<�8�3��4��1��9>����c?ld�!�|�ԧ��LWl6�c����!���.m���h����M}m?iL��Cd��cd�F�by��?9y��8밦����%�s� H7ltJ
�� �$%�Q�V�I���)%���lt�������{<�����v���}^������(�y�]�x��sS�/���P�éTm��O�Xܣ�x�uD��������w�����VGʑ�ux}�xD�.A��������#�I]��80#�/о��F��g׽-�£<T#y�x�G�	�Yې �Ƙk=8<zC,[�(�8�����'-��Hd�G��a+���ru}T��x���ǴVؠz��������|=�D��C�tE}�f�B�|�.��l�;�t) 0���"����γ`h�X�nH ��8���K��3��e�I濋n��B����4��᪒<Տ�H���Wul��>ڋ��\�����ba;=����0Ix�����0���ɛb`R�w̒`�f��c��0*YN1 � 1o�,���B���PG޳I�uQE�";����3��v�IZG��Bz`�}�.9aހ�����l� �t�_�_���.��n�_�ޡ���Ow��7j.+Tp+���4R���������ƪ���8�pIF[+��l�~ܟ6^qD9_&�
� 0,���Kfw�������)� �t��򈂛ѣVH)�<oB�������#��:Y�k�R�C�m�� ��؎�<���\�P+D���C��0�,b�e�~�����o8V-T�4:04�_v�E�g��G^�*
/�}��h�i'z�<�?�&����R&$ˡz��-F���m�:��l(C �H_�xR5���2�Rx�>��!�p��as'��ݣOt(8M�ঢ`�S�$2Q C�M|Y⥧�����~�s(s��c�c��O�o�
�H�6���^tG$��lػ&��]H��/B��ʠ���y[����"~��'��^�"��Ť�E�5{��[ˊB'�;�� �]�:'F�,E
�D���kn�k�:}'Zp�^�~�����{.|�P�ᐹM~��r��v�µy/�{*�B�u��;�Q�<#���z�p��9j��r�=��n��S�3$�ĵϔy ����z����O;���Ld	�D 8��	� 0�_��	�+�?�j��*�-d�li�2��EB������� �����Ǚ�S����o���fw�N�N�'v泚�m�1�JW=�-�3�Aׂ��G=����_���M}�ra}'uw���Z�s��)O�|��?�&9f�Q�(%I:b&}�6)�J߁5ؘ4ș��,g�[�~�v���7A�{�8ة6�$�[S��k��z@���b���a�����q-=Di2�m:�\6�1HǌK
B�l�f��x�jL�!�������-�7�>`��f*C�/�/"�3O'�[�������&������9'*�B]L���Qo�b=Q�R0�gAP��Щ_�4<�a�������ڌr0�J@;���=ij�:�IC��Q�����q�ٙ_� `�P*:�9H���f�-xJ:0:י	�l̂ᒑ��K�����c���!������&(��ʅ�\�Xl���+q�{�U�&�FmY�������G
Dp�wdЫ�������.J�����,��s I��[����PA���aK5T��.�U����xRk���=����R��N�)�ŃC�sל��������(�������~g�oZ�d�)�EZ\�o���J���`@~U.i�ϟ��I�
����Fv��իRxs'^��ͪm>���d��v����P7�ե>D��v��F�<*�
�^�f�������j=���0�8}�}���������8�
�j�sε����
�?���Q�V�WNCG�B��~�6��4�I�a��+��w"w�LC�q %ׅȗ������ۅl�s�H����p�#��¼ǟ>9z׶N?��Ҟn�p�?�;k�Pz�`�"[�~_2nb�*��"��aj��Wf̄a��A��iL�u��:	��"���8���&�b��O��:���m�f�g�L�뚧�wU1v�H� ����m�)��?;b�@8��K@�OY�z(.�ux	��0���͜=�^����%�6�[�{�R���S�����6^�j�
���d�61���v��J�ݣ�G�����+1�2%��?�؅��y�F����)Zo�y�m-%`��R�JA�A��Ƀ����⦠���b��G�#0�R�i���":�
�����#�
��(��?s�������b9h�
	Zݼ�LzU������r�v�.޻,��H�T�%
��؀r
3�A���)�eW.�-!��5�mg�����i��1�_B~�
*��[���a~�Z���l%�u\o��e�}�ne=dw�{���|�����Iv�8a������@��M~�Nk���җ8^�h��(o?R�t�0�0�J�}���ݒ���3�8���A�xVA6��1����ڦ/��:aԋ.	f����l�ꈾ�k:^-�j{�33ݘ���z�ü�z�iXy`��*y�pޓz������f�t�z��"t��(��p(�͑�7[��oSr�`��M:�����%��M�A���⮳��l�Z�t�  �w���XZ����_I�M��g���CE��'�!�1�5�=ޢP����}2��*x])����r�t�Չ��ݘ��=ܨ�d�`���3���&��K!�J%_�xN�0mɿ�k\ւ��w�*E�1!���ėC6�gD�%Z��U��k���wMӐ�or��II�Ջ�J$�%�ո�329����漨r_A�V�רcd�t*޾yjC=)�G2�G��g�Ӏ|:.�z.�:n�/t=[����v&Z�復�����ț��<�w��'6�+�5��,��w(���43Q1��=��v�;K�7��#s�� �}�ގ�>H�79P���V���,y���=�%���R�Eh�т�(��RZ'��Rr����\��0�A.�y3���7���Q�MQ]�H��2����g���Շڎr�b����<���P��{䴆R�f��h[��;�ޅ$^Ц�=�0����D�tx��1�(T�w�2j����,V	�!�h'7�C{�jgQ=���*��^!���a�Oo����]�S���'7���Ǣ�[ԃ2�D�:� �
g�!�,�8�Z�J� Ŋ�dU�f�l�z>�NU��$�&�=U?�D�t�8|6'c�Y�"��72p$�������mP(a! ��Ef��jq,�w��Xy�Y��ބM�,�+�.�����y�=�kiEn� �)��o�e�o&��?��.}����뙬	�X��z�%�x� &�"k�7A{�am.�_�Χ�1k�{&uK����)��w��G�~�KJ� 2�[���{�ԃ�K��<ϘwL¤k��-Xܧ�0�eJ�lr8P%�_�6茺����bIa��-�IT�e�6T�ZOfuyFAw���ⅲ,&0�k��[�v��z�ef!W/ꀪ8ܝZ��=�|���d������1��;�77���޷�+_]VX�l9���^�zcKj�������D#�I��g�6���%��e�ߪI��Xȱ���+4���7�?���+TO\nbn�>� I��|�*�wUtU���P�{�W�b�jY�!e!�o6��2c��ǻ8��G��[��x3�op���2.�����d�%�>���#�Z�/rH�LY#_]G�q���|w�[�i������
9G-�q�	�]r�U��:��G'$��{4��UvE\Y��| У@�](�o������k��̝'"�����x�'�"����G/�C,��.7��ܻHԤ�:�>bU
:��cQh|]0�䂝� c��xP�3�a*�Ț%a^�^"�-D���[S�<��9X����,��:@�Jh�	���x�������E��ױ�"���9�e���A����3������cuU�*1WB}�"����F��k�o$PS`:�o]n�e���ۉL�0��C�V�b�#���;&"6�Q�J�Q\s�}��؄إ �^u2>o�!��e��~�`�Ia�`m$k�;s|�t�&�V*g_+P �\���j��!�����1��W`1~�ycR�h枘O�L-�c��fb��6.M�R-�ez4�� ���ok�ӊ]ߡy�g���U��d@K���#��>=����'�!����vP5=A�-R�]����ұ��C��O)���c*>��7p��K���2�ƍ�4����%f��o��ik/	K�׊��� �R-^��Fp�t|
�pE����վ ����]�u����>�y����4����%��9s�X<<"�ϡ��]y�l�ߎɩf5�
��i����)m�;�1�-pG��I��ݯke�30.d��Z����N �@H�L8���ko�����H��|���j��F���&.=������P�o�n�ů'��x��uz��{a�ۮ�o�v��k��2��4oK��=���˃�36�6	�㞲�9��S�����z�}A��ƙ�+H s���s�7X3�`ħ�u�\��3�z8��ײE��	�Dj���w�TV��\�:DCᶲ�4 .��j( �#���7�V��Ǩ�%�WM�ȃ�xf�^@�*�+�������L��=����Q �9�+�Z.�o5->~���bP���N_i0lr1S�O��@���l,���4�iA�n[�����)7��32��B
d�⢏+�o���t�|��M���+��T�F� څ�~0�?#�!a��p[4�����%Ӏ"�-�/�QD��8��Y!��܈:!�t�6��rR���n;�W}#�mZG#ŷ'��Gv~ǂ�Tяa]�c�8uFh[>���cYX�
��y�_���f�0�_�`=Ŋ���'hY�%�dPz�\�b�F,VS&W \�$�� ��a��뀧�"&�B��?���よI��х�K�y\D󏢵���Ը~���K?{O�^�����2��7��D˯��Z����B���n54;���h�,� �q��#f��/2�**�ѲM��0J��t5�G�6�����y��I�$He5
�j"dC�	�r����ڱ�N�j+�u��~�bk��hY��g�ĖO����FZ*�yuF��K�ò��<.��D��@eW17J�g�z��Ǳ�	n��b(I�2!s��z���[�~a�޾"�Y�sTz���U�˷����1)cg%��3���-K�k�H+�"���>�cF6*t��[|	��CIo�^����>���JC����bq��i�t*��U)���xSJ��N�k���5��_F�R���G��W��С�����O]n��eo'x#B/�+��P��[�?=mq9�4qO�;'AHP��Ȅ
-]U���r)�fͺ�:�뗯Zd��_�,h�3��%3E}]��G"<k&j�����a\�#(�\qq[���?��T��w�X�ؓ�w�����P狃)�lU����q9EXJ�k���`�8�/��T@�@r��� b뮜��Lk���ؗ�yVyk_�l9��9p���0�i�b�t�;�Q�|-e�lPh�]j�ku���%���x}��o^&)��M^�`�E��9�ve7�$Vͺ���8�� Q��U��C��6�L�w��r�pu&9VJLj������Ǆ8��$�����oBqpB��(�bUg��g�0��=3)������R+[�ѰF��wdս|zf��*<��NK^9����ӵݻ�>��ܭ��"G��:V徭��q����W�/t���#'P��4ޒBY�	,�N�����>-�+��Hi�?�Fwx�0�C��$˄^�Wm��K��W�ݱ��_0���
Ȧ��(���tU�G�U�{1W��M@��Q�5ù�k���<)�W��7��M�L{6D�L$1+�s�l4���,v�'�����XX� �!�b���y:ӫ�+�/�=Fh�z~�8�AIE	�]�@[CE�*�����!{�+���
���#<�[1R Q=�C�������Ն��R�}Hv���,ʵ2���;@���z�voR�^)����@BnΜ۫?��f�N�9�����g�l��RB-�O}�$�y��ݮV���3�V����N��O������5�=+[  q}��Dw���t�l�ja���#������bYG7�!d��^�OJ���.�Mt_A��Ӎ�%��o�}�&2��`zG1fu�r����?�6�~7�`����J�5^��_�6�||�^��O�i���\���x˚��{����몫�EtV_�iܘ�kQ[�(>������I~.6�f�jG@1^���x��2>,c:�B�~�S�B��j��w�u	��������6t��4F�I�xU	�r�ؚ�h�)���@�jPoC{��>Ϻo�wy����mJ�-��]����%<�OOn��:�g�������+wFDm���+�2ŗ��`�I���bF�"�
��������,��,��4��m�������~sw��
��= ���u�Ӏ�Z����T}mM�HC[�[C�dTb>WI�r�g}��QH��o��Xw�@��!],m_%%4!��S
|�|r��l����L�����b,/������GP.~�ʛ��s�BՖl�-^EW�ǿ^u"c$yK�z�:�6Ҩ�����o�TA�A�^�6%<��#�ݿ,`!�쵯���.��o��AP������E��iˌ�.
��k�4��j�������b�dEH�.=X��]!~�I�hze��&���+ɾ��� M�l�ײ��#;���Ժ�����?����Xn���];�ZV����%������dS��F�L9�zx�У��&;�,e;�EV���x=IZeE�`��S"�U��%�̝��Ǎ9D V��]�zZp�XE<�9]��t���g�C���a�?��ωO�&�8傳�-����L�>�B��+��N^������1f'�����~0}���䡤����mۑ�����q^H�ʣ�J��ݑ[�'�5�o����
mt�|(U��[��{j���bRz�ˎ�Q�|y�������=q\78~}FP���~����������}�Nc�͛ŧ�$T�_�h�������f�;������M�����3�������!]��ˊ䚫��(p����Kv�U���b���BW�qA\P���ϛwt�FX�}�f�]�	PT�/�@�!��A'بǆQ�*8	��H�#"5`�fm�Hp1�Ռfd�����ɡ��Y���Xe������P��]�e���x�;:�S��L�m�f��J�Pݩ֦���Ĥ��T#Xs��W�=�S,.+���Oû4�~̳�W;�R�@���	����ֱglcq,9���L)��`�bg��-*����_���h��a��H 13��xƫ }�ډ×Q�'P����-�S(�	ɞ��wʁ�{�{��^�k/T�w�|��}�����q����f(L��pR����g �a�R2H8��D�vI���ZqFdU>���c�Q��ߦ�O�A���G9@��;9a5e<ʿu�L�X<���+X	<���Eu��|�>_V�3���%} ��F-5���e� �i3Vgz#����؟�v��-�@���Js!�e��~�i$��
���ڎ?�~�6_YM"���&� Ǧq�w󑘌31p���H�/QT�5�06Z��N<Q�!�
�i�����:l%��#�]�@^o5NxV>n�wi�	KuF�:E�~��^D���Dg��܉N��d�)��'~�hږG]����+#�3[ͯ��Hp_����1�G��iA22�w�%<��W�r�:��M���2x)�A)���!�Q��S�O���:=<7��/��ʿ~*�e[��z� =;uW	�E��L�E�_sk�36��ɧ�9����%TWMK��EM���������{b�c��/������xE 3[l ��e�+(W�"�k��k���s�{wP��`�跱�M-��᧳��@���*���T���Ҳ1ؾ4�b���kD���\6FF�Z���~P����>��ӲT���S�Åu�W2첿7~��8���[.�OB�/���h����0شj�?����D�]������#�4��@l��#�a{2���ӑ�Ou��B�6Q*S�V�T���3�'��k��KD'a���<�����,^?�/]�Wy� �ݡ�K?g�+���(
iX�����B�C�Z?���ޅ�˨p������s�~�����K�>wOf�W�NL���?>=�	7� ?���������� �o�]ˆ�~+�ѯ���>���� [������>�6�#9�K� �ۣ��e\H�4�H�>uw�ȶȹK�m3I�K>*�W�gj}�V����5�c�ATe!��$��:�B/�]D����2%Ծ��Ww���J��?��j�һ�U�͙Ȣ٧qE��Z�p�ћ����Z��xq�|p�}ڜ��˔�d�{0v�ƅaE���Q��3�	glK~�3��E�Q�c���7�s>�P��[��[.�:s�D���6��l #���BM߼���t��W �[R����}��I}@���@�Yb��?D��/��Lt�q4��y�ȳ
�x�f�K��xT�u��3��q� �R�~��V�łY<���÷���O��6=� {(h�ݩ�+�'�^��?+�Qv<��f�Du���aгv^�+u��eI%���Ĩ�
?�Ku+�\���
����Ԃ�{�F|���/P"4~��"v�o�(Vf"�C/�#E�Ɓv�_Ȉa�_��� ,�3���l�1��������M�jM�L�8k�u����{��:y9��,gz��X�� R:�ۋ~'�;_�;j[�li2�Z��R��u�pH�׃��8	y���_MԮ����
Bar�D��Rod��ޭ�j�S��V�د�r�[�|��H�v����!(�����Qܹ�1�y�v2���j�y�w�`�sP���ā��!�a��7Mq*�p���w/o��,i�:��F�3�*��N	�Enk@�J�<Pb8.�ꙇy�(������ͨQ�i-��-G�UǼ�+�^��������?U�A������@��H:� 
�;�@Uh%;�:��&"H+�ٛ~y����3��]_�͢Ѻj��X�S�j^���y�V7��y�x@n�Q�- ����'�
���U���������|?$$�	�u3�*�]P ��w	�����=Y{���	�b�[��<;�lE�6;�.##EP;�����:���G�sxm��o�G]�!�v���Gq��u&o����z_�s��?��L�Swig}�� �G�x܉�u���>����%=k!�Ҷ��r�LZh|�W7�_�-$�ܫk����@ѣ����aG}���ƪ]��kP/����_/I���B��2���B�I��v�ܟ|�P|��z�a��U������Z�ܿ�rYݻ6��G���yl�)�lq�K�hl�R���|����	���v��&�ӷ�\�B,�3r���ے)f�6葾Bk`^�}���LEZ5���gf�Ԕ2]�����9k|XY�K1Q�V�be��f�L9������ψ�cn]ղ��5JY�=o��{�"uW4�l:<�)����JJ������w�U��R�1��I������_�7y�L����c`]��&x�h���Bh�<- r�m��	_Y��"��~v���b�xN&n�.a��\ɓ)���c��%��7ǣ�b)�t/�,0iuM���p���|��#�	0$e��T�b�<�-G;7�I�aAi5�׉��UT͵<m�u����)��3(��C�O�n���ߗ)e�5)Z��-p*�o�X2r�ّ����ұ���_���s�_߽����W'���[�+�ۃ�q'I�'�*!6f!A.��"i�W�^PT��1q��u�-r{�P������!v�@/���,Q�������[�;����t��?��@TZ�*��C�hs�5.���&VQ�J�� ք��jk�n�r^�iSw�����@��Aٖw���<tu�&�F��eU.D��.	;��_�����;��'4;3�J�_���_#TtC��s����5�_�jl��-F�؈OIO�Sw܄屆�(�S����u���z�/4�ͻ�k���6��7�� 0�0{i0�{E��egr�k�@vOG���N���Y�hg��V�����:d����'9#�*1��i�/����>Ფ�:��9%Js+�(��i���"m��Gׂ^Z�k��+h^�;�`0
5�N����+�")�&��R�'on��h���A��^f��D�@>a�����s���|�ξ�[.YZ���)`�!�֤�G\��^�uH�NU3b�v��x:�' �@��D��ae؞0�$�¹���ؤ�$�X8A���F�J��9U�=��0tU�e�e<�t����x2����oa~�,+��:��*T�_֞�ַ-�ft$%��t[()�kW�w����	Y��9�dl-�< �05��9��X��֘1��)��-�Ǉ&#���b�g�6�BS(S�udz50D�C���ȵ�����f�iC��Jdp�w�J� S[��kG��g�A�_����v���eй��Ӭ�(��[-��-B�z��^�U�,΄��V��k�"��6��4���wľ[Z�h.�R��z��K��b0��߉gE�֮]���X��,2WwKi=Wncz�?]�����X$��������sz���S�0����M�)��^K�7�Ia_���C>-�
6*�{�^2�6��X�:m�:m�l=����=Κ�0y�);�%��'��i��?����Y���>iф�勁�4*�-�Zv����s;�4xr�� {��DJw �vڝ��#.i6�}���?,۬�G�[�iG$1.�$'f<��P`ty&"��3������I>Za�I�~�3���b����f�#aQ���+���ڇITW.��_��W�3�B��mѸ�S
?R�͹���H]�������P_}w۟�>꿰�����ŷطC���N���vW��Y�����M��/s�j�;��Q`�e\D��T�K�۹3�݅� ��b��?+�xo�2�)�1��U��;T�ϗl�0J�T��E���|�Q:�3!�~�qc���D>(��q��S.5cs���c�,�{bqa��z�Y��]����R���3�Z��k9�ê�b��fv+��<̣�yɸD���4j̶�!��9�`��A!Ƀ) �R<x�P1����1���錟uP����Ԡ���2F�<�+���|��h�r��!VPW:�~7�y�/=u�P���\7��<q�29�k����i \5R2[��ۦ=H���Dr��� &��Pɩ�O#]�
m5�`�=E�[�	o��KrK�������t�N1�,F��"�.m6��R�K��,�
vT�5Q���ư��ǥ2t
����h������>Vh��+��7qg�QA�[�wl�g�>����ߍ�=
~6FM��_���>#Q\�����ؑ�)cnK�F�Z���P�ͬ�3��|fe-�4�W�� ��8���䠝�!�[�΀]��gt0LJ�܇�H�fD��������f�����@��ƕ����w�s���e�[7�;�r�ӝ��u��7�m���.\tn�.l�^��m�~�"��&��Y��h��$���4���Hn�E�� ��u�ȫEfu�e�2���d^9��:���#�ωhVw�Ci�8me��t�	��R���:ӧVl��*@�y���GP6��[�U ���*�u�,n�u��<Ln����`���Hc�dQ(�J:�č�T�BYX�]^����UYH�\tni�����/	���,�w����9���|!jkt���2���|����'���+c�v��y^b#�8,C���g�����qx��kx��Q�"��d�"�|�&�	þ��Au�k/��ַ��Z^����ߴ(��m��Ky�w���w�:�m/S<�0z��I�(�|�g���C�B����H��yØU��k�@*�\'��M0�k~��}G��K�t��-O�G���ξ{�Ut�ǭ�_i@%9cc���D�6��ʯ�t��0��KJ�2�:�(*7�ji7j�	2�g��rTkF@�����D�@�w��q ����4Q��*��)I�m���	�3�*�Ė���������F^|^r�bf��Ȫ������
�܏H�&�������B٭���*����/n�TF�`rW�݊-k��n��6��3�D������S�f�?��D�U�*��]e嶔��q��"L3-$\��:0�7`߹[�^�
b�[z���Ѭ�d��s�o��s�8(?�\�~Md"8���v�y�cw����uFv�:6��?}��C��!��#P�����e����8+D��z��0�.��F�gI�>f4�ˮ��I��/C�;y��9�5}q�����<��M3�B`C���ɓ�jڣ��c#�?e��&5/<'�G>�Л\�鿼�<Lw'F�N�k���9�n|�Jٛ7*{Wq'��0ӽ�w�J�֥�r�ӀA��$
�0.2���E��Z)�K����b�F��׹
Ꚉ;��?DR��/����Lp���P��_M4^kM��T�J���:�B�~ؗ�|ם� (&][{��O8V0h��ddY�xE�	ͷ6s}��%�J$��(���X�ܽ���ʜ�LYt�����"8��
���m�i�e�T���j)��C���so99�}o��oI�m�����=�������� 6/hcZ%EХ˂t�E7�z�h��#n=�a�}P]j��!�4�]t�3�����[�؞�D���u�W:0�KNV/���6M�<,y�S*�yNxHC!j�F*�S�q�O��[B<�y�<"Q��H�B<-k�𔘅���Է���D��2"� ��ݸas�~�	�t��2��UD��]vD$����L��Ӗh�ቩ,�K%A�q�KՐ�,v���f���7�ATv��]�.?
2���؇XǱ딒e���	%3Qa5Y�sUN��E��x*�������a]&��
�Rk�V���8���;��>��?�p$��I��u_�a�O��.���Jl^��k�eA���~�
%���>l�G��R�y�������`�7��7�ĉ��w��P�LJ�e�7 
Ъ©���L{���v*yRǺ��PO�ڕE�4�H��"����k�k}M#4G�V�r�v;k��\���)����qrM��?�j7$p���u��ەKT[��i}���z�),�����Tc<�����v�n?�΁0\�ǱE�}Yajn�8�Z��$e	�����2o;���c�w�|� a4>��q�*�e��;�oB�N�]�(,[S�Y�¿�%^�����y��r���	!N�A/��M�R־u�l2��35ئ�NX3��7�R�/"�8B5%�W���w��;em�H���v����Nk%�.�RJ�Br��^�mZ�F��\|S��(v��&�d?��ٲ���)`b$j�T	i������.��ł:��.��l���W��"���Cr�)� �����?�<����y���A-����nDH�c`.m2���:�5��U�{�jE��mx����G�˖f�EbkS�]E���f�;_�[�V/K�}���dj�~�v��Q�J�n��J�[/q�m���]�����*N��cs�`Tlns��m��L=�2�
�ܬl�7[qB*��e�kyS.���^���iA�(��@Dyd��jzDd�n��AA0�`ܮ���Gm�_ڡ���?i2��O���m?����Wųh���|�c!�&����Xt�����e�tla�(U<��gG(��\T�y=�v���O\�5�~I�W]E��S]���ߋu�J�y�O�2L%�jگ����F~d� �U/����1�0���Q#�6�T�΅,;�>��0��ؠ���[B��Oi�I�I�a��y�_�\}P�����C�f_	�1�pg�5�ҋ<�Cu1�uJ��X�v҈���ָ~�ӿ���X��6PU��ꟷڶu����Z=�(֊Ǚ��:�E�T4Y̧KgȤ�&��6��Cn�����0�PU�g*���@���O*%�y��
�i,̉b%�I;�_�����8 ����lQE]rm�G���)��(�>��=:g��#hV�)��A�t_|��Դ��!Q{m�{��W���,NK�u�p+�Q �� �;9���5��a��ա�Kt6RNU@ � '�NJ�i]:���&��W%��X76Ĥ�t�m��%����{MS~7��բJN�l��{t��E���~���Z�)�����ɞ��9nOx�<�����=w}c�Z��{�K����{
�����A�nO��P�A7Mמ
�W���;��x��kl�<"[�`�ҕ7�}�k�G�ǡ�x}bD�D�c�q�t❜h2JUE���'��V�{��X�o�� �P�E�51(cF���)�����Z�6�>ǲ��yj������!�{=foZ3f��� Q���Z))�)�>����.^M��3�*�TZݼ�����N�}>�z���E��t����� ���.��@�|�~ ���K��&�
�3���d�|7zj�V�
uz�����\�~��߶o��9�}��{.H�:�9fօ��Y9�HB�E��ү��f�vg�`h��#9wi[i���'w�z3�ל��ޠ�;�0��ktnc�88�ph.�ѭAkb`N�����d��H�
��jy��ފ����=�-�~b�ʟ��
��X��^�.+j?e�*A����͡MA ��5	��s�.��}b8�B8N�Uq���c�C�6��T�����O2���k
�x��;#�!����)���J�!����en�9Pm���7v�0muh/�K�0ő��A�C�K)E(�����/l_*�<i��,1�6r�L�}~�^w:��nX�ȟ+���tsu��L��� ��R(֝�����!?��P"Xozc�@��1�Ĳõ�L=��r�(�]?�����0�}�eBg���G��oHLp-�
���cW���Op�)
����ӿ��[�2�\	��E'h��p
Ç�_�T��n[uD��|��F��:�= 
h{��"��N�۹6�;�3���}ҾO|LP'F_�狓���;�7�l����s[�>~|�����1υ��m�H�>;X��{�*���Ձ<������"w8�ZH#<ˈe��3�����0�L�ൺf݀��ڵ���޿
�S�'�A��H�8r�j�ڨߣq����ļg8�%K�o�{��P��X�5��U�J���>%
��]������v>`a� ;Z��[w{:-����p�`\��K�F��X��'�c���8��qx�2e���UK��_�j��rjS!�i�iu����M�u�&.�Y)����1�����3�㆗Ѥ�<V�[f*��W�N��i�'[z+�]6l�/\�s��M��~�b�_Û#�>��/�-�*�]��L��Dˆ���v]��8D��l��߹���,�
�t�vo9QS�P�T{G������ۇ�s]:�� �Gv(��ւa�"�[$N��� W����ŐIO�,w��xr��X�ŋ�\�ܧ�x�Qw��B�i@�Pe�I�܎���>��mz����6��Lqm.��s�E������ai�z�F��Wr�a]�e]�O|������?�(Y2��m�|H��X�Hj`�q�݋����O�K��p��ǊlPK5����"L��G;->�[���N�L�y5����c���2����l���DY�������� hU�HU�
���f�Z�S����Z�
��p�O�����&�M�f�[ht;\D�^�H���b)��ö֖�Ν��B����l9�D	���f��N�t�(��ew����դ}��3%�������9�������a0+l���w��"M�^���HR���go�b���c:�@Ω%��A��� �ۑ�S[V%��!��4����5k�z��#�m?�Oz��|�E ���wqZ�h6��Z�q�����p�&��yʋ��(�!�4<�Cw(G�U1�b�s�|͢oĲ�Q��f�+���jR,'�������Q���;����9W�["�7v}���~x�>�9�(x*<��<x$6��t٣w���Cp�����s� P-=��ؚ2��b��kk��=�:���?�sJk�6���G�ݳ���d�M��g�j�ۼz�jLf�߃��E!.?��fG��'���r����1d:[�]J����Z����TwB�fΥ����W�)��K��$�Q��*@[H7m��VE2�]ZJ�HY���Ȫ���M\%c7�Jo%q;�:�Ry]�ot;Ӹ	#�DE��U��p���L]XP�sh��7^Kph��]�l����.���P@�0TL>��'��H�{��g��r��&�jj�
m�0���0O֐ȫ���K����������ˉ��˥�Ϸ~�!x���%�������.�ܕ�+�{�r��<n���od���r7an�}�Æ\�\��J��B�5��urK3׹�!�RJ��{,ג{R�-�z������׶��<�s���x��貃����������K3��@���'�#�E*�+j
�]����S��L ��wm`���0�U�
7����E
X�sمs��۸��Ht��������\�s B���3pq�{l.�;�@4��myn�p��Qĳ�x�����c�{(EΕME�����z��/�T5�k,�̺)�;��A���ydY �L�mI��&[{+��$T.��W��_W�f�Uv1�<���o�Ϟ\̈�\}�SJ���o9����g�sb��wk�1~_�)���g-F^�%i�.IۮP�>j��6'�2W��u�Y��F�{�(V�l�f�dW��o�lq�D�mI����fFE*����۽'smqE��I�JԊ������r�')ݞ���������y;�l�e1�9!]���jw�E����O*c���ÿX�el̮�a�5��mN�/�x���Y�0�l��a��30�oB<I~��$���������Q�`���(_0�O>�Pz�)GM��󃫇��Ön|g��}C�5a��_�=����"���ʨ��&�7�Jq1�O�+�U�NU�da�lJy�ݭ]`tEf��>Ӹ��l����>����F����S⻌&��q��' ��o�YS�D��"�h3��v�<T)@f�P>�lCF~�?1�}ms�C5r<����#ݳ�����]��(�WO��,�W��`4}d����Y��au�!����ᯤ�*]�R�F!�Ľ�����I��]q|�DQS_J���ڣ��������sL�.�Mˎ
���5�W�A�Q;]M'~�;�8�k��~l��y,iC�}Z��\4g�>��1�;��e<J�6[�:Z[U�u���H錱�Z���A��a���3Y1��.o�����Oo��=���x����P\�ѫ�a�v�m�������]M��ݟ"��z�^C��~z�O��<�CZ5�rkZj���?��K���<yڹ�[��jw����O���tL�.�aQMԓ ����>�s����E��|� ����us�oS�������L��	��؁�����f�X���E�	�^�{�m���.z^E��`q-�D�z6��!���҄`ǜ3�����_�x{�����˔��&���\j?��~���XC��F��^&�^�URY�:��P�������CbH�Z�!h>u���:"��\�����I���э>?y4�_��U�8+�]�z��aK�an����*����EZv�.��5p���@@���)�(k��[�߯�4I�ƾr�'A�@W�8�V?���I��DN?"���>**�~���w���J�t]`>�E8�]0�Y8��|i"pA�1��`�#]����k
����s:9��>k��e�^�;������y�?+^/꘣?�=����k(N�Ȧz��Y=���<r�J��{�j)�=�7LU����\�Ye��9��٘��FX��P©;�Y!��f�|4B�t�誀�n"��y���-��z��5Vr��etF6�T�mg+�7���H�e��f���c(.I�<D[s.m�<{�J\��"2ץF��誆\����.�#o��U�e�QhK�ơ�wf\�mQ����� ��%�>F�LK䆡p�m�?�wg+E�Q>%��A]��E�D��P�<�V�s��B�<��㈝,�����?x2q�QO-H���^�����)oޛH��b'�c}3��xՠ\����X�*����_.ӕ;�������.5�-q�-sM���b�b�����W��=���!�c�S����FH�������V��z��<-z�7�����[��ɝ�P��+p>����S?����	��⛗x%��I��EP�
���K�6��'��ɸ����XH�E��(��������������#�O�in�3��0�jy�'�,�Ҭ׽⤧����&�_yX'W5_��Xs]q ��R�xf�����M�A�vf���\�򇣭[;�I=]��OKZW��F�˖DFK���fW#'�)�f�����p �R�m���Ki	�6��N���(R���#��>��t��r	i���f�΃�Ug��s��?�tT)����?��sy�3�φo&M�o�X�YM׿�y��}q��X���#���9p~���y�GM���1�<�[.>�;-��K��h�l&\H]�����o2f�e��I�CO�!B'ke7q�@�2���鑖���ۛ���̀D�rf�\��'�U�al ���@bp����TL���v��l�>Mt���ŝ��[u�Pw��J�-Ԗ�PQ���g"��]���<!o6�h�\��8��H���@�t2;��M�H���D&�)�l��a�����\���nz�ō?ŵ:2���Z��'�E$O,������xv�6k"m�օ��:F��b�B_8C�}⏄��"�n����F��(��T�#����e�*�_�- Es���/d��t� ��(~�@H���s�����l��Ac�cT�`"0�b\��aq�b���K�Z��}ܒQ�^\]r1���o�� v.1ƺ|�ؐK;7V�/��R��4�.�T��7������T��d�QA�����\��eQ���s(����U�/1T��D��Z���s�۳dYT��4�(�DE�c��.�̝w���������1Og�gG ��W��"E*P�F�L¸�mӱhߖ����k�	��	|�cV�B�ȳ�&d����-?��b�bѤk�ql\���1�M2�]���BE�M���&�v��V$lW��`Fa<Z�F+�Gf�*р�1�q'���8-;��f�͔"��䉫'p�$ERR��
�L�tGqV\�-9c�=�U37/v2���w{�=�����)��᳍�o������Q&(K�_��3�2��Y��n��H��pL��r�CKg!һ��{9Tw�rj����>�|�GH�I����o����np�p�U �dm�����5�Jli�����@����媤aiy�+���m�Q��5�G'�eA�iǠN�79�~�'��p""���;,�6{[�����=Ќ�.�[7P��-�F�5�ˆ�1pT�H��� ��	\o�V��~�T�Q�a ���P�#eIZI�� <���>8x�OJ5P��@�H8UZKܠǋF��a3��+?�=�/Ķ<s{#x���) >i�`ܥ�s��i�$D�I޾'��D�Dq��e �@@���h��-��Y��ٿX[�vt�'�����[����5D��=������C���8�%�c�J�)N���v�Dj��:H�LGF�.r���1��bW>5#��B5���6�;�ע54)ek�̍9)<����
��y��P0~ E*3�M���d�8���f���i�Ƙb%�|��ϟޙ�;5�D��҆���Of��_07Ȯ���sҺ3�tX�����̐|�O�I$�Z~[ph^��l���W��������e���p�U�eb��)��~��RMiR�p�nJ��n����1#J�~<s3��d&`L5�USHKbL��?�>f��X���X��"F�'��5ud��k�D}d��Ǻ�������3�qU���vU��"��Ydb���ū����]���>��(����ȁ{h?G��K;D��>���PF<�r��YRC���wr��������ي���@���.�fO�J����9d�Ʃ��$��7u�)���z�`�33��]BFd�ŗT����MN�Ni�K��e��G-���Z紁&.�<��]7M�->���A�\��zQ��Z�Ha����n���A��͌g�ҍ���<�rs��'4\݈��{=�?��t���hٝ<�N�aq�����4F>�a�%�oU&}��/�\轆da?�G���QE� �a�7S��f'�Bɇ,p`:�<�P�&��C���8��{���ݻݓ~��F�^�:�N��f�h��~K�.��^T6B���ͱ����*~甶��x��:������n��N�a>R�:�c^���טJr��)ev���
�Q�W:�g�CzRS�
�o^�C�����ÁCl���ik���m��_�I����&���B��b �Jh'r
��ۈ]U^4jK�+���̉ZM�t7c�In��S�b�ؔ ^$��Sq���_���@�)@�o���C����M��ߤJ�Ϯ���1#z��P3Y�홹�&2�^�u�xt\�����:2Z�k�k|J���y��L�n�R��'7E�^g�4#����-w�*C�]�:����%��I[ky�C��(DS�>=]ߍX��eaS6i���U�Ϳ���0���!R�7:�h�}ԟ�H��t��Ȧ�p�����Rg/��J�p�����l�-����o���w߷���%���*�1<��C�6)S�@�2�^ǖC��.���S=����ǴR�i��7<�	@����(���;�E��fnk^}$ȍO����	�3����'+L��W/u��4�3������XLn"�?� g.����c���OT�TDG�~�A����`/ȇ���dk��g�c�dn��1����/�0���p�i�o��N~�s��Ň��Y�F��cH�)4���?t ���ז�tQ�(��G���3�6x,��oH��`Y��
-Dǖ˞%B^S,�����_�:���`��� ��
�}a��Ӕ:�@S"[\��8_�<��K_�4^���q/����aZۏyW5���Ct��G�CN�/z(��`�LDl֦9�;ݚ�E��'�rKa��H��:݁
|�Uh���)��g��>1~��J9�|������1��&��}{O��ѕ{��1
3��%���\�]�x�!�y�$6���)�u�)�>3X�&��n�`���?�qH�᷼yR2�5�g�SeZ{��_�$�/�I��)��
�����v\�^
�E4���f�K�Nf�&�ǒ��s�ⷠ:�&tKYt������w��.����d�)-b��-F^�����;c�����;כ����"�C�"h&f'�f����]d����s�����÷ˠ�&k�؈�� ��jszc/m\8ƃus�)o�\�o�6ܟ�jo�/���{�U��e��ub�O�J)�f�UIҽTm�e�����`g2�aSr������{f��IO��b��[�O?��
.����dfO��/H�S���|�O��W�z5,?�DLG�����u,H���[+cY�D2���&Fvc]��F��x��HD ��0��
n�\@��4��Е�=��Y!�:�TY^t�s���܈�x�n���,1:R�盳�(����DZ�BI�˒����diD?�u�39��7�gwG�vIO��~������$�m}�~��A#��\�e�􇭘���N��E�'��'�" �_��Q��䞗��2�ֈ7ŝ� >�y��0-��l7"��5�Hϰ��P`״i,Ye�j��l���)���"�>����8�3<��}�vJP����FF�j.��;F6gĭ�_ʈIJH�
��bd5w�X\�^��s���d�K��qoL��^�\���Ι%�}�c�"��y���ER�S�L�7z��I���h^�T���C0s���Ms�ts$�������T��2P��tˋ�a�q����鱳�M�O6�v�����$�*� O���]����P\�O�D��o�6}��q=���f=����U|ޮ	_S�ߦ4�%��m��f�^��n|��U�c��.K�cw[���~�N�h�m7@��٨�J  ����|�i��j15A1i?�ELp���;J�;���~��^m��6V�;l�����q���R����W&�
n�F�����Un�U�?+�/ΒI�&��s�m1׻-#���͏��Z"R���/��c�Hp�2�O���j$��
�/�px�W�Q�ڶ옎��%��}�u��^�?�Y��+P�S���\��`\�*����w�){:���C�ꂊ�D���$��+����	���4�o�+9Hn)x�T���z�@)�1�M� )Us�b"��,�@k���:l�-���0Ǹ�I��z���K��d(H%��?o�����G�[#�D��7�e��z�,Ċ����-�7`8;��L��ʲA��ƨI �u��=��fƐ��a�^��O[<Ŕ�)�8V��C�s���Р���
�S�-R�sw��>rc�x�����(-ig,����͍�d�m�	�ВB9Ab�W82B|N{�(��A2�}z�ʳ����%� ;�o{σ/���8A�U�æ���F]叁����T���z�]��"�Н��1y��^���k/�@����ȹ�;�	)^GpkTpI�� zb�L�@=��
��L	o��ɖ��bݮI���9��I6��I���R��oE�S}���&k�����]�@9��;�Y.�:cm�Z�Ph�?c���V�o���u��~��f�NL��Z,�c;�Ʌ��oE�7�����2m��^��_���:{��V�u�)���a�nɹ��ֲ��ӘY���}(K��P���|���:BZ(���M}�j#%�.@p�{~dO�E��Շ���;���PA318�wz������̷`v]Q�8�����"�(��n�'��q0�1>�5���P�����uS���Tw���.����2�h�T�q~��u�X���S�o����O��(KVf@W�7Wo��l��K�t�O)��J6��,
^i�s���S��aU:Sf4��Bx��U�V?=��X��~���iϫ�Հ���]8�N�18�rG8{�0�[�����C�7OH;��;������ih("?�s|0~2(��*�/ իmX���$�3,�J;C�R�x�O�u��q����yhq���m�0ͱ�w���
�J�1��$?u�1M��Ÿ������e=�I�ߺ[,�}h"�0bSo�a���Ƒ�n"�yVD |+#��U4`]����J��ߌ��Q���9��v =䎖���ʬ|��a=1�w�+�_��{4CÉb�+��\W��e��.�MQG�0|�EW8�Tf���`嚣ս�Ǳ�e���zA�n������*�5��	���چ��3�A_���t_�faG�Ab�g�1��	9-�r�V�Q���]���#tT8;p�sӼҢ#.��#�ޫ@(_��&/��nx�`��Sa��D�T����*�ϪzD�l����t�F.�?�Ο�Y%$�B���Y����o��#�y4�M�rrN��G޵O/�쐣~/#�E��g7�,�ܒs/n��_ˇ�b�e�������W��N��-�9+I<�g�<^�K]r������x����]g�b'zٞ~&W}���yi(^�v�W�)q�0��0��Z�XlX~�l��7h΍#� �~�!%PX~K�������A�%�$~�x�`��I��Σq�:ܟ��_r���1eͿ�➹%��H�m��(*�C�ykp;qo��UF/Jl6�cq�<�[0L���$!IdO����K�5�%�Z1���`0�kR�i���@�b�%A��Fg����rf���t�u�Ϛ4	�O���A/Z�	יO��WID�.�����f��%S^�؅���G�Z{����&�`�>�n>��0���e�jCk��S2Oc�9��w�E뷯އx���L������3����6��_^�_f������l�������}�os��o���}���~���/	��UN������T��=`[Wot�����Nh[�5�xkq������N�[�yǅLb(��(i�V�R`Ql�JD�N;[��ϖW��D\��v��K c���R����M3d�Aa��.";�����.�j~+o{������A���W���v�C!7��o?Pun�I�{.NPB�:����x�{���z�bl�hH"!���W54.�)e�(C� �����ћ:B��*Dm��+�8m�hǈ���c�v��s�����`�e6.L�8���������Ӕ`��m `{�t��KeN�V���҂�b��;�����*���9�h��.W�sǊ#�݊kͮ�q�d���LMT�|@��`�����&�a�*CJ~,w�.δ���Òxw�N�<�m�tME�:�F�%Q��:Ơ�n���~)���T㴼8�|$�B�8!�V�ХDٵJ����0h>İ1�G�Z���ǅ�(K����'Ak��O��B"9�W��a��P���F����p�K�p� ����0����d¾~��kt��FK3�N�p�X\�u�>�����%jgD�����7�tvڮSZFI�տ���ɷ�Qr��1`Z�]����<�:m�
�.����UB���K��R��C�a	�3�+�X1Z�Ѻ�3h���5;�U-��{/V8�$��4���iuŭ�&Vrĳ�n����i@�Q���UC��Te���䧴����&~I�+��y5�HU��<��>�$<�����xt>����Q�7�O���i(���c�F����/ﱯݛ�����^Gu�?�l��V�V����;;�_�b")<}��\m�蛵�Z ���z�m�	w/�L!���.�P�F;U	�3�h�i���x ,P�GE��l�e䦞��� ���M,�o �)�h ��@�Ww��b�g���%I2��uZd(���W�� 
z���w{�H3��bPu+i�Xo�7��cAeʾqkZNfw�u]�{\!��mj\Μ������.�
)��ܞQ_����U]o��Q� ��a<�P�֔�`W�� �Z:A��{[ S�I�7Gv���%VlG��94@)
nz��T�a-�E":����%�C7d���RI��KPg>�ޕ$�ݨ�4�/������sDz�Z�2\��}�!&���G�u�a �E� ��6�w� �s%��H}�m�]�9��*�!^VrOI4���U��F������l=Q�9�K�� �b�$ 8�d"��XӁ�����,�WZ�w(P�������kLכ��y��t�*7�"�g���eр�_M�u�����)G������|E� _L�#��.ɤ
Ș�����0`]��B@ N?�߃� P�F�	)����2��w�n2Y#�hb�<��:���F���xa1T�Zy���S���_���t<����5�qK(��5���鼕����E?�;�f��E�rk(
��(���G���&��N/�Y5JƯ���v�Ŝ!��M�����R���y����+�Ze5��</��t���!&�;d��r��LhZ8́1ڰ�9�L�3�������-8�ܼ^n������b���:��������u���_�+�*gn6����B;����S�*u���믋X�9��:h_���Z �7�`*q�&(��i]q�������ƬݍR3�nT���tG�
��Y�������%�$l���K��9��Y��F��%k�ujU����N���p�q�~7�$�wP.���q��vjT޲,{p�t�ˮ!�[�� kaV�����O�~&�u�u9ao?.��s�)&o3�����M��1��&V��lI��d|��\0̓���F�}�n�U�t���;;�bu�Ь�����$l�^�j�� ]y���	��z ��3�iԚ��|9|	�=�L�`��/%�%� V}�&���S�vk<�*�l�7��S�v�ך�W��@�� H�G7�r�{�7
:��h�4��'չ�=b�z�������H.RDԳ�:����_�_���!q3��O�c���iX���W���@�͘~�c��
�C��*�R�b]`��!���q2vt
g�P,�+r6�©��ӼO.�3Yᥖ1���LV|�������ڵ���)@��^7���QJ�g�.6b�͂W��2�ʷ���t�������B���dIY�F�ˆ-���'~��黽����,��<��K��.OW��.1梒�?H�t��@<*@l�����v�猝m�ao�k<�:dC�*_.�H��q�հ�T]xbf6pdW�rm���[l@D���!��2�8������w�橴EoT5���W�Zm�)�����}:�+NN��ӎX�~�Jkh�j��8�z�w�>�0�>X�$��]V�����GK��P"�lتم����+_ZDp@s���k���C�_���d��~s�����Ȳ�%+�ƿ�Ɣ�Um_��ӫ�u�䴕�|���I�y�����;5>�[��CV|�3xKZͥ���Bm��gˡ����14��T��B����*?�~:kqO��w=�!b�%q�4�I�%�$G^���I.�!l��|%A"[���*�㮔B3�U�U��^uj	z >���ԏǋ��*���}�yS��I����^
�%�9.,5�Z�L��7O��e� ���)��\Q=�ldw�D��	�,R$��v	-�8�A�B=��=�=��܀�'���j���+��\���z�-�D���)���i�#~�y
��q|���F�NA�z��7/���J�wVP�ҥQKM@�د�	�6��R�"&g��*��P�T�> �	&z��s�On���CNn�;&�5�l�*��֘��h��j<�Kh�{qϮjk�u�D���?ɻ��DwH�R.<#\H�F�z����E��[�B�'	3)]m�mj�@XN����֓ė�eKG��Dd�̀)�2{g�F���o�ec���nTOS����yyQ�(6�)�C�)���ב!��ؚ�a���,��Os�+*:�L�e������+�1�%-��Yn��A��_
�7e-�jM��̢rf�	�RV��S����rRJ&������\�|2�zK�Ӳ�\m����ˈQ��	W�O�ݿ����܁�\�^f*N��<rfVhU�}���V|�N~T���dl�0�������T����^�m+I�Y���+vx��K���*OLX�#�6�SqaѺ����{�C�bL���Ŝ��߮�U�y�Ej�5�]_~�<���g�e��AZW �J����І�9w(�<��t;�'�ռP�˨1���Ն7�Ls�����ug1j����7V�(�qv\z���L���L�7���Ey���x0��a�Z3$3`��H:���a/�F&j��X�`�	G����_�y�ms��A�5CbPK��{7Y~��j�܊�ɇ,���Ȕ7�O�k��>?h���R�����RN�!�6�zyNwr4216����-�wq?kb� �?t$���r ��&��S�1�
��ݻ�^��$y'>��%f�Smm� ��tei��(�ɿmA�I;P\���94X�q���p��y\�o\�\���#u�������i�V�Z�n��/�7�#ߊ6�xcn��b��{k� �'�@��	��3&��������:��*�f��VW���!��=O��1?�V$���'�p��~0p�W�$n����$���=�h�>�, ��EçQ��3.�������cqu���W�p�0�^*[�P��;��NA�.�pU��b7 S.�s���U���#��t�I��CY�	ǋ�J��G-�D�7P��5�J����y"�1�������:4�W���߳�)��鈁
�����	��Ow3�S��.z`fm�5��m�����<RO�qG��!���E�1SY۬�>�i����~��R2[�T�8���fX �)]IJ����j��|�-���Zs��:�Ճ�I����P�����rf����׼��%Q�>�w��7�h��E�P���MJ���m}�ٛFUr_>���0|K����oW�^����|� �}L�;��{�b1�/���XK��xjx6qԚJ$ǹ��_[+�Άq�����o�q��x�zX�f�;~�}6��$�[��:�{���,>.��}���iN>x�1�e� ���kĲ%v��k��?Z&[�s�|��萳��'͏�O���Lr��Dh�K��m|�~���*�����+�akv�ޒ�i��<1*E[�g}_wQ����`?`l��v1�#�yx~��/�����N�Т5c����+We*V�3�ec��.�>�r��KO#��~�`4� � K��Eª/�D#����""��H5]zͣ!N�{�I�:�e��k)���v�}2�b���3hD�'!�Eq��(�Ҧy̾"{��ۤ��ذ)� 6��	�����D�|�� �'W_	+�5�A|b��+R�t[w0Q���W
���b�q��8��i
����C��/�M�P�'�ny!w��5!+;��e����4��a�7H�i��%ʒ1u��R�=e��]Ϯ����ğ'7VN���^Q��z�c2����;=��<EOK���B�!.k"}��uWy���Zc�L
�s�y�Ւ�760�'�&�O�u4R���j�º�����1�����=JjI�r�%=f0��qD���kB�3Y���F ���qwKO'_Ç���p�.:�HD���"��R���\W'x�C~�(��B�`���=���}s@Ӱ�e\�n��W�;m�[�u�G��ސ���
O��[A2:wE`]s:�?I:�{H3�� '�$��͌�ГD�V��<�90����ٹ[-��a�ƿl��)�d�y$2�L����a�`��b��t�iQ�β������F����bN�����f��n��	3�ol�Xa�1�#(E�%䫏��~��&cU��e�<�ɠ�I�0���!o��c��� s�/�{s$��xH����d�xj�\ƭ�� ]��Ѱmm]u��-�o}�q֕piBF������,ò�F�T����9���j�qs���3�nU�u/<��ّ��O��힘O�Q�ϥh��X�3᭙��MEJ7��!?^����Fٍ|W�0\.�������R㜡d�~C��k�ZJ�o�i�  k9�<�<�e/|�k1��.��p����B�<���$Lkq2�=�! %)��1b]A�\�d�M�je��
�9�M>��9��۱.���=(ߔP|��U�!�y�������m䯛r���h�	�؉�⬒&�'T�9ox�0�#=�,�O�����,)�@U��V�{�Q��H}��5Qb�-2�����+�I�0�Tl
�rf|S���r��|�눲����y�q�Dr+9!�-?ߜt�h�<��YG9��|�6����e�lS@�����U>�BAS��L����H6�(��c>�33\QM���á��ɒOK�����p^r���K��s񤾦�tk�8<x����~Ð�-���L�iP��:��gu���擉H��k�%�t�ן��?d�����{0�d�ȣ�^���T�X�_*=�x� �8Ơ7��4ٌZ�_N������jS�u�+�b�6:�]G����C�M� a�F�ur%t���+RV��
E\%W.3൥F���ȴ/9�y0@8�������eW4k%%f/�f>6)� �X��T)���S�ɓ��y��,�d}H���ڽ���4O���f~p"��z��������*���?��U��f�_׽�
tݙ~�����s.x����Ϛ���z� xBk{����j�d_M�i-�'�,`���?h�/Ԫ��v[���_S�㵈l����_#�f1�~g!Ϫ"ԯ��H���>+��yg�8��,\�@S�c�,�n�:�!d��xMU�+���9�FO;S��}� `�Ɣ�f��ȍ�n�a�z����'�{��i��W��ү���[���-p,�d�(�����z�|��pxp��tG��BB�@�SSB��@����ᵐ�٭&�$�2��/Biϓ�]yH��rK�3NM"t��
߸��d��T�������K�0�����b/ﲩ<�8�U?Ȯz^S;�ݡ��\��Y7�#�[��Av��ǘ�Tǥ=������|R4�F��K\�K�Mx;��%�ħZ�8��tHG���w7]
Yx�vP��ߗ����)��>�կ6�/�k��L���x��3O��ȃ.yЈ�d��k_7&�r�MRn,���8��@�~�%�zAh��X=Dn�W-x�bD��\(�]V�����4��?ֺ�\����$��d��2�ê�Ϥb:3/��^N��-��3َ��`�g,#���Y,l��s��gn�N8J�e{&���@g�T���O���^�xO�T&��N@Y�Z�=P��Q�����-�<����_��:^��[�Y��ӌ,ڛ2I���i��ۚ`�??`�c�^��ߛ�xI�A�}�#�g��5QzZ��7��<���������
�5)�H�G��V���{�RFz��>I�j�f�����0�gL����'%��g/��;��XR�a���,x��fξ���}��,�fc\<C9�^��Vޔ3ߒ�c�H����4d�������iȖ�~��/�Von��.1i��Wn2�?!�.�I/�4==��4�����m]ݞ��]����՗s
��s%�ˤX�V2��y��D~S\��康Ǹ�N\��96tW�>	 ,A&�m�u1Ѕ4�CHlL�ԋ�t�__a^��V�8\����4?zU�Xv�O��L�<��=�� 31p�*�q���|�p�1�e�N���)r��rD`B��y��q����<:W{M��@۟l���1|�U���<��l[�˝�+|;���dBJ��3��|A�m��5�_Hsq3z�n�r�Y^�X�IXR�����hw{���^K�Q}��Z�uH�W{P䊛V�|3Y�u�U!R��*L���8rru�UmV@�t�#A�Sӥ���e��s{��X#3Fǧ8���5�O�0qB��A�ME(�E�#:+��'�h��؅�����e?��"�{�@���q5�v��5����
��꯰ڕ��Ԧ9�1�Ĕ"F/�w�CәK~ñ�]���z�
X��+�������t^�SX==3��+�!�d�C��q�q'MR�*ec��ˍH�r��E�w��7��ɀ��/on��.M���.�:gUS4��Q��j�~��T:I�L�J�T�+�@9oԬV��g�wU���n�w�(�!�]�������.R^A�%$�JNz�ԇz���8	
���0�ɋ�"AW3*1���0��4kj����/c����鄅���2�f��	3@�B�;b
�7羍�Jk��N�-����p�+`GXf���f�%��� aߩai��|N�M�p�)�P[�f>Cٹ��pa�*v�nl$���7��[��էB��TI�Z�t�Ɗ�`c-��N�T=����Mt[��|E|�?mGu �d����V1`�0S�1?�-��k����~�1���{l�;���v{����%1pZ��!��3����3�"���0�,� }���I��ŷ.��{��v�C�R�8徉��������s�Ff��!�9?��ו�O6?�>��3�D7�=#�~P���&���ɸ��ן�L�W�����\~��5��\-�^}����#�!�ƿ6�v&��.
IK����K#(����RA��!� ϥ�{O#t*�(��Ӳ���e�{ m`���4K�����z�~b'm�|P�z�3r��Y�!�S\��r�{���7J�B-�f}�hΗs8�a���3�:?�O��&��g��/a�"�2	�1�ﺼyd���á{3��IÝ9��O8���b���G�0�kiע4t�ڜ��}��i�^0�+;�Ѯ�U����/&�ݘ2�}]�Q�/��3{��8���ꌹQ#�n&a�6oY�ޱdR+�����=<I�<�Q�8ǐI���Z�������r&:�ŝD�����(jQX�����T�@�P�^9+���o$3�1v���TG���ȕ ���i��+��L̗B� !0/	\�P��$g�W�aX�%@�\<�L�Q�!�Ù+�Q�����I�	*���I ��P|8�`熌���v��\Ws{���rϑ+�Q��~�@%kV�N�Q���7F� ?2b<�ҷ�@��9�ؒh��F��_'��ms =HRp�hz'?Ӭ#U	]�>�?�阃�ϲe[�&��,7uB�E�Hi,Ze��I�S.�S=��&EƼ�3�J�]{�\�N���d�K���ɬ���Nu]���0r�-Y�̼Je%�l������	�S�a�e�l�� �g�C�.͈���;]_�,f�{R:@��&O��MU���N�0w��_�H�P7d鶞��d��B�;S Kd���ۋC�-�(7�V�`�������Y�US���h:��ݣ���|?e��<Y�3�z�lΛ��[t"��$>��d���"�u�@�j���W�_��Zl�	�\� j閸q�w!��}�� '�h�&N�-����VB�S 7����lށ���e i��נdk4�+��)!�͆�n�Y?��%0\�'s�T�@�r�6msMF����RrfP�k�$}a�5Sɝ�����RGL���*֑�%�Z�J<6����F���uH@��"h����YF��|�A
�ݭxp	hp)����k)��@qw+���ݡ@���š@/���u�͚�·93{?�oϬ9�i��N�}o�Fx>�OW��Ti�?}���^�!�Z>�k��Ȣ����	)�)p�%�층jX�g�����VEHJ� �J��q+@ŭ�*Bؤ��.���
ʢ��*�Żب��Z�}�����#��)��@B�y�Bz�>*�H����Y�K/.����[�����
��1:(�����s��`�Lx��ۘ+��i�݋��6�����,���!���7�͛����^��F��!R�! c!�L3��5�̈́�r>'�%J]j<��Fr����M��X�aJ%��_�����w����4W�g�?'�}�F�X��!<Op{qp��x�N�֏"��5����D����o�t��	�Vmi��\�+�J?�p��'�bz[�xg�G�R�����6���D���K�o�W���(ڌ/��7)����7��/�[��ı���Cִ�2(��)��c��C:-�sv�3k�Q8�J�v�y�����'?����R@m9�}����A�Nf7Ӎ��)�.��"�$\��x��h2��PS��G���Wxq� E	P+b�uȲ��EJ�Y�tn��L��������R��W3<�@�A��_�Ħ�;�k�;[�+|��?�N�n��ף7O�;Wk��"�|���$��%�2��{y%���Xz�q�8��Q�i�'�@�^���U^C>��*O����E���	��ce�N8���f{�(�Wo���2�2�<����B��+ �y~����ͱɼRSm/��\�'� ������	.�S��d�O$i[�"��N���9T���3L��dh����7�����/nj��"X�{�|���� �Ί6�0��;��ʖ�ėɗ��Ʃ"�4��x	��a�����ٵ0̂��ޢ��FE�8�z�B`�u=&�� �z�W�v��=���M|"����� 凎�U�.�O�ȪW���2�� ���D�f ��c�B�LI�ߨ��g;�}�,M6��G�n.�ρiD���cu~W� ��Jc@�nHYQWD�2����������Jt�A�=��2{���l��D��k�)����7|n�l�8�����v�H�����4���Z��7�M���3�-��QX�t\ =�� ���uXc���
��?;�tx���O�ȫ���*���lo���������É��W{6	"hֽl�q����ŶZ&����T-�F�X!�2�$(�\�l\���u�t)��[�xá6��}��+d�(�B� #�/F�{F�-�������������R�}�yW��4ą�mi���_պh���k*�����,g��%u���g�.8$�;י���D��B,}�$���?܏�~Ǹ������W�!�7�<��SL���Sj�w�/��x���X>��mC�M��Α]_g��߼U�{�������s�܎��<�3N�Fܫh�P��,�s�y�u�>�Z��L���_���{���r��x��`q�'�|�~��I&<g�I�1�q�*�ʺ)�O�G���yU(�C�}�BtD�W$FIVPHӶ�E���j�� E���A�%�&���z._�F�G���$�^�7�c�z��
�ڟ]��
ŵ����L��%R�����D��JzڴmgL$���ز�Y�g&���V�s�MX�W��������2� �=�� 8Kϊ�I(�kp�g�FOРyi�����yS��e�'nD�\+d�X��#���gi<K*8J!��r)��	C�V}�E2�Lꓞ�Wh�[ ɫd���c��?Q	z�A���5�����d�G���O�;R�8�E�8s��7����Sz z��+,�0�_�w#�	M��>%�0��}���Ff�N�*q�1�I�q�>��a�nY�JV~<L����g/��X�z�o��>J��$����C`�F��C�F��A��J_pj��`�P�-�X�/��a�yW���t�=+��t(�zǔ���;2�U�.��1"��Q{u�eo�mRoĐƈڅzgw�%���z|z��3{l:^���S �e��:g�Ֆ�JȞyD�*�q􋐐��@����ρ��8��K�Y��ˆ�h*������e�%���ߡLjB�y�2�(@wAT�^k�ď�u�0��tu�?��DK\�Ť������Â4�j	ܕ�������;X�����$-�u�l�_�����4K8ټ�zr����i�������y<@���>x�~�TJl��b��{XT ��6Yf����@���E�"έ���?.�9O�`���$|x����U�ޘ�d��ӥ��u-�ǲ1�qc����� ���^�)���=��5eyu�#���B������qC���1Z^D�����ߐ��9{5�܃��<M0�|*.胃qss�@��&�/lC�kUܷ� _�/��s��M�q��kg�_w�-�?����=��Mxi�u.e=��O�6/�Gng�|�Ǆt[QBHk�l����_I�Jԟ��>�m�k��j� ;�v4���L~�h��ۀz���[CixU�H�3lh3�b?���"v��M�� �Y�u�G��m�jd��l�ζ�'>��i�S����e����������˖�G\K�;��ɡ�G�s.J�O�}h���s�iʊ(Gi�os0s���UY��IX���X���+c�#op�/G�T��b�g�&^��,=�׋Y����b��t�4�x���햤@��o��?i����s����
nv��d�"G�]^����OS��r������uv&����k��E�DSȞ_u���ܗ})T�ƛ_�^��d<�#x�N�l��u�M�ӣ��6�]vW�;@�Pv�M8C�e{����5�	b"�� =�,R޽��.b�6c��t���[{�������M�U�P��}D��q�J�4@(���7�z:?j]e�2)p�$�Y���΄} �1��VK8�/,! �h���)���2;�)����Sq��?Ζ��tE�f�0���oʤ��@j�겐B��Z$�Z�7G6Z��p�e�D~v+�cu<��֕�7ؘ�~�>E��\�:ĝ姪�h[afQ!y���� ���0���ѩ�?�[����ͤ��V�4��$��G����������w�5�.4�,��8~<[.�zW��M��Fy�����z��!�]9
��Vt3� 8;��mZ��<d9���\4QKn4䘙��e[֧q���l_�Q��l��8�L��*{�J����1)�o��-D�5М��ɚ(�fL�h�f=�� ؚ�g�i���;/m1�_ܗ��hZ�u�L����8�˗#��%�`��iqa,n��,)�lTJ9I��W���B�!Z�2y�"&��o�})!���_h���Z�ApO\��0GT��P�e�ɠh����W�%S�����pGI�!�H6O] Ul5F~�ֽ���vGRw�W�יh�DNև�>�	���EP�dԵfX!-�*I; �X�gi���Jq:�&@��P��+��W(F��+,@�V���+7�Yf-ϻW��Ôd۵����>w�^ �j2���뺔�-mqx�YVҤ���%+�YL�ܵs:Z�Ȱ��S$�@ X>
���%4Oh�x3S�Ͽ� �Ĩ�L^Q�Q����;��f˦�4��.��=!��f���!�|�h��� �e!��d߳���๵qt�q�Sb����վ+�^+�K+D��7�?B��18�&U1C7UX"^�G��\ e�*F*�V���bY�@[.]�D�2�0,��O0�"���D�<J�9��	�U<u�G��G�ԉ�u�����Qӱt�=�����zu���2A�/��f�MǇ-��������ʗ�ZHK1;hp=�7֫S��O�׏?�-�ˈ��=�S�F�Lmn�5˭+ϥ���������?l��g`��� ��"�ؒf�5�7�;���RX��Ḅ�A��rj�T�,h��s��g��L^z��I��FH��[�<2�����˥����EL^e��Ok�����,<>�T<��#�?n��kl�*��51U/ü�c체:�;L����7W�Ww�� ��h���d�?Z�M�p)x_l֊�_2�=4}o��  �r\-�}�Q8N/�:����FM'���*p�o�G�L���jIӨJ�(__<��G
��Q7:.@ę!�ȯ�Nt%O���͉��׌��,[ջ�����v�@
�
���XVV�UA���Ɔ���(���2�;��2�m`�< vӁk�7�d`���kg�k�ʤ2�������{��at�9'��O���ֳ$n��c6�� �@�	QIJm�X?�	��fA�����QgXgdKE���""pX��,��P���x:p��S�P��{�8��&vTOS���d��6}u�$�Tx�:a�?;=�����0�	<���#	����dk�܄��(�F������?8_�I�e�UCD�o��]:����T������I���:�H1i��gJ1�� ]1���J;>�m�e��FN2#IH�H����=Xq�>am2�?�7 �"�SM����4�E� ������e�xǳ��� F�>嶑�<&���վ��>C�"������r��G
X��}Ⅰ}s0k]�"(�{ی�Ә|�p;d�$�H�C���@]�Dq�d�l3oU@�ـ|Zò֑v{����ˮ8k���?~n�������e����DM/�k(QF'�O2-�����F��@!*, �ӡ���sU�s"�'��l�_��3�s�B��3�z��+#�#3�_�6c:�+̈́�!�8y�u�Z���K�ݘ�/oK�g�!(@\��5��ay��iT���yݳ����"����/nt�2�r�L���$�_��[��[7x��Gх�G�&qtiEg=��<#���w΋�oK�D�Q�z㡑wS@z�߅����s�'���N�-���N���F�ϗù�q}��i�9?z��g��=y�����z��<q�P(�U,hT���}֙���&�U���t2涒Q>���4��X1\�Z��@rʗ,2��OX���^Z�d�;f�i+UF�L�������$��؎����N�"�:y�edS�*I�����%H�Y�U�S��+T>�a?������Q�"&�x�w��4՗��ۨ���F�Y���l��"$SS�MP�m���C#�d��n� �špG!b4���;�ىo�fxχ�	p�4� -���ɉOn/#��(�,'�+��Ic�%:R�]N�#~��p��<:�6T��T�ց�I\~�/t�Xء0
�a��� !�-'�i��,?�y�Lnk{�;S���z\�ua�����
�@_���c=�:���r��ȜPM\9����6���]�
�X�+�AgH.�<<�e�7���N%�Q� GЃ+�8���Ͻ�D������f_>FE$Y�FX~�����O/�Zr=�	�U	�m�C�
��e�F�,�*�5
����)�XP���Sk�Rh�L!��,��k��5��3-�dH,��s�O�c����b Y�d�l��y��s
7O�,G����M��$���ZG(
��0�`�=+�5��W�(P���ٓ��(��)��_J��ğr�)lq
%�lc��z4�Ӣƭ�<?�D��1�3�pڵ��ӓ8@(~lou�)ԅ���e�Y$����x�/\7�L$_Ϸ���V���<��~go�QY��ѨItt?6����%WW�Etk���Q�VͫZ�k�/;?j���`����yz��h�Ǳz�A�k���S/�֗˚�-���M�Ij����i�z��F�_�ӿ����`wX����4l_�v�(���g���C2�@+Gg�KW�'S�k�n�3�'��D1cֿ)+��x��O��J�8�3?�J��I�}�i%�%��M�a�n��V�3�S�\R��Vh�K��k��e���Bm�~�^X�&ؓ��� �+R�����_/�ܹ@Z�K���އѳ�ַ�U���k,�Q�"��,�Vx�I���)083���{��LS���C�c0ܓ�r���8g���$��k���\����?�\H�9�Q�w�@��M�й��t/������y%��e~h�����H�Jא(p���@�T~$��5}����2��ͅ�U�0r�ߣB��F���"�|�q�U*���g	;��ʀ�$M߼;�L+bc� ~q�o3�Pe��� Nׂ������bm�sD	�����R!BH��Xo�v�Ub�)/��'�^®��^�}2�����i�H�0�G�ng�ìQ;E7�Q^������ι��z� �Sl��,�{��5��Ɖ���5���U�y�VC��;F�.��?�E��������½l���d����AL��#B�������l5���cԞ��9WF���)}�:w
�䭪����W{���I��]��O��5]�z�2!�c��@��U���
'��nkr��O�{�Nԡ���s�(����L|���H��9�WI������Ӗ��a��c��VF��{5H@�d�
��(����}�<9A�/ĥ-f:�czd(Ua���d'jeG��&�Gv組MB� �Mz�ȴ�R��߰? ��n�f���Bn���r�����|hj�$|�20����M�o�_�P��M�`��u
�������Y�!A��\L���2"~�/Z� ���X6�~�>F+�+*�uޫ����T����1?�p��,x��m��˔!g�1V�M7E7�4�]kz������;�"����ij�Rgb߷cm?n/E7�j?����^y���LK��U�)�C� ��$j	�@'���8�Ӱ�W��3Q2/Q}���� Co׺̗�3ޘ���ZS�����p�J�7e䇁�x�!w.����˵��i����S&Z'V�m�dOm��c�JE8Y��|Ib���`�D/T/6�;\��p�uL?��D�8M�/H�����޸|�c�ޓg�\ޟ`�}_KR�k���^7���F�B�M�Z �d���TQz>�F"W�Ͻ�G,%?�7�"�C1-=��(F�΅�A=�Aɀ2��HpyB규g(�Jɔ� ]釾7i�V��l��:x�2/�hjh-,|��N5����>��q;�Ub��3������- q/���hhϘy�������f�%@g�N$jM�u$���=ђz�������җ��0ؑ�xeۂ����0G�Mx�Lh���
��m}?R�܅��A�<F�1-(8@:�ɼ|[�E���l���qE�/q3�n�lH4Lh"�M�B;�����$�d��oX�P5�n.ykRQ[����f3�(-ؙ��Z���Y�ر���wd,F�ކ��ς[��0n>sm1�#;��G����!4�L��νΕ�>
����4u��B�C	D��dRfM��i8�ѝum���!��9[�L�K�%Ns�mK�W�V�f��k9�#Z��c������(�B�deg�ɯ���'�;�vl�K���^x�᪕h��Ҽ6�¤x��8����a,��P�#͌�9sU���aǵ�,qc�	[�^py;���Q)�tX�]hݎ�tʈ���c��%���IU� � ��-���P�!D�1�?����i~�Q�������$�xq�� ���^F��p��ӱ�!�������A��[蟿��tS՟c/s���[]Ŏ�=���j��)�_��o}P�4�63��I��(B��u�]�����w|X����klv�8��e�Vq0�{�����A�y;�����'�sM�Vt]�:}�ߣ����d��Dg��2�S� fa,8F����/e2cW+�Bs�/�/��9k��҆�{�z��;C���ί�S��^H������y��tC �@X�x���D�;�������a����3��6n�Xlg���m���8��-����FJL~Bٹ����Q����h�Ε��:�]OL�I�w\��s61���W{tב������������ML�@��fFrWW�J��}��1�	���1e��A�f:���~���ڕwV�R��i�,�V[� &g�A�c-����Y\�m6��)<W�\l���Ӳ��]ku��{������6
s�8[���\�l`�<v��x�>t�<܌Del��6�,�J�I���4��|�ƭ���T��_� k��ne���Y%��Z{J�@�����<�ઽ�t�4T�,y>�\R��"�7*�s�"��݋+�o[���%l4�XU�`\�[�b��l�ݭ &�o�P�vd���&S��Z����r��5z�?�Fo���2���3bd����ʉ(�&LљbB�r���+'L�[�}��U�Df��q�R��4D�&������������-�ޕ�3=�U�}6�8��M�� �b}�,�so�r�����3�y�G�mI�ŵ�\��:����H[H��8ww��ܻc��\g��yE-EK.��b���i�R�����g(�	Ax)�J��_��E�wj��0I�ax��⢓@�e!V-[��>��/P
&��@Q�W:Fc[����VܝV�����co��6�~s�i�M�`���G�g�O���WEh�vY@N-�U·KO�Wd���%V�rzk�r��/�'����vE�uY����i(-�b��L zJ��*i���@X�����A�L� [��&CH�Y��[
�*dA5�y�bd���{�b��S�}��9���ʭ��*D�%�c��k��t������-�scs���L���Ҝ�j�j/��/P%
�Y#����K��C�#�.��,E�vM��C��Z\y�H8����1L��߯�J���#"Aw��?�Zf���O��׎�?aZ4)�vhaӾbЄ=��	���������4�)��9�p�"4}�̘?�z�׊y�dld��2�;��|��UT��+p_Y���ʥ�3>X3n��B�0�k挘�e��O���f��u����z"M{�9}e��,J�
I~�1i�hML�%���g[k������0bz���7M��-ln� �q��g2
�J�� ��qe��?(�l�Z��C!��z���=��63�H���-[^$�vHP��H�#��|vS��&Pl�'�e�_`$�ҁ�;�������x�|��urM��`ʭ��g
A��+I�����o��w�c:(1��ñX��k�����:��-ۢ���s�T��o��o��]��#�t^)�K���۷>�'+f �?dQ0�Z�TQ(�@�o*s������"���f\P�:�-(P믡� ���>��h@�(�@��ݡ\�<{P��ܗp˭(]P�ҰM�͘�'���-���(DŜ��Ӳ�� 0�C'`$sT|E�n�ER�ƭ\_��NS]N�ӟ�q�DՉ���v�ykUUߊ��o	��3��C؝�lRgPTP/��᜛!��%7έ���]��G��EY'h+�I�k��:��<����oCˁ��'P�	rz߆a+?�q[�u�]o�ds�o[�rz~�����"?��9nYQ��zI~�Y+�������*]�_h�/��Po��ER���G�o��\L��W���3�'W���+W�]#.��M��M�!ś�HӇ�ڷɁ/�������Ա��Wա���v���5�0���_����=cƿ����}kQ8��B3�J�+6L0:F�_W�l����@�_Gԉ����Nx��5c�6\z�ʰh�XX����f���M¬��A��? e��J�Q�� �h�w��zoL�p�ۤ �L%5!)�v௼�I%.��gA�*���U�W�󢉾�d�{$�sn��'�{�b��9�zj�]k�� %nv�kk�LȽhة1��	h���8�p,<��)$(�H��.=�"E?xu -Z~˾����a�y��ٟ9j��ZAҳ*قg	��C��_�~�J�/��{0j"O��:���eB�P�
#�F�`:��~�Dv*��hkP�s�� ���i0�S#�o�9����������1���;�K����z-\�<��2�۝D*ܳ	�����8��M�[�쏱�N�x"N��*��hA�uᾪ~;�^6P����n� ��;�v>�0aXL�S��f�f���?�3(��]Hom�Wte]�+E�g�]�Wu����J9�vW>8��|�rʆ��.�Q����C�D�Dz
���p���*�P��3p�bX\�1�|�S���Y4��6�.j�Wg1� �&1~���<�]uA��m����孚�[��\��Jѣ\C��Z��q��BޝxZI�ϩ�*8	+�5c/}F5�ȱj�*G��y��/�j�����D|�K� �4�J�v������</"3y�Z��v��ΖB� �ΰ�Gc��/'&ׯ�i,a���~�>��0��"M?ޣcu����鐦��a����w:7�ᠦ�y����t���=��&���䯂��ꁌ�1
'��Wv1v��������z�)!�l3);� ����<�yVWƁ]S���p��(v�D��&����S1���}��0./ؗ�ė�j�Z�i��
6'�G����:>�6�U��j���W;�����N��s�Y�� _y+�aXA���{̷Y迧���y�k�����^̦���7Y_XY�[q�y�����M)~��R��F���f����B�ꧠ�2��~��'� �'��ˠ��(�C�ӯԏ���QGx�������cq���_�P�b�d��[�6�@�l�2NB^�P�v�� �qg2��Q(�ա�X��/�]���mhl����D���/1�Z/��l��+��/��D~��#C�ĥ��yDO1%����l�ũ���L�����f#ds�pH���d.6�-�F��ܕ9�X�>�hc�\���;1|Q�A y� �seh��I���hI����[K<�;�(�}�������h��oD�y<pR�i���ν�Ix�`�'l[죣 ���p)��PX @⿘��M �w��!^�������{�Ǵ3��~���0���5^����\wᦅP��CY�Z��~���db񪦪�&@B���-��1�.Zi��o!�T)݈K3��G;�� ���S�OY[���+��Se���<����,<,���&��#[Z��V�5�ӫ��A:A�AM[�����"� Y�;�{�㳩��dk�BE��y��p��S�V�1���Q�"^I�h����v݋�t��\)��p��O�0���U�<{G���"�o��;y8ڣ'W�|G�]�˂º��4l�FD���u���!Ԭ��e��df���^���(���F(�#�����]��W��Ʃ�#J� ����O��D�d��H�F�/��D����R�t>}mے�����n��zi�K'��Xx���:������$���W�Ӧv�c=?䤧������ϛa�������$xІ���C�G�N��uI��<k���6
k˭��go�8�{��^��<�6w��k�Κ�����o]CP�h�9���~�&�b�?�`Ǝ��v�׊�nu>�g�y��~��5���|z��GՅ �h��$�LLH�&oNq.�7��]�0�wl�=}6���1�������P���z��P�0J=T�������]4K�,�e�d����mLU;���B�{��W��9���|d��A�4��� n�;�;<�����3��R��#*��qÒrz������_l�O���3��&���~�!PdF-<gG��$�q,g���t�F]��`���K��݃Ao/ �����1�G�T�#"֜����P����xk;�;�3l�2��8�׌�!w���6��4�v��������_��DǺ܄RE���0�7�'����:|�W���Gׂx�'1�i	�<~�"��Q�oE��G4�8k����uPi�wy�U����I챐�=�ގ�*.���=^���G����^I�u-���9���҉���[F����Ց�8Ë���n^��c�5�ڳa�gf��w���Y�c��`A�"$�﨟���"����UE�G@pi����F�6��:<vAiN}�;���n�v�$�A6�lޱ!ʓ�r�[�?q�^�нhD������L7$G��*7k��RYR�5w�Ž��M��9�dľ��k�'K��{���K��t���yHʁo
#� �X�fW�JU~N�=g��L��D�����X�#&�y%�Y��a���A	��zT�E��T_w��n����N���m�ާ7*F����3����	y�,I����a�7�z��b�X�������v�*F��{:�a����o]/8���p��g���0	�1z9�Ґ3Qڡ���&�I�뚼eBZG�P�w������V.k�X�\<3C*�ƨ�g���Hx��k����Z��=�pP��Ɲ�G�_Bԃ Jk�q�X	��+l[%	D�N��`;�M8'�0WO��{R�*��0��,�Af��xP�Z�8��"ۄ�utY�u��K�	qgwv2��.��0á���bjI�b �(�KI�<��/����PIW~���q|������M�=b$l��y>2����J��O�+{e������5C������=QPKh�r+�?
N�=j��sf$Fo�0��PK�L��.��Z��8˝�)�\����#�a< ���u����׃�|�7{�o���9v|F��T��x�=�|r��rYc�x���ߎ�Q�<5~����ݣi_��J�1�E�^?a�,��3r����C�K�s�L��r�>��~W	�<�hɄ��h�-�l�'��f�I<��<4r�SV����a^�W�m�M��4,Px�� ���5C�8�p<
��nW���X�Pz���?��J�TH���U��������#��N݅v��̅�/�$�\��;TK`�G���kA�w�E����Yx7Ba+�%��\���ŏ�+ο}%8F���� 0�T	
F��*&�	�g�� a�X����'+�O�D*&�c[�le���1tM��=�Þ9p&�C���ɳ�K�"�Ľ�xz�:����hN}c0͇<�¤*/nK�(P�q����\����r:tj��",�Hl�<���2�}b� 2ۧ��S�F/�����MM`��� x�cM�(k���@2}��t9ߏ$t���0[��X\r^]|+���ԛ��X��`�?V)f��b)%p��f�4GB���;C�Q��K���>�`=E��a��s���r�;��,]]�i������Z���1�B�v�&�}��l��(2&��8�Eq*t
7u��Ǩڑƣ�uBwr�p:�?�s���b��F�R#�pf�V�9\�LVF�0>AqQ0e�lE�.��G����x��;���$Q{bjW��~[M��x��?���wb隵PhFUĿ�><G�;�0�t@��x��e����FJ܁fGw�%_��B��!O\���0h�]=[�_�c��y��ҷov4p0���ݖ�/O�)S��j�g�n�\�}�(�c������O{��t
��̲���Jȴ6[�;�>�E�o�C_p�y�(2M�n�S��|���+���Ѹ��$W9� ����ZH%9x���'��9Գ�v ^JF�,=(��Qۙ��I�`K$�u�Ǚ����92$(G;B��·Ū�P.鱃U5A�#K[�$ٛ�P�;ح�Z���-u��]�b��@Rژ:��_i�ʱ�s	�YD'4�~�]� ������ ܋Iȗ\^�ٽ_�T����H�F�����ȅD��s��߫�QP��S`�3�:�*u����5)T��x��(3No�xT���݁�m���iV���������{��������8�tr��a���`ϓP߬~�ed�P[�xm�t��*�%\��!]�B���wt��O�Ί��;�t}6%`Ln�a�-���q%��D�U�6��lZ4�~�"=�FT�Vd��B��z�'��ŤQq�7����[}�+]�c�&�y]��Ȕ��/W��6pp(�~B%��������ׯ;Η�=��b��8�jB'��kSd/ޯ�|� ���f��{s�O�FNr�4�s�*���� aU��E���B�`�P�Y�������#�����8{!�AdX`n�@#�j��7��s��TP�'���\����3��÷�N1be;W�c��8���� {����#�awN�v���'���1�EƷY�o9;K��oY�`��/@���И=�qyq����;��Fe�>�RoU�XU�R��,+Tŋ�I8����y�0l����bQA�����iR�+��w��������qOK���p������*����:Q~@���H����%5 fWgIERG�'��dJ�sK��	�H�\����Eg� 
���%7�t[j���^wo(�	~h�v����]�t�&�Z#�l�q�)D�1i�Mb���wru���b�о��c$�}��苜=AP#�^�Z�	'z:yrӻ�Nȓ��r@ⶒ���'+�j�o8�(yu<L���QCV�gr����ʡnU8�Xb&��Ʈn}N��I���Xo����9�ayLd��E�+S�hp�]�����ǰ��30#V2�л���Iw���&�B�!`|7��d|�[�q�G'J�A��9c�Grq田�hRA�'����h�ocI�n�|'�����0�1d��~],�_�IB�ђ;O(f����pt���s1m�r��,#�@5��؊���t�bi����';�_��ۤ'�)���vq��ŵ� z&���x7�C�z~$�|�Q�L���+O*��V�M]���OY�W�X������V�>�x�ν�B�h��C���a�P���\��֋t���f����L��Oo;0j)>��b�e���`�~!���Y��]d�i'Î����a�h��k�|2�8Sw?���!��_:P�/QK�l�W'��!D�#��F�Y�YY��fƑ ���ON���R[��,�Di�?��r�x�d���`�vԗ��-�R������p��yZD����5�FF�5\�ox:+���p�:	,z��-�N����b��:�2ʱ���ŶF�gW���6����aHʲ�G�3��Fc����؎�	��Ǫ	�u�A�@M�C���'v\(��#�@�� �y������l�u�t���V'c���0�b:�Rnq���]�ޡ1��t2T�Q�=�-5 �Ñ�B ��)KX��L´�VbzY�g�eq��x���f���ҀA�3��.����CIZw2�Ӗ�������{l������?�f��΅� �E�,:&�֔J<7 �K f�/����~�W�"��Wn��{�:�='s';so4�:�.p H��~�h�d_���v�R���R����6A._��P�z�2��;��'��B�qn�҄�1�C�������L�?��}�S�M�mv~�Z��L�U:�W(Y�J�,-2��l��&l�j��}��;�m��<�[m�0�RKϡC%>��wo-���L 	�� q�X��wy�0z\�#YXU����|���}z2�:�Q��=۩FO����_Se�z�'�YQ|G�U�$c��5��<�=���;s@=������_������=!9/��٦}��Ad�,�$��ðǴm��9���F��je�Brl�Z�N�� ��D�9�8���I�
�7��XR�	ʟ%(v̳���g*�]�<aUu��5����X(_1*�[7��x����w�8_�&r�u��vڑ<%/�WmZx��\(����k?��a� -]���L)���E����*���
�]���oV�'�o��W�v���֦N�x��lO!6�uk�J�(�� K���W����bv�8k�>��A�G���<�m��{�{M�=}��� \ᅷ�-��`��6A],��t�{���9����$o㭋Ô��¦?F �مs� �^�<0�#?<E�X�̰�s�f
͋��c�b,<p��u�����.��qI�м����6BQ=�6�V�0Q�q.<���KJ���Q�pe�3�V˖�<-rdNq�c�b���蠪��m�ӏb������1�n�-}I�Hʩ��B(�Fxr��n9=��Gl�??�J��k�~�>Sp��c�if��Rd�W�V_�3�pO�%��q�yO�l�@��B��M�P���~��ȆveB�������OR�=������q���U�RD�Ċ�-��Րg����Q��򧹫�
�n$�����2��Tڟ����׶�����o�L�;E�����>��#A�e��4d��`{ʁ��ၚ�"�b���5�A��y�c�@�أ(R�>�O�S������޹�)f2�t��۰��N��.�l8�L���|����?5;�����~V}�>�#!�AUBc��#� ��<��W���b����#'��'�}�-�Ø=��ta�h9��!6�#$��^��Z��@����!	3K�Se��d`���-#S���$�|/�td������M��Vf�х1�p����ЇvF1!�J�7den �g�c3}Qol��̀T�N�!L��wB��R�l�L^)-�
n��e�n_7�N���I$\2����HN�߆im��R-��0-KzN�Hh��煄&:1,�)��m8#�̉�1<�|2y����?,|n�@~1��!��m�ǞW-0���C1���)X=��9����n�n�d��s����*urq 3߇na�(n+	5x����y��І��D*	���Ig�_��/�F,�[��^y��}��j�5��|?u�J���E�zN0�Ge��dtu����Ԁ{?���O��,�*�ib�l&��G	�=�Lk�:7bw�z�|�6�n�d#|{����nj���7��#�2�Z��f����nq"7��A`Ԩw4��_\����N��xI�$��.g�I,�|�djti�C������:�溨}Pi��k�؃�0)�", F���ӎ�}�;Vr4���f�3��#IԚ���ݲ���o��Բ��u.:i��M�1^��$�wn��֩)>m��k|c��?��s�W�mDԠr!�� ��M0�X��q|$��1����p�ad׆Q6a* ���n�i���"!N$� �IЀ�h��Oj�,��i��IO6T>�_9.N��_x���>���x2�e�m*5�g�1|�&:zŉ�v$���\膆.�GG&20܎$8x�\,�5������y�<�G���j�-�M����*�L��O��h�:3���	�v��LO`�wi�w��������Z����~��_�NWj�Pa��9�.c�L����������u��    IEND�B`�PK   t�>V����  l
     jsons/user_defined.json��M��0��J�3 c��sk��CW�n�K��0[K,P]EQ�{�Ii�M��	����#�g���4
-P�*�BW*G��L��
8�A+m�Z�-�o�?�ɋ�}X~x"��%�z��\�W�[��=�spL��"�����p�K&�i��,��c�C��հ�J���Mw�6�z��D|�T����*j�آ�Y�)�Ͳ.�x�� s)�������&"�C2�J��ABu�?vF�f�V[��t	+��q�2�^(�b��=�n�Wُ�@��e�*�v�yzx��E/����'��O�\|䪧�vxz��♋�#����3���șt���3;t~C������MMx�dO�l6�L������nў���ݢ%ÓϦ�5ݐ�,�!ݭX1$~��q+v������]}9��Wm���`�ԍ2��7uۣ�����Z��}Ӕ�)� �	OY^�J�ԇsP?�a��Ƃ༐��3��)�	�@D���up��۵� 	�A<{��]>ޯ��(���?���ry�E����z�PK
   t�>V����V  &�                   cirkitFile.jsonPK
   ]�'V�cŌ ~ �� /             �  images/40a6b5df-e714-4004-b865-d48720df955d.pngPK
   �>VS'49߈/ q�/ /             Џ images/a09c37b2-5d65-4269-9e69-57a504bc5c33.pngPK
   t�>V����  l
               �1 jsons/user_defined.jsonPK      <  B1   