PK   ��'Vph�(  ��    cirkitFile.json՝Os��vſ�+���B���K�*/^�*����"A+qBQ;.��)�D�������c	}/��9h ��?&����~:[�����a����(w5�ج�_����W�����f5�e�|�8��#�^l~���էϫ��~3m�.�
E��g��ա�ݭ/�mB9S:�L��ͻW�+Y���Y����.�%���K�.���n:[̍��y1[SXn�[���mk�A�t�r�����]�^n~/��_&��x� �d�P�R	5��"VB+����ŧ��SB�)���PZ:�
�����B�i���PZ�?-ԟ���g��3ғ�PF�?#ԟ���g��3B����:�%��\i|Y�]4�m�eQyUN�֋��ƨ�����ZIv�E�֒]Ѯ�dוh��c�
�5+<֬�X��c�
�5'��p�w¹�	�z'�e��	���sB�9���P^�?/ԟ������B�y���P^�� �_�/���B�����h�/���������������������7�/�/��V���/�z�gE9+����o�W��[�,�!�렞(aOʗ�|^=��$��ѷ�.�|
�V������>�F�7'�A����/�A��z�/�A�B�C7(����ݠ���.�Ç�[�]{Ѯ�d�A�k-�u%ڵ���u*�v�r�3�r���m淫f=<�D��@��g$�'��C`���J�K'ǗN�H��w���O�O���/=��.&	��1>�U��z��(vhT:42ꏯ���ʰ��Е�S,>��K/]�p��gY����O����d�X�˟�b�)_��mv��{�?��'ŧX|��W&���?���/��I�)�b�����x��W��I�)�b����x��W��I�)�b���ܬ���a>��_n߰�L���`�i��p �vq`'y���Q����JQ��L���`�aOF�����!*b�~�r���Ό��1DCT0�2�H��M�*���lGe��ˇ(@n�(��Q��#��`�
�X�����#,&F���� �&;:*3:B�}"E
v��Q�����F����!*��!��G�� [F���Q���S�F��4l�!*��!����:��l�!*��!�iقF��4l�!*��!�i�F��4l�!*��!�i	�F~�Gö���!*b�R�`�a�Gö���!*b����`�a�G����!*��!�iQ�F�n4�݈!*��!�ii'Y�@�����Y��
 �}��Q�����6a��9[ݭ��Z����۟���Y�E#Y��"Y�S��DY<җ�d��,5�:H��z#_��W1V�I�HX1V���bͨXCs0�bͨX3*֌�5�bͨX3*֌��bè�@����bè�0*6���bè�nU\+UUsI�����V�f��Ţ6���٪��AM#Iè�2*���-�b˨�2*v�\옹�1s�c�b��1*v���bǨ�1*���=�bϨ�3*���=�bϨ�3*���=����80*������80*��ƨ80*��+F���QqŨ�bT\����HO;�C+�N���w�}Z�4���@�,�JfhiP ˫�Z(����-
dyut���׌��eAO� C+|����<���yz~\237�\T�2Ƕ��e�{����^Tǒ ���ĳb�{g*y�K<+�4:-|�g��9�ȫa�Y�Aχ�d8tZ�a��//~�g�itZ�
2�sU&/��g��@��3� �=���xV�itZe�
2�c��Ko�YA�!�i=N<+�t��)/҉g��@��;� �=����'�d���ĳ�L�<��ĳ�LC��j�xV�9�L��~&��4O0�lܙ�ߜU6�W6�Yƹe#�e��e}_ eG��$ߘg6
�LIR�o�6K�w�iI�1�lܙ�ߘy����Ӓ|c��(�3eN!�1-���<�L�{B|c.Z7���3Ғ��|Z�o�Kw��)�7f�%�>���#N
w��)���3Ւ |Z���|�Qpg�B|c�ZRB�OK�k���TP��W�����(��)�ʧ%�����,)�����F����
�ͽ�6�i��k�L�V>-�7�%�N��$ߘ�6
�L�W�o�_K���iI�1mܙ��ߘ���O�Ӓ|c��(�3�c!�1-)�ʧ%����Qpg��B|c�ZR��OK��k���T�������x+�����F���]��kI�V>-��母�;S��9�K�ڇM�i�k���ͺ����k�Y4�� Y,��!Y<�% Y*$Kͨ/�^��W1�U���`�HX1V���bͨXCs0�bͨX3*֌�5�bͨX3*֌��bè�@����bè�0*6���bè�2*���-�b]3*���-�b˨�2*����bǨ�1*v��tcǨ�1*v���bǨ�3*���=�bϨ�3*��?���3*���=����80*������80*��ƨ80*��+F���QqŨ�bT\����k�Y^�ip�Zy�/�Jfp�Zy�W3�b�<˫�;�b�<˫�;�b�<˫G�����,��QW��gy�|2�bm&�ek3����t֧G� ��I�XKg�@��T@�Z:+�4:S���
2�s6*��YA�!Й��tV��3>P���
2��T����L�\�k� ��L�Z:+�tϕ3P���
2��T����L��� k� ��L�Z:+�t�(P���
2��T����L��@�Z:+�4:S���
2��� k� ��L�Z:+�`&YZ�OK�'�O6
�\�Z�o�*�+�,�ܲ��q���/���xZ�o�3w�b-�7f���[�$ߘs6
�\�Z�o�<K+��iI�1�lܹ��ߘ��Vn�Ӓ|c.�(�sk�1#-�܊�%�Ƽ�Qp�*�2|cvZZ�OK�9j���U�e��L��r+�����F���X���Yki�V<-�7殍�;W��y_���ʭxZ��_w�b-�7毥�[�$ߘ�6
�\�Z�o��H�4�^J�_�+^AT��Ӓ|c��(�sk�1-�܊�%����Qp�*�2|c�ZZ�OK��k���U�e�����r+�����F���X����ki�V<-�7母�;W������ʭxZ�o�_w�b-�7毥�[�$ߘ�6
�\�گi�������t��[����o���j�e�n���Y;�.匿��]On޽{��٥R� ���N��Pz1/l����z^Tƫ�,��{�~�����o��t0v��׺��2E�t],B[߶�ֆ2����z�+Jؕ���AW��d}�N����ߕ�����z`)�(�a�XC֕a��E�f�u9n������V;_����~�7��. Ĉv$�֢]�Qd8h�N��o�K6�����cp=�h�\���f\+�iZ�c�M_,חZ�͝����ez�Iߙq`O�AB]p_x�6��s�k oٗ�W)�8�/|-�Ç�������������n'�u�����_�ul��/���A(�D�~�A�#�y���f@�o3b���1B��y#���9ك7�r�=����O��΃o#cq��2~���&���RgF��A#�ԧ�W����c��P �X����W�ob��{0�|�M[y��@�ܾ�?8ި?�т��.����~�o�OͲo3>��":ե������y���(#�vio�#���F�O����x^襏yF<�]��g������z��9�x���G�R�z���_M6ͦ��<��Z,�v7ݬ�����揋�����Tpɫ��Zo��V��)$w^؝ ����TNb=J���TRI*�&�ŏD	�2TR*��T�Z�D-��J�R%j��T�Z�D-U��*QK�h�J4R%�YZ�D#U��*�H�h�J4R%��k�]��$��y�I>ѣ>��S�|R[���T�V�b+U����I�S'�O�t>u��ԉ�{�JtR%:��T�N�D/U��*�K��J�R%z��T�^�D/U��*1H��JR%��T�A�� ��JR%�+�+�+�+�+��J���хo)H��η�t�W��A7xxI�	�^�]B��{�ğ��k�K�O���u�%�ӿ�6x�������>�&x�b�����~���ŷ�˿�;x��u��!~V}z����2� Vrę�߹| �̔%zK��Y�]Ȣbfiw.�br��ׂ��ԍ=u�t�Z�BXę�ۅ�&g��IHj�r��CS1�B;�a1��:ԓʯ\>�E1����\>�����QO�r��3+�s���QO��r��3��s�/��QOj�r��3+�s�C��QO*�r��3��s�W��QO�r��3+�s� �v������ �90����R.	G�tpO�0upW��u�w�/z��IWܖr	x90�ܺ�R.;']SL�p	8:0�ܚ�R.S']/L�p	�:0��z�R.k']�ԓ7Y~�Z��IA�	j�']�L�p	X>0�ܲ�R.�']�L�}�U	�| tno)����^&dS��Q�V�r	B���`B�K��Q�Vޖ�T �B��`B�K9����`B�K�JW�2\��2�b��K�m�u���̭�&d�\�t%h0!�%�
�(s+]K�\�t�g0!�%�
�(s�XK�\�tg0!�%`�(s+TK�l�tuf0!�%`�(s�OK�l�t�e0!�%���(s+KK�|�tUe0!�%���(s�FK�|�t�d0a֞uBj�[ z��~�|l9���=<���C>��ܼ���5��m��^�R+_��/>݊Nw,���A�bK���V��*�V����UP1B���#t��1B�#t��1B�#L�0���#L�01��#L��1��#�A��1��#l��1��#\�p1�mA�#\�p1��#|��1��#�v�b��>F�bD�!F�bD�a;�1"Ĉ#�Qň*FT1����|�������.`�W�y���!�!�)��R�z�n�>�]�n_ɇ�7o��k���7�U`�Od�/�~�+�x�����|o�dE���WA��EB�Se�so�nh�~�@e���c`A���/S��m3�knۻ8ӦS��?��ߢ���n�I���n�I7��&�n*w��t��m��&����Ma�)���ݦ*^5wwӽ���b5�[>l"_���Ǣ��\?��?fz�.6�1c��H�ݴ����3]/���r��"��gi>�[���}l���z��]o���������O�c7�������}�)��^M~m��o��e>��x���<������������,������Ю^>,o��翭��y\����f�u�#�Ss��hf��u\r�����z�T$�Iו�0_n��n�Z��z�'��������3v��.nR�z��Eǌ�fH�:Κ���s�ꪶ���:�]�o���S̠K��j��k��3y��cr��ݵ;�ƅkwU�򰯵�p��Q������1�y�͗��Yw"�fU���Q`���<������gu�h�>H{��QEZ}П����ZU{���m�D����h��˦���fo �Q��~��8ۯ�����VA_�M�dȴ��"�.�$m���Yv8�fO��YF�vyv3��5�`�a^ƙ���!�0Hef��L��8a/��$p��w�����|�k�� wsaݷ���n����9*�9l��NC��@T�U鎍��W�z���o�uO���"|_��q���b[����N�-e�٢�zc|o��1�1�7�싩�B2莦����]�tf�e�ͷK�ηK�Ϸ{�B~[F����ft�m��Q�aFU����f4�o��`�aF����ff��m��o���������6�����v��t���u���e�\/�CwR�ݏUO9�U7�Vu�]����_�۲�n�(ڠ�S��k[�m���E��x_��c���?'��A�L}��WQh�!8��ښ�o~�6o����o���cL����Y�uǺ1O���B��5�~҇?������U��X�l���o�P�Ean�ʩff��p,�An��:��a�3�s_��.s;�o7m��u��2ORW�q���f��
8���������#����u��+�n���oԼ���v7������E��u��v���igǃ?�iŀc1�����2*�?~7b��\z+�k�ݠfǷ1=��4��na�q^�]3A���v�]�Ciͮ]<,���څ��*z۰���N���Ә-�9䫎v�tYW��VO8��U�{�B7���_%���uiuU�����u�黛��scC�\��+��$����|;AnV�<2)��]Ft��z����˘�o_���ǘ�ƹ�u��?~l�kw�ۗ�ߎC?��6�����.ߏ�v����e�忺)�!Z}������������u��������,ڬ7?.￟o7]�Pl�����L5��6׺��ٷ.߿����Z�o~l6���x���$ڪ?,~�~ڞ��_o���>+w;!M�T[\m���C[uw�{�?��B�d�����)�P�EmBK�#��а8+}�8��?�D����L�9�sX�C�_I��8���YK�Ã�P�8<+u�8v'Q�����L��������G�,/�Z�����p�8JX�Gy�8�Wb~G��U�3���2�ա%�/��Y����c�'�!}�b�V��j�V�ޞ)��)�£:��_4q���{n�p~��f[YA��;�~~��v;�A�j��5X���`���j�L9[_*���V�.n{�*T^]��yrH+s| ��ף�y��p"<���D���*|z�O�9�N��|���kX�)�pj�*�趍��6�d8�M8T�G/���o
?'��{��ܳ!�t'xhF� G���n}t�6���ذ�Y�g�3�JJ'��s���y�H���|��Q3�=�j{(�A�z�h�.��~X��ٴ�es�R�����e�������cs��է�7��ß�?�PK   u�'Vׁ��( �' /   images/31de6c7e-4b9d-42ac-b555-28e4a5bb4aec.png :@ſ�PNG

   IHDR  D  +   )*m   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��`Ƕ���9g�ﾛ޽�m�lPiFa4Y�l@q43�H8��䤀��焍��6Nl���E $����2������Դ:TWׯ�Z�իF��v��ܦ7�nY�t�[W/�����k���d��%[WG�,��f��7"���k��^A�겦i۪�e���l	Y�ue��W �\v�k��ŀ,��:���W��]M�l��4m~}ٶ��D�q����+�Y��M��KOzY��bG����r�����Y�c���/���?%��0�&r���
�L���+/9�O	�Ű�{����VK����ͯ��KN����°F�se���դ~㪺+��n��AfX�g�UOm^S��ˋ7����4�x'}j˛�o|��I߈w��mo�]X�Q�U֖Jj�2�VV��Ta��׈Ðtci*�2��:�U��U��#\QRkՐKV^�P1 iz-�?U��
v��ʰd��j��q.9�OJ�Z��A�#\[.�=,i��t#
��Fa���iX��D2C�,s� H��ݰ�� sc�ae�4����`GQU!;�u���npay,Y��l�k�T�ɨ.�.(V��d��t=-eU���)�6�zD�;[�qEV�NR[�l���DkI��8�R�d)F>�V�p�K�h�ƚ��l�[K6����J:��
K[�,?������]��2R�x�_IǼRy�!�
�NWd�ę��3��k�a�V���W���[��#k��׿�a����l���[�"g֒����k��j�ˏs�����d/v]�_���/�a9������Z[Ry�<�<5$�-a%���%�L�hSj���J�h���$}��P�S�[�����HU�I3����J�������zM��0G�ұ�o)r��MyBx.J�
�őe���Kzj\u)���a����~�;��%��J����\��w��$:��XF2C�z�_iY(��L�S�Ys��HT�+���ՉȆ^�Sg�t��6���0�̕���K�+�`I5<��k���e�-|EhHC�s�r���G���/_F�9fd9揖WiW�,�يPWX�5������%nJ�	�Gq�S��ě��������oGtr}p��%"�:�Z�T�����ȏ�/������L�*���?!���
m�����$;�D>KK^�� ��/�K\�ĥ�|��ߗ��#g�N��k^xi)��L���3T��,S 2Hj��5E�jZJk�y�ZU��W+jK�zm`PKj
#������7�3�XV],�ө/_B�W�K)�Q�5�/IId9�X�N4�G*��_?jC~bˡrٟ�p,qw��D�b��-��D�ms=K��8�q�����-�jr�0�"��Kx%sqw��a;;];&�~��\�$��]A���#ς�<K�1�{�\q����>`X���� ��P��5�X�n�)�7�����6nZ	ߘ�� m���BKq������?!H���������2�L"��6P�$��x;m��8;۞W�l��]W�Z�(�(3o&�%�+�/�]�͒�l.�-��q#�������۟������è����������?#oG�����w�������b���1�.�W��3�Ț�������/�/��;���?��8���<[�Ϙ۱/�X�?�(�m��6�3"8N�?b���c���c��_1�y�=�oN�3^.�sNb�AcS���������o%_!|��*jH�U#�G�J#��g��Z��c"ѬN�
-2�^����_�g�ߩaȐ�N�+�Wv�p	����;�-��cY��Ʒ�K��C�/���5YL��F�E��D���[��u�5���M�A��^�L��+|�8M�GJ�  aU����i�X� g����?��8x��+���*��\�+\J�z��5n��G�2b��F���-7���?��������q����#�򏿏��Q���?��,�����bbbb������(>EGG�OHȌ9������F�A��;�D�/�˟���?�	��������8������	�sdTl\B�095U,�H3ryZZ\fJ��,�^�jVf�M��|������p���b?Q{��Ax�Z-����} c/⠻�;˪���858�Qt=8��+
+�eB7��G@.��'��I��6�7:�=���!gW 2Xê��_]��"/c�+3�A��RW���t�w����ͫ�3{�B�㮰"���i"�6ƾt��[�~�A�"������$rRv^V`�*$t�X�f-��g�1���bĈ[nqۭ��_�cSbE�II"al�@ ����I$�������%VHF#�$F2#��;����������s\\\bb"
x4 �t�$&'&
QD`,��d2p,W*dr�$67-�2c���8E֢h���������j)�3"l%4 �ԃ�V���c3��`֬/9��	���	�a�Z2=���\Bx�_G�)X������+�Ȏ��J��Ȋ싽�ĥQ�ו`�i͌�G9�G�QؠZ��B�b̊Ȱ���#źd3��?���s$r.VV�H��!�b���?�#n�݈[o��&��o���;���D)�0Y"K�$3tYJNNNOO�J�X����4����<�#��'hǟ����2�����'
��C���I�(J�JN����d�B�e2�\)�-�#��(��/bw�I��@Xu]r��O|����kdGl�`&%O0���aD/�s����YH���Vd$3���cx�_M��e�u�?����EH�O�#6���vau����0+*t<ߑfnڲ��y�Z�,R2=�����:�eݞ	�?���z9K�D|�#_,9�+2jc`f� �R�U3`�����Iq���Ba\� )1.!>Q �x5|�
��b1t2��*(2b'�ef3~�^�	y�m���4��h���L�4?N(�0>	%%ũ� Y�̀^��%�4jtZ��<ʮ�Z��(�N�n�&l�G�:d�Dc��f��G�Ek�^�%�2r�_E�څJ��E���x�$��H� �.� �E
֠���HuA�/h{L�:W��~Ax&�ɻ���~sf͌���#z�����X���W�""'��
�朰�`G�����+;�'�2�s�b�z��_�����~�t���Ia�A��<̿��vh�ajb2h���(�Z	�j�-(Rfcfhf6�efHQ��,�#$#1K�� H#��3�K�����!%19=M�"�IS%�b�dTn�D?3ΤK���Z��})��=��:�Zb2����F:�F:�[+�zŋ�-��:ڮf�ǉx�Ƭ�����,��1v��H��<̫D��c��a�y����_OX]Ej���	U;�Q{����d��U ��q]W�3�������}��aFV��zv���6���h�f�bԤ
~2���
�t<P9�X�h�_U��"A~������b'�ti���LX:q��y�3T�2�i�d(ȸx���ʙ���|fP�<g`�H��e�4s�������$3'	��-�$T������I(]\<�;i)b��43$]!��gT�L՗�juR�&E�N5kĆ�U[�챊b�@d�W���2r� �n'M�]�`�
�Z��ny��D���ش׹��P�˗W��g�o�-+@_ �F����0ϼ�{�W�t!�����YilC�1���Ô	Z`a�*�����h���0K�|����v�T��W�3���j��fO(10�sKku�j8ߺ�*MV�.�R�SAKe55�?H���\l�<�Y=⤑*f��B#F!Qx��e����ʲqgIu��#�t�M#n�����B�ɲ�f���e��<�d(R$�<3��a^tJJ
6 ~111��d������`f,A;�@e��,���'�P@a2|f�޲B&���J�2%�Ψ(�]T�[�SU�6iT�Y-i3�
�@��"���P�q��mersY��,�0�i��2��0͆�f���m��c��a��2��2O2�8�$�P~�(��
��*3I�a��R����O�!جU���W�X��"�	~�@���)՗��5��;L��2]�Y�g�ƴ
�h���{�̾�)�B;����%e���\��83��Ha(�^��gi�;������#ߟr8����[6�_Y?�0[�H�Z]�f��]��Z_g)�5�%)u�(�T~�ӯ(t�at/�AJ)�>�tټuO�S�����u��W<�X���faM���*�/��Ӊ�F����A��$����[ڀ
�E��a�p���2����Ҁ�4փa0����׿B'�8�}x��@���`����1����Js�C5�4U�_Wq�s�����/o|2��Ah��x�$s��2EO[��V�i��*�1�;��upg�r ]��N�����z��$�+;����e\�z\9�݆��n�i��r}��yqv�{�����&�i�k	�Vg�Wjf��$��XKa|�.�N����!(�-ז�fd-RO��_���wm�����Z�u�}��C;퟼X�4_��Xb(M҃A~��Se��"�f����0�_M]f������Q��(�/:�DzM�~f���|�}����Nqg�в���Ǎ��Ά�>�������ʪ42K��qxNr�(�So*H�G}����]3�S-�0���!'5i�r����EK��֚Fs�b��v�Ӹ�^W稷Z[r��z�-���6��ɎM
�`�� i�At���Vb�����f<C[�'�Xm������e@5t546�e���"��g?�^I�df��a���m�:�~��r�WZ�h\�d��T��2����d�RX��m%�X�f)	�[|B@4Ƹe~���?��s� ǝ�.���/�����y��[9l�@Ǥ��8���{�7[�|,�����v�� w�N����3�3�(�DcBq�q!���i��P33��Q�clE#��f�U?N��X���K�<S���<�ܩn���;��������o��uP�TE�y��2#�Pc.N\\[_r�9O[�^����PX��i��ԊbͲ�;:���pg�]8{���s���q�}��i~	9�tQY���qU��\��8�"_d��Z�N�j����������yT�g�\�iM�T˽�덍Fg���Y�l�z�ىVoop8���:�'�ea���K`���&>>66Z~/��BpJ���O���4�ɠ0C!3�̌m��Rf�+1�c�qB�Y�R*
�Ŋ���	ׇ�M�m����&K�S�����ep�̩�"1�af&"�*��|
��<w��A�.�������`<����<���~/[��>,���<X����6c	 x�~����F�Y�LE���w�jI���k�f̋�.48����/��m`��B���3�,��3}�Opgi=��}�|�n���l��A=ʐӠ��q��3�4�P(6i�=����L����z"B���Y��in���4���.\�|����v�c��l(I��`0�"�Fd*J�ǚ��_V��\�ͷ>P��dq�l�z��a�;�d�������&��43���K��3��q1q�w�y'<[X���_��R�Ы@�h�x��A�aclP��H>a6V�Dv����!�)�b~���j��r��1e�c�Yg���Vo57�$1��Wk3�:�)�B�|5��.���N�"m������Ab�+��Ϝ�9A
����|���{�XY�`o�N���鲉穾����dS×�	u4u8]7STQ4�v��wGϷ�lx�>����;�%�����	v �����
�H*���rhA܎�3trl����b8�>[�N��Yh_�.���O�^$��.`-l���{����sgN���B\�K6H+KĶ2!�r����d���Ņ�����Y��J�,���mT�\g���N(���F���iw@�uǎ��!�����&̂��Q��1�N�q$A��!�C0��"���2� �O$��J�1���(g<k�A	S�i�n��k�Q_��U�g�����fqZ�N���`��hY���� ͅ�(櫎H@�ɩ��ʝ��̓�6 nq
�C����-��9y�8"^�K0�2]=3Kl{����q�'����-���I�p��1�D�6ͦK�QO���u_k;w����Ν��;�<��c�,�Bd�]�ɝ?{�̙s����?�*�?���$��x���~��Y.�,�5<��N���KUm̌+�Y�O��F�g��%��WE��Ӭ�	���D�qhE���`�U�9F����&�Pr�����0;�����`�k�6�	Z��p����O��$�����b��	��~2����2,�Y"�Sd�72�����p�t1��
��j�6��n'K�y�)��%�+�2�Mon�gN5��#����4߉J�9�bF9P3���ۀ	�S:���WXf�:���av�1�O�X�W��h[~BCI4��,��uV����;XѮ����J�x������-��r�ˠ~�ƫ�f_�0Rl�����B\����wO���i(a$ ~��rj�z�K���5���8�&�^{'�;��_Cp	���T��۵�v�c��M��&[���pV��A��:�l�o�54`��c@��#n
3P�=|���Cwhb�G���^���'2��ȟ��qID�0{5�C���LX��	O(c���Φ���۫L��/H7����k�O���aN�Q�4�.����녭��:%D�!�W�P:�w�сN�覮�A�0���t�����������1N��!�H�����b����Fۋ���q�����k�q�Y:%�S\]��{�w/w�ǝvl{-�����{��9ѩ�߷B�N�;�p5�͟>�89�S_�.vs���4�R�b+���G9K�a+���
���δ�.mZ0�:o�u�}慳l�s��U��z��xۭv[NN�̷�~;`���<�	q�_�Lv5�ƌa$�4�`֏E�o��xB/��X"K�����G�n%	��ib8�0��f��Nz��h�i��s�/�m�?�<o��I��E��Ezw�j���b0G�l( �f��]����_G�����W�K�~�pK��,�k�S����!�7�� s5����1����}����L�F�K[�/(h]����z�E��/��}蜿�;.�58�$��:�C�4�p����݇�8���$����������/�F5�/·
���WO̧��� �dTt��j�����_W8��䯔L�4#��Ւ��a��l�-x�Vm�76��t*d�����[F���o�b�M�K	����Q��;�`c3�/��B
��+'愣�q:����?	b�E��IUU&�P��ZY�Ze�J�T	 O���	��YI1��h���l��6 �;}��O=]ݐ���;���/,u�t���bB�t��tu�Nt�Nwt�j�����!O(�	ɝ^w����A�;�ּ�M�_l����Y�yf��`��S����f���"sa�� ��d��-ʺaE'�?����J�ˠ�ͮ&07���-��R匳���"�����|���y���b8�T��7�����i�k�9�QG�Ś~u�gX��^Fu�=M��uv�ɨ7d)U�z� ��'�g��Y$H��3���{M�2ð��dlC-3���I2�		���t�R��ۼ`��x,�r�;k�r>�f-E����1E}N���*�|�/�*�o~�	�;��I`�x��`(�;�P��"��pt��|����τ6��[�5=>��	bMK0����A?\ׂ�<TY�i����|�Ì�%W��
L�����̎�����׵�>s�$#�wC�vD冯��8�lp��1̆qt�0C}��u��Q�����s�3���(1i���}���y��������x҂�F��:h欌�[F�����;.�Z�b�c�b�l�{Q;::D1�����`	�9-��@3�{��z粥��YeU����L�Ǜj�n�`>0E4'�[0�#�&1����2~����1����+p�i�v�?�z��P���ˀ���=�F�Ė8\��o����Vͅ"{q��O��u�q��P<���I �w:�%�|�`n�NOw>Nq���W�Q���7NQ��YB�z�a���Ar�0�p�[�a-�Z���7~T���[a(��?M��l��d�Z�3�nq˭#n�"Af��񉰣٧N@	Z:**
:����g�OzBb� >sFF��c�|�q��}U��3���0�eSh�Ƚ�>��0�{OBpp=����}���69��H��o����_}�F�B?�I�CG�{�v�9���C���Ì5=]'�Կ�!t.�D�DhP�>�0D#C��lE<�|n�W�X1@�~M���L��Fa�Ԗ�ul�	ju��E�����R�(:�O%��a��+l�bl�xS����y��%��m������O����ǿ���iP3''
�3�iSo	���2�P���y�)���n�IYMK���7n�]wO��)*t�f�$>��'ti%\C�󙓽0��ff0�7z����*H�kD�'�� ����.{k��%j�C��Dt05�Ov��`���E1vz��毩GI�q�ו���E�v!t5T�g���5o/��A73��J�g�)2��s�����f��fl��6<��N0�sZ��B�zm✉#��� Fo�n��[���3G`��0�%ddp�`�y
�Ț�C4�D��3[���0�4u�L���o(�?��Gj
�U�5��033��u�5�ـ���AW3���M�`3h]R�x��ݡ��x΁ �\����Fvx�o��z�H�t��f���}�����������D?�2��¹�a�k?fE����;��Ɓq�~:����l��y�!�L�Pց w*�q/���)�M	`N����O�	n�#܄�h؟�㏀Y�� H��̈́3S�CY�0��,�O���]����B�[J%X�a�$�c$Y�Y����*���뾴�!ף�	�A�3�i]����23��"�������v���D*	�������`Ɩ�;��mȊ��O?�a��/e�C�N�QW��t��!����u&\�	�K��&�qQ�w���0���ړ�YӀZz?�N�D|^�ZF:�����q]�jS�F���:�k�`6���L�#n�r�����n�����O��a"�O�N\�0���˓��?��	�>Θ�$����˥P�bIJ�Xi�5��kc�8���_��&s8����>?�,�+����n[<{~�)��t�����顎�v�����t�u��:�.����ƃ�C���tG�of~�HA�C'�(�����o��irQ�?�'45�4]����{V��`x֏^D����$����ov+�ֈ`�Ѡ���� f��4�|������z��[٫��>s�0C���F���
��f�Z�Hdi��Y �١���4��%5pm�I3�i��a�!�H�1o0��P��� ̞��'���:w�ة���֣��=���ͧڎ��?�j>�n�i���V�H��ni�������I�|&t	W����mˏ�C��L2�i�Μ�r>�e����p��NM�?p��pt�kw�)�������2}uc(�8w���.g�mCa,�(0�o攚�3��[ �M����;�����qI;� 3�f�vR
�$.&6-%UFK33UJh�\q�iN����fg�z�?)73�=3�kf����A��C'���{��;�mn����q`��Ж�:6}���q��=��6(pO�	w�����M�I�/IpP��2ku[}{��v��L� �<L��p@~�+������fN�ҫ���ҍ�}��)���7̄��7tsg�ܙ�%OJL�xSQ��$ƒ7�"�����6;V�K0��e�7����E`��m��'��r�J�J���NOO���f�Ό7�[��KP��lo�U`&�s���.��Kʹ����`�w�����ov��z��sqW��SOu4.	56���:����{�������uü�Y�ݞ�������'N�ꅜ:��~z�w����G�e�O�+�IlY�2oՆ_��H�4���m{U\K���sX3��z|��J�p=������p�{���e"�������<�>aq�@֡�_.�9��8e�Ģ�Tͯ��|?��Y;f���o�$�q"�'@3K���ܜ��f�TV-�X��&u��o*�[ޥ�p�a���2�=A���\��@���m��cO=���w��Z�5/�Ӓ�ϊ�wL�L��aae`՚�}��=._�����n��6Lv:Y�F�QW���	�	̄?]��A5Lv�=x!���2n �sNp}G���{��������[G�9����=!�|/w!���p҉��x�q���ǉ`�
��Xsޯl���RV�F?\\�4����z���v�-�c��0�裎d�H�.A�)��n�<���ӂ���F��^
'N��������ρf�/�v����t�;��~ݮc�-�\�K?�r�G�'������ߓ��t�ҩ���4���ի�8��q�c9}^��;���1�����<���_s��0�8]�Pm*Z��՚������@���Ý����ZruaҼ����A�c�����2cZ��G�������;��N�mY�ZQ�j/�1
�8E������h��E%�OZۚ�u�\*��ۘfN
��a�Ȝ�gc��B�9%�t��
�r���uN��T[�hk�0�Ѿi��.���3�*u�y>������p�;��7z�3����7�L|s���Ksw�-���1C�w�ʁ��w�Z=hf�Z9�#�53$�RG&������Z�{��g�7�6ws�׷�k���PwU�as�fn;ҿ��a�q���+����Vfg?���`��D߰�c�׿ޘ�P'��8�#Myq΢���8���u�_.h�w��.x�b��,v���
�0�~��`-���"̉��ilZ"43R**-�f��F�vj�����"K��9є������`�����n�w�4"�^5c�����jX�.gLSJ��y�53rV�T�k2�>Z��}���
������}�����!7?�3�w]~h���٬��P��
f��Hd/�1��(ca"�J�$ý�|�Xn���C��Y�z�~�5��=Q�ޑ��̾�f���4h�*���{�x��p*|��H��-=����<a�,E�jAP_�PG�Z���t�aa���G������_.�]�I|�tE0VVScE��~p����l��lÒ����,4r�mf�3�&3��M%hfO�$�I(lv�TRQ�����;+����5O��/�ԨjJ3j���|��<1����**v0&>��̃<�9�f�0��_���w<>/��w����3K>;f�2�B�*]���G����St̰Ȼj4s��5��*�B����5,�<�%D���\Xm\q&�-�,E1���%�F�N֗%Z4B4��Ғ�'�M���a-��Ʋ(�������0��4������J�:�Bu���ۿR��p���һ��4x��Ġa$��Mq���r[?z9s�VVˇ��[_T����iп'_+�(	���〳mX�����C�9V��cv(����.����P<�y�c�6�k�)�n����i�w؝��:
3{ܘ�7����x�)"'S}3ߝ�[��w�QD!��W*$
�16�nvZ��&{U��b�uQ�e��ͳ���u�	���h1�L�8E;G�ь�T�|cH�h�3[^m��LQr�^��@���t�@���g[��X�љ�O�3&ˮ��H��.��b��|Ձ��_�W��0�e͊�#�w�[���`{����y�����~:�HK��^X����GB���Ly�=��(c�ezl=��h{Q���B�Y�(J6N��N��ID�5ę�E6
�#1h��3^:�����s}'�#g�Q���Ν�o�RW1}�������.*J3�uM���^����A#X��f(Yt�d�Vᘑ�� W_f�����? i����}|$�����zu�'E����JL:F)���*���)(F�E�Y�a03A�`��WU�X�װCѭ��?al���L�QtN�ü��h�8��:;�����s���X����Ą�0��RR�h(��r��b�CRРFG�bGC���t�Z�p(p.ģ6�RmA�/I1����:��H5�Oc�>������ɀ����r;��>_W[���������dm���퉣�榿p����fn/�R=�������W�=|���J�L}n��#�o�f���z4�`̐��l��(I��S@��p0v	5�v
? �)��S�R�9�M�nM�[�U35��4���3�I0�Z���b��6��8��i>�8�������������ɣeOU��ޓZ��^)ue��hSa���g�̺�Q,����ZKR�u���9/�v��޷gw�{_�o�Y�f��W�|��j�d�0�Ʋ4s�4j|�H�%���g��*f[^"�L;�pp�4#	2�ءd۳[Y����d����%���d��a�;��[�P�v��r�<f���ۆ3,m���p��8l�:�!��ٙ�aw�̍��)eIVm{9$���q����G�5s���^M��N���ӎ]�vwg����き77�RX����o�f}���mt��lknֺ��V,p�Zٷ��[�
��<ސ/
�;,�̚���a�
����.0&�i��th�s���kI���CQ��0ɀJ�H�傚B�E+v�H��⌅1�B�!��+�6��J�r��S-��?x��C�}�s��>��/N6�{�s˺����<Y �֤�'�&�+ʢRH��6CT�]lB"�j��r�c�H�U�%�R�a��B#��'V���e�gdXfᡒX�!�۸�A�2�$Æ�xC0��d��?���!��`%v�fv��i/�PX���V"#7�
lB3�����F�����
H�֏�>~�8�<�F0�/�~�05�il�Lf�X�
�����;IQ[�l��}u��R��;7� N�C��1怏\��	ϰ���M]_��6��]�����%������]����Vk�TV**�����WUkZ�z���?�py�*��;���y�~�HV���������xk|L(X���NV8Ţ!��WS������֔�W+�3DU�h�RkY��D��������hC�52}�X۽��R�B����U��5:��L��Tj��j���x�t�b��z�ЌѶ��7 s"?��� {8Ř���|5��h� ��TT73�9Sdӡ�q��8CQ�C�XOA�h�O,a��xv??����G��8�;S�|��]��������']�afE�4�큊�̆��a�Z�&��Xg��;�0J��O0�L�F 3�x�2��o*%�;3�,K�r�LA�ƍN�	��vY�l��X��4�n~z��"�ٱkAr$>�=T_{jw�0C	�g�Föh�)g����;�ڼ�n������'�|o�y|�ʖ�W�V��[��o�K�o�>�j��7V�v}�}�x�7�w�B�>�;\���r�4&���|A���ih�0�Ѱ���le�Z
����L��抚���-���+�7�<����7���}�>�z/��7�TU��/�G�4QÌgi���P�	Fh]���<�Y�`����p��k��<���8�(�9_`�g�m��v0'��Jq%1�|x4��S�����k��tj�Jc�ڿ���nȇN�whcl�Q��(��N���%�'b��Y�ìFHl��C�5v*X�yvpvLv?�}�\sJu�]�{�?g�Yf6/����Mv�Gm��T�{��`7���#����ۇ9C�PJev~F��(���n��BLM6��~���Y��a^�1�[h�8ff㦰:Gu��`1���~Ã��j?}�xo�9�!��`<鮠�������=t�����?������9}d���#ݭǻ}~�e�Q��Ѐ���~̬��ȟX�:��@�'u��-��
U�uO�>��{����;Ɲ��T���m�_�n9�۸3�ܩ���^���0)[��DsI�Yg��gc���4?�q�]���N��9��u� �Ao-�7�%Z���,�af��`�'G1�"���ء�7L��;��Qe�(�2�fk�(�]T��.Ѧ|<�Vb�� ��(�ȃ4$�(���O ���'���X�B�g��q�D,�����p&8��ٚG��,Xn\����r�KM[j�4ٔ�|�1���m3�ֿm���"��(�l�L�i�8x�p���:6��h�?�d�O�lxhY�v�<������Sh����ލ�����tS7Hny�!R�@�>�
����ؼ��=�q�q�u�wOk�}�����9h;��=��o�
��`0��[��A��3C+٥���6Q�B!qಚ���dH+*Ջ>X��p���߷|�k����^^ܸ��ů?W��r�ӎڧ�uk��p߶f�s/�]�����@:�TUC������0���:��?})D>ږ��M�,Nt�U��9ܼ�3�]�"yu���I��on��IQ���N-o,�� '���+"k����VD����4��qF&2b��/��3<�4$ͨ��""|p\���%�Ȃ	��R=	.���v";;[Io�̺���N���3ܛ�����i5�?�Ը��bk��luZm��9W�92��o*��OILωI"1�B"5�V��5��ǚ��'�k�^{d�����{�[f'���������M��UǷ�1�����m�3x���e���y}/)�6���mBno{��������qX�FvO��D5-��{�0C�U�A��1�m0�Y^X_��p�c;�ss�W����%���zc��޺���vm��Ŷ�_n���歟o��Ŷ��m|���/o~��s��8σ�-*�Nl��L�a������My �z�lEdT�j[AB=�>c/�F����mp�y��`f�ĄV��6�s�O�9�
3���ˏ�������م��^�{~Q���y�0{yŽ�<�񾧫f=[5���=O���T���5�=U3����g*f._4��E�?S}ﳕ�<[9�
͊
��<����a1s!:x��b�&�Ov�H��Јe�NQ�ˬ,�Z}���������Z23�#n�y��7�~�� ���ǎ��6��u'!?	;�Ȱ�al["a��|\1��u&�̦���iR����aa�f�r��>ot�\&M1_[�WU��HU�{ͿW�A�����a&3�"�!�[��Sʙb4���`#a}����B�C�^پ��5�ݝ�'{N��9�{�{�$��>יi���o�� Ww	̑6	�3�T�	�
E�=�RS,�,^�v�A�sW�5�ٗ����/�l�jۮ�_~��VW����zZ�Z�z=-�����]�|���-�~�����ݟ������6�����9t���J֏A����ݑ��@������o~��@���V����%0��o+���$���1z5}��;�M��Nwr�!�?����/z��%�xi��� ��N�sg�p���A��(w���|��&�I�qc�`Zr�쎢�X��݂u`$C ]�]5�h���&��WӦT�裩[�d �afI$���?���+V�x��^z�%d^�Ӌ/��r�J��^P*���/f� 1!.>��dy�0?�p���Q�|��F�˃��2�A�n��ЦԸ�'�Dr�����H��PW7�ƆmҘj���� � ���"A��o�;��.���E��3��@	��t�����3k��MF.Y�� �X�P���Π)f6�p��\��Z�s�����������kn;���i���
�����sw�ԞVO�1�}����{?_�㣗֮����8�����0��E�Vt>��2�<}<�$<�?fv/VAa�"�sP?֕ܒ���p��~s���l˺��u��?�������}����_#��|ೖ��n���>?��燾�ݲ���c��������G�:C\��֧,�7�dsAG�����D� L@���*&���T1g�BKU����ge�F�z�[`f̢�$,��-�y]�sll�T*�H$�����Ξ�0���L?�`9q���nח��槧�%%Kę
enf�c�48-z�Y��L��D�&^	�	7�5&� ��ȍ*�����j��d
�a��`�`R�>���Qr�hu(gB��3>��u�a��E�Fk��s$G�Ə-1�,���u϶q��۲�a��-�l�z�WG����4S�����j�uz(�Y��{]G!~S+�?�r`��+>YS�JCwru��L}�pQ>xfg�ċ��a�mH</	VM��Z�,�q ��N����#�8"{��~�q]�����Q-(������g*�e�g+�9$�H�T��*Q�J8Z�>&C�#O�HgK�&�L.�>�A��'K�4�/@Q�=�UR��7��N��
@��:6y*�d��LX6.J�0ft���?�����aN�R�~.����0��Ǣݙ��ѣGgfff�)+++##��� �������0N�O�'Ĉs�T��ȊKԚ�e�:Y�xiu�����P�e̓WvI�@X�1������`� 9mDXb���0��3�L/��G �9��"0��f;��bt�N]|�4�E�2h�X��I^��3������aEw=A_������=(O��jm�Z�f���{<h�ey}�o���z���O�z����|����9v��2�H�3��!z�DH
� ����A��?��T&t���IL�����1��m3�}=D����O�:�g/�1z�̬9�)�R�J.U*"��o�*-C�������"K)˒����I����&U�R֖?��� ���7k��^*�/�k�
�`%
6X�p�q�bc�`����`ٷ�;)>ح�D`ƒ���I���Æ9&&&..�4�����ao3�����b��}�	0�A��ɤ��T��R��ry�2:'UZ[��,���:�Q��8�Vuea�4��c�p53O&�Z�P����3�MC��++�ӛ�z��ȴ���y���l}0#�$������''5���DSa��Da�L���f��ミ.~���_n�s`wkˑ���x�����8}���ӧz:`8x�``�����f&>����}�ݞ�G�o�f��-�-��5�<�����}k�j�e���ml9��/3���q(̑���-/�9�����k]1K~o^�dU���*�4S���$!e�̂�2��Y�T�*S������Ӧ���LSUͨ���N�o݁m�]�Uc.���xf���Y��Kο��z�A#�w҈��z��dc�<�0̩�?�Y$�)چ����>�� 3 Fހ<-- �d������T��u&&9���bS��rI�\�%�)dr�$M"K��J��,u���h�t��A?y�fuń�Au� ��O,�<��x&J#��_}K�'������]�����O d�����A}�~vqg�3k?R���QւD'�y!۪M[8m�����ʧ-|��7?|�r�!W`�Z>u��M;@_�;s�Dg��r��|G|�c��h���ccHk��������7�����W}.�"�3B2�gVլ�����T�_��_��ɘ�s�q���+%�/%|�㧽=���U�O�L�+��c�
u�ʥ�˒+s��T)��I���P¡Ud��IST���?{���d�&���$��'6��s�x��]�o𠳐�`�O�ѻ�$S�șc(:'���l�<洄0��	ĮX�b```�ر`�B?3������sԨQ��y�	����8Q"Abzj�D1&]�)�)�Б$�ɫ�	v�l�� Wk�al���+&�����&k���]D Aɑ����4�O�[�_�n�Ex�u����\�HK`W�5��	*�N5��j�z� �����om[��w�n>�s7w�=���΀�v���u�������I_OO 8�	��}ǃ��v_k����q�Z[Nt�Z�}������d
pUk�E������	2�2I�ʧ�Ce�ea���`�O���c9i�h�g{�@ sˀ��?�ҿ�'����(�2�2i�B���f+�����R�D�t���91��f(�U�L����eˢ&�=�8��n�zK�~���d��	�&���*�H��ri��Q�Ǝ��7�����}�-P��;�`ff�����l$�k0��l6f$X07��N�\.G^&��w��D�9!1E��"��A-f�D�U�t�h�t��BX��6ޝh�Ktij.����ő�Y9\�<3�ִ����F56��S��nw�ǅ��v�Z@���v�_ql�&�:H!�y�I3ә/���t�1�$��r�^p���qO�d.J7?���������]��?��2Y�-� s����z��!W�T���h�
��������!��%�>����t9���0����][W�g�w;�8�*6���H�Y�L�n�O��͝�I���:����#���˒�Jݡ���|�DI0c/lSD�4���6�&?�Q���t|�: K�W�� �Y�?mbF�EjutI�*���|Ij^Jb~� ?]P(�&�b�������Ly�s�28�pј��کx@nܽYY�Z5g?�ƅ�t-�� "j�Z,�Sh�$�F��eFԌ1�V��&��������ĤQ<��'�5+���stt4�g����N����w��H,�t�ܹ����nח sj� 5Q�� �UY��2�J�4!'EU����94"gQL��T']u����A�1	�N<�QB���C��F`�{��p����M.��
�
��;�u;\�.�����;zv�����3p��sG��:����=��}G�t��:;�]no���R|��~�s��2Xq0�Np}9�{�(Ot��,�p���;�!nvu�� ���[�dS���'�R�X���^c.P8��p�U;�z��{�}9�k�~�1<n�������6��x��H{����>��w�w�F�������s<l�zIK�y�ښ�p����~fy���;��b!!��)��4�T � Cm�'�P���j������0��/<�����T`�
��h6}�R���$���(KP�G;�k�����B_x��r��(:���0�ꑖ�1�<�Y�a���e��U��Ly���NO�O$| )�aa����#��'�O�~X,(�&MQ��eyF�4�vZnք��8Ժ�6�j)n����I.��l�H�ds�%�JR��l~F�ߑ��o7������7���w�%A�"�a0)�q|<u7�A���SRR`igee-^�xժUo����իW�\	�?_}���^{k��û]_�iq�([\�@��e�22���,--E*�e'gՖ�@��J���4�c����O%G��L�Wn�4�!�.4,�3H�a��#ݮ`�0�[��m>O(�s��=ݭޮ��l��kM˚mo���2�����_����Ъ՞o����}Pс�ΰ�#0�"�)��P�
��C��eI5EB}�a��DP_��C{ ?"[I\�T��@H�b���%EoԶq��O�7�����0�yI�B�f���/p��oq�1���t�.�=�ϝ�Ŗ�pT���>��b����ow�^_ۺ�z{�\{����N������bW��8��N��L�sX3_#�.���K�FY�F�a�$�KE-�gf4��M�M��$G��������v�)vM�}��X�P��4����K������?x�P�ɒeR�V�R���M���ML��8��քxc�(gtlcTܒ�x{����X�H8E"�/�+��P��f����b�f\K,�B�Ѱ����_$����pۨ_��R���*7���ro����[�?��?����-7��91������;�LKK���&7t5�Hl��Ì%��f+�313;)>aT|,4�B"U�K�49?o��i�D���%�*�/U�wm��J�[�JB�����Kl�専D`y���<�4��݁&�y�=����6�g;����ו��n��]]�V]q\_y�Pݬ7�4.k{����G�dTA��#��n��`3��R03�/�~@�I�@��?m�*�k�y�gJ�ܥ��B�6�� �:�:�qf�	vYAz}�$��'>{����۾�����rk���<�������G]�w3\蓝��O��xil9ۘ`��AL%�l�j���>��핝_�7��5���R
2\�/�ڽ�f�0Ai�7�\��(_\Y�i��I�=�A�K��2K��X[��e��T1i C��P(�̗�u���������r�D��ьTz5����#π�L0g+e��i�bg��uU��I�6�O�d�-wM�9�ϦL�`�h� q�H8],ɕ��J����5�$������iFM�����Wt��xi�BF��E;��E�9
��h\�}y�T=jo�-v��Ȕ�v�m�9���Au�0�Rp�%�f03�������E"27֛-NN���a�B�@�2�|�Q��n�[4OܓS33�V�TW:�Z��P�U�Z���O��:$<y�υ���0�4���Cf�/@f6�jo�������ٲ�PS�:MɺiӶ�m�~����6�ݵaꔝ�E�ִ������]<Bm�_ʹ�����$�/�����k����:�fu�y��=�ul��nغR�d���\Z]*��;gEW���O2�0�5K�2�k^��֧�~��}m�g|���P���P
���3��yCA�g�fy����ydz�jkv7�f�sx�G_n)�?����'Ƃ#�����8�0=�l�����*k���%?H��;�֯η�B�pm����S� U����ͯX�җeXfeT��ߵ���Iy2�ֲ��/�����G�bEreaRm!qn.���][�;ӎ;��=j0�;��dI�		5�F�PJޝ��~�TȦ�i�j���|g��ք؇�NOɑKG+�2���jJq>������X�6��c�%�d��j\?,jT�^�C!�F��Hu����V�@���^�R;E �9��
�o�����O�"�����A)�e�Ԍ^X��'{�<r�H,�,~�᥄����x4"���*�b�cO4�74,��Z1^or�Vd/����[y�&��uZ<����0'��Xok=������D0S�42L9�=�m7���K]Y��.o�TkK��Mm�ߙ2a�8Շ�)�S6�&o*��ә�_�J�j��U�����$,t�7��1����M�LCa�t�����,�k�k�r�����a��N����������o������jQEtR��L`./�'��0��|��v�����u�����>�����=^��3,m����:̓���ma0C3f�̰�C��'PE��}�|��֙�'em�����F��J��.̙53�gn�N9?Yq5͌�D�)�襅��V?��5?wbŞ��WܳƬ0he�Ғ��� w�.���E���{�q���cßRj
_]X��ˍ��<Ν,}j��V+���yW;<g�j�g:P���c�]��Le�J�)�(K~$Eh���4�yU���7�9oe�+{�͖�	�#�47a��ta�J��W;+##+� ��`��t��<�̗�LߔQE��'�PD}A�"��N���p���h�;̀y�*�B��v`�MAE��� �NF���_|��v>�ܹs׮]��޽���?�ꫯ>���m۶mܸ�:�qp��I�J�RI��+�-��5�a�SW�PZQ�V[�f��M��B�ţ���t�6Ѯ]�E�o@��Î63�m��r�{���F��k(��n=޵eCG��w��,�ů.��@3�ݢ���1{-�?[wl��5+���J�9��|gzNѩ�ì��B�a0���2��,�P2�ro�;����|�k��nw7��8�u�o�g���%�im(��렮s�x��o���:��*��!�Q��>�X�L�23�Lq_2 �{i������6w�!�|&���Pˡ�_m{�9sZu:�����0U���M�nAD�{qU�y�{��@����3�֝�|�{��̪�2�� wz�Kz��U�+�5�U��73�3�a���P�1�SS,Z���y |�sUr�#NA�*��B�Yr{�s��3�e���%����䇅�ؑϦ'.O��:����wՙ�gL8�`������`j�x�H�����A�g��_����*��%ص�3���+�Y�D2�V��K�ĤUt��R�Q�����y�K����:�u��.[�OOs��Ca�q�`��-`<c�r�ʁ��'Ntww�������bĲ���$����v�7��5�/H��ũ��\��Z��n�P��e��.5N��W��rE]x��Tb��F�e� f����=�:q��;h�O�K��O�O�6��'��5`��=��ܵqݩ��k�d-UĿ��z�$�B�{Ū��kݫm�z»���G��|G�����'�'{hڗ���3�,3������]�j�����6��q��ܾ�h�}��>�Դ�/���v��)1�`��ԗ'J�W��������r��N�̞�|�6�þ!0���@Q���]� 32H��L�]���㮶��=�7~��gM*Ky"oA�3Ӏy~�H�ls5�%��k��"3{��5W�9�N�,L�+K�**����N�^�N5�&R`��$�V��6��Y�g�n.4F?��� �սi����Ģ����c���g*ҍ����Dg)�;�Ӥ&m[�Af�X�$��,��k��zQ��\<�m����o��?���L�Q;�r�s��s�q�X���� ͜��̀Y`��[.v��������v���L����-~��~�L��Y��9U-��֛/�����;|N�̼��`��y��S73�aX�/��"�]nn.�sv5�p�cbb����(��6��"&�$�ɥR��Yi��i�#~UY�UK�,��t,���r�}ެ���ǧ8���``�����+�*�=�9w�0è����O~o Ļ��`����:ޱ�#������]��J�?(�y�$������w��o{��c{;B�͡�֎��=����0	���p�)Xob$[�RGy�^=�<'�����&�ϯm��(������C\���7<��]X]50�Z,��M���������u����>��n�������gPJT�]��P�V�����ێizM�㕳�^Vu�	�z��sA3��VhfI-}@�V��Ou��@X�̾vX�]e̓�!6i���z����+��3cjRgř��//�rg�5պ���5K���[`f��효/D%���-{��;=c�´M��O�(���DR�vt��?�=v�"+7]���ɒd�C3�M�7�E=-Nz)K��0su��]M�����W���e���CI1�����4�T�����O�����9�Ub*��Uh'��O�"q-tQ`��ׁi�n��]�У/Z�-1V7�pM���h3/vX�lN���J�yҘq6������E�ʇ\�0�7� ��C^�bߘ1c 0�sc��bJ��4�¤�t�DA���V���a�;��,�C��[�آo�V/6�_V;k��TEnC[���P�?l�5#�u��F.���0�A���zg�~���YM�yʷ�c���/������k�U=�~��S���x�v�[�	 �餙/�T�s4���NCm��ick�%�c��.)h|�n�Kp	�6�V���}m��}\��(4S(h!�֠�I�6Ѩm������s<� j �%��t���xi�&���2��f6ۆ�gױ�������n�wxߦ�;�3��P�x�0cj���pa��`�Nm�)?ڮ��
,�zf�6'��B'�KVպ ���5_~�ó��	�,[mHw�����t�&o�cXy��E0e3���L4q�HK>���s�.��K���hfd���)�ԇ-�����U9�7�g�>=���Y�MQ}Z8q���1Q�
'�S��2�J���g)����r�o��Ȍ%z�¿/��ߗ2��E���{<�:w�S}��Qg��ۜv����r48쀹��0f,�3t�0c/(^��EVV�l%���L Y��FJK�+���f���X�����8�N���4��6�ˮ��o���h����\8�� .Ҍ�H~&̌d3M����?�n��8����I^����ٯO�Yu�b�4%n��"��ֽ��3G��Zܝ�N�����1
r�Y�����)6]�I��-Y��=֛��uo춬{���1y�FXr��e���h�a���˚b�d��������z��3����	�}-;��W�9��%0ï�T��Ou���Zێl;���m�#Js��ߒ���n�_�XC�I��I�������-�z��;xZ�R	�[j~��%�A�߼����5�T;���du��-}��;��s�%;_�����p��+��-��;�;FJT䌑g����R�$��/�e�e��3�+����5r�r�+����ɓ�S3T��
�2+sJ��30��m��Q<��fi�vhF�����Of<�u�湕K�MB;�X���uu6
^	�u��������á�x�Aˍz���.�=:bf������ L��ا�%�J9�b��~������
�Qe�-�Y�fc��!���պ4=jG-�%	줙	f>n6o�����o�`QG`���G�6�����\۶[�|댙kv��uwOY;m�Sǿ9)w���GV�W�<s`_���1����a�-�5��Rs9�t�k��B����O=u��'�-�1�ˍZ�A�`R�Z�MG�M��\H���f�;��OW׽�|���|-oi6���s���0�S�`��C:�x�Y���Xg�������[?lڴ���P���4����)�_fH�M��,�F]h�;m�0��ܚf�E�W����uOL�_���矷|��N>�N]RM��1�P2��Aw��%ի��pGρ,C�Ȫ��5Ͽ�s4hD1.W���9f�,k�<sjr��ؤ'��X�)&����).�*6�&U476�,9m�D��P�J3r�
���}\���7�L3��A�ai�I�0�,�k	��p�l�m�"�S�l+����ƌ�妛ai��A����0�L���9��?���`f��.���`�s8��롖̖FR�6�p�8�,�u�s��̥0�a��;����>�q(k73�����/7�E0��l�ut�=�=��׬:XW�kXjX޹dYpI���&ϲ�@}c���?����].4����C�@�������f� 3�����3C٦Օ������E��D3�/�G-p�D6-0N3���Ih�~~�%OШ�g}#�z�2Ӧ/�j9��[ێ�F(�P��u$_����`���<�]��U�������Y�=2�z�S�	�(��nÿ��U`ו������
4��к��q(jt�ڒ��B�^3�5=��|�}c�i*V�wq�:���j��jb��PY0$�M��ӏ�-|}��_�)��n(5��]��~���*x��9Ҭ1��y�T^&N���<'E8K�8;9iV�hvZJYR|yZrAj�]R�h�*W�=VF�\,I�/-8��~�g�T��3S<���O����c��\h<����[����h�7�A���F'��⠸ّ ���Q�o��?�/�
�,��0C�I������?�<ڝB� �iiix4����S�e�Y���V���e;�}�������$��V��{/P֖�G����-&��ٔ��?�C���lI�`ގv_'��li	|��s�����'�<k�k���o������]�u�{����w ��
��=]�($2%����eZg㾏��珪ӌt��괂Ʋ�:M���< #4��h��ZL1Ii`/�_�,T�sڸ���e�[���h�].ב���#��.��q��h�ߍ����-_�hz�6���瞤��Nmt-��^�&���̐���)�b����?���C�\�γ�֝��x�]�+rcI�O��
�=�Q]��P�թcm܉�WZ���iƒ�_��A��]\��oOwq��|�'[��̚;+��j8Ý�Q�-�!�g(%�UN�R�#����ǋ�wI����NHO�(I�;=e�$m�\���T*�Tʜ\Yv�"S���=n/w�}���0#��Ff%�;i�/�������<���b�Ѱ�V����2�e6sMg��r�ر7S�׈;n�O�ߟ�D"�233s֬Y�0�K��H(��D"�b��b6®6��:[]��Vo�YlY����r���MO<m��d��T[f�M���΍3��3kU7�N���a�)�.$�����uw�=��?r��u�x�@k˙�c]�#'��ζp��q@���wu��8�����u)��s�	��L��(a�f���(��\k�&0���,�h��>c��d����`85��7~�z����l�g{w8����`��Ͼ����f_��O����ݭGwo��!��>���g��������:g�>T~��g���MEūj�߾Q�ݻ�]k�����o�z����|"����/_��%0Q'��.���Ć�P�iz�=:�}˲ke����6�yo�ێ���d;�W�4͜��;5�Y��$�9rE�,#G���\�)W��c���d�bE�J9N)ϒ����fg�fd��r�YnN�v�筝\�ۇ6%i�<��lա	�r(`9چ���k���љ�G�s̟i�WR7�̹��i�Z�P�fN���ɷ���?^�9�h8	F5{�|jj*4��3�$AR"L�D�����&�Xz��b�3[۬u����9��:�|u����'J��O�{$Ѥ��Bs�RJ2AM���)�|4��Ͱ_M��c�0�dW[���f���
yz��`xO�����	�?�a�vx�@�;.(dX歁�t��}�N�E�)�5s�u6� ��7Τ�z�&�^�bW';h.@KCel��(@kE��z
&]*��x�e���[�lݧv�����X����v03��f�$��� �����rǗ;��~�˝�}������f��/kQ�a�� �.��,Q�-�U)6�$��=�^C�a���<=��H8�M�ӌ�,��D5�R}��\�}��	�"#�ᔍ&��bo>�=���9�e=�M�:6mt�83C��g��f�$3K��b�R��+Ik�d�$;+mtnJN�0'+e\N�qc�,7�b��}��$CQ,�>v9��90�~ZT��P�m�e.,]�ͬ��jʲ�f>X_]Sgv,�s���l���,�|� �0�D53|��&��vJJ
���v�/O�Q4�Y!Kҍ5�v�	��lO8�Օss�)�h�0\��B�4�Ӱ��R����M�i�0e��b7�� ����l��vX�4Ƴ��tw�|]�m��`�"��>r{Z��[<�����z�B��@�t��3���	u ����$M᯦2-��C�zW$�-[u����K�%̿����G@9�+4���B�]_?�]b��ն�G����H�fR�s�+�_IK`��2�:T39���/��^���#_��6���^"}�
�̠��|fo��d���lX�l~X;����l��z�hL�C���?��M�Ε�f�����)�L�,K*ϔ�\�����*C�R)�Pؙ��^�����KƎ�����]���;�����f,%�8"\a�4�e�%�-oF��{�^�48�%��P���[�3�l��ؤ��d�Y�O��t�<��!P�H�3��HX�~ޠ���oOBo�(U�_ W�f7��
��*3S��Ds	�og�w���tS����8U�S�Ɔ�=31��@A?IKS@w����7�(���5l�66��o~�W2 �c%�����l��Q���+���Y��P�l ��PѸvE�r��Z�ۛL\�ιXb/�T?��۟�{�͗6}����CAOˑ��^��i��f3�[�^�Q�����q�؁V��#�Ұm_�O7��t����ʝz���Z�*e���[2�Cž�٭�k�a�_<6�Cyf��@��%�8RYC+e�%�3E��7��-��yE걲\�^�,���P)���K�ժ�E&l�x�<C7I�Daʢ"qUI��g	��7��0����:\���`����)��|b���F��an�oȒ+oq��o���?����a���Ç GGG�s�=���ǎkkkknnv�\---Ǐ�멧��dfϞ���X���i)�b�.��'�5:˖6�w֌���:��ـ'�g?��K$RW���3�%�)���=�vX����� '�5��7�)lx���f~Ko�0���]f
���e8l��+*�ndd�3�i ��/|wI�뷾��m~��������p7Z��!���(��C��;-�փ���>�n=�t��!�����g_o�������\��/��4���C�qm��Y03]����P�١��ĺI�<����c�]��<l�Cg�A�o�҇c͚TKYVm�����I��ƨ&�˞8n��	�&dO�����(?y�l|�lZ��u����ZM�����ߪ�����k��P��#��i�w�Ĺ5OXlF��1&;�6�4�0߀f�]VV��W_������;t�О={����=������ׇVy�ܹ�~8��u�$����"��222�&,x�I��0�u��ʪ*�u�v�BԌ����J��7���(�0�!�鋶�)i�/�ڂho��E�iC���3l� v��~�$�L!�a�����%_T����m\_�k+6�����������hok�t�u{�'��`l����>r��j;��v�_}���_n�p���ז�o�>W�jcN7�"�.+��7��a��Őf�KF&~���_�?d��W��ӌ%�8��;3��d[y��4���nr��h�2ut��:���9iV~��s�p�����q�d͸�y%����]źg"0�Ljz�8��K�f��b���Q�����?�����������W����l�e(gX�P����u�����J�����NF��[�n��!q4�M<x��d8�I��N�4m�D�8�|�7�z��8���P�������o$���H!�{F4/�;;/l�p8?���U`F� ��3���*ӌ�=����__��ݗ�|�sǗۛ[C'�-��=-�������փ��s�A~��΀�����o�z��[߯y�z����b��6�Qc��v�/|+�03!��Q�1�D�P�+#y&�2!��B��[�� �;����8S5�D�'��dI�r3$����Le.$C���*�B��Ks��q�	3&f��VT�W�}�ϝz}�Fq-�9�z~�@�+%�#���%���:�_G��������~���n�{�ow���Y����`���İϕG�����rrr^x�6��ɓ�O�0[���nח@�(%��sR�L"��̄��R��i)���8Ebf�6�ZJ��P!��ȽZKL"5T�3�J�G�d���e���m��>W�CsP�"���i�{:i�J������ �NCAi3;�ayF5� 0�HL��o�m�N��g�c�E�m�pݧ���#{[�-� }	nC�ֶ�áv����ñ}�>ߴuצ�l_��S�ny�˝~��S��\d�o3Sό��N�[�π�a̓L�3$���x,�C�������|��|=\���x�:�nR�Xib���l��͒gd�Bo�p�Ǩ�r�L���+���c�,i���g����{����Zu�C�(���)<��"g��a�� �ʢ���Y@��܌t��3�0`���?f�L�e���P(���e˖��~4C `2��Rizz:�z�w��nם��Q<$<
�T.ÃO�� �I�i�5e�V-]�S-t&�)��"REZQ�a�y|f�L�#�+d�P*��\X��c�H:��P�?�O�LK(d`L����q��ך�b�0C"3M+���ԦY������U�c\��~O�;�_j|u�[�|�퓯��ߵ�~�o��}�s�N��䋍�wo[��%+�r���U����b�S8��Y�w�����.���7ן��!�aC��G��2`��|q{�����1s����jMs��,�?c��≒q�dezZ�\66S��TeʳU$�D��_����͔�ɐ��P=��,Y�Y�8yf�T�K��\߇�7Q@?����(�H]0�e2a?�K�l�uf�̱#�_>0�ͤ����;s��Ѓ�Æv/�4�|��c��s����h��Ux��$����X�f�D&�˥
�D�H�J�
`�D����8�t���%�4VQ7sX-�@S
#��I1x������j�nk���>���_J-�-�<;<m����N3�l(�]�4J䗀����\o�G�H6���*��壛��D��+>}o�RS���eo��܇+_���[_�f��M�bzyq����￼�T��<_N}�Ix�4&\O�P�lE��<<R#'��-�Y0c� �P�
�99�G�H��Ҿ�hc�[�n��؞e�1̾s}��L�N(Ҕ���`,Q�g+�c���ie)�e)��)�)c))cŉ���*�J�.�T��d��q��'L{�?�n��F����ݚ�/�Xs��?�HbciT���F�9)��M#n�����ɉ���3#�0��j��g�@����y饗-ZTYY	�,XP[[�裏VTT̛7/��pR�����AZJ�\No�3�H��tie	�xb�.ʖ��8��Ǆ\A"���ŭ����~��`F���p  ����q�?z���g8x���'��>�����N����}�}��
�܀0�� >�/����l���{&���)F��\�^U2���߼��9���?�umj�����o~���m�q`�z�wχ|\3׳b����ŵ�"K)���/C���X��gq�iZ���l�0_#:'!g�L��@fv�6kQ� M7j�k��eB#�(�U-]�@�2On/O�鐗YJ�j��b�N霉�*KYJu!��"ZJ�՚�����y鸜�lE�S�T*
�;E��NiE�3ҒJ���gJD%)��)q%Raqz�]i���G�U��)ͦ-X�]<#Pl�٣x��(V#T��������s�c�����&�3�|f2�I/_f��a���˗/G�c�X�Xb�]TT���Fo�q:�l><�L,I��$��"�iF��(֩�kP��N�tRtNfa�f���DU`�HK��y=LõH�h~Vޮfnt������k�9������^?����/��|��Ы/u��b׫/��Zٲ�Ў�g=��OO�a>s�/��D ��RH#O�r�`"1��k���R�~F�3U����<��V���Ǿ?�������O��|������f��ҋ�Z��^m+����NgQ\M�.�%�A^r�kn��`��ِxS��~��ݯ��<_r-�.�s�;8�S�Mb�&լ)z�rײ�ysJE��V�k��n��}J8��h�k�7�I�W\���^�}���`;�6��eG�u��8�ђ��\y�h��/K/OK}P��� f� ��;���s� z� �qa�é��$%j�)S%�Ѱ�����S���b_����G`ƅ08|Q�0GY
ج `c�v��V�^�8s<�����l�|��Hr�7��`ff�ĉ�̙�Y��͚5��3g��� SZZ�<Rqq�X�q|l@a�@�.�fN�J`��D?*ɝ�$I��*�ic�����γʇ��(��_f����P�p�)�};��Jf��|性���X��;۞�E�P�ɻ��X�f�"W���k��j[��y������~��N'������a�1D����APU�5VS"1�I�3ҫu5�F�̙R}�}����/�?�X=�>oₙ�kh^{Ü�*�Р�2G�i��F7���85��$ɐ�Fp^z�kn�Ohf�����B�F`(�����^i��j׽l���>[��EP�'���=7���m�z�/~8�F;�0��;�}N�+�]2w��:���޴=�����ۿM�*�K��iݡ�'̙ٹ��12U�Bvwz�#�BS�`�8��tM�b�R��\��B�"C�L&]'�?AT,��le�B�!�Θ���B�*jx���h]��0C�^^(�v�[Y0@5���q����c'N�����f��b(̃�Fn���XBy�����k{�d_D"φ|���?A�c��D�͆fVef�5%��7g֜�l�$emy"��9MZ0X9����pm��0S|\����:�H9�C޶3mǂ��{�n�+Z����/�V7~}����r��L۳���5��:����"����o����W�W-i�	�Ca�-�dk��6;�ZJ| 7@ȿ��[�w�����>�X'�3��{��-����W���J�f�-��E;4#�4��N�t<FE��h�����~���Ei�28���"�.�ăoڥF���(�Z�j�jWT�q'��5?��9��)�e�y�f�)MO�aK��,�J3f���O����̠M�hFY�Sj5G·5�,�"���)O�
�b�Vg�>�k��y��L�U0񫂻�.��h�xKB�#�i�re�*[��-�Κ��~���Yd��V�_��`�Е����h���FvUi�}yO�7حv�TI�vo���K`-�	7sBB�p��\�K�y��;g���#G�d{]��L����,�J3��{�1�#0�=���Ή����ap����B��Hh)� ~V�т��/��b߷{y��݀�v��A�`�@��u��ڱ�㮦�>��&S��f�ڙ�/��\6��Yw};[}̰���kg��y����`��<��)���EFm��,�9�i��o��V��g�C��z�gV,s<����Rd,�5<��+ۏ�vq�����/U'JӜ����-����Q��0��+�V�	��fC���v]���`6���z�/V$.��@S[j�K^��q��o,��󎫙Q`��8wr�;6�sVZEa�e���@a*ͪ�N�,]��߈kKbM����2����"c�h �-�Ε�2T�����LQ#��W�M��l��I�h��(���#���w��
SӒ����lhus/?�EV�^=�&�w��ui��gƂDSa��8��թ�BIea�����G�78�&0�P)G�D�`w��f���^MA�FGG3��mjj*t)�X�^,�O,KF�RB�����0�e2�R�1���κ�uΚ:�ݖ�D��c/���,3���%�֒>\6<CV.���H�݈����`�h�5Բ���&H�<�wK��������?�AN���1��=c��r�.g��y�f��,��~��{;\��}�N�r�����a���Ck�[�U5��/���9�zq���W���z�o�o�j�'[�m�t�/v��l��_���O_���K��>^�i���\難�fT��ר��v-,��zM\]ɰ��[p5��jgҌ��.��]�x[Ij��;�ᦗ(L�B㽀y���R*0��%i����-�q��[?�u�{qi���s|ؐZ],YP0�vςM�,��B���j?yf����]�	��.��	w������R�䙲I��y�I樑M��Ū�5%9o�r�,�\W2��ce�J&���| )�.qr�B����23���a_˥5R��Ц�4h��&�̠��J�:�Z3�jV��V���`�4��+3Tp�/�9E@#�n f$ ���/G�������������AaaaGGǴi���\_��O���Ix
�a�ɕr�rѓ��F�ݾ����BQMKɪ4��E0aR����dcS��!"�z���/��)��P��s�����l��n>�:Z����֎�]��j��5]�k�:M�\^�Y�]�������:��� ����_�n��:9�V=�9ws�.��K�r���������Ѷݟ�>�g���Zێ���cۚ;����}�}���v}��zh��5��=�}h�m��^����q���D�/=�Յo�W�9}^�ǿ�ɝ�����`�sh��Ţ�2�����ǸβՆd+�e[o,Q��p��1<�d���_O����s�)��c*�ko���������}tz�;�ϡ��E�u��,�R�/�\S9��L�*[�Rɲ�	�u���S�)c�Ҏy�|����~x�dkɸ��??"��&N�RH32���L)3\���'��7���gWh�h��ڼ}a��X�/�W*+
����ViXR�ʪ��l�Z�u�ͷ�|�-��N#�~����֬Y�v�v��7�x������֯_����y��a�9s������	1�qP�)i��t�����R��Zg��~������ܚ�܅�q�r��O4�@&��DD�c'.��ކ3H��������/����a�{ZNz�|Թ�i턱O)D��e�R���,�#m����P{k���W:���x�!9�3�W���nXK��E��-�����:l|����nٹi��_�ڎ�|n��5��}mm����v�=��.o�#��}����[�غ�奛��h�:^a�0�
j��i��Nz�-����?�3�(KQr�(}~JMQ�}.�a�k5�]��(�nF�EW@>�i��Ɇ9G��O��;���zͤ���,P�~ݴ睌Z��V�^U���j�:�8�����a�zf)`~2>�Eq���G�Y����`�\2�裺�ډ�1y,%aZ�0K!�� �0�������a+�%�jc�0���/j0�n+�4W����+������y�iC�rk���饋�&X�cǎ�ǎ�
3�of�
[z�ʕ�ƹ���	�Y(�in޼�6����`�4���u�	0� 8Nzz�\����Pkl��/u�덆�g�y�6�����,�<mz�i���*�-yXn-K2������e�7Vc����8������|;�hW�������X��O�L�D"xmZ��ѯ�d}\������35ǫ*ܫ^=s� lhf
�ľ�'�/����i����٥1��]2[���\�4��ozr?ױ5���yǺ]>�rG��C���W[��-�n�� ����$g���Aa�]ǿٽk��_{��v}��z*�>�a��/�	t�q=��0���~2n6l 洵Tf*�`���~q��\&6iŶ2 9��E���)�*�W߶����;9��Ū
M�q��ݻ~ 7� �z��J�$9h��cQNm)`�p�lvnE�V)(2_�d�Lx_B�9>�E�荜�7�*�(�z� �����f�^2����D�S��ivrEv�tt���;����PV�`�$Y4�#XH3��c�4�$�h�K-��yq]u����i�sZ,d`�,V��6a��[�}��0�A<R�@H>�0�������^��=f�
0Cè޴i��'�|���V&���@��*SH�J��f�;��R�068j�MNH�bGu��f������j-?�� 0o��G�A�6���?`fC�@r��<�����cb���t���}���N��z���i�w��>�"_?)����j����5��=��d��Gc�]m�(��n����(
����9�L$f�����8��wA����G�ɦ�DKA�⒑΂xSA��줛uS-|s���A󋍛�������4��'�g�h��[|�6������U�������!����{����ֆ�Wn{�����P%6R�5��s��NK���q9c��穉O%��|A�r�z��b�T�Le�����:y����ZQE��V>�Պ/���/.Wi����u��'W�K�,P�����vɁ2j��
�da�ԤM5kby(�ȡ�T�B�̹crd*�%���ʂf���OZ��W��og�ߘ���.ժI���ek'f�?>�6f�#)��baN�\�T*2�ҳU㊧vrkl�T�a;���g�ꂏ@@u���<�馲��G,1[�lp)�ڛ�F������8749����y(̃�9of�b,Y|�}�j*66����ر$�gƲ��
�?���l��L��;!>9!�\.�(�F�$[�V��N������h}��Q�BUM)?��ˢf0�����1�Z`�WS�
��h�E����-�վ�>����<O?�e�̷��}P4���c6L�u�uwMX�U^����5�?|w�C_�;�F�t�{�����fF�%m�-]�9֜��L�
y%L '4�4K����{ޝN�T5Ŧ�J�5�����N�,�m�j�7����Z[�!kw�����}'O�t���*]�㰴�W���:�妱� x��G߿s���������m�JD���?e�{ Cz�\3
��`�u
��
kY���纎p'�r'������5��T�T_R�҂o��+���U�m��&y��FU�7���o��A��NBc�z�oݨl�9J?�	m�z�s�;�5:W�T�&���̑K���NU�	�Ɖ^H=�,\���D(X��$1�1U�DL̜��	i�rY�2K����ΚR8�׿fߦ�u�]_��g�uQ-���'7���h4:��F�u����\������VGCC�4;�a��9f���'�[��^x/''kpX �s��� �ԾP��O�;w�43x����ib�-�X,&>���i�4�m���&����ش��\gz���]�`f��z�/��6\��|4����@B�|>�/�9Hf8!�k���5�7�=��zI���cq�%KC�M�%�=�����t���.����������N>nv��� 3�-�i�2��B.Jt'�i��8[A�-��֢h�c��B��MB���VMJUQ��g\��%�ز��m��s�������n9uz�r���3}'��C��3�I���\6Xfl���km;�;/>��S�+M���+G��+�)��i�E�#�O9�dO%�ς���jE5�S�z���yǹ�%�>Y���/.��ҤpJ����5�5ř������|�0~�CJ��f�T]�n����k��f}�{���j���4�V}�|��sgY���1ي��t��R�*����(VX-X� �d^\��1�$	f$%��ǦK2��1��*EFff攼�O�`xF�Pldu�Sþ�f�`�E�F`Y��Zb�o�5YmK)pe]]�)-"�v��#n�)�3�0��ȫV�Bۛ0aw��tu+�����^��޻w����D�$�X�,�I�fS�þ��9:,��V��	b����-�5.£-�J�9�Nf643
0ff6_u3�pa&���G��I�a�hAl
�(P����:vn?�c{��Oz7n8�񺾏�]�dc���>�ܰ���ç]�N7Tz{ ��`D�=]����D��s�e��ǵ(ƒGs��l��>r�_�k���X�Kl	�	��=�R�`,g�w�9�������J�e��-���{��(���(4�@�)�����3]�A��J����f�d1��בP�_���ۺr	3�����:i�%`������O�o����tB�`�F�9�RL%��y�d#�)M0G���˱%6H�&�䧛�b�.�&+���e*I�*�T��T���f/�ïy��ԅ�ܻ��i��r���̬�J��rYIj�.Y�N�
�ŢiJ�$yzz�d�d�\>F���d�Q�U0��K������ 3SX�$sQ�]���9�r.��wl�WM7�;I�e���0�f#Z}����4;)H��f�w�Q��"`p����2��P(%%lCc=u�K�O����o��a%z;�H����������F��^�9��v<�uVx�&k�r��%4�_��$>�C�\44�ȣ����`�{1������z�M����}A߉��[�O���nk�k9�w�ع���-m}�m'[�'|��.o����ti���w�)]�a>Q>��X��*���x�i�D��T����C�x���� ��,���Bc!�kʸ�Ew��|��/�~wd�'��=�l>z�3��з��';���2��	u��T�خc�]{��5��
�gK��]{>}���w�ǽ+����W�'������{~�z�0�:`�F�iDKg�2�5̠c�a��:'4��i)���W���R�=_DEgqt��4C)�Bg)�X����*�ױ��Jci���>������q�EJ�,#[�=Z:])W(%�e����Rq�\���T�,�4S)Q*�J�ev�,�KT*���Gz����oH7�� ��ܹ�|E���������<S�h����P�dz�ɸp����fl$�	0��M���r0�# ihN`��	�k�|JXXBc��)��T� ���Ke6��fҲ��uVs�����r��r�i�S��V�,y2�`�����H��:��^"�U �f�>3x��^$ԡ�����؏PH���y�':����n����P���cM_Vth�f H�z�t�B/��{N�S�	�[퓂�֑��[7-'T��.�ЬKbb�Ě��4�M�A-�������9����U������m�
ć9�t?MK�<-����+�? ����@� f�g0mL]b��@��`�����o>ݸk�s���NOX� S3	F��zf1:�L�_f<��4�������<F?�,X�������-�ba�~*4�0�a���^�7gaTCɝ��Q��"�[�����%q��,C���^n���A����I���LYn�8C����d�����Pe��J�lY�B�R��ʌ�
z��Yr��ѳlo<�͝~�M�C��x�o���\N�d�Q��X 1j&���e�s�ុ�sǛ������Օ���z{}=Lml�||��z�&̴;� y`�9555����HP�Í4���ӤT�4]b0�Zlf�b��cMz��i5�N5�;�|���iֹs��;����R_�8�|c
���a�{��C�??(���I�&��=@F3�m�o?��Q�A���v{)�6~RL����<f�;��E��$fXڀ9�6GP_� ��p�Y�2�D"����I&m���I��E+s΀	�Z[��/����G�nǪe��ڶ��^o�������@�fX�,ή��6�l�|����3�fl���i��`��.ב_mmX������b"M�D#䓝Z6����D�f�3�l�� N w��4�W�X$��K�f�<?��skAb���i��x@7�8 �JcS��j/E+�5��z;����G�j椖�7N����\Ϣ�_Y*U&M\��&Τx`�ʜ��L�"3#S�!�ʈ���3=wA�s�+!���̺(2�'3�["0� tE�"�px����4����O4�6�l��T
%H
3�������5B)����%�	T#��;=܄�D`���kk�V����cF�ц��
u�^#����Kd�*SY���&@���4�:��f��B5����`�
mQ�>w��f3�P�@7������}!��u���7H�yG������4�����As{<n҇P�='ث�A�)���~�����+�3�~��U���4��k3W�f�f���R���l��앚��5j�n�Z��Wq=��wmns7� ��E�������"��*h� �d����	��?p�4v�����n�ث����7��c��7ַ|�z�W��t��~�!/��f�c�^"���A���.�\L���oz����_�?���f6����p����bQؠ�������)Ʋ�ڙ�9�� ��P!e)2��ʇ�*S&��2��܌��t�DU��%�rph��B7���^�8.ڡ�Ӯ���W�9f�5#_x*	��	W�����y���N��l��� �o�����D�+��x҂�L�[���S��yyyZ�ˢ�",5MAA���ӱh�v�)!��%&� s�\Y�h���V�4.Xf��!5��!�q���`����|~R.V'춆��E��������vA�80l��Am�V�'��0���������sux<���m���wx������I��K^2�w�4d�e6�n��Q����!��w����N�=\_��ws}�$�\���UV�S�Ũ�����e�S��ܾ{'l�p+�r��^;�d(硚����|�4�ŏ��S|3x����zX�_��bӷ��_��襅�-��p�A��ll�F���?��0���[@f�%?����0ӎ�{<�P�r��N�n��dզV�]�_29+��=���ƅA#gɕ92�e&oU�R�+��We̾[Z[&0ka5-X���;��W�eU�giLC)?�c�9FZ'���1��B3�HEU�K9jmv������L v343�,���_f6|�� [yyyoo/�}�̳pb1	X��n��N�J>Y���,IMS�%��=am�:��ϵ�SU�8�<<���A���VV0�X`uŪ��_KÆy����5��&��f�M_%�S�����Pk �}���§X7�~��c�l�������7����Ll��ʫ�hQ�Y��)y���~.T��S5랶}���;?�����j���g-�^2����С ם�/����i�2ռ��>��=�̞֐�-�:�`�3a���H�ԂF�0n�4=?E���(ml�{��u�l��0/�:�}����\����=�@?)��a:Z9d` 	��� s�;1z�}�v-ܕ��3�1V�5.+klN��ѐ�qLr���@U��de�f�b�j��r�L��4�>�������>ٽIY�Z��.��l�����m4|���a��#F�/M�1yꌢ���hޓ2i:�|[X3S�{������3��u���&}�e��f3��uuuV���7��`>��u'A,��q)�ir�茬�9�?�HU͢�pҬ<�|����R\2}��:��G�**���Ї3@e��'E!B~&|��@�7����B~hi'�Ӵ4,P>���;p����O )�gwW���c��җ�p�jyE����w�_;3��H���� w���
�B
�U����� דi�%�ÁTK٘������Ձ��Rw`��Ϳm:���d���|fڒw������?��f�=K�V�[&�L}RT��H5�vDX[�௿��fGn9v���?�����0���돽��7&��	S�����N��8罩�R�Q>4Uv�J�Q"Q�$*�8C���H͒�e�ę�L8�p��d��|�DV���x��R�n�5�ç������2�H0�b��N�l�qU�/�e��Ek�G�~Ŀ��m�r�-0�i�ȭ7��(%������_���3f�(V���E��쫩�{z�����wF�f��bD��4[��D٪�4=+[)#ͬ,Í���A[a�%�]x����b�u�`��뙏L@0���C>�b�"�����p><8�������y	�*h펐��N{?���]83��� �0�il6t��Tn/�-*�����������Nd/�����s�xCY3Sb�)]�^�� �+^�/�k���k'�g�ݳe���}ԏ{|2�/����&�`0����,m8������fϑ��8��/�eԗN]٨a�����Ϭ�2aw�ݔ�s�@�C3a+�[n�����'��l�ȟ�^��h�|�?���Os<�Q[�xh�p�L�!����X�|�B?�5�L���f+����daa���٢R��W���~ؑn*���c�T
;/�v�S��Ul�Q��S|]PL�v��/�gf0c�353`�h{�'O��F���QQQ�+������?����L^@B��D�P*�Ueg�e9��Y������c�-0'��4�A��Q3LXEE�����EIft�Ka���ϛ��.�)�m3�wz��I]�Al������h�`�{`a���ۃ�N/�w��	�9������a��L`�$��+�J�w���g��J��j�}����*��Y\�ɪ-���N��r�&�P Z2;�\2z���wd0SLl�����f�/2$q�`fk.����O���@������Z:9ɦ�0�c��ѝz~�������G�m�`���Z��f���#C9�����(9�-���v�73kf}kf�����5\�+� 9�HdI�EřY �cQ2g��ٲeɖ,��,f[���"1����8Y咮�+�����bm�"�"#O�8���>��A[���6�<�8��Ĝ��JAj���L�)TJ�21�_pJ�"/Z�P�R�h�s�^�D�����MK�,ǹsm3�t����:̩�q�D[(.4~�%����xv��g�k~�.�'�0����{��(aB�����իW?{�,--ܲm��8 ��㲉'�p�;�}�76�D�8`N���d�3����JMT�
����4؈��bo��;�xY,�:ܢךh�`�
y���`�(B�|��`��7n�������z�x�z��{�6�<��=hl����mj�"�Ul��|�S}�.�̄�!E<�7�G
˰0�:ʥ���l,��_u���W5CQ�I-�n�|���C����Ӿ��3��rm��N�؇E��Cm��%�Nw��)jߢe��A�<��$�`�I�k��2��LxO� E}�si���#�̌+��d5eC'#�������[�RJ�M�kz#�I�13�y�;tX�UE��	c���eb5��Пxr�+R�����{��a������Rԫ'����0���*htt3J�
:��,94-�yB�"%��U�;��?�O0P�>�3+�4�W>/����SE�o���B��L0���^�9R��03[���l���=�ek�/��f~����5E�#i�cXB�P.�VC�B&�I�
�B�S_��p�S�-+̞�h��3����������gΛ��(7��Q4?��oz��<-M^�R�W��ݮ��s���CGn��{��;����K�����{��=��&4vS fwc���Zo��l��0�q���a=����Jss�<õ4r��߾Z�5���v���Q�������K�����ņ\�������G,?�����>=h��+o�3H��_��,pOx�G��v]�}����P�+�M���g.pO�f��j0L�ȭ�v4����؎�����9D��&�0�1�0��E����(�:܆�Ь.����˘��7؇`֫�?�q��R�	���d�L.��$�z�}�����!	���ҁ"����%��Ri_�"�(��R�S��e��ԔD�|hA
�7�il6*9�5+�L+���;g
;~��P-��ω�a����?���{�@A�� M�<�T��nL�Ι3��={���?|�0�ǎ;t�Б#Gp|���K�.�|���l�'!F ����EJ�
<˥p7A��O�P��Q�{س�0�3$,[�/e�L����0���L�ZC0�O4���[-�ͭ-��Μ�o�T7qp���ŋ!-�2i^��a�
��=7.]����D���tz���ߐ�v3��Pqv
,)*�T9qM���j:����>����g�֋���p�`�Qh�L4f��%}�~6r�޾q�3�fX�D�����.��3c�`���3����Oͭ&��z��<����QUE�L�Z�a�y���uJ�"����‮�E�;n����?�7~��93��=s}�n��)���^UW�%1i{9GM��1|�>B��&���|eY�	fu�9g��IӾq�m�(�P>�+��/�=M	�4%^�}����se�^*eZ/i/�J	U��(��0!*zjx��ݧ�DM����1.��'�a�$q�g7)5I����HN��f?�~f-`-4�'ǳ���h��u��G��N�jLL��u�Ot��i�)������{�D���?G	��0&6{A�����ڄ��ݻ��s�nݺ���͛ط����۷o�#�[�n���̰���b�<�\��&N���''��
��/����ponw[f�='��,��4f�j�g����Ca`*TwT�($�;��	>6�[�`j���Z��͍��v4-Zt}ZQ�ԙuE�5�3�̘�X:50kJ`������W.�������l�A#,�Q2�ܓ$�(�&�ށ�Fy`��"Փ�����	�@.���{�^�n�Xd�}|_m�5����_�5�����Sb��_�����g��$p�V��Sw��������9t����W�p�㺴)�"E�X��K���Ы��YU���7���Mt�ϩ�}�k�s���G׸�W�{���*�â��./�rN>���G�d�ag���v̎�QX)��oj��ܭF�?���[�f��ݒ!1�^����{��3-E��[҇��K.-%N��2�w��j��o����������Gw��t���R|UZ�<5Y�S���Q���܃�?��aVǚP�Oς��:�;`f3ݐ�EMF���G�ì�����;�����_��_�������w@���̑B! ��GG	���7X��911lH6�w��Fn����pW��0�,��c���8A�JL��Qև��X8@�����gE��a��_?�t���CQ'���3kA�0�� f-�Hs-(l�3?���9@]P���&ϝ`m�����s�'��C��������xf�K��L�ռ��<���MAz�@��
�Y���#�H��*�(l�A{$Ғ��]\�V/�y��c�|��S����f�<gO-�-�m������`n�Ap�;�L07��7���k|��>��?8}h��%>���`�A2#�Q͎_��7`�A���ؓ�[�./�d�z���6T)J4�`Pe
KA����m���Re��铫܃��:��0ڔiʐX�	eY"]��(k�[�<��z1��r%e�5�}��I�i�s�UI�d�&t����mRv���20m�G=w껳�bC�L1R �/��Iɽd��ĞI}Ճ�q6]܅��ERK,r�y���fօƛ�T+�:'�D--͋�a~�S��m�A����T4��10�����X3c��Of ������p �.c_y��DD�p�r�"��c'8��2}q�dZ�9ƘU�ף<;ڙ-�e�[�_�*蠩l+���F�@'w�̔3��7��Fzu��?C�LAh�羷�ƾmN��>}�蹥�-�?�nd���{�1�JANsi�oݚ�W/�@3C��i�f���v;�̺NYyw��[�T|lU�v׭K۪���b��3G��_��|޺[-��~���"���!�y��y����|�V{�P���X�{swu7�Q@=/�: ����4�zk�.�y�#X�;^�PZ��Z��S/,�1��gA̬���5���[/m��L��I׏�����7D	@a���Z��2�߲��¢�D���J�S�����JV�JNR�TIltl�1��U��A�GF:X�������d:�>&6��\"Q(SR�HU!��p������"s�ó9���Zx w���J9�Ȃ�L7�K�nX������*{�ӑ*�����v2�ccb�1Q��MHH ����ݻw���l� �ѣ���3���9Y�+I�**��t��y.w弊	����]vk��PG�,4b#��=�2k�D��3_�I~��/��ss����C#B���7\��w���9[z�U����n(L�X��Q�:9>��(u}�4�k�\��DC���qZ<�&Z��!0�aF��pf�Q�siИ.GV���}Q#��h����ÇN�o�hj��
������R���3�^���v�$ ��f⭻z�f�R�0�]+�6<nYvrK|Yh�+J/@��,�߀�okf`�Ւ�j[P1,�4;�6��{8l�Yh���ۮ���^0����y�Q�mr��3�;b֐hS��|��8��!�W�6uz�ֆc^�[�ʆF���I�O�Ӥ^_��&OJ�'+���?��û-E/QE��L٘��mF�ެ��c5Gr>���ild_y�D!OK���蜃r�6_ح��l��둦4SAd�{s�+�điO�pf��2��U�����6�4�e��V[�T�.��J0c(ώ�8��y��)a�ڿ�ѣG�1b���|�I!��c~~�رcq��u>�ֆ�&F!���r�X�P4i��j1�L�f[�Q�9>3�8�ȡ��-9��H3���DQ�q�� ��(��׌4B0St�`��S�f��h�yo|O����������@�>]�!G�)O�9?����?ͭ�ͨ_��V��`���45�(�X�;�_f�R����[�fXgȍ8C�Ġ�iy�q���G�+f:{����禠�����<ꋂ��0�y�yM����ۀ* ~����;��p��/�l��n����Pˬ�b0C?�%�s(n��Q���3�NWο�,ڏ���G9+K���(w>xN�h�ˋ<�=m����K_�:�l|�{0b�El/�;o��_[v�k8���p���m��LQՈH]FJ�������W�ԋ$9M���/M�(�"�H�sd_�}=��M�}��?��P��c�"?P$Ȓ�1�RȒ�)�2�<��*��j�U�Ö�ͩ�x
<r���jb�cmY0���pY<7�>Gc����T8�N[�˝�PR��{�2�Cq9ۧ[@O���`6lسg��H����c߱=~����ק�����jMf���G
���II�$��TT\&�<�'�>2"ө�9|�:^�-0R�w�<X� �4�
e��Y;3
��
N�3�M��-���� �{^_}k��ەs���=_�}�`�,�7ٲ�ڤ�3/��^/�
�y��f�3��a���`f<�[�a��zL�<������=����b������xж�<�������`楃d�e3��7���G��}���%vw׵{%�? a�d�H��W�0��f}[s��Z��䨿�kr���YF�s�יb����m�\��N_��f�`�jA����3��G}e�7kbMԜ�o�Y�/��g����7li<&��E;4=��\�������~2UIR�v���c�=��ˢ�kzo��`}f���W���|X�����)�U�rX"MNJJ�1�'�Ɏs���.�߆����3"�����g���Y�5��4�$1~�6��Qn�U�,6��3��M��������Q��i�f|~M�a9C�/\��nΜ93f�0�M�2����h4Μ9��󡯽چĄ	���	fQ<M�KͳJ]FS���t�tn�h�DM���Q��OG�}�f��R�PX��c�!b� Q�P�k���LA�:�Lv2��k[ ��k����PӶ}k����Y �f�򻜴M��m�'�d_;���f��+��]�4��z����b1�^��Qy�s�=+ŷ'ì�1f'Z�:�+{x?װ��.��5�W	�z2�;K�<�4��FTX0@��]>����Y�~
��#H�eïa �Z�g�0�AX�~���K����#\����9��z�ǦO s�J]�����K�|�b�u�n�u��Y�W��5�A��٦
�ԡ~	i3-��*R�:���Kq:R�kE����&���W�J#�����I�s�+%��%ћrzS�����y^�R�7��.���">��R�9M�S��28#��/�L�gDHP^e�`��sg͚g(�җUt�FC��Zn��- ���f��O߷�}0��0�`R�Ttxl$��ׅ6��U�V=}�455`3s'�B3����}�
槯7;L����5h
�T�2Zf�]n��f2V�;lN���j���f�f��MY�ϭ���D���gM ��@Q�0���!����`��o_��������n���@��-[7`����$��� ��c�Ɓi��d����u�\����s����t�Ks&��̯kf� 3뭤{v�i���:܄JM-�i��9�L��\w�Nx��Ȏ'^���<
�H�~r�ކZ�1f074�!����9ul��}���v{���q�{��J+"���̨F%��8H#�o�3�� ���xx�hL�����?Yc������1����_�\�����U�Wyp]�O�~�����	&M�Ui����g�M��Ͳ��޹�hT�:�B�F^��y؂7��3M�Lc6�
�R�8D?!�Gy���	����o?T~�ls?��~�S�d~d��mr��BLR�\*��
��|�5�l���I�yp׻۲���ި��f�iA�4���ԅ������p�m6����,UN7�3x���h�������P��3nzY�]x�`����O8�q&L��;6�	�����Q1R�L!Sb����n�HH.��;lV�Ֆ�Ң�mS>-Y��S���$5E��/:d�@p��D���03�)��	c3��V��f��Nõ��O�Wn6r]�>���ٔ��u�ԯ>콶w��3�������'�O]��@��`K��w��F/K«��$�t���|�T�!��D�ǕNr�cw�ǹfm�~��{N�x,��h�zj���6���o�Ֆ ��4�4фϹ����<��䁉�ң7�_�nf-�)��ٵ�7T&_M�7�0��`tƩ�^���������_{����Ҷ�}K�ז�bNy��M?��2g��D=�9��������F�|�j��#KJN����n�������E��n��hSf�^�yL�Ӥ�N�+e)JE�eZ�h@|�T��<&v�(��d��>����뾊/Sd��Tw�6!>�#Q\
��$�4-5�WJ�ܡ������QX�S�"��1sc,p5��M�k�Uؠ�*��6W� 6@ɿ���֟a�۷/�������H:�l�hfl���,:g�>}��A2�0��1���q��� ;���xal� 2V."�����4��r8��\�lsX�.x�;u�m�S��q9��E�Ø�B1 �du�1��v�0�A2!݄�Ne�%��s�������V���r��e+�\q�σ+��X���7[o:���ll�A��C�ݽ��`L��xfV��W�.y�1����}\{�~��f˪�]'��ڿ����o-���`#�@c흛0:j=55�׏�=v�����,ڴf�<�۵�9��ʉP$����ڎļ� ���0sF�K�?���9��,8�ys�%��e��%?�����gЈ��UwyZ7z[�1*{��MǸ��?�1�?p��w.�n��τ�X�//�jx��{�ү�4I�R�{&)R�$�������"�ᑖ�]d���/
��Y���(	�F��L��/�%)�J%'�}��3w�C���ӻeZ�L�S)(X=�-4.t�U-2�t��0�TVi3���
��{�0hf�_���,�3��b�xѢE(w����G����`f�H4q�����A|a� !:A)���rY�H�4�]F��h�l63��5�!]�l�c�u�kV��<�Y�ꯇ[�ݑս����*A�%���F���4t�W�$�h0o�������5>���{����{�Ǉ�ݿp���s�{���<w�VCm[�֭�ɇ{�^��{���;���ς3����y�Ζ+�j��aIfǨ�������Y&/�v�7��8�s�]���|�<ؾ|�3�O9���S�:w���GlZ5}�i�ޯ<ܓ�7/~���5Jh�x��(2��5˫R��4�>zF�!+ٔ��˓M�P����Z�.[bQG�(05��xSn�!+Τ����eQ4�t�!=^��*��g��]�A��3S-���?	���$���ͻ�+���OU*(X�B�$룐�&�G	���M��ĎD�Ǝ��)����
�D��$�$�895LG�V��0��� ��LԐ@��	f^H3���?u�E_I��M�Ҹ\�
X�v���i�U:\��~@qFx�i�H��0G��}}������bA��{���K�R�|>_ss���iiiy��.x��0��D�2�"Y,W����rW��pA9��dv8�f��\a�W�ڧ&���)�[˺�B��a�o3 3�t����� �����C�[���	xn��|������7�kn��MN��F���=����.���Ş�}$TBE��L��(q&�s���&��5�q7מ�>u�q�l��-k�ٹi��m��st�ûwۻ|�ڲy���K�����s��]�c��T��Ĕe�;�Ȍ�мo�h������.�#,�nM�!#�hH���I���̊�!�ҡ���nf̴�s�M#�ic�ىf->R�b�w�7e'�+^�?s�̬Eu�e����?w��O�eC>�왜���L�)OIQ�������$�D����!"�@�h�4�Y|?�����RA�;ac�(�{ʇ��>�l;�Gnȏ����R2t��'؊0)eE���x�
��av�m.���KW��U������}띷���3猊�N) �wMEFc��S�)))�֭;~��իWO�:u�����ϳ��ӧ���s�2���66�%F��(�"S�M3�ֲ������;����R2�<j�,�Ak���Ԭ� �X���dV�Pk�^k65e�cL�Bx�)X.���M-�A��'��@�ƻ��� �h�o�m�F���h�~h���w[o��< ���|�'��D�Z ��R������G��3��F�,9����=8s�~��-󶬴.//v�-��/�l>��D�u��"wøe?�2�Zfɋ.M����R������f6��c�)������}��U�rJ@���|c�i��ͤ��aH7{z7�P�Cm�
3g	�y�6�Т�n�Ù���y�t��>�8"6�_T�"1I%KK�+Ti�Ԟ��TU��d�,U*K�H�ŒdX�I2Z+6�@���R���M�m|�=�rzg�N��
��2x�P�����͹I���α�͘��U�+�0N+�Ϛm�Un4϶��v��
5�AZ��ޢP�����L�͡A#o8���0/�*�3س�p�_c�ǥE���	���B�+-�t8�l�JX.��i*v�x�Is��/�Y0Cf+@E��CM�欎�=_*(a�.���K<S�6�ԂLv�?L�5��h�{}7=�;��ݭ-�����10��B��OKA��4�l_k�%�U`f���Cp�=&���I���6ʘ_��t�b�F���e1b�n�٭���^�n6s��m܃��f���;u�/잸ޕj,��Rk�m��ʣ/f�U7�9�d�� m��8gnW�G���D,��]X��ƌ���㝹���sGu-G�s�,�{>.��ڮ��� >�44֥�����H����3�������;ܓL�D����Ai�d�,Y�����U�
�*��IPe�RRӒ�Uؒhq�$er�,	:jY��?y�ֲu����ڮd�BŞ��,�B���q:��uU�Faʃ�/�ڧ����nZa�m��T�hJ3sx�0����`�>���l�^x�l��l���
���ĕ�[�����h!�%�̲d�X)-*�ewZ,n������(]7�W��$�0�qDB���R����c���`�YɤBq���J��N�,�.�0��4����� �B�=������`7 Z�������@K+�e>@}������n c�(�8f���vZؓ'��(GV7�@ا�.��J�%��!;��М�/H+���U8�9�h�C��rly��3F��^�2S++��d�
&�;�9�%�0L��;���|u�+xs���oÖ�Q��7[z��Z��n�\�8�:ƒ�M�K��)W`��k��C`B��d�Bd�5x�U�CcG�s��YBkVRI��y�-�� �)����A�q�by�\�,��(ũ*���d�Oo�\���
�J���J00-u�VYT�ߵ����ty��Y��֬rN��L�3{y=X`#�4�@��6gG:5�;r#-���Nt���t:�.�%E.�0`o����W������B��h�*��c��&N1E�;3�Arbb"�������z� .!^��SH�M7;Lx��s͚�i
}atIV�E�(��h��Ñ��M��aH��D��_k�/��_>3����y	f�
: _��D�|�6OK[-�so5�h�4475��4��=ܷf8�������90�?K	3?�e�Q��0�;x�e��!��uP�i��ؕ}H��L���6�}^q�{�6sO���~������|�����	�O����H�P�'�5q��p���=��j��`��'�cWW�_ܡgf��=�ag�a�c\�ʁ�B�w���&n�ZS �F���>����=)�1,�$[5K+�X)�)���h�f~SB'+Di
q�"%%I��ɒ��)baZbbV�tZ�H���w.m��n�q/�,k �bW��eA�A
�B�A� ��yfB�тL�J"����ï	u��4�c�
��?k*..�����h4�>L���q���H$2�LR�4��W�psa� �Y&�l��/**�{l��Ot�$��Y�M90�c��qp���c*.��wʨPAG��ޖ�a���:���\2�scsk}k3�1.�Ɇ�f|���o��7���M7o4���o�/�7��Ya,��O�R��b�sx�� U�cGn7k�V���Ęҡ9#���};�Ax�d�%��$���Ӎ4m[z���ݿ��i��n^��|�ey�q�۾b�ܯ�o8����� ��
wsΉo�����t4�y���0�'�k���H�K�^Ag���� ��ʺ9����=�1>2N؋gbY�c�<�9�I��|o}$ի�'=+>s@1&[���,ꛜ�+�OZϾ�=�%�N�}��� 0�Ꙝ�7U��B2$���dK!́D�v���-܃o��V�Q JꝂs�N2K6���s_bǫ�f��\�!��FϞS^�v�o��[�v��?�%]�c#�i(��|�כ8ŦI�X������{��
�֭�I�bfx��I�&�T~��'�����)�j���&�T
eJR�̙3�VS�I�_<~D�Ue�h��8�-��ۅ�#���7��/��<��=�֑"�)�=�Lw����g�J���	�7����F��������s�}�)�fZ̕��,3�;^�{V2Y���ұgg�ݚp�إ&������ ��5+\�����+���~�k�q�7��c]Vi��X��Wۏ��u���3�w߻��}�m�~W��y�\�U�6]{�R�=p}�e�'pj�4,�b��� _�y����~�����e/{&8f���~�=��$�1�=�f��J|
�rF>��� 4s/���Pl*T����.�%��(`Z�1NQ�O��גL�$Px�qI�����QC�J�K5c���s��.���O@�M���)��g	�i'�Y�Ԙ���_����������������.o��w��a�5�k
���W�Z�B������\__�r�J\ ��C���G0'ƅ	c"��$�H"�|��G���~q�R��0��â����@GVt�.�!��� �-�iƥD6.o��L����nc������~bƶ���^���m�o��	`�f�͌�	u��ˑ�=]GI��8�&̔�ָ�VA�O�ئ���u��+/����rl��x�������9{�<��ճW}׏_<y����G�?p��/v~cY^9���ܽ��2�O��ȏ���Q��I�+�,����0S��߅/�/ܗ�a'�+�I��3��q+��I�h3|0�/2���g~��}��2B9S��@60-^%�sj�2U�L�C�%'�Ҕ��R��$�H�J>�\<,E7�x�B����^�QOXh�@aE��;됎G�S˞���L!GJ��G���Q�2�������.���#�ѡ*j�~m�Q �իW�б�ٸ-x�w�ށ��P�ӦM{���j�k��f8=�#q@
r-�,�&�D�����
�hW~Za<6����l�R���_���]S.�Ů)F)�����~�uf=X��x�����"o��7|�y-�i���_K��FK��6�|��ӳg?=}����Ϟ���3�`�"a�&{"<&{d�p1�G�����-TǠ �2�l�A3�b{���[�U�7��{�СӇO_8}��ZC���_W����Vn��=�����K���s|��=��K�?���./��g�6�D<w��a���t��Q
�8�D���f7��Z�*�}��6��+L-C@2|o��|���0��orr\�Sg��G��HH��S���deJrJRjO��E�3M�S�J��R)=i}��TA�2���)#2?��_�ݚ w�սb3�LTX�ڷ��m�eHX�I5���ڥ˻]�zD�Ɔ�����wZ8�fJ���H~=����e˖=~���f�	�ܹs��a'��ӧO_W3cC�����(�L.��Ȋ�K���)�������ݭ9]9a��pgV�����:��aŠ#s ��^f~%�v��aC��:=MAﭠ�N��=�"f�����7^�׷�h2q�� ��=���Fu��A�r��Gi,�!����/Ί(�.�_2����x��a����n�|�<4#,ϋ���Jr���{T�v��J��3��~��Y_��뫇�����<�:�No���j}����z�[���T_>z�Ю���lX�������֨�Ůal(D�PRSp͛�wX�!�-,*�!fv���if|�ܐif��7�����.�5O���'����?JJ�)KP��iI�$�B%GIL���dL�)r%��U�L�D�+I	*��oj_���_-��=���.(��(V���I�v��2;��G�K����3�%x���3�)?���Ifzx�ڵ �o߾�>3NB3�۷�G���"����}�7�J�;J�(�'�U�<1Q))����(i���%�4Oyv�;3�InC�ɯ��r	/�ua&�iL�[l�d�do� �h���6ܫ�v��Ż5w�?�������F�'�������M�u1�m|��݃��߆�'�Ǵ��g�����S���DH���Ҍ>e���]?s��t�m��[�n��� ���VK0詯�v���ikѵ�����s�lFET�TG)o�7����M{6U������܍��Sd�¨�'J�o
�ys����47�Y�Z�{��N�3+�|��0�* 7G���?�z��L]�(���D���:Y�"KLK���Yr�,M%륒���짐�J���ԅ��%N+����=�0�v�[���W6Ņn�� /�K�[l�Me0���0���-���f~<v������Ç#F��������z=�@A���<t�P����u�fc������GD'�e=�*X9���R�J&��4OpP����C#lC���;	cҙgd�'�%��D��m;[��������7nj^������Xs{��k�����j]`�W���|���	�*݊��{�t��0���57=I��a�<Y1�e��Y�n��M�xW~�9'J��d-Xv�[w�d�����N\8�r# ��p����X���-����7ZZ�T54)�	Ȩ�~��n5���{�5W[��?^:���>˚�-�=o�e%5�����\>Q�D��yc�>��Td��-y�Y� _�k�K�+�a�� �\l ��2��1�q��07?枋���&KR�RS�U�$�J)�'��$ǧ������A�Y�:�Fw��{%%%�RTR%�q�R1$g�]����{$���X��[袇bґ|��2���Q�)Ѡ��i�#�i,g���}��̀9*�g��n�׆�3f���P��b?���|�A�;���Ǝ��DD�D�
�B$�i��咸�D���Xg�v�ZN����,bw����++�s;�0��2yþ �����Uw%p���U�/Z�~���`�a0��~��k�4����
���/^���m���׎k��b���/�;��]3��
��3�qd����AX�Ѻ��`�Zc�{�^;w��N���Z_w�-�ᇏ�@$?}���<?�s��P��fO�Wh�����o��v7�mi�inn<v����Lk�.>,=�-�4/��
�o��M�j����΍-ǿm:�-p|����7O�}�Bfɏ(��)[|��X�(Α�r��yu;z��g�Ɣe,��]o��hR��
Oh�P5a��~�bM��6�_�i�TZ���L�S! �}%�W9���E�E��E�����&�D�%�IR�W()f���ͼ��^�^m��9��G�QH��2֜�Qj��U�a����^3�K�Լ�-�3Hop��u��˫�����N�Z�2d��`�={vEE�����������jk ��D�D�$b�J� JLMI�����G)b��	ԛ��,Di6��f�?��Ꚃ���#�X���aو��uaf�1��Z�x]�l�Y���7<n�iڳӳh馌���wg}�7��Ό�d��2�ߞ!�kYp�+��56��ڼ�� ���#�03�P݀Y�ˋu���h�$�99iTLkv�#��%#�\��3�/����"�C��9ae�.�A |�U#6kU���k�\;�t��w��|$ݶ���4�ݽ����3�{���;7����3	xfQ;�ڑ7߯�S}�o�yU�$�59Q�C�l��a�`ۇ�3�H�v��X��7�nC��p���E��n��;����=��Ҷq߸�r����5����5��N�i���]����B�#th{�{��5z�]%'W'rpi�;�SJ���=�8y�^�ZW��L�K.��W�5�*J�X�P;_U^�8!�<^0)&2;.��B$K�ʓT

����{ኣrE����CXee�E���=�1B�ge��JN�=�o��?���W֮�`�lf��f����1o|�sbb"�p������73������J�D����^8|X^ʐ>I��B�MVꁏ6�|����:��;��\6��T�� Q$^f>1�0�P��0���yC͍]���o���=%�s��-�;�>�>�<��YSR��bͣ��n{�p����f�a���%��3��F��BK8�s�L�1̜���ةq��,����]�+�Xdˑص	N-`�tj����K�-�s�m˫��q��⵺+MAtoc�U�4���֦��nq?=��w?}��.N��A�`=�h����p�V�h�_����Ў%_�:�����Ҝmʌwh�F sש���W`�m�_�9��|��_���6Ү(�r�:��i5�4n�IV��r�/M��j�蛹��}Ӟ����%�j��1��D�s���ܽ1�JdM���ܽ��c�K���F��Q���hUNe�>�$~e)�*E)�X?M����^�R�����!{�mW�W;�Pz�o�$��~�xE���y��NN�9�>�dӅ�2`�D���²�Fya�dw!�4F�֚����r�N�N�M���N�K�J������%��~����� >>0�^P�``�c��}���+o�h�4$^,JPʤ�I�M��l�r۰�q)��[>�O�aZ����
�ڠ�5�Ͱ��
���%�_��0{��{�3�fB�&�g��ߵ�+7��=[��l�演o�Jȩ�Y�Ff��f6|����m�F�;�!&��$3��`�8��eX�qNB<'��`�A�D�p2���+�vd�>#A�U26Z�S�c�ْҜ����;1�%�O$���%4�=�%y]l�ܹ����}��'���{7�'����_ߪ�H�+o�����=�����Z�u}�{ЯrL���P�P�g0褁�c&�߂�o��*������{��#W������t�3?ʤV���{���<�y��4�#j�;�vʭ�q�B�k���7u�1�D��t���@�XX�᦬xG^��0�L$��iIJ�LA�?��M���t�L���l���w���ߛ�a͸�C,qa����TR|��]$���YQF0G��pM2J*i![6M�r���X�:�(/_?�5�E-�Iɩ���~�_��Au�>l|쁎!��������a0��K��������!R�U�)�f8�*��)���ֱ�z5*Y�+��rmj��F�����6+=���s(xP'��W[�]�醷�Y}���o����A��&C�6[�^#_�+>9)����Fc`�[}!h���0��z��lD2Y<��ny��#��i}V<�SeH�6�5?�$+ڨ����gʒZ�2�Z�*��eC�E��As'Vsw����������j=�-�~��t,Òp��y����֧�����#\���<���@�����A] �|��ʾ����k��ڷ��D��(�Z�P���0���
���ݳo_��0�s6-���J,�L�'�nΒ�|�M\��0]43�4c��:w{�R}�sB#�_c���'�ɳG{��U����_X-�U51��n�FƉKr=�i!?hf	-���<�Ӣ�]aaKD1˔�2R�Q�ܜ�ص�ڽY}�"��Ә�A��^JyOUj�<%YE�:`FDC#�����^)��{x�μ�&�i�D�'��/�d=�\W^�p��6��43����l �`��@��u��=##c���S�L��dl����_��{2�A{���ـqB5e�G����\� �M�1�l��n2�sj����|�!Gb+�%*��тip7�9�H��f��%�����6�f�����V_+hl�7>�T���+���g�8l]�r�Z�iX�����s~,���	��5���6Z��ҏ|��V;����Wo{�,�a|���է��j�=?A3OQ�/)��@i̓�U,��f��2d�h��C�0�_v��[��|�} ���%�[��꠯������|�z����m��������[���k������𷛛������~��u�O/k�'����Ԡze66�b�0�givx�vi��m۲_�9ڝs�/���%�Y�O�ܽ��&�=/ґ�ݜ͜��,�=i������yO��@{��`�9h�.E��F��٣�̚�e98ϛ;yf̊ri�Fm�֟��޽:`�'�H㦄E���X(��#[���Q�g�����'iv�~P����CE	��^rZn*I��qV:�y�K���7Z�H�,�p]�$�)_b��{M���
z��*3�w��g��<%%�˻�A3��?� 3�������Y1v�ػw�>���ӧ?��cUU���f��Y�����[��1�i���hq�H�P����R��Zi�I�c������1�����U��V��]�U�fK�2�����m<�N�(��	+@�f
<l�����> on
z�jZ�l�Q^��w������i̓���MY�sc2.�e��g�g�[})�����Gg���3̨2.��$����U�(�hɕ��¦|��1j����/�ޫ���=���G�.�T��/"�ih!Ag~��`��i�6�vmZ���]P�-�>oCu[�$z�/�5�7�/���ײe"�o4�ik�{jA~S����M1�A��`c��6PW�?�����������K����N��k�i���TP��j��l�z{���j )1�&�� fs�aTw;k]Y�M��7���õ�>�᧖)����e+l؏����M��2g\=� N5N�ig]���@�*x߂�S���)�T�'ML�R�0ό�-��X �M�\��Eq�3Ҿ��{yJ�퇥��7T$�)U�(����Դ~��7�'_]ګ,���b�T4��|7r(kXv$s��C�'�XP:~�~�l��J]i����TRe6T�]FS��Zaw'��~�B�fZ)��1o4vu�nݠ~���g̘q��P*��l~��7�>.c��kojr��'J��Tb��l�TY\K��9V�~�m�\Ӥ��)�3*Jf�+�lQIn��ޖ�1�*�N�_4D�̬<����`�'N�`���<�M�62���Ձ}�[gW�0`]�⛁�7N^������g��0xP�̢�����3������|���hf����2�f6JL���������W]~���=��y��������{9�����M�e�0eu��v7dK�}ʆ�<���˧=�5A_}k���oj���m	�6��خ楖��)�_��!���ꛂ���?0n�������yOs��s��ʱ���Ԩn���2Be��/����+�Z��o,��v7fD��$F�P�콜�e�&�Ig+�I3�q����LVn�����F����1�,��Bk~���ySGΝ5}�&��j�D�iȊ���sj�5?�a��0�T*Y���,nrd��{����M���3S7���S��Y���K�̃E�)y`N��`��=e0'�)6(������s�!2P<�۸)�����l�v��e5WP,��NW��>�]ջw�w��S���}��|��3C��Z�� ����e˖y�^ֽ������ϛL&����^mÑ��֜�"����[�B�c��nw�,Uv����9MF��t�)�=!�TW���T��r
�7���3�`����g~�6os�/�x�S�ۿ3�d��̬o?���~?�iP��{n���@���%F�/^����P�8��Z���!f���mf�N[^ā�3s`��)��ƫ��?��+�V��\���r���:��i�!s��lw~�UgҪfj�<����3�����F��&fo�- ���\�MMu4��m�h��{����H�S��M?���khj������s��v]<6bv�� ��d�7m9��0s�āe>�&��_����b,j�Y���A�鎱��
��(u�^W�)֫�0\�|T>VU����<@���܌��:򺛳�M9�k��jϬ��eΞ�X�)��w3d�ʽ��%C��,KV%%���垊>��H{d���-i�-T�>R}�r[?ő�i����D�����X���ќ*�\��ξ�=�|� �oQ�	[`��8>h�����xu~6s>E�w:,�.��a�8�.��a�V��{���>�����{o���4�9����s�hZ8�F��x�$�N�#G���f��R���r�#[�`gee�o���ZUD"���r��n��fv��j��NlV��␖���q�3������$QK�?�F_hX¢y�����lң��(:�S�����ͷZ�w�����bå����y��U�������9��5s7n�~����p�Css�Z����Cn`O���{Sl#�R6�^�-O^��u��u�u��Tcp�g%X5���$���m�\�O��2VM�5/���T��͕�g��i���$7�+0�`�z�w��<���G�д�����f�Rl�@���7����P��6���+�N훼�*3�|��BX��/N�b���os�>Sj/�~h�w�/w�G�x����.��nH��r?^2�4w�y�E�ٽ�7���Rf�GE�Ԇ;4af*+9�K�pm��ŕbk>,m�^[��9�W�2%9YE��`f��%|g�,׈W)���)˔�Չ1k�݇�E�R�0Xª��Դ^�B�����>B�M�w	�! �5�๘�N0����Q�3;�����B�@�%��ęrWE�������@'���)n�������p ���:h�3�={��v���E�6�]�Z�K0�d2+��p٨��lxH
��p���S�y|y����+ҡ�eAKĘh�9�Ki������<τ.������8C��U7�����ۗ�5>��nW�7�om��Άo �6nn�z��ڭ;���p����RS6�zk�͛mwBQ��<��ߓ6~֔������+Jr��T执Oq>lih?�����FGv�%'�Z����f([h�Mt�-��k���;�\9���W�[��͞��:fc����qp���d�Ug�i)v��WZ��^_M��������3���]u�@2�����
����^��SΘ����u�kۉ�mG�̿�����O��'�s�9��3N�Y��&T���۝߯:R�>}����PG��a�J��%'V�*HB->(.��>k}�=IJNJU��ȓT*E�$?.abTlQx�."�(*lFd��Qݦ����}�(�062G"�e*�<%�'9�i=���>�d�=�e�.ڡ��R�6<���hLQKM�,Ǹ��&g��m3϶S鶻]�6��"f����f��]�~�?f6������Ͽ}�6~��ɣG��=ZVVֻwo\�G�ƾ�����(�H�
�Bn�Z�N�c�j�Ѣ�x@��
3�貖U�Ɣϒ�P{���l�X��0������!������s�B@�w����چ�׫zk��?��<i�}�X��������F������V�ܾy�~�m8 �����`����ly�pyi���׿�W�:K�bI�(lp��Q�QHP8��n�=��n%���eb�O����SWN�˅!�� E���C3���Kj��+�|#P�o���n*oS�u��5a��P<g8xqlm lF�K���o3tZ�13�L�J�ZiYN���]-Ei$�w���M��f�E�#D<��Z`��p�xW~��A,:'�g�I2����<{�0�_/�J�R$�LJKIII�K��Ҽ��Ⴘ�х�Q��at~bln<0�"�����*�ErR/yRj�R10/��`㥽xք�݆�H0�:`f�).�l�d��2s���0�[�;����6��t��|�]�;fff�`�@�̰��g����7o�<nܸ���jp�->>�3ΰo���#1=�����K�2�<LF�`TRp�i���+��l[�\���3�:m�9�;o� ���,fi��0�����0�$cc0S`�N���L!���z���G�����fO��bh��Ҽ�
_��z��[(�A���N�(d�u��7��)���MY(l0�qu'8�|-�g���a�*��Ģ��f_#w7r��D��8�&g�⼵ǿ=��_�����4�|�[~	f��y]�t2������[���|>[��Γ���bfa c�!�(��Y0���!p�e�<�5?�h��;�8�@;�[s.�mǘg�]�>֜������\T�48�0�2Y��?pܓ�tQ��\�T%+RS�I4���L�O.�'�(��d��JQOi|o	�'���%ь�^���T�X��f�Ά+{P�t6��-3�HjQ��t����9z]��8�V4�\4�VRe��q����t����睷�m�򙱽1�� j߾}a��%f�n�olS����x�=�Qq�8�V�\���J̶
�@J+M3�ӪS皦,0N���Ι.5��"�^ 6����B��=0�pmC��Yc�ɍ-$^Q(�o��B>�oh��v�s�!~?�(�_[Ss[ p�����&~��>m횙b��#-d��<�[V�k:�2�����A�D��2f��c���p�ě5�2�#�������j˲ݧ��*�`ׁC��[�����*���n�Ҋ�8`$��	x3���zh�d�����s�O3�d��l�)$	����6H���c]y1vM�>ƶؑ��Ht�]�yȅhw^wy��%�b�z�e���cf<8�PL����Q�pw.��f����tf����1�${Ƨr����~�4���+�!QAhQ9|P(SQ@e)re�4����\�,JN��*������f>8�Ȁ��/?n�3�x.*��L�MiR���֏�*�c=�0:�4~B���gv��iw��S��~�ݷ���X����P(�'����ç��{`��1>�D"f��������BA|b�
��Pς�mq�M����Q��gY�q���[�@��h���f-�PP���v������5̌g:���`nh@��[�eR�����lE�hm�����R���&P�[��;��m����J��r�53�ӳ[��T��XG^�SM�dK�y2S��8Ch�0MHEݔ�BH�W�ACGf��ʇ*�E��-���-��9���[�	R��`���	�h�H���W���Ar'�af�d��Gf��S�f����W	�H��2E/��_	_��,2.~I�P�n�ǻ�af�']�-�o͢�f��� �ak�B���PH�H-K��]��\��U��L��e�?���Ɋi���������'E�����M��K��[��[�S�HQ��B���N��&�%V*���k���gݶ��{�Օ=b=0=��Z�!t�nc3?0����4k�e���lE��B��i�l���6��t�\�Y�Dc���`���`~�H#�./i�Y� �Ğ�gTxli��W�1���a�@��T�d�3��I�u�<�9��~T�L��D#)�ėdɊ��e�SȖ��;�xe�g�#3��u�s�f6�j��$������2����滬�� T�������(1�g�	� �0#~�n
ܾu��3~if�����ص�PơP?1z
 $u���Qh�GY��3��d7sfWغ���%�깻ƕ�mGv]��������wS��a���� 3�a���s��P��r`{Ś�^���婢.lUffS�ܯ�����a����J�q�y�d
�⠘T��_r���� ��gQ�)���d�9q=�e��:�#�C��:�(�$���N΍W���@�G��J1�d�d(&�TiJ��P&Ao�R�@Z,�(�Rz)�r���5,U?r�����n����þf&xF$ �ݖfJ�L4dv�)uZi������pٝ�B�y�hE���̀��H�P�9�Fhi�<�$43.�e8`��}����8(�&Ƨ*TIR�̩S�j�Ya�pN���7���s��Z5	�\C}����t��LC��:,mRο� ���3`fʙ�p0D5��$  ��IDAT2�
:�����lk��MM-�&�㇋���x������7x�	f$���ÜfaΡ�W5���5Ӏ�>h&��`ʤ���,1Xڰ=߷d
玀�))�>����?�^���C�_��B�<�)�4�E�C�4ޗ��e��m�zffC�=�{��v�k����f��e�q��}I��s�{A�{��}>� ��ٷ�	t/����(q7M��E��p�W�>����f�QϪ� W@���<��@1=7>���D����RAOib/�4M.I�ŧI���=���$1������>R�PK��b}����닻i֔�O��`ic��"m��D�')

�ʹ��\}��U�t���f~�����7��Q:lذ�ׯ���x<���z���UWW766�|-��.}��6�)���%�@�R,-�1�n3�g���MH--�3h�x�1�=`s��K��ct�~���X�3���0͂�S(����3`n癐&���W�!�A�-�5���6�p��9h��&o3]Æg߼}����O���)��6Zqe)�D�؃�$�Y�(����޷��x��l���������x�oM[�4��{�|�Ԭ�%�KӧBC�@���jkS}�G�]CnR���O��f�����S���>���A���3���佊�����'I�'��t�� $�w��3+���Tf��mܣ�9��5Bk�Ԩ�����P<����qAy�I�)
?�P<�c鈏#�G�`��ӏT�3E&�#�3i��������iy�i��)BɃ�\@
;'��B��P��#>�H;dVѴ���8����owy�=sTL$<��3S��|��?�p�ҥ.�;w���p�p���˗A5
�ĉٷ^}K��Gڄ�1��D��iI��&M4��&M?h�&�0,ޑg�U�+��)F�"�;�fd����`�K���a~t�>�́ -:C���)5q1��rҰ��@��z��؊���r���ko��8��nݺ�_f0���`F�!����nx�ْ�����~��g���t�j��=��]��J*�C�'�?���!��@M0X��T��n	��f���K�Vo��5���<���56Ws7s*�%������K����]"�C�O�X0���H�T���|�{�w���V�D��h���'���iI�A�`�u������D��[̯�
�B3�q��a�5kc,4��se�� �3x��O˲"{Q0Z����3��	\Z3�~3���ݵk���D|ıH$ڴi�",m�l�)S���D�$�>:J'�{"�H`���P�����)Nˌ2��������΄��3�
j�l_f���[0������w�����ۗ`�0�ϼ�H�]V|��4���@#����z=��g��_�V���4�3w��6���$�8ND����/�a���v�w��q�ٞ�qHt��p���܄��;�{�e�oo?p� xnn�g(X��!�|3�?P��_�z��iUl�3�u5T�� ?T��W{���]��W�_�Z�ج(R��,z�L������̐�3��/I�՗`�<����{�r�{2�jR?�0N�N��cY4Mf�m�հ�3����dEZ�ƚ��Z�ɰ�g�V��c������t�(����$w$��t�^'~�CP|��O�w�;b�0��^�w�������Ϭŋ��m۶�O��`MHH7n
��.����!��&Q'sRJ���RȤ�a*��,9�`�����\!PY�����c9Ê;�'[3C���O��t�gO�p������?dz��{��S�s^X��gϟ?{��s��?=�����fS���`���@f��f��f��Sy뀙���b��8[���4�� ʹl�ȮQ9�%ٛ�\�4�U�����N]���4�.��L	6QGt��*F5���?E����ם�xzۑ�/n�|�7�l�T��, �#e�e3a�!��K׳?u�9���	��r")݇B̥GZ3P;�ӠV� p��f��>�����
����n
���)�n�-f�^K�x��#,����g�M$"[~ׂT���;](���f~�=�L�^�3�3v�۔��h�A����o��̝����I�&={�l�ԩ���چ	Eq��6H���͜����)V�FE�0�͚HC:�uG�*��C�4����1vE��0?{�?�DH=��|���?Kh�%ӟ|���=c!� ��;wn�r���B��gn_тn�`Ʒ�$�f��=]�-O�R�`�NR�X�Nu�KۣtP�]������<7��x��G.�\{)�⅊nn�U���녙]��Dvu�������������W7\;r���G�n[��ǽW�[�*'Jy�VZ�������w�̞�����ga׳?�t�%�8�n%ի럵���p��1�_mψpR��aZ�����2j���F��s�wfW7a�뙭�Z�}1��o�/2h��dF�$u~��t>�x��Y5=F���wy�ɟ��'>>uM����Z�q���p64����Q
ax�Or��[�n���83z����^y����D	b%�`�"%%E&�&+����J��0�}�YF��D�f��ff7!+�i�y��#NR��o��������
�3�L:]�~7�����[�Q��0����;�0��%
0S�(>�#��!�Tl/�젣��d}Qƌw^��xW~Bq�f���m&�.����='�_��c]�u�Ԯ��.6�	߸�����̾`Cc���k?��p������^8p�����`V:k�`���¿��35�0aq>����=Ԉ�/$��B�`���c����~޿||���ů�p�EMȖfʍ0��-Q��ߢ�h'L�B�PԦf
��oP���8�14����sJXR�8�~�X��p^3���]�ʼ��6-O�/������`�peq0��fl���C)^�reYY����õk��ݻ����.xō��b�!ёQ��	R�$��4�=I*�N�-#��wo�
M����Z�Q,@2�Jd�3�f0�rƩN'I��ܒ�<3��x~�ZB��:��7��oj�������� M�޼}#��f<�1�o0wV6b���8[n�1�.MX��;���@8}H��c��ܺ6e�~�/w�s���KW~l�{L�8[�f_�e�d�3����zMc�W�qh�փ;J�̧�W�;��0��8
{����AEB�����0� ���W&!4�T���Ӧ�c\���F�W���ߦ��":�����`f_{��f�L��2�\鰢Ý9�6M�9On��>&�rJn����)���B��.5e����� \��⶿���}'3�K�ۍ(�P�,.{�LnJ��]���߽K0C9wtM�>s�7�̰�ٲ��6>�n2��T�9�ɓ'���^�j.}��6�,��J@����b1� ��A�R*�I�Q=Ec!4��Fq�ݚ�j��rF.��kd�p�W|a��b0� /1�(�����<]X��;0���y�h?O�<o<�D5���;�̟P�b���{^^w�L�s(����-�L7���6�)P�����x�����I���-j١��Ԯ�n4�77Ѣ�/���|�����󷯙U��j���w>���3GO�p����\��z����S?�����S7���^5~r#w�����鲢\���kj]�|�$��г�1�����[��N�j8�������7����X'���~��{lᱍ	����<eI��ݽ�#A;u�2&~i������#���o���2�����ӕ����-����?�1��j!�3�L�آ��O&.4[>�_�n��5K�]f�|Q�sf�����x=��5��`f�g�[�B���=g	����Vw7j��~���
�5��w@4	�s����9<�FJ���LfA��g�!�=0ƍ�8��;''g�ر0�G�ѷo_f��o���"c⣅0 �R�J� JLIVɤ��4����4�0d~�)=�B��6���T�BkN�9'�BsX�A(Ө�#�5]�Q۷xdw���>��(|�h�]�$H�����ya�A�<�}evMg�&�����{�S��zd�6Ͳh
z�>��q�&��O�����OOq����xR 4m�����,��C';�f�t\ ��q�\�ϑ�����n_|�]�s��*�u�{ӑ��O��vf����>��۳���;��؎y_/�U�,>�����:��Ê1���8c�Т�w�h�I�Ы��_���B�F�3e�a��^~q������^vy��͕�Fd�|�k�n4rm]�����a�ܽ)۪t����qv�m���y��}k��]}u��U��;ձ�Eq��_r��`���Z�0�b�2�YGN^d�X�p����W�X�x��+�^a_>o�\}jI���`�&�P��Y�#�y� �C�3�=?/�z�33ʑ����<���.2Č���O��&�5L��,L ��޻����s�xaxllL�P���	X� �к���̚�q�4���q�}�7^3���@�@*%)�{�M;��t���)�G��.�HM�WY��0��Hw��������b�MYqF�ʬ*d+��I>3�0yzN��roQ_�c�C��Qɫ����G���Ҽ��|E�6~�={��񣟞<x����o������z�Z��t�����7Q�W��c����ܣf�A�!?�B0�Ff*�<3T:��?/a�!��,qyA�M���K����-8��:w���q����}_�VUN����R7m�c�BK險��VA�5p��۟W�M�=AiRG�37�C%��v�u�Ы��k0��s�F0T��T�	}���iM���c��%e�$�'�|��!�=h��������7������sc�.+�� ̩��m�	�AY�M,S�ͅ]6LYrKC�����r�8?�����d�{Ғ�O�U|�d����\�x��e z�j,�j�����c�� �?p��@3��3�� �k����Ì�-�P�����rųr���Κm6;L�+zI候i永��S _?h��2�e��*�3���GPݵkWF5��+nsd�06.&.>N"���r��I�f�;�s]��zOS+�y��lɌp�� j�Ce�ބX3!�7^t.�T�CPH>�5��݇Sz��fy���= ��Ǐ�����yy���'���<�7�Y��jh�ַx�h�p��w+���F��>�=�=���x�{)<�H943�;{���:���u�J�t\���3gt7�.M��)��au�2�(޶`�����ݚ�'��� �?��\�n�O�+h˔ArK���f��i>�flE5X�=�^E���0�w�Γ�]���_����mW!j�!�O�ܣ��f���,p�Z��5��+�?m�UR���ӫ܃	��e���6su������N;<�,S<{T���PV�d���3r|쾦�ҵ�_.[�d��eK��X�t�e�V�x��e�/�[���)�*TJ�3� �y�<�K03VY���32\t��P�^-6j��F��S6rLe�n���8��4����}����o�3 ��# ���b�u6�,��w�6c�cfN]�$rX�� ��ۢxg>V(��e
9|�Y'9���ZTe�5�O��]G�r�]�Q����r�4ވ���"�`r� W{�f� �S��k���\{tG݉�u�T�<���Ѻ�����o8�����|_Gr��܁�א=�'�֝b����Ϗm��ݚ�o��޺�j�
����]_���k8��E4���9�m��ܨX�Hw���;��JZ'a�0����O /ʥ�ۅ0��>]��ϖ�rRgh?*�1M�<�h\Q�_R>s�%O?��#��H*�S�
U�ᱺ�(}&�u��d��}ߚ����+
_���B2�}�o�6/�5��IّQ1,�1l�u\�[6+ڬ��c���ծ,Fm4}�	�������ۣ��$�����Ԯ�˯<��YT6f�哕F�NݭdH�3'�B#�gy����r}�s�9S��je_[�l���K�]�jՊ����X�t�ꕫ,]X�f�a�\Ei�АeH����0�J�<�Tn�b��Ț�P/F�� X����a5�����Ys�%�{vy�Ù$���ܥ�?��?E	b�bX;6�)v ���`lL�����n�_�~����7o�|���ݻwoܸ�w�޼�<\ֽ{w�Q�o����h��P�*�2Y���(r�)��a�}b��όBEI^\qv�9?^���H(��ɦE��j�ݨ�h�/_�Y�_�X٠�G��La�她��<EI�hz��,W��EfBp��8�58~u����A�d.��5�l$�	>�<��@eʗ�j�y�2�FQ�_D��&�V>�q`T�څa@:ΰ�"sQcj{��0�*��U{�h��9BX�����;˱c��ˇԜ9�\w����3{��Z���Q�i��2����rPD�6Z+���W[FD9A��S��_�Y:#wk�ɿ��iƲ-��M�eY-c�Gy�-B{A��F>J3�V��ґ�^?��s*�9�*ww��N� 5k�;{�;�Q=����5���8��/�%1��?o��=����� �B��i�����U��~�lɗ+V�X��y�r�y���U�/�o�#-ʔX����f���W��h`��f)��^����G�1�F4�`?�<~�\���fr��������-���-�af��o3Hl�G��8����~��[�lٶm��ÇY!�.H�o��qBje��'��<Q��U�X�NG��T2ב��e�4�4��u� ��!�����1uW���[�>?��3�̴aeH0����P�û��^`��shAEw!�n��q���y��cm�h�k�v�P4K�BV☝�1���{���k͋��>ƛq�#yQ�H����OBž��T���ݬY�
�&�\c���=�Ҏ�O�G��ͣ�{/�y��ƽ[�p�D���O��ܓ���%Wvg,���H���F+�ǡ*�(|��W��7|f2�;�n�)B�f��j�N�j}�QK�my"}��Ue�9�0z�2sw�x�)����[;��4+��|z�e#֜��u�E��H���q�D�U�SK��_�g���0Z�h���ͫ+��Z�z���K�/]��۲e��YR�n���z��b�U��_�٬&N�(�L9S1�-F�%5ȧsJ��6����*�%��%U6K��h3�*+X�������m���k�M���	���kn �XNKK�c̢������c}T{���Ÿ2��W�P�@PHŒdyR�Le3Z�N
jf�[�s*�+����>�g�l�a�R�s��V�ͩ��ʥ)�&�������CW�`ay��M�N����6�/O�?�=_��=�8Ʒ^}O����},,Gq��{�5�-uab�*�v`���A�Lv���6�5P1����t\F%�v%�����Hh+)�>�Q��om��]x�[{�[��ys�/]�}����������w~�}��-뜫��ߺ��#o-wg����9&-�<S�2�_���W>���+uM	�H]���'07r��2H��DEJ,I�_Y�ʩ�=����c���������/���F
�Bazu�1M��گN���;W�c�`J���k�s?h����%~�jf��֪5��Z�|�%K�Z�jђ��W,���2�s����\�h�\��ˌ[�a��`��qx���#p����O�m�̶�`wq��k���V��������o�.o��-��^�9"���l ��e�i�팿��M�6=}��ĉ�G3'��+%4�j���N���t��A��iї��v�U�Ms��l������X�4)ҜO
�g�Ar�Ę������vЕ͆I�J&8���{�	f���VQ5� ���[F�e(����$�2^(�̗U^��1*�Π�Of�gvοtο(�QvM�!+Ѭ��?��E.X�<����s���{b��S�v�y��.�=~��Wϟ�|�ԏ�ۿ�Ȟ��ܲ�j�������W�Y�A�Q�<}Jc����W>��
3�̿3���x�J��q5��Q��z��Z��x]F�eW�[��)�y�7V�p�� ��f�)/�8#}єO�[�?��Y2r멝ǚ.�#�'���9fhf����O���2:��X�ڰ|���sW-��|��5��_f�jѸ%z��%`��B�� �b3���Q8~���:��������r?���:�d��[���i��n��BX:)2�W����0]h�+V f�T��A����fdd�f0v�=p�@v海�hhf�L)��mv'����b���.�Q�N��lw'�g�Jrb���L@�(��`�i��//��$l�MgTBŎWq���w�����y���K�TvK!�:����^�"��H3���Wǖ�L������~<4gŜ��;qt����k�_�5�Є� ��n��R5?̮��v��g��q��W.ޱ��k�y�|?�H�6�IǵՍ4�ﾚ�	�]�YkȘ�g���㛛N�p�����t�||�f�]�Ѫ���*�@���=�x���6�'�d�ه/���w�
w��{��ש���N�A�/{��ꠚk���v;�i`�DKLڏ���,4꿜��fY冥�/���6���n���]��K0�j�`��ǎ��kf�Q��?s��\e�;�<�N���[5Y���ݷ`��3of��c������ +�����Y�f�	&0��5q��o06����r�T����p�,��b�vuTY�-��6�\��j�MtL�e�������i��ej��X���P	i'�A�8�
���'I�dt�P��x��X�v�%��dJ*g�,��ɇ"�aF
ɢ0�/��]5w�j��/�~q���O	�^mm���m����(�(�G�/d��ѝAO���zC��K��>y�#;,+\�
�s�#�hQ)��Ot�����i~S�I��S��d�kIݮ���.��ݒk;\�6~{%^9�������RWa�#/ڔ3vK������d���3?Fn���a9��r櫪K[MG?�p2�v�m�����ϛnr�:?�5�Oco%Z�S�Z?:gZ��O�G-(�tON�K,�L0��n-��2�����0?��#�3��f��U�D?>#���5yqN�y̬*��e.��f[,�&��
;ԆR�=E�v���������l����k���3�Gq��a8������ϋ���'(g�أG|�#F�}핷X�E�S|�l�D�4[lTK�\����m����r��i1X���]Ӓ��@ Өd�i��	+���E��}�ݾ}츆]�N�g~��Ѹld�_ܴ�G$$�C-3�gO�>v\�cx�K.:���V��$ǰd}A屍5�׆E[�|w���8M+�{�|��ǁ�Z腰�~-��`�V�
6y����9����k�^xذ��ej�w�覣���.|�����8�e�}�r�9'���i��X\f���t��}�X򢋆�T�T���}�!�Qc�D���̙p�dfuó����t�68�#��bB-��V��z�U�|�.�I���3�wfu���6�g�c�;`főnE!DByAv̥�Cl�����XlVw%�Jꌵ������NW��}�~����L��	�m��a��6�؀+x޺u+pe�O?�4u�T�g#����>��gϞegg���jH�0#��R�4)	<�fZ�������d���f�6��P6�8z��$�5)�[�A�p�Ȯ		�7�a̝I�,�<�Η�'�Q>�6ficHCp	ƃ@p@�����cF2��L'���a�N-��DC�J������=��m��=�����wn63tۚ}�n6Cn��ۂ^b�S�W�`�=~�I�A�d���'�9�ۺ�������Nai�!z���ᓍ�Ծ6��|(��م2J�� CߐP��4�ݝӣ�6�=(�nN�1[�,���q:Z��t��b�	-�X����rhcM9����֡�Ń�~f�5�ݣа]n��I�9��p�U-4� �fM�U+�愛���0W�a>(��G�Bm`�5��:r��'u��[����Ee��M\h7W?y��h��<��v�-p,����ow�o�s���p�G�
#	�(R�!�^}c���p�R��*��ǃf&7γˠ������W� 3s죅qq�,Y%U*�e�r�k�W8Kg[�V&��OY`�6�8yn�ȪiYd�w�܆�b�W��~�< o�}d�>B�_;_��g���{����� y(���7Iu�,�!�����7��
̌d:���n��~�HnȐZ�rC�@��+\��{�lZs����k�մ�+���ݶgܣ��'Ϟ?|x���� ���S�Φ�@s]c�փ� ������u|���y�ܣQ_:�ဓ%�U�O�����n���5 F�&���aQ��(�t(��
ml��v�B�AP�A3��0ӐHS�,\�.��u5gE��P�P,,C�,j��������]��o%q�Ro�0g):h�Kzې����fMm_��=���A�>f��v�g�Я��cu�2�V�S+Jr�t��Rm���1��esl���a-7[ҔJ>r�2��l5s��0�[0��b1`Nó���c�jl�{p�/��/�3��շ�0ǈE,�i�̢
��n��-*ʲ̟�*)L.��*��Y��i*L���T\�	�tОo����@$w��������q��=��"8����������f0w�Ύ;`�5���W��0��Y�YC����I��r��c{�|���g�Բ��篿y��	���<?���wZ| ��F�9��|A`���@u���ز���kܝ���̵|E���0әr-��=L>
�-����Єokƿ��l�/��M"���<x��8, ��LS-�cΊ4��n��B���4kj40�)R�{E
�]bQ��%{ޚ�ÞA=���(GV�;+ܝ��>`C���0��	(��ODY -���~*Xc6�2��>GQ��4��\^fp�*��
�,���t��YS�91J�N{8����?ܒ�	�pBB�fv5k��N*
��ƾ���� ���%�ry��iUV��i�UZFT�1��+ˍ5�&Xȴ���0����KE��p�P�ۋ	`�yn��m�I&8fw��Yݩ�g�q�nN���<�A�"��@���oV:��>b���J+�Yբ����3��U���~���g=p��j��-��7^����q����{���������;-�:����w=��`1������&oC��s���PA�{����D���G��Qi�6�_�x~�
9̞���~��_h9qYv�]e�y�l`��|��֡�
E�H����ƌx�:�<;�d`n�����?�B��ECrP�&(�v4�"����g�q7ˠ�!�I�����%/�L�����c��~��H�ƂB��|�rRg��O/q�*]�J�5M�$3���� ��̴3�Y��e-a@�a��8��1�����[�1q�f�B^<yZ���v�f�t�m��d8D�n-�\�[aQ;��%S~�3��%=���P�g03a��sN�3|�a��t����?C����ʅ�䰊&��W�0fN5�A����}p�-�2�R�EݾS7/�^����u�7�7}^�|X�_����[���"�Iݺ�6�5��Bj�"l7�ƾ���7R���g�n;����[�;���0�Y�Zz�Nj �	�󨼻��#]������0���L1,m>Z �a�:�<��ٙ!��?A�GjP-�>ok垴kfR�@W`�Rؔ&|�L'��2GJ�FϧG؆DZ��J��b=Ea�	D-�e~��s|)|Q�Idjt((�Y5��_����l�(�s������y�M������T3��m�962*A�Ϝ�TH��3��(��\�̝<"��Iwsnw����&��"c%�r���w�ae��D��~M~����vu�Bp����]�PBTn� �B�.� ̔NS�*��*�yf��gPC��ex#w{ٖ5�}��b�@�*���Դy�����Z�����k�[|��ޠ �dr?lj�%#o�@{��>� �)6���z�������{�G�_��u�~,|�ɣI��Uag���.�a'æ�{Lն	���H�S��:$�:a�ڌ��5��=t������_�ǧ��?�2�\�� �f�<`��rG��6���-���@��dFӺ�vr̴>3'���iك��t�̐fT��s���#��A���x�+��៩,��-�۴��0#m�j�RY�J� �i4��#�����6�_`���4τB�Ҕ@mga$3�G\���'��t�#R���ba?���SC6�D�䋬ZTaa�����]�x�y"[~|Y�ܘ�h�
e����e�k��=Wk/�� lI�V_MK��/^Q����+��|��6yΏn�$�����6��@5�Ty�)����Ss�쑕���}}�� 
y����wqcO�������<��)��E�`���̿�uC�������f��Ϩfpq\9���&��Am����O�t/�ܞ��x�f����0'	�Z;Cn=�=3�I��p%�^hc6�f�A�Y���w;�Z��N�7k��t�/Է��[�a��A��O��i�?2��1qQ�11��T�Ra������JU�cz�E%�(:4�+�{/�KY�3���G��ЋtV�P)��)���5�t�Ic>����EqNBq�جI��	mZ�� ޖ'6j�e93v�YڸK`���<r����C�_/9p�Pm�5�LN�����O0�U��(���7[w�ݸ`��Q mo��3>�`#����m=�׹e�����N
	jnΈ���9�Y�g|S����Nj+�1�ݫa��H?Z��Ȋ�PC�v5�6g;�;Ec��4J>���K�K�(S7������p2�#�P"�$0�(Z�%'����az8�Ü|7���`t��g��zf\�r���S�.J|�ۍ3���pAl��[o���w 30�Y�3����	��@�����J�X��d�qѩ�2>�Sa�Z3��YD�צ��+/�E=	L�xW~�E�bv���Oj>[a�d�~䗦a��_�[�G�6��P����U�v�!�4�]+��ՍX���#?�@�=���zQlu��|v�����U�h�HZ��WU��f��:oc׵zjo��>s��Γ
�SҜ#�uCD0
@=�N�b����;`&�ޚ�`�I0�HLZ���O!��q�����0��6u40M�`���~0���PT9�`_L��le)�|�o��4q��	�pf�&dQ[(s�p�=�:�-��5 �n�!�E�C�׃F:`�q;ϡ�f�`9�ꃺ�CKdeG�2��������=���rv猦YSd��aa���`SA`�(�JU2`NU(TRQ\O��TK�����/cB��+43�!�s�e��3A"Y�����5�o�SHLeY��L�Q-����䆟�����pw���Aw�M(�{��!�i��3�՜��T��l���ɋ�h��_�L�Kk�`5Hj$�&/��)򮯎���qA-`&���7��Z��ݧwN����EB���>�z���LH�C�`� SK�D��4�f_$��"�JY���
3d����&�·+�n�9}�5(�r=O_�ꑡ���7ިr:�<�S�ˍ6�3Ե;�,|X�v�K�9�.���A:��!��@������i�!K�������{�&Z���战?"� 9�:���b�T��2�8M%O���i��bM���D92����̝�S��w���� ��1'����mR�%3ѦU��=K4'V_z���r���
���E���wO__Y��ʱ��rUŅ��^�n\YzT���K͑:C��䎳��P/q�P3�X�D��O�O@��hh'��,���o��ӕ~����0�:x�����N��Ģ�03��d�0��~1�q���5�t�Ȑ�b&+QK�s�-Ñ�]v�>S���^6D�/��}��Xk^�!3ޑ��ԞTJ��Ԭŕ�!T(K"K%~E��e��#7��f6�	��x��J]�J����O))H*-H2��{,�S�$��A���Ͽ<6�`���dt���g��	c�2�F�:��>�/�����2�[]����Nq�٨�?�f���
�c�b3��J�8Q�$�(��؞��?��/	�'�^�_��	��u���#�N~FW���`��y�%�}������;���WL��@9&���Cu��8�T߯o�nHf�3��Rsއ������KgI'���Z�l�8��3�r��״z�I҂r��|l~�H��Q fx�Ԡ�xm���S�Z%:��,�9����_�m���)�|�pv�]=l�}�����]xu��=s���א��M^t}G��2��8E�/;�y�qp��e93vϯ����b$��f��^�9�N���'�	����*R4�>�d�jǴ5�V�2\Sz�FIJs���Z<n��0#��Y�׎�mώ�af��;�Ƌ�/Ɋ�1����}��~���~��׏�����HHE�G�D�B%S%���`�bz%��FƢ����C#��Y�,:�˨��(���$3��T8����Ć�d�v�r}=w��{��ظ/��q�Fe�^V��ս|���+Ҭ�}F������6���	�R��o;��}f�ᤷ=�<�2ll�f���V�D-�X��iMA���K�N��@��*ˡ�
�p'�Z	5h�Rn�/�w��T�H���E���mg�r6���p�l�U���~s֕]��\�n%���i���{ڍ�8]��T��ֹO/��3�0�j��g�j �͜.5i�y��&Ě���B��b[^����g�Я�pmX�^�صn�c�"ˆ�SV�>���Q\�w^�~H���fw���5���ᆌg�|�d��c3�����Ǚs��(m�?'t��Q���=��o��J����� s��(>|/�m�T.U���,u��#G~2L�q
E�r�٨���3N
r&�J��,�"\�:�}��	�Y��/U�9p �90���+��ǁ��{p����7	\�s�j�ۻn�0le�ܘ��@=�Nm�.&��c�O_=멿~��O�9�Fu��s��f�N�ИM|��PO>�O��Ss��㯹r���7������
�Si~�C�2��f����t�׹Ϳ�_�9��7b��%7[�Ƽ�,�^��|��=�(;�6LP��`Vg�(��\��=���
��^����D��|8���q���d�yQF�C�g����ϩ��ff���z)��ơ��5����W�Z�`풅�/��f��/�Z�-����22QG:V
`�#��� f4¿cvC}|1_� C퇖�1�h��L3M��iO���=l��Â�Lf���f�PGm`�3+U�ϦL29lF�I3������:�H���J'��] ����ppx�;�Dw�#�����r_���;(>Y�)Gl/�-ˊ���j9|i٦��-ܣ �`G�4��$[b��٨��+ܔ��z���{N�on���\�fn���&~��a����3�3�-3����M�cN|w�`�q,<��4�E�Q��D/>,�#K3��4*Ӓo�Cҫ8��{�^V"1�	K2i�'K�fyq�`ۥ�T����k���{��7��✴Y�;Z�,�a�R������O0��8���r@�I4������=�g@*y�H#0�'���۰|��%���_�bd�%��.���r�W�
���d�(�k�6�`~A��=/d�C"j!DB�#�fj2f��.p��[\�B��N�.樘�(!�!�c�x0���Qщ�b�L.NN�8k����rW�?�"���LpR�]�X(��X΀��,x��� �M�d�5��)��?Y��L�C�#-��C��F�����hƠ%3D���츊aȍp��]"�:f֐I�U}81e�i�}���&'�5�8���|���س3`�Ml��W���W{����:���w��o֝�<�	߇����#���Z��JH3���ڊ�����|�ب�r��k�"c��V�&'�,m�/0]��^l�7���n�m��X�:={߭W\�!+���{���X�����aK�0?�3~�n�y�n�٫�\�d���k�,]�d���+��\1Ւ���L^a�g�L9�6m�!���afw���0��1&aa�)�	�=;ڔ#0k�l1��\�7��E+�P̝a������~���3;N ����I��NT)��n�ج�*��1-Y7B^��`/%�x)�zZ�T���A2!��_0f*0�W���,�lH8��Mn�i\���ʋv�G�i*.�S�� ʪ�n�yߞ��4�ע�C,Y2�v�&������>}�TS����C��{�eJ�U`nmj��M�M�uޚmGv�?_P�=(:��Kk�95��n���0�I3���4��7����"�ق������_�#u��� [h��[Y���4���x櫫ߏ�L�r�?��!7����� 6@ɿ�9��즤��Ĳ�4���u��8=A-貫��V�!�l������8F[6/�Z>o��%_,_�f�勗�\�jŲ��/�\���*yq���������f�A�'+�=��?�|�)+ʴ���^E#m�Kg[����]ʴ�b0� ����1o����&� fad�$!Q,W$(3�:��U�pZ���s,���3��OqaZQ~�./I���\*
��mowH�!_������z��\XYmJ'��6a+Mw��Ú�ݖ��D�{a�����e �Wa,@s���Ȃ��$s�.�|�k��?|�hC��{Q�2��ۚ�I�$!����̨��`e��'8���>��Gi�O��;M#g��H3�!�/=�o�,���m���Z�{���dDXs�fM�utw7sMYB��;����-�\�̖�c���S+˚�G�m����fiv����������w�k;�����U��1��q0�?{f����S�楋?_�r��K��^�$/_���+W��bi�J��~���B?�o���ÆM��1�jbF��\��sJ�}�H봒y6��\��&�Þܻ'P~�]��x����рY�菲EE��c�"��x�L!R(JM&��9�Qi7[��+FYg��Le�1�1]c��S9a��yYV"\����L��Ӓ�|^�ǿX��u@Ҋ��;�L�d� �f��v��'����C�y��ؒ�Zh��2�LC#\�J�{2T��/�����x�y���k~�5{�����*��$����a�5� 0����+ߟ9�p��c��[��ILZqy`�4�)�:��@3���k�����8cΊ�Qp����Q�ܽ�ue�2��4a��m�vm��{0�6��Լ��;���{4�[|���n���c=G'}]1r�e����c��NIgf����$r���/���8�X8cMŒ/W@3�Z�l��e+W}����k��Z�<f^����� '@7k��|�k�'��2�qs(�}�!���1���eS�f�5�U��UVK��Xn19Ms�n�������4��w�9\Nfv4���ǃC\LtbT����HJ��a�:f�f���YRe�͵���J�X��5L^�+�7%�,Wf�% {��p�_���']��
_/S�Ig�Y:����j�����:�T_�iH�3'�En*�	�Բ����քY�v��s�2�8?k�n/����oV<{�Z�ՖV/��\k�V��B0��L~�6_S.�;q���c�\�������:��G��9֖3��ua~�A#8F.@�IM�˘j���sC�cFlE`�ZYT��S[>K��-ٲ0@M�w�l,��4[�Ϭ��/uJv�bM�Ԭ��6�u!�8Gb��]|fh�ܴ<�2(�H1{��"���\��,Y�r�*�W-�X�ذv�`�����XQ�53���t�~f��y�!!�ņ\eIn�}��y���e��L���f�Z�n��P�tX�>�������?�w���㢙���'��43�f������'ʠ��R��鶕W�K*��,S��R�(��uN#�}Ƽ���S�rd��+�����K;
{#L:N�A��6�)�|�J�F���	�l��,(7%��M�ID4��F�w�]h��FR�����:���
���{����_ [���j��Rl]&�a$�m��&Kz�՗��;t��}yŹ�u{?&MW�L�� fW�
0�s�~?��H����a`m�O�umn:��w*��9�|nS��Ěx�&Ƙ����:wo��Sy�&�8쇟|����n+V��m��\`G����G7���Կ�錪�@��Aló�������vTCV��pԼ"�yK�/]�|��%�[R����_���NI2j�t|�*'�Kc�w,�Q����#�~΅���&Z)�:�h���2�,�9Vg��9�ꮰ؝fk��e���i�����o���?�c��i��-H�C	m����`fǉ�v��jv@�8����C��!͕��9�ѕ3U3)J2�%J� S�FB/�	�#� �43y��_�o����T"_�o��ɖ³�|��?Κg�zt��g�oC��@CKC�M��B�x��j0�o��뚚�l�6�77ֱX�AM��Tsq��=������w׹��9Ӕ:TKG�� �o�������ֽ�Ҷ��lk<����V_�5nk��9,Ґ%w�p�ߘb�	b��h�?l�]^�0�թ��������ٽ'��z�k�u{�$��AQv�ܐ���̨5Ph ,�0~�\o��asf�ָ+�ϟ��<�ڊ�V���Ln̥fX
��CC ������p�7^��3=6{ӝ�p�\Z��zu�},�2����t[��vw�����v������@����fMQ\�鋇�B�E����Z�)���*U�\�r9�N���p�W�d���r8�v
)�����i�,�,Z�o6�?�x���Z�4;�3�G���c����ؖ7|�����t����sv�9x���o�����&?�	h�{�x�5���#n��Cp�9����k���.��}|���_Ω����:OVD�,PJ;��o���9֕i��S�̎/�L,�,9�Ho�+����3p?�2����������u��8�d���.����Q�p��,Yt��H2�cF��b��Lb�����(��_5#�N��&ٽ�����2���鮮������ HY �����ڳ�2w�ԻP�J'����㞃��w��E�c�HYy�`�&�1*�>*�44ܔ	!M+	4H��G̾6܃�0��`����'[+O��3[;۬/4Z�l�B��خ+4��&{���͆��	ԢΏ�P��{N�����"���0D���9@6���`�e.tX�F��h3�m3֢B��Ē;�8|N.?O�	�ن6g/�Ab�p�z����ݲ���3���3ͬi5�����Ê�+rJ�kvn�ulס��@_�t���3`u߻y��M��{���;��]�to�y����.�?��Ⱦ�]�ek���.��^��Iá/�䳷 ����?̘�{�� ?6I�] v��@? ɿH�3$#�K!xp_�I]@�-li/��ߪ�0�����)R��ӽ���:������f���Jip� go4*|
���r�YF`��mP2-��[����/@9)0���0�H��A.���/5�\;��FT�|�Թ�i�l�皧�,���V��~���>��@R;�{ց�f�
��׉�n���L����:ciѬ���"��0ۑ]l�u���0c�v�|CƜ�\-�@�60��]0���-�f�Q�Ԫ��Y��O �w��P��rǆ��~����Ԙ�ar}Z� �۷��ϝ?y���'�v��Ҳ��^?wΦ�S�)�|����)D����-D�3\��bܽl�\
5�c�,�+�8��᝸�8$ƨ}`�9T�"�M4���á�(T!9�C
�90K�����hv�L4�Ab�zCq3�]����+������&%���eĝ��ȡ�ބ�W�m�|�v��,�~	�d�� �4ؖ%�5QY<IY8Y]<]V4U]2cĜ����a����q�ߗ6���o��\���}}���q��+p�_$(5,����d2<���;r���&Θ4i��cfhf�2sFF�d�̩�S��I��:��	O!�p�\N/��Q�����`�T����N���l�MNO�=:�ng�-ݲ�e��-���9u��K� �×.�����c'������ۚv����g�Yf�y�u{#��[��M��ɕ^��ۉ�g��0c:�����.��~ �	��6`��(�p7�����b��nWy��+[��M��gY�o�� �l� ��TVN�77̑��!�{��E� �3�80⧻��y���ibN�<�j p�F�~�P�<I_��	#{�A�����O�d�de���i�_�c}&���|��O�Lo���e0f�=�L�������Ϥ�|�"�y|��NV2�T�57O�֫�2
ҪE�t?�/����؂_3��:kJ�(��?Fz�����Möf���)󧬺��<ѵ�Ц	������{ڶ�޹�c󎎝���lo�zp{Ǿ-�[V�ʊ>+�/k[v�x���!uz�ɠ����gf�%/ޣ|��/~��p0�
��l���Z���F�*�)C��"q���:[���v<�SB/GZ�'��q5(��q`�2�`������.�W^�|@�٨~�� C�ٜ�b#�I���x��qG��C�U��ڜ�� fFq������	���"s���j�t��_��(�t�Q	 ���?�ƿ�@_��	f�'�9����6��K�?w_�A�^<6?<���2��@6��c�Gp������%�:����Kc�0�t��)�=L��V��������D��@�`,�t.H�#
�^�ի�n����x���tyoњ��J�ƙ�N/�7̳X�sf'8r�;r͋�]�w�x���բ�K�98l9��0���)܋tԇ��8�qիC>�*����Q1�ah{�4�``�ҼJT�?q��~&�jI��Ka�T~� �H`8�i=�q���E�*H���f� �u
� C��dL�Tv�? �"�P
�������l��wI0�}/�IϹ[�@����yS�PB��� ���$��d8�����O�M x��'���g����ǝ���w�L ��_��p�xp��`!��<sD<.���d�k<�I�j���,g�%�'w���"���*Ў��t��F���`�F��f�oS�S	R�K���c �)歼���%����C]��>�~q��'� �^&^^ �7�;��~~�m�A<�&Ѐ[�h�p!Az�T;�R�
f�B�t��J��$�	fP��g[Z�Y�~%��@2ζ�5�Y��{��x.&`	�`���$�Ӹz9h�_�?�ybw���$Q�7yT����T
�B�f$
��z�D2Y�n�dT/��׬q`��OP3����� �?�[�O@ ���>^t�{` ��������Ay�>�@/,)���s1���
xA<�o]P��mQ���~f����:;�5�O�������H�`P��(�����Dڇg��5�k8ӱ������,��W4�����S0t�
�F�{욒CR�3�.D����fhc���ܶ�,N����e���'�N%
�b��6��[(0�� ̠�!��*�cL���5�EB�I����]�u0��#��E
<D�C� ��2�q��]�_!7�@�����Ǻ�������Ո����'�:��5<������}~F���	��� _<���ۓ���I��~�g��+��O����o ���3 �\>���nf�3���U��b ��9���)> ���_�ɷ�?! Q�H���~R��q�I�f�+���k�d2�Z0|����c2�w�������f Ƕ�<�_���$uы�����0�v�7������eWc��"��A �K�cf^Ejh��0���P�_-0*Ͼ�y�x>{�����@T@]C0���}�M���`�Y����X��⍐����z�
�ե{gD�_=f�?���������p�3ָ��=����.�?n�����|�h�ށn^PN�jY���x�����#�mF�-#К�kS�����O�A���F5��z�I�9�g/7P��Ӭ�@�:�������Ӛ��,*?;N aܒ�Y��r����#A�f��t������2u{8�l���&XU� ��R��Ր
b
��q	$ r�Z��S ZWn�6H8�6��f(f�i��1D	(m��Q
E�?Aۃ���`r�Y�; F�K�^_9�C0�0�����>�ɘ~8����q�ss�p	����Ks�������>����{{1}���@�?����:�0�9
����:A7rCԽ�Q@� �=��K���!
Ɉ0RH>P�]�"x+褘�@� ��;�W��ϔF*܀��C���H��e�k^2�:!Fa��Q
=t9�.D�.0�*F-��H��]�X7o��Ǫ���"w��H�l�z���h�,�2�wm6�C��	W��#t� ���������6�@Y�,�&���`�~i���f���{�Cx`f�cb������}���/��A��?��۠8��$�?-�_�-q�y)�}�p�oEniW	�-U��*��k
�5����JrU���fe�?��$u�+�.�c@��QRi���$B�P�� �'8�VA�PDB �E��xbYO��Gz��|�CUG"�k_�F"_��`�J����[&W�d�˘�@ח�{hW���t�7|�]�p�p�
q�L�+�T��Lo��U'�ڂ��7����P��z�1pNpb��b��~yb\+j���&	`��:��:�Z��������{��)0CMy�L�l1W�d�H�yݳ���7�������Wq�8W�oEl#F8��Ӝ/��	�l)=7==�
�j��9Po� F��.�`� u��B��w�O|�8�D��y�J�po� �YŮ�Ts
`��TΔ����w!h�
�V�Wգ�5^�\v���ꞥG�V^ؚ���eRC.���jϷ:�yR '�N�ᕡE#�z]���^�p�sͅ�.�Zq�}���E��
�Y�`x���<��b ��$T
�Y�� ��Ć�ěF$�G�3E&à�Ar�>�2���w�`$�(�)V��9M�	C��#u��Ԕ���J��}u�
�@3��e����똊�j����XCf��I��Pti$hL��eR1-���\���$�S�zt�����{�L��[�����+6ݬ !M�1��&"���c�3π�(�V����y�%��R�"����w� ި,���o!l���Y�#�8]ܼ������-�-?�%ku�Vư���d_ ��"�&�Fsgȣ�Yg�'#�Zx5����֝ą�_�->�i��O��8����`?Lݻ�H0���I�koG+�� 1d�J�N��ۗ�//�,�?�Ɯ�G�p�2��� ���5G;{��z�3T��=���d�b��3)0�A_�·��~W��ޅ����"#�g��%��{���r��C�\=9V�KT[�=���*�����{햃i�2��Ab<�>����}I	�5TFߵ�A� 9���&�2�Xl���#R0���Oz���^���d��X�vAo�x/��{��D%��ɨ<����zS�~�*�WR��n5`>�j�i���&� ��������'�d��ÒoQ�R�ד'4\w����'����1-���֫$�1�G�:ǜ	�wPXT�E���#@���!$;#�8�4�5v���+t�s�
�9�?�6��~ߺ-�����fp���������|h	��SJ�s��7Vͯ�k���ٍ5�Ʋ����i:9境�O3�F�{���G̤�]�:�s����5��|�<"U70D,�RG�¯
��١v��th<$FH�0�z[�~9�.մ����V��Y�fM�pdzj��jwrvj��L)~�T�)�n3�x���rn6��U�l��=RgK��%�Ǒ�nN��MkRQ�En)������@��O�p$�	{ЉX�k�R��V�
�E��dUw�(�|Q�HJ��D�������7��_�? Ѝ2H$��@ώ'��D�'3�μ�0ï��K_� Wx��tQD�J|��^���@�ب� ��G�.ƻR���>�C N�W�TԻ�ԓ�;�	(��u0ct�Gīo	����E*Г�zE�e�y�K�����_�+VT��&�:�ع��RL��D�ȳD��%Vp�q��w_��k@������;�Q3��T�AI��펛�N,nӁ�0t��YS������TWVUUT�4,,��.��[�PWP]2�8�mT���(�b��M����{����w�ɀ;@X}s��%LP`fhZ��T��>�ס���=.��vs�|2Mb�!��K��ⅺXA^p�68RoM1�ɭ���1�g& ��"S������|A�6(Bj�
��q��,S,Ǟ�t ���)P/ط��?��N3��i�IB�#t7b(��#٥�L.��n�3$��w'`E �=�0z��xC	Oob�]�TT&���=<������'� @B��B�fޓ?6���3�u|�zs��C�)'��`�>���q�"*s��%�ܨ�������O`�a-�I3;�}�C�K�f�XǞ$�+t�o��Þ���0��3] ��(3���]&53K� ����ܴ�Nkj�OO�]�N�M�7`p�ECi��8�O�#�Λ,H���XX��
�H���.�_XZ[_YUS�P7kyu֜���W$�
���fh�^F|�Z�T0�>4��I-�&����
E�O@]1^D��5�ߌ�|�d6I�9�g��q����:��0h~Y̺�I[֋u���1��Ρ�e�ߪ>�Yui��Ҏ�K��^�3���!����E�T��
���鴘nPA]ʜ�r��R�mxʌ��:Ê�|H��n�[d���}�iq�����6�B��^�����N����[�z��.U��Rv�����	�@T7xxH�n���!z_��z�<��Q��O��	��=E7�{�P	�Ex
�3�@~�$��dy����+�0w�;��uC�7��*ҧW�e����t�Z9�&�M�\2�T��uW���{�y�u�k�r�,9X�4��=mÜ�ē�[���C�vܰA/�R'Z �A��<bd1���s����\WS�_][Y�������j��Uf�^���o9�"���Hw0l�f�xzR�������(��l9�x}�
��L[��9+��NӋs#���=kH!�Q�ac��-���%�f[�����	�:�^�G�h�A�G�n	�)��Ɛ'M�OZ��t�?�L��U|iG���㷷�.�Ot�I�!�p�6*�K+��K\�`~'��+$��%�5�";�47�<��
��0Qx��v��W8�È$
9������Ⱥ/�B�����Je�`R����Sْ��R���^�}Be|�{��K�!������=�S0�0c��s�$�л��	��M`�e�6^���6�ľ���!a�x�� H�N!���Dt��l���2� ��IUչW��#SF�X�O���&�*������]�Ubr�x���VХ`N���С�<I0?{��/�^oa[]>�z~Ue���:��[UW]��P]_QU>{Qy��B���H���������a`~�C&�R����Z���F���\�j��kS�ӄ��-�^��~}��݊;�7��o�'�mO|�9���g��O[#�ZB�Z����h	z�*z���=�E{��pH�5�~[��ք�[�w�(�v(/lr�}xy]�P7�(0{Xb}Kd��JOrͬ�C�e���d���n'��ݚ�eQC������d�'�jh]����!��U��I��Q�Z@�(�Ջꯤ�dPZ@�"�s�;���C������c�RY�dS�M~�}�
 ?Q�,!=f�4EpOȒw��Z�[��R��}0�=ܼ�տ����}0���t� �̳;�}0[��O����`άӳ�*�<1��mV��r/��9yS囻δ��V�����-rn�Y;k�y����<I`Q����;W/��f����wf64à7eW��-���(���u�⮬���.�����bZ��`��KYҩ-���Yd�ll�
��'dw=j3K7���ɠ;�1�y�ʶ���$�6r�%J�Hմs��;3�o?��ܾh�x��tok�Ӷ0@�Έ�["�l}�&z��<�lz�x~�
��#���(x�eG�����1O[��wJ.n��=z�*i��0A>���dX��Lɮ�4�9C�l D���Los��Y� K������y��GJH7Q(�%�!���D7��'ꋐ��*@2�Ad�^䐰��O��7���A�.)���dԵ��OHF�Yw�(�L�)T��v羚ս�s��y��sA���ȯ�}0d��8����F��
:��$@
͚�(�Ǭ�f�y�on*ìP4�!�$�G�r�9��o��]C��c�9ͦ����7�<�dxe��^��H�/�8$��̗P`�B�B���b(1G�[c���������jaE�����򪪚������2fO���Y�ў#]�3Y��;^�CB!�{�C��YI�1B��(͜H����u�+|�ilk
_���*cvl~���)�;v�=m�z��Y��UD����x��~����U��#�egpW��)���5�YK0��v�m��u{�͡:�n�G��H��#�X���q��'��2����$ΜC���4}f���?9�ۖH�Di�8�@�?��)'�(���}���D�f��	?Q��PJIgO�A�<0*x~EJ�M����P%�wŀ(�#Q%�����~�2���C�'�Y���3��$�S�'=ƭ�T����,��3?G�r��MM��V���\\g��[{�]�o�\�p��UL������ǉ����A����q��)�ΈuE��bG �^=w�ⱺlF�Y�nQ�$�Y`�I�:f*8`�fh0`�_�4�x��a������ڪ����J�K+��48"
���7�>��o�҉T��v}ǋ�B=*����\P�v?H��qx�Q<.+����؃jW�O�μ�=��%�uSț���͑]���iy�, �x@�o$zˀ�p�@o������0R��U[��֠7-�W-��§�  �뎨�QϷ(���i�jꬰ�\��@$,L���h���1�j�7<z@ib�D p`x{Y4������Q�~(�~��H	��0�,��^�Ki]x�L��!%����DN���#�W9H${�]I �^�
L��ʊD�W1��9FvX��"N���{\koFPE�J�{��n��OYο�o�g���v�f�c�K�k϶U_�{�e��20q�
�=����P�0�1��UN[=�d߲���&�nڔt�԰�.~���֓$��z43fP)�8�|L
�)+�dF~�̒�����֕�i(���j|�!�4llo;y@,N��-���;��F=9�3C�����&�rы��>6��6�_��Ú>/��]qq_��-�/�B����o7�m�z���-���gMA�V��^���9�EK�������3����G��]�/[C�u��/ۢ��=��ږ�y�j�X�Lf��/Z@/ೊ�R�t2� �-@��b/{"�hw��i���J���H���4�����w�`��eR��el��aP��`@��� POuhZ�)�{(0�K�R��f���8n���@��YqU�U쉳t���.�ds�O�O�5�By���Q�0a�X_�\�g�c���)(�H�&�T&	�+\�|9/�*Т�ɓ�[��Zಢ"h&o="�}���2�0��E#1�U��oQ�
���r��4�mP�`B��^�\X8$P+u�KeZ3Yy�p�p-���-V����u�-
�I퓓�'\�nH0)I͌���53�8A���cUHy٪$Ӹ��g,��S_�Y2=�<R����p�����C⯃��]]��q�s �l���jܭxЩ'pä�vdy�#P(氧��on�^߯���2�B4��M@AD{TW[�㖘'-����z�6 ���%
�h[�>�!MW[��Ψ;[�vF=m�|��M���a�{?m�|ڙ�3�Zk����k��s��y�`1lR�Y�O�f�Ǒ�aOŵ+6J�����{v)��^58�#���r�\1#O*�W��G�i����%ˠB,,��D��"��Ô�i�x�V��NA+Pp4"mf\T�I`^*�"��p�Η;����Q�T3<8z�",H��Ӡ0k\s:�
�&� ��|��3|�Ӑ�GX�ޜ^!�g�놆�g���)�� �ТʲB�HS�]y��D�� 3���:|��t��N��8W"�)�ˊ��Џ�W�/���g�"�3�w��0 �Y��g�m�^f\��[(g�/��y�=����<��L����|E�#`�!�f���@+�p�)N���� �g���"��� G��aH0k<�j�S�p�(ݭ���L�0s�P+{g��ږ�G;�O:�o ���$o䃫��3�I{ȣM�ǫ鏗��XN#���`P����Ekx/�����)�����m1uH���Oo�"_��#w �?mz��}c5o���n�!���W���f�*��H{P���^����D��Ǣ��B2�b`���u�u��x�n�Lˢ����.��gM �G ��yp!m�@��$@�pe~R�Q������7?_ll�x��i�T����[��٘J!907-�4T5w��R�iY�qѼE���Ѻ!�������u�x�+d9��"2M���x�8Ϡ�,�63���Ĳh~^��1զĒ	�9]+�Y���k0��80B���{� *Fw���h��@Ǫ=���f�0��O�2��ڱ��Mi�Eg� �5`n����sb�8����
 ͉'_[TGÞ�g���+�kPC�-V:؍N�7,0y<95���������N��b*f�9@�]�	O0�J��-��dR쌀�d��)�o>l{�5��r#���/��[���=i�<\�p��ӥ��W���P��=�}��Z��<o�#u7��
?=o���:"�v�>�z�!$�3�/��]-ض"rz�`�A�i��*J�7��d�R�*�$�M����3����� A�
��et�:ܴ�I�km�%f7�ͩ�?�aAђ2��9�+񶱁� �X�ȍ.��AЧ��J�Uퟟ��k�sg�4Κ��z^m���yՍU��eWY�>c��xd�7�W��ex��,\�5�\gZQ6ke�܅�sj,X^c[2r�UR<�����u@2�Q>p��J�8Q aΐ�fO�Ve�������jq͂�U3�W��R�f�b��׿5��Nv����A&��,�:0�����ηD���i�cb�ROڽ�8[%�lP��voS��17S
P�%�+`���.��r�йr�~�*u6�q��C��G{��#�ņ&nr� �_3)���h��a���ZH�OR����R�I�exX2!� d��}v��[�qDG��Ȯ��nU�,x�%�m�����U�����_��t%�M�hG���-�$�E�C��]R?�i�I4E��m�3��Г6���#u���G��W�-_��lb��C\I��FM��H.#�:z��x��ʄo&��0��}fp��]�̕6����Z��r���ꅵյU�uU���˖�--5�@��/xK��?�<��!ױi�`)�L�-_0wi킪�%�˫W�T7T�[^]�hNg�pC�zJH��,��#��W�Wm�.+���z������r(@ѱ�tB�1ԐᝍJ�@��r��a�%�G�f�_\U�XWV���tAUeyYu9<�//M�5��+g��5��C�]$��)\��LP��jд���.ť��2���=�U��UE��� ��Ӻ�R�o����c��	E�����7��w�
�_���V�p+y�gّl�K��3��wMu� �gF���`Ƒ^���3���@{��q��-�ä�K�rX7I�mI~k�z�����5-ގPP�D�����K��,�|����:��e��=���Hn��n�9Id�6@r0(�78���)
�u3�������!�o��~���9��aW���Dig�Hg[�gQ��%�f�L��q	t�PAP�P/�K_��7�ޠ$Q9 YeХB+�4`[-(] �(--��V�TUU @1��fif��&�(̔qY!�1ʯ���c6��>sYUi]uuyE���ť5������՗�^U3����;�,Edy��[�gT0�i%�m��f-�*���,�X\Y�XYW]Y5���x��#�tCz���C{,m��P�b����5�+��c�����u���k����]��*��8�p,Ө���_O�,��\��fv3��1x�!�B5��{����uI�����̤p3b	���1�A͢:%�wa,�ԫ}fn��M��+�jZ��h��q�pZR|L$�0³�7�J��䠍�7�F
̔:%��;��p��
N��F�9@ZcM����4)���T�쁡�6	���6��4�^t� ���D�n�}�QD�����{�������<AK�!�:rAI��HS��`�X�M�`l�O�z��Z�����m~��3�eG䳎�7���|�tНe�uu�q�pW�x`�ĥ0�fNd����23����g�W��2D�JR�=�i�@����_<���� Oc#���V��\Pe���f/*?_��&�3�6��#;Phn_���W�K&��WV,�_�PV��aqC�ª���5�s+f.*SYƳ�ݦ%����g���<�z[�Ҋ9եuU�K��̭\T��^X?��,����l9G��	�E(	�'fU��N*<Ocn��uMu%V�����faE��Ҫ��5�j�WVh*�
��
�?A(���A��W�BQ8�`Ó���#Vq��!͌��K�ĀO�
t/ >С���| ��zQ:4�봈y�+�n?!^��&��
r��_�^ �TB���'�槉��J �Z%��l������R�V���1��|B�\x �+td��Ďo'�8��$�a��'��cv�M��b�F͏��C���Z9�6�����=�Es��MQD{��M��+��.uFZ��f��֌�j�s�~�6�{��`&��{����=�qG��v��ָWM�/7E���Z�����f���O�/��fQ��	�<��;��J䁖DP�^���=`N���y��XD�G��II
N��x��XedAf�2pqA�?���eUu5�kk*�K+j+��jkf�)��{��9P`�~���Y93W�*K��+��*k�+k�U�.ZTZW;���䡎��ѹ%�[t�6�0-J�9�3�*jjj�����+k�Π��t~EuM��yK�m+�G�k@��1m�ŀ����l�I�(�L�����������4sMUm}mCMy��ʆŕ�`,/,]gcq��'��O���P����S7�������ψWO=~D��Jt�%�_$^!\&�]!]%�"��&����#�[ģ�����	�>�����3��5��3/?�ۢ+ �����DPe�43jc܇�+
���gk��:J/�e��T�pikګ�W`T���l�{�!�٦�o�S^l�|�B��.r~�xЋENO��i�Bʧma�I ��Q�Rc]��3&��Ll��2�����j�|^tK9��8�4�v�U�ϖ {�i$�Ӡ�R��,r �\ݙ��'��~͌�٦�2op�5.v�A�sb�}hI}em����J�����VV�VՖͯ�_��a~y�����{��p�ɝ�����h� ����>�<waCu������:�P��Ҋ�E��+j�UTT�X�)��0��0�� �׀�4P���N�8Z�D�+�5�.���[P�XW[Q����lɲ����UÃF���/�Ѫ����~����,^��j�Rh��F�,++�)]XY����vA)P�r�������l\M![���8Wj����q)�a��#�
YX��CȢ����/'~��ޛ.� ���� �׈�w����緉�w���W� ����%�d@��W��K ������ě+��YF�X�g{�%����F����fҕB;�ݖB���M�-	#gG\ޙ�%]�MB0�ߴſj��9�醐7�!D+���WK\^.v�Z���Y�#�		濃������3� �_���Bxw-a ��$�{�z�"��x��.Ϫ]X��cxٓ��7�4VМ�kʄz�YpUY� f���Wூ��f���(=m�]��������fYeeuM qIeE]}}mu��U��u�N�[�ԧ������K�(�݆�#��T�]E3�8C��9�-)���^U5��rnÒ���C,llXR^]e���,���y�,T�*f��M.�;TmV��#��#�\j�_� @俲TrUEY���`�Wה�5T,�\�Xm]>��-��X�fU��>��=��U�����p�P��ҹ����UV,�F �7,�n�쏪��������"�݄�gq�j�2{\KR�(����2�vhqn�yl�ud�mx�ux�yh�ex�ud�yt�yt�	�#��P���h �����6��1����G6-�Itu^=�֧C��_`�^�Ji�n0���ņ�@I��Ӛ�a��,kb�Yxl����_l��{�*z�"�a玈���Oۅ/۹�Wzt-s{����r_�I�
g��r8��] �W��7�,퇛��o	~��������7�T�ȗmQ@��Z`�f��k����<�,ܾ,>Z�w�$����[�ݸ%�����($����d�}�h�x�rIr/J���JgΫ_^V��X���j��9����**A?ϯ�t��e��o
0�@���K�D��.Nm2�I7gF�ǘ��Ϋ�_^?��qAE�����*�W�.�W��ܸ��Mc��mI�'�)g�Bw@r3�5����������*�.�F�������5�U.��[X��:�,�e�w��ˬ�3i�r����6��ʀAN��'�(��0���}����A��Օ�/�aA����Yb�(r�L��8�k���Q�Ÿ���H_��?�k0�����۷�Wq�Q�<5��3�Q>t8��%����!{1p/�`�qH ]8ݨ
0�Ӎ�|����:�rѱ6�|��O+�F�&���|�iolH4#q:����,�YA���脫��o�R=���6ы�<����o��=n�h�>^��t�۳%�/���Y�{�0��+I�u��& 0��|gk���`�#H0w/�`O���
��)����%�.�1n���`]��)��!��3�c��d��%U !(F�`3gV�E��P����k�&Y�Y-�]�e]Uy(Rp���W5�te�gU��yCX2�Iΰg�K�K�)��.�iMc�p �a���7gU��E �Y�5.��l��_WU��vN�<լ���D���ќh�*��.h�0+�v,Ô��[W>{�����,i�����_�,]\?��Xh���1�u�}�6%ʡ����,�ڗ�;|��y�u��������K�J��jX0{���s���,��[/�ܨ�q f�A�|�@��4�����o�E-)���K${Rh�P)�U0|)Fl��b�3�Ab�pU�	w��S���s/���h�2�Joc2��k���*�Ȣ苁G��KA���[�R�-���$	҇�ϋ<�s���hP���^n
��
�h+�m;����K]_4��l�z��	J�mktbA���QHq�>�~�d T���^�B���uK0Ы!��7�E���)��:ΣEN�W�;�$�0����6	(g�I��l_�$lZ 65!�U&|!g��.j0�l���LI^�h_[��)���ʜ��W��5�UU����z�����W̙\���ֻ@죗���}��@c*�,�[%~�@�`� �Pr-CG��̍��V�)[UZSY���za��t�W1N"��O��è��)|��t3�j���F�N)��_[�`ѬʆY��fWϮ�//_V�Wk�&�t�31�A�ŵO {��$7s��Q�]�v-�{ꓳ�fXfbwPY[ZY��p�l��S�u��u)�0m*�-���.y������T+ �'��g3[q��{�x�lK��~f/��&��8((Xt��h�'��ꔑ.V����V0���_#�,=�B����I�Tm���o'�I8�H�ܹ^0C����M2�q�D�_�V	�����'�	DG��MϚ�^�
߶�f�˕�/{�l�{�8�r�
Ш� u����H�gLC%{��Ն+7��a&ׁ���Lѫ6�����U�ig6E��E���O�M�b�`Rc�C'�f܌�}�	ň\qY���èmV9M�̷˙:	� ]0#=�djA�aNEq}ce��]�cbY~�A����-�B�2��-�kJ�05�4'��)`�����#�h�e�����[U��:gA�vZ�vW楹�[)���J��x^͚ζi躴@�\�@kk�Rb3}V��¹5%����&�Ӧ�F������G�������ծv��z����<i4GhH#2�3�&��6/��*���ZR�+����kJg�'��4�4�@�0(-*j"�r�ɒ�D���"�ɀ~�c�3��ӊq�i%J?h+Ί�Ę��Ol깏�K|l��H��9�i�M�Ɋ�-�-�X�.T���fFSj��o���p%6� �kN�[��bQA����䏶��mJ~�1�M� ����j	y��|}г5�g���kh o�9�]H�?�	'T�=�kNȟЮ=���M��;�i;E��qG(��O;D/:D�[��V�n-8�J��!Tb���A�Ж)��Xpi*N��Z����/���.��3������A9�i� �hVN�pzz�g���sj�
�*�3ƅM�2x��9r�TY�6�Q���'W+K���~�it�`tӺ?��-V�*$;#~r�y�����`�U�3.6{|����-_���R��=�JW��T�NdЄ�������iCC������6���r^͂�S�B��s��}g�,�1�{z2u^
�y�e0Ώ�Դ)ת���3�3FL��*���sf*�ǅNW2'%�A&�@�gk��)D�2� {�g�������ԋ� �h�Hd�W�9��A\�A�nmL�*��=R��9.V�&�+ǒ>m���ģ�_�A��q�M�ዿ��o%JXQq�	`���foc�,��{���e�g���#�Y�w���&{ڜ�|.�z���9����g-�]C�V�-���o�/����E@$�)Hw�Q��0&��i^�S`&i���H��Ig���(��vE�i��^pdUТj��<?�!8@�bX|`�2�}���� a��C��������h8֑e';��/9�n*/�Xp�eչm+���_��tU�򃛗��Qsv����v,:ѹ���i��L7�حD����Cԟn)=����s�k�n�<޴�d��KWVֵ4,;�i��֚��/n�9Ӿ�|G��u�u9�x��+CJPڦm�'��No.=�e��}O�?�y���E�k/�]��i�]U'�W��Q{fG���On�<�V�W1�
]��һHΛ5��T���ғͥګ.t�kY�c��%���5�8���Ԗڳ��O�U�i�:�\}�e�B�=�U'�� qD��e�'5��[���3'��p�+���n6	�hL�j��/бBz#��A�$�B)�U��]�)�*�"c�9�@3w-���B�u=�w�w`F�a��n0��K*��8YE,cBX7�|�Ρ�vg< �x��MG��qg��خ�ؗ�`?��z������V1���h69��j�9��Aj�����Q��`���tu��Y� Wq����-�~K��}͒�ˣ�e|q�o�6r6Y)Ka�3�j���
�#��B���\�	�C�8���`��ǉ�W��W��ǉ�G�{�q��������ܰ���q�:�u�x~�xW��F<^z��oT�)�j������*��k��9�8C��@������#�>��i��CZn��w.O����// ���S:��Ge�Ȳ)6���xr�xpOhx�/]7���55\xt��ޅL.o./@�$s�=.����,��?�2��6A����<�����ŭ};ڗnn^�xr�xy�xs�xu�xs��t���t= ��Ϩ,��ID
$r�w���x�-D���`���	�g���*Ͽ�s�}0S�Vl�$�"�(�'F<�Q���T8v4�<HE�ΕV��)�7οEt�8���$���V��<$�p��ی>3��@@0��l�#�0���H;o�z����;1w��w �AmF=!u�֐�-��Gm�W8X��%�U3\�ߴ�	?k~�5�Us�˦`p��	gPѯZ�/�8/��/Z�:B�F�mO��Es�9��<f����K�1����@s2Y}���J��Y`�2i\���q�Y���,��3Ϥ�W�^y��j<�2x�*�@��;%I1%�j������lĤ��i���i������̓ĕU7���%<���C��6d�/��A���O��NIO����Qg�KX^���<��bR�䘤�q1S��s�D�aZU}�x0e�,�%o}
8h�V	X�o�9J\�*�y��Y�����O��h_9s���z��ԑ1ʼ��32�'*�e�r�q=8/�mJ��`�3�Ϛr� �lk��,#%oh����1�	�3��XYضr���i�ǧ�M͌�2cX�n�E�Y����;0��e ���^0c��j0w����~��`�(/���IB�g�=�5�ԈÀg�y��18	� ���4���Hn�2��$���ux���c�6�p���3�dR_����݂8x�F>��8��Pqr(\l)�IC�X/(�M8�c������[/�D/�0l��Έ7��W�'͂���g��r#�Z7#hq8�5�yShWS �Ugԛ-1�뫶�ם!��Eo�DDG���#��v�ѝYuk�W0���5+�sR�lX0;X��`S��Y�������~f��=�ÑHV�}|+��b�@��	�`����[�D�V~�x��������Iq����Zs�Ț���o(j�4��ސ>]�X�ɕ�>K:Eܫ��B�Iᙆ�u�}zd����i+�Tq�u�|�/���qp����]늚7�LL�I2d2s�g4νB���z>���Ke��Xq�V�q��1�:_+1�"�DN�5�c��/��vd偖Y�[�XS4N�719B���Yz�	�Z�^`��S�v�挄9S/��nj���DNIL���q�ɣu���\�W�u���uެ�<q�,� =p�$i��K�Ӫ�k�Z3n"�3�b�#7�`���������[�����|����$�}�Ԇu�������e�� �՞ `��^��oSql�:�v4`h6e�Y��
��u���k��G�������#���|2�����Ҷğ(���P��K\�$�V����4BϮ��8�C}e[ʽ�	�;�5G>j��^8e���-�i{ԳΘ�ѯ���[�����u\�"��?$�r���ꈸ�~�%�NgʕͲc��k7(>+���s���4o��אI+�l�X����6�)I�L3(A� �n��oR�
0����Dr&tp��?��4s"ː*Ȗ�!^6���L1C�aK���N�X|y{��ݵ��[6�2��-j�Z>jfF������A��v�%����ϕ2
�zi��y׈'CʧF�%���}����k��\t���D��]+,[�9��)Zj-��5�es�/G-��}��n��
d����7�8���`FZX^�cI��W>_wa����.�߱Ұ}SẦ��|�� _�t��I�>ǀ;��b�"����ٓ���l
���=�eo��k�喝����֢�,k��-�Zf�C�,j(�U�i�^ 3
3	f��A3#��d(Bl�9�YSek���_�� �ċ��	^�{{]0KbKF[a񵩽�4�V�%�#?5Ц���r��LW3n�r��⡍`e���@t�?�.���)��O��W>��Dr �J�C>G���yujo�[�£P�K�ύ�#��t�JS�ܥ�֖�+�2�>j�~�z�=����Ǜ�O�b7�?��lSX�oZCހ����<o���@ڢ���iK��U}~�����_�5/>��2��h6<�:p��a���oЈ�������Ϥ�7j Ơ���|w�� O�8����H��#�D���?Ӕ7O�]ti��;���[i���G6���5l�dZ�jL/H�����.�!�hAk�P����`�b]bv\�������_{y_��KN�/��2�}��s���c�c�6aj���|�x8r������Щ1-�9ö_�t���ԜaSL>x����E綔���pco͑����Wk�n4-k�e.�Uo���q�n��\��n�(��ƃ_ӱ6n��r�ܓ��<����֚�W^�\t���웛l�3�V�"f$��F�"���Y�. 59 �����|*�( N
�R3w�}��4���/'�Vq��ċ����4v\u�;Z�&颋��dZ5�y)\�&�tr̼qq&$�NJ��hQA��h<r<k/��W��|��Zs�L�@<�c8u��;�b�8i��c�H�B�PO ���4��mWr,� ��G�J�'�jåzn����*d_����!g��b���f��-�[ew���ݜ|�s�����7'<�|�#�Ng��-����׶+/mO?�Ssr��C�,��)u�0m��eJB8i��s7H�x�b�g1�f�#�k`E�D
���%�H�s�'�8P��!��1�[��g��߄'r��zuH�H ��d�ć�̾s�qo���Mg�&�isp��d�cmc��)o�O��&^�]���0����,}s��볪�KF�:�u�|��恂k��OwN۵aԑΩG7|�o���S?���]a�N<���oU������هs��u�;�œ��l-�p�~g���>�]�7w�oj���U��-c�m���5;zFd��-���,��,�B��|L�9���Z5����f��c~t�����W�Y�o�Z>���aG�F�\;b�v}n�P�V��xԸk=��]E��N��2�����f��6�o< ��`Ƶ�`�B�:�9����8�Ұ��SV�$�!A�;E<<M<�Mȓ0�Jj����f7�#�[��"%����Ǆ#C��$�����8C��A^�(9�O��&���> c���Brt�%Nh��ԅ�hEY���q%���F�o�k��C{�}�o�{F��5�Ԯ!_l��bg։�#��wp����֬W֮��%��lE��u�"�`�)�_�Ƌ�Q�d!ϝ��!%ަx�1�iJ��Rӿ8X]�-����H���_J̙�$}o$�KAq#4f x��ϕ�"n���*{f��#�yt4��!�͝��'�ol�_�»�Kti��lG���tR�1�f��}�H��͐��$׮��N��Ui�w�=�O~wO�ˣQ����<8q~3���[[�.n�b_\� �K���Yf����c�~-P+k���:q&}:���i��=��u$����om��¼�H��樝G��s�_w���Ӄ��
����9cn��w�*mL9v��C	���>;�|���A�v���]�puK�ѭ��;��0Fw������x�:���Z0�4��يK�n�'�ŕ`p�^'�,�ˮ-��k5���(i�s(�t�l�ѕg��չ|���C'֫O�0Oo��455�S�w�
�������?s�3o]Lz�� ���Fº�|���0ݑ��6�V$��v�+�z��e���q �]����l�*�3D�e�Mp�g�Λ�='hJ�`��=L��hY�<�$���	5Dr�qtS��%�ϒ�c���0L�C_�l�B�w�ҬI��eL���Y���.��h���ָ�2�U�3�8��h�Vz����d��"��^q�~���~O��?<�`?��>ڣ���h�r�<�[���=G�m�������Z4I�5�U��_Y���kZ ۱s���/�=������������<���t?��.��C!��m\1s�K��Qkgy�2�%.���v{ǹ�ԓ��1��ި���G����}v�{o����컻��pn�:z(+��:zr���g�o�ǒA�e���⡷�[�[�K��x4��~n���/w�����b�g���/z<;���/�cψ���g��E=`�|f\���3����r���Q�[� ���3�0`4xʍgP\"8֗g�C�T�K
7��/2i }r���cemN@>�����$�=e7��$�����u�fV�gڙz�o�=U Z��tg38�j�7H��P���<X���XFY�h�����W0[�� ��D���N$�� {�I�0%���\}�@�*�&$
uq|C4��2Ek�装�X|�O���Dx�fJ4��(��{l ��?AYx�v4�ޞ���i��9���e�V�NLeKv^�B��O =$p�&�%	�ex�����/0/9Y;�$��	�˟�J|�3�ၸ�{#o�/�����;"�P�7^:�{���xy';/�cP���l�>;��!q�<��S���<<�|�@НC�GB��|�7������cn�M��W�a�lv]�5���E�zz73�#nw��q��!���'�W�e�ۑ�����8 �n���3�������N�P�=rj���C��DD+�� �<u��;ĝu��V�O�z�����{c��!w������#|�?�̎���3��#w����|f0<�݇�S$�����[���&0�[,9���-�|fh
̠��&�Y�q徕�MY����Xryk@Aݢ�.u�x�X��)� �rw��^�A�+�E<0s�[�j��Xyrҋ�A�v f��tW���(q�Cũ�k�rQ)��"0��C43�#�s������R�L��1�!Ep����sd���]_�+|^�(D�9@�S�M�pP�J&��C$�8��	�Q_���>A}�K_����]���)��gR��ҽ���_���;5'��4��9�Ɏ1�����w��Y��ӎoH:ٔx�)eW[��xJ�i�֢K�y9Y|���� ��L����$�l�u���q���îJ�u4�����m�s�R�4���$>�A��sd�.�Ѡ��yy]�`�ؑ�1i���\yqB>��nی�G�o�ww��'�'<�?��Ɣ�mi���?oJ�ݪ�k���}��lQN� �=mp�4g,8nKZ�&�~q�pa��{Fv��tϨۻ���9���{�G�U����ă�=�Zb��*@A�R��> �5$
߅H��7��׸h�:l�R C�*uW7� }A<>�+x�vT�>0+CC�cKǁ�L��P�Z䞆4f�W~��`��̨�@RJ�@-{��
�酙�60M�ʐ�/K��7?��p!$Z�$jy	�ES��d�{B��)	2�8�����i�ӏ<�Lh��dnT�PT��� �(s�j�����^�ʯ@_M�^��_��L~�ڏA�у8pۧ�Њ�����T�,=�y'����"rcWt��-����h����{;f�X�wp�gG�}��yjk{�g��)������g����Ǡ��k�.��V�q����������;�l�����6L;�f���ڍى�Q9�̐��n0�?X:u�ç_\�-HȮ�:�Ŝ{��v������8���c�Z3���	�[�'�ķ\�y���2��Fn��3I��?G��ڱ6jRĦ��.�{���f��9���Ck�j��o��c�������J����C�>�Ww=���r}�@�Q����g�2yxڣ�IF��D�,?��ט�^�`Wz@�B���������`�}v�_I�؃�<$�Y��u��琻;� 9�������"����`�j-Pn ��r�"Uz�B�oy8��ER�b�K1f�A�4��n�-{��z�� u�Ir_7�u����ګc{^De���ۈJI���U޽�]`�[�{��0�J�c��{XRh&�2�f�W��r�xQvvsD�2o����n�-�9����qK��%Eg��ά��[m\�Ѣ���0Yq�x	`�g��3��}�"������S7�+|th������럶/�����E���N/+<�inN������3ēQ�mL� �E��e�27_?u��MA~�Ěrt��G;Ko+}���Ag��UEgV�O.5]Zc߲ޖR����.��x 5r��q�Т7>f���ī���u����E�k�o^��u���UgV�<��rd�����e���&��0�2��?�8��+�^�O�!���C 4	��d"}��@dL�X�
5�	<����6%@�2Fu(L��I�3�'���X7�!���w���?�e��<���mLcg���hHOx����h���
9�7�����Ǩ*ɵk�P���� ��N�J�GAzz��iF�@��"箁 %�q5
Z�t�O�M�S�"�9ִ�W�������H�EEQs��7�j��+������W��y�d�5G��J��mȌ�q�xQsb{�t�fRJ���cv��7cخIM�ĝc��c$��,�<.<a���tѥ=�<5�0���M����<�`�
}tn�ۘ��]y��Msx���Ǯ�^=J�6>�fJ�Pc&`�`q�u���%V^�h�m�@C���珿��̗�祬�;m�ԌC�G�1�@Ψ�q�Må�cǦ��j"�%LC��KO�`��Q`�1Kc�M�H��ܵN��2Ԫ^c�wʨ#�'�<i���#2���� [<Yfɓ��'e\�Os��P��Q�H ľ6[��dK��i�w:�'��*�85οPŘ�����i�3��� ���w�f�n�H��f*`���*��]�坝�1hX��6�������hx��.�_�橃��*�Ws�H�%<�4܂L�V�	6*%(���G cIRC�0�|%G�$�k�EA^fPn�07����f�����	_apU8�@�~B�Y���"(����3�~����J=�[x����-��Xl�F�e�
��+Xz��
7�9�0�ݖ�Q,a�d��;��`oGeg\"^,9�/vJ�|�`E��>�����u�ѿ�3�}����#~�G��>C2�⩱��$'��Wv��.�R�0��ڵ�.��,Ώ��T0Y�����c~��	?������d}�㑿� �O?O�i�EE��NXjck�`L����P��:��9���@���WGd|����ḣ?�_}2?�ב�T��>#B��s��|E˅����t���&������N�N�,߲���,�,q�����|�O<��/�|����S��8�O?���={�4���`�)� �!�90o|���ˁ!#��Az5߈��\Lb����nF1�ӓ��D5��~�Ɋ|�t��C�
�gŴ�`ېm�ŋ������y���m�����ۇ��>�����Hp�;��ko_���@<�HܹLܺNܼ���5��e��Y<�����s����_!�x��z�,��,��"��ʛg����~�x|�x9_D�<�l�a�ҷ�$o������@��s�
QoQ������`��"�K~�1E���/�}p���$�#�m�yL`V���y�ޅJ�"�_�B�#�D<Yr~{��jb�:�/�Of����_���>� �?�3�}���L�H��-9F<���������C�fZ_�ͪɋ˖L����f������G�~�9�u����d��O�'?����׫r��\"�[� 38��~&M��'�]����y�s�������~4�X�a��3�X�����囒#�f�m9��q�k�xZSi�PTɳ&�"^Vn^*�Ksd~���e}�%�a��?�3����?���ÇE�f'F����_ܢ��!|� H��H0P�C��k�$�6m|�[~<����{cLS�38x�`�6Z�="��p��W���ݑ�6P�����n]�q���
��ۯ�}����Ǐ�=~��qד�@����z�����{�Pz���[���~}�� �͋��3ĭ��Fx��i��O>�n ��/��z��ƫg�_�����î�=����ݗ����H�l�x���Ç�Ç�t=}��Y/=����H�B!��>��z�t�u��O�۳�O��
� u��k%zԅD~���Ӈ@o߼:��zP��I���C:�0�ӚZ �����13�T�+��l��?{�A���e`ٶ��o�j/o����J�mg(�`���,NA�aU�5���zst�b�gI�q;c�N�<�3l�����Mc��&���椀���d��e��"/�0�e;bX�׏�~~��������.O�]?n�vԞ�dp���Ó6LL�=M>%^�Sm>`��3���)�4k:C�J+0�B�l�D��/�5a[��}�����Ҝ��9"m�U�T��lux�4�:���?̯n�rΒ	��r8���"��>��4*�_ٶ�8Ǵ��,i>v�853��Jf�g����$;�=�/���Ʌ���sĝ���luX�:f�&f�L���䱣E�(QP�(,4828844�̈	�ń3�D�H!O9"-~�**[������|S�1dEOMQ�
	
���D���(�!�ʎ
�E�#��"~�0L?N1�`h�N#�&�N(�z2�}<=���=���}=�<�ݼ��=�<=�<<]ܽ�)rs������#Sc�H�GȢ��A��G�"�Ib��%�Ŧų�LH��6��s��3d��������{��z��yz�xy���L�-q��M�����;�R�ɑ3R���i��NM��ew��-�;m���^yb��c��h��c}Y����⃨������3�d�n�P����1��8(O)�����u�v-|�������4f�]���ļ}M�h�`�us�̹L����czb� �r�A��ҡ3/�r�RN~x����G�\�~�s���5_�-�|q�U�/+�;oJt%zŦK�N7����TM�)PȊ�o�u�`�A��{����Yw}Gō���:�^n;�`=�l��e�r3E�����׈��`������г�� rT)���s4����w� .�S���pE4�Uv(��S��(��}3�*<Ԩ��{�DՑ�>pd�,"��S�T� W���O�Kzӹ1��p=�����<~���~A\ $+*�;��?X2.-X�A�cd9/�:fd+XC����|��'�B�@���Y!Bf���>/�ˌత��Ib�I-Ц��~����ۭ������@�AN�;��r�AnN�\�9�pq���o�K���?��'����@���������� H0ȩ��S?7��nN���MN����ݽo�~:pvT�yy�40��xKg�6��˖�0�F�J��ϴ��ʔ��6�<ܺ�ek�ֺ�k�N4�=�������3�7Lg�'
��G���W���dl���(������U�	"��*�&�Z8���ګ��O۫��_[Wr~��̢��Kl{W'j�\y�� ��K�og���f���)�^?q��K���oZg��i��m����l�9�l��e���<�tnuY.+'�ߨ�t��i�6WQ`V2u��noʶ����	���<h){����7Z�[l�����¢�u{�dp4��#��'���w{�s�("UJ:Ѫp��d�������ߞ�4O�b���~%�~�X��O��fh��|�)�Q�X���bq�o�&`�C��#��� t�lA8G 䋸B+H�	8�\=����'�Y�t_3��c��&���l�  ��	� � rqD �5H(r��_$'Pɜ�����W�O��ͭ/ ��2�����ǀ��<��tq��<��i���������k?�A���[N�t�� ��O\}�< ~rr�r���A$AV.���\�tu4������ˀO���k?�@N�k�8��&GG��U�@7X
f��#ן�=1m�������G#~�gү<�}����a�$����C���2).a��,qo��N^��eI�6cH`�Qa�P�Ɉ���I��)2�'?�>��g\�>�~������A��?�(mLl�>4��ըe%Ё��dáS�g�q�؅緂�d�ӓ&G�������>� J2�����ϲ~�g���	7=-�4d����l�|f�?���$M�;��aˊ��Y�E+��g�O���Ϙ����>��g���d|�'�Ͽ��6=9b����f6G�8�����8�Hj\�>�To��|�ܞ�a.À��zC/nCoy�1�l��.T{��~�����18��`&�߁�=��}	�<�!���I|���J��0�`&72((<���pB �~��C
��_XX����p��EA�|�`�gZ�3��8���N��(�� `$}��$�r���@2�m@�(X��z����1!U��Џ}}���<ȳ��ǀA��
��r�5����������������{��7�RgW � W���V����wq��7��@ �3&v�tq�vq��L +���=@Q�����@g�}�?�9p���/��A�|zT��lCT#C���lO���:N������g�~������اϴ��x,��?U~�'��w�g�iS��/m��1,os�ٔ�6�]#�Y�OK��@������d�G���h���>}���ϔ_�I�M�cG����|��ˊ�������iv^?u��f�t�db���#>���>}����?�є��t�/>��q����l���mg�]"�?\`����xY��(����Q���L�E��?��M����|����G��SBY��`&�f㑮���$�qY�ehZ���I�ɓ
dF��)�fOw׉K4``��v��.���+�fx���`>LܼD�
ɒ�c�"���<NH� 8�' �X&2�e�;���<n4������!.K���z%
C�����q"��|!��P!/X��K��(����q�688�(�F��Rh1a�t��뀿� ���sw�����s_���`]h���us @t+��@��T:�2�
���px��:���}���K?�ᮐ#�dg�J�O��7׾���}�'N�H%���b �O=�&�O0@�dVP��3�牗 ��I��I�q,[���17�s^��\�g1˵���8<�w���Ϥ�qjj7�@�0�pE�MhTg��u�x2�>7iZ��`S\@I����>��7��(	����x����#b���E������,#t(� ��=�U��e�|�Ȱ��	g���BY�Jn6΀���Sc�eك#�[��9�`F{� ��`>O<nh^���2yj�%�6�5b�h%!l��W�w��y��c�s%q�#�s�z��X4.Ѐ�C(0c�9m2yD��<�_�4���P��y)x*�C�W�"��0O� ��s~���u��t�#�A� �(0�!�g�����`nH��`
~�Y�es�Y�86+�ˈ�1b9��,F2����&�xQlN0���k��$E�"� 6�dD2���D�V���w��4�Ŋ�c��~����B�A�^<�_���x�x��������|��\�,������n�ß�{|������g�������X��O��~N?!{���W��W>�/;�/�?Cb��_�] �$����=���W����1��1�1�Όn0C�)038�:]y�x^wnK�d��=Ko�]�hg�íUOwU�n�s�:��2����k��o(���8Y����F��e�S#(0[j�F7�O*{�P�m��vW?س�k��˫*ή�z��S����JV��ɕ��-up
́&qC���u�ċA�kv��Z~g[��ݍw;*tT�_i�b���2����;����Fd� ��w�zɰ�=m0v��kī�;6(��s��Ҟ������?ܼ�zsÁ����Vj?_in[i�P1!ڔq�?vj��x
�����p�b`�������6�+���ե��3�V�g�~5��䮩w`�*��w�L.����7/���	��p�H^������#�Y�y3'{~��?���3_�����c'38Q����Y!\f0�s�0i���ֵ�H�aq$l�0Z�X�	�~�|��z�M�����?2���b%s��\v�*�>��~
��Ӏ�}����w�n���\��X39qӤ�։Q��ö��:�mb؆���֤�ي�2��
��
��2�²�E����U�u�����������9QmC��C��!��	-��O�I��J?R��׾�ȵ�_������@C3��
SO��� �G0
����'g�t҃��?\z�М#Gf><���ҶV��N[�MM�m;g�Y����z�xXe7;O�3��A�R0��W�]'�V�3s�aϾ����������궴�lX�ۺձqS��-���L�7L��~�x>|�� �F�M��W�}z&)_��̢'�O�w����� @꿫��޶uֆ&�����M�ֵ��윝�-!��@���1��0�Ϝ8w�e�Uyk����s��Δ�?<����ˇ��Q��fk�e\�:e�V}˞Y�˲�,Y����Bܐ9����|�(��n�q�6Ί4r�n�P?��{w��QL�)�f̈́��l����O��*Rck��gm6�N��TT�(�"��
�����C� 0NܼE<�DX�(�(�Ǐ�r�LM``�w������avw�{"=\��Xr&;���8�`7�/	"BBÄA�f�\�`Ndq3h�\o/����l�p��9�]�\��Z/�1~�ì#Ƕ�q2a�?�6�������,��K�ƶ�]+�ݘ�ݜ�ђ�Җ2�#i����ړ\�J���d,�Q_]����Ĕ9��ڢ����]VV��"/z�$nOr�6x��$̡-٥%�cS���TߍY�����_�������`r��xA�9�� ��
���`uG僙����z�����YMeg�-��&������/�ѓ��٩�����c���+;�yJ�A`H�I�qM�m�k|Ŵ�#2���� ��!�ҥF���K)�C>���X�x^��0�`��<d��ׄ>��7�Cw><v��Ʉ��I�������F�.@e���OK2�s������xm��s�@32��Ҧ
0J玽H�(ݼpL���&n���(b+rYC�E��Dˌ)p�w�zΦ�Y��l�����=`�p��m(��]H��n;��ޗ�^�~�:����`~@�(nm��`"��z�XXn����\{w����B�Ҩ�)( efӌx|Q�MƲ�?'�_b�תC]-JW�p��T���D�x�g�� ���"�����)�y�5G;9x�:���{�Uf��Ty�d��4��W秃f�A<��	�B��0aH���d��xy��ߚ��-+iKz�M���L��Ȉ\o�,lo��N5�� ���p�(�'�Q.0�9),������ے#;�[��24qkf▬�6��j.{�������r���AL&s����n8��<ȅ��+G�va�u? �ܓ�#3rs�h���}���(�������t��g��'T�&仄�zDE��NA��"��O*�y�_��_���������ޞ�/#a�,zm��6�o�8Z�߁/����������x����`y�{KH��A��KN�O.��Q��7�?��W����4��_��q����_|4��2�/���Cs#n,����#g�t<�=��M��#�LX�3;���������>��?�����|�_�~���?���_�v�o;��|KH�2�%�Ũ���*p���rg�$��j�}���S�����v�����_�?��g�fT�ߍ��F���?��g��hį~?��3�g��t��q�����+=�R��8Eʸ9#�����6�B�+�/�8����o�>��菠`��_���������j�ۧ@]�`nصt�s(�lR8i"!�bOJ ��"���O�^},$A���H#��o��@䓿K�e������!�� r���$�|���Tp<�Q�a�U�5��&d/����дj�9�m���T�2M�3��!5AVݮ�Ak��r ���^0��ust�O����H���C�ӏ; �yǈ�$�Å `np� �� ��ֹZ�gT��I����OM��#o�Ů2����Ǳ���!�cc^DHp��0��L�D�� �=	�Ʀ�I?<E~l���D�����lF�����f^�0�3p�K�~��;�w�d������Y���GIGF)O��?]z`�l�*ycTh%�kA�pdxx$O ݁H �	��`4�YP<�����r��x�4��Ĉ�Y���OW��udt�I�&���4����}���w��"��}���ǻ��tÄ܅�S�`=�䥃�����Ds��#�z�G���F��7Y}>���g����4�׿��'#���DQ����7v��2M/�ˬK��&�d�N�-S�;����;�����a}~���Oc��1������x�?���8���ĳ!K��N��cƓiFE�탧�s��� }�o������>��O�~��Q�~䇿��?�����#�-	-W;�7q��=�ߡ		�H�J��!��_U���a��!�W������?�N󓏇��OY}>������_�?�4�/����bM/��lT�p���PR�PA� @���#P� �AM/��~3�Q3�#���w3�L����Qz���t�'�yoV�͌SSfr��,�ΕgN�B<9����ĝω{�����G�+'��`	�!��u����^z1�$���2 ��A3w�
�_����̢�pX�<X� �Tm�����i}��U�A.jJv�B:��	����gp���!\/�ˆ��p�"^��/<��D�(6[N�O�����ڟա�]%�(	j���H��Ƅ.f�u.��4�(=T���.�>��pr���G�����8��~�(殡��B��ȣ7)"V����sWh�+���Y�C��2C�i�q<� !B�]p-4B6|��>!��ah��H��Ԡ���5*�
5wMz�ZI���0��2���!�?����ɵ��K_���~��W��^����hfj�!
o���d�)y�Y���T�>5w�~���%��66M]�i����Kw��M��9�A3�Y+�n�؆��
�4K/3�+���0g�]�tiۡ�G��s�<jkٕ��}ʢ�i��d���0m̉����z�x6bU!�ph����aUq?������)����n;:���ǋw�5o�[�4myӴE͹�[-����'�\�8I\ȓ�ZԮ�* ! ����˺�e	9���v��ۼo��}Ż��o�o_�>�qӄEm�W��m��,]�=�k�Z��΅:
ll�n0��45"p@2��;L�=�E
>$��?�f����o3�ET�Q��v/��}�M��r|%HL���]2:'|bl:��:�����5�����T?�������\�神�^!���\(s���`���r��n0cn$����gF�,��,
��� �Q��f7�����a	�҃WK�$����bf��~>)�0�/� ��s0sB\!t�HSN�M����/-�#3q�<l�,rcj���!kb��|��78�1lf8W���.��fvr�t�G�~�8#�W�b��2�u�&f�&r�&xIwyQ"gyT�򰏷���H�g�vd`������0���Ā-�������Tv�&
��D�Z��R�*��"�u�ҥuZ�π����5������`�o����ă�_��ϐ����c����^�_y~�K;K�79�l2o�d\��X�lzXn|�^	�T��t]��V>��]�0+r�λDt]l�4ʧ-�����ӧ��1�ʁ�c��ݭ����37���(T���V�K8k��^ (�M2����y��%�n�tI�Ę��j<s�������o��Z���d߼mN���XS�0g�櫻����wsƠB�yR���� ��b�Q�s�#K��?�����9�7�t�Y[6�,j�O��ɉ�/v�3� kf6t
�)�g]�! �a��}>=v���z_�����U0���֟���f���]>@E-��R�Q��l�Ot��«;w����� �n6��]�1��%Vn^m���o��)�"�.e�Y&5ːγafzQ���<1�à$#��\�9���簪�w)��C0�ڿG<�3[(��A�n"�6<����11b}Ft���(=xef�E�ڤеa����@�� �E\�X	�P3��&��3i�l6ۿI�:+n�&j�,l�,�I��<.��-�s���cŸ0�L���� W�9�1��q�HѶa���36�G,����+3D+R�Vf6���}�h��'�{	��<�'ذG	��\XB��}�'�,��xS�#+v���(c,W� �W欌�jWz�L�������.N�nP'w__��'��pt���7��E��������["s�a9�iFٚ���,9���܎����M-ō�gMl�͏ei��S��Op?s��i�(�%�k���s��V��t2�Q9i�����S�V��Q{�u޶���;�f.�ʋ5<�,0?m�"�Y�k�R�P����ˁc��p���7W��A!6���f�9��K.�nܻ�p{�5m3��&��$�D�^������-Q�c��=íP�z�����9�BID�����5��;���]U���l-Z�l+m/V>*H���%&�0/ޱ����P�ɸK ~ i 
��<���^� ���'E�	�	���,��->��s��}�P	�ez�dn�ӻ���|�s��q$�����-�S�?0rN�Mmu"S���0�j���UH��H����w�^� G��ؽ���`������ӈ(3��! Dn<�64�O��ܔӢIX�
]�	kT�,J-���>�����2F�8a��*�x���+�>3����ݒ�V�X�J�<9dYR�ذj� ��ǢG�pq
�vQ�����\���\ �KG�n�]�]�Q�B*\*c��V�VFЖ�~�>>t�\,���A�+A� 	AgÏ�Oh��2�_s2o�2z�T�\�^#]%	Z��[�٢�o�����w�0����7�-����+x���*%��M
^���r�m�9��9�Ҥ		��q��ܸfyQ�c�dj|LNBH�8gv�����ޠ�L�i��U�dN�3I���$�F֙E�,�N���}&�_��{S��s�˲?˗K�ű���$�yX���3ă�K���F��A�j��p��yp﫫 ��tфdi�jT^F}��Pk�楳�/�64G������Ҋ�u����~y+8'3@�q7��
3|����̕{VC&��iR]�||��x|���Z*��ڇ+���qP~Z�A�S���k	f ����F���pp0F��N�QC���B��Q��~�����1�ý��%��$쳿L���� �3�F0'��a3����c�=+�A��1������d4J���F��C��FJwc���4S`�/;�ρ���HPe�C~H�Hȏ�0�{�m���Z���������V��V	��.�h~���.7�d���
�#c;�3���3O��_��#)fQ8c&cP%�k>ݭ��2!����v�������h6t�`~ �>�e� ���:;�g���ґᛇ	���7�7��s��3���<V�BX+�n3=:� D���D�p.;���s�B>�)І�2�GE��pٖ�)X�s�`,�V<���VF�5+iMSi�>�5a��s���ě��	�q����%v.DY3O��@�;���ܾ�3;�^ܳ�x��=�7��h�Tw��}';vo�}fǖ�ۛ�m��w텽��t��K�RǷ�M+��#��%�u�ص����'�<�o��[mn���h<~z۾۶���y�pӹ}���w��ы����@��V��/��ke�w��"�����rj���?����#_lݵiqӲ��{��=�mץ���n�va��S��]��g��,�/��ۂ�Xf��J��O��8�o׹#ۿ��9�Ŷ={�:V��nYu��ۏ��vz�s[/�����D��V���GF��s/hqu#�a8P�I��}��$uc�}}�E��;n6���>L��D���������eO���sb�8��:�5K@���`#Ѵ�9�m��Η�;T�%/�*��-�K��.��2J{���N�}� �ω�Т��f��`��qlΐ@�a��j^�".w^��}>�^J�d0�B����f���.�Zn�5(<t2��
Fn8�#�3'����^�g�p|JٞU����B�ls�P4�53�9�����8��ǥ�u0pv����	��GKF���
��ʙ�֋�q>�g~�$�y%�u��o���촰0�#��I2�e��007BB�A�K��&p[FG6Źox��;����ׯ�?��շ��\)�Q��8-���W����f0<�}A3�}|M�>3�0*���~ڴ���3�3Peg��g�޼@ܺ����k��u�ܴmՕ�w�[��޸AܾJܽL<�D<�=���f���Y�U��I��ϹF<��o��<�~���w��:ڷ�����ۯo�|u�꛻��g����gg����v5�emJ�CE�˗_�u�xz��{�xt��s/o��v�����延o8q��ח��μ����{`��|}�>Ch��4�m�C� �S���3������p�қ;�ܱ�isۺ;/��!� s� ��'��<���(��+A��`������� ���Q�ً
J�=������X3�+��ǌ�ኁ�0~ Ɣ,A_ W.�4Hif9ݮ�6��[��v9��l��
oӻ��T��[@ �so���1�-@�,�_fU�ex�ux��ݐЂ,z��gΐv��^4s4̈́qv����<b�C����|��=kp|4��0!G��s�J+ۓav�7�yx��x#xx�{zN���d2��H� �'7�,F�pBD\a0J�CY�:g��w�t�8<x�����4��m���$?�14%�9��@ߛ�q8�<>�on.�^n�~�����O�x|L�ؐJz�"�Y�צ�ꔻo���{m���Jk��-�� �p?4�.���G��H=+Գ3'aK���T�)n[$�mi.�R��R�Ҁ����Q�U��������e� g�����O��g׹p��g����Amc����t��Q�h3�y�lYDN���Y53-�g��d�J�r�j�\]�i�O�2))���EhV5t�,���/1gp���%��s�sJ�/�FO��(��Cx�*v������]JZv�L8�ķf榁�&0�P90��g)��WV7Wa/�f�*���y(c*i�qSr1����@n\�<sN�|r �IT^�P�乍�
�fF�P
���|<�mP2tr&��&��CEh	���ǆ!���Or�&��Q��]j����� e�6�M^��!������@�#�M�A	�'�l�C2�3�:��4�@�yjK��Z��-ĥ�&�O�O`f�[ ߙ�XI��cR�%]�>��i��y�qG}���nVӜ�N\�/Ҳ�JrS�� �:�?gS��M�����}G0%n_'^p�#�����p^h8�*/�����M��7��wx �h?���2�3��lA,7��
���H!;2H�� ��^pG ��xyN�.��}���� �,�w�t2t�N4�>sx0� <����c��:�iР�}]\�r=?��Lܔ'�45|ڦi�-�"ۧ�wL	�2)�('aMAZvz\|X��x|��CB¸<���eGq�'p7�y�['Gm��95�mZD봘�i��Ӓ6MOi5(�*Y���}����:9�:�{��ġ��~B�T�Y�|� ���(�+�I��e�#�F�gN՗:f�/p���@�8s
 �7_�kL�&�x�k)�_(R�����y�'s-��⑪93l���j��g$�'rHc�����)y�!:��2}��U�yJ�n�d�����U���O�=�c�m�x���L��F$q] eN�ȕ�R�s�6-�2TU25����a�cѼ�9�ư�rm*9�uA������c�@& �x^�EP���+ s�-�2�����5p����Qh��/T���?f� .y��y�V��9�Ü���=6�o��.T��{۔�f��M��5lt֣P�d;[%>���!Z�d'(
i�1�"�pX5��3|�cI?M<��oը�������g���B�Fh"�W'�Ʈ/���5���Q`�R���;��0�XW�9�#������lN<���dĳi�\�i�c���ف��}#�h7�ɏb�B��P�G8�)���1�@rxhEP��H��TF`
30�n6�˥��67�ɍ`	ùA�	��,`�����nn΃\�<<9���|׏�}�����М~��g���s�C�?0����g�����%����w��ߜ���w���wXᖪ�����W��_1��� ����7���L��s��u�=����9}�����,pwqrwr��`<C�|���O8�o�Δ���:�<J�}�jN�*�2jZ���0���bA���%�E����9Y3s"���� �Z0݁�=\J�H��+�e�9�C�N���J��ͯ�.k��WWWR_����V�M'�2��c\qP��EhYhShq�
td�
ȑ$�ǌ��56�)i(-�ZP�P5����0oL�%�:>0OM3���N^�P1 H�l��F9C���?�-�9�K4ԕ��ϯ�)Z\�S_��9E�9@��}�%f�����4�]�8Y�+�� x��t� ��M�H���CP�T@�a� �@��+,II��`�*����%n�ǀ[�
0��M�j����ަ�u��=m*(�+%�"U?c2�Q�f���@q���y�cl to�?� �Y4'�'c���,�����o�g�OJ�Q"nO�8���j%>�q��"���F�����C��s�Ӱ�RNZ���`F��CC�|N`��|] �	����>�*Dh�A<�;��&
�V�3㘑� lv6_��s��`;#�q١<v0�#�@u�
�(䇂�+�������������}:�_�~�U�{� ���+���7'��[�~n���O��?uw����e��@wg/H�����|���O������.����\<]��W�A� q?�^���ny�����t��1�?�A��q�kࠁrr	`�p��ӛ܂LЫ�lD�z�P���U��ʯ),]VY���������������ri}��#�j� ?2�?)�#@&=`�	*PJ\�B�mo(�^ZQ�PUZYQU������XT��)<s�W~*��@(v���@���I���妒�Ҋ�u�kK�kʪk���jj��ZR=��jA��� P(��wk��1� u��Ani��U�PӰpQUe]]mcYye�º��u����%���Y�As��QD�v �2�@��� ���fnw(=j �$��
@��)���Z�!i@=�O��wrD��p����v���RO��Ϥ�;2�,�6Ӑ�+�^�e��6�<M2�b�N���	�Y+
̏���cɅx�5
�@h֜"�k��uC��̢�ƍ7�2s���!��牮��m��ɼ��įP妗P`��3�%��P�^`>K<���)� �E҂p�5?|g�H$�A��p"��BB\C���D�O�U�7#�m�Q%�J�	�r��!°�Wq�W
� �(m�(X���A!~!|�X!-3!b��'��W�O]}�@��q�z��� '7��9p�������@g�~����z������;r��������������pu���i@O�=��.�(�5ؐ�i���.�9��׊���������i"�[�����������H�)`R�J��,�rD��Ɗښ�����ꪪ������R vŒ]����?�R�^���឴i�p��-��֗�V��VV5�.���*/�����h��Tc������!DZ�2�:�'�{)��l�u�X3:�ƪ�*Ȳ��������8_97#�X c�@0�	z���1|�aՆy��隊򚚪�j�,�u�`��C�*��|�W�h� 0%{8L�}��Ϟ`K�#J�*���ח��2�/�_����gPx��p�È�fx�;�lR0{�	0~��K+�Ã�K�ϝ2��0n�m�BKFiN�iDH�&9pB.Z_
] �+`��ŕ�
0�	�L7Ƀ��g�'�:hZېY�eq���AZ5/G>Eq����R4���9���k﻿�:�u�x﮷����q ������c���AB�1��6A�snID�&�8���6���6ƀ��$	%�y߮�}Ԉ(�����6��:U�vU���s����`00�+��@?����9������'�ӕ��gf��fL��O��tl��5%O���h�rv�ENv���r����^�d���nՔ
m����OW̤a9S��`R=%�ͣm�`B��� ���sON���Yz�)b���;���5���y��%����#򮈸�qtN�.�Ϙ;#�|W4`��Ȼa��uGT�_�����;��&O��������3���֝�q�~�_�\1�pD�]Q`+����wa�����w�ǿG���&��bZ�ei���cN2?��ބI�K�g1z�70����;[��[�`[�a��`a$������'�/� � ��3+#�t�2�M�?�vKSK[c}3���-f���mSSs{G3��E�G�mPn���[ɖ�	N�i�F��-� ���mm-͝ sSOK{gCsk{��--Ou��`�9�WWɤ!b}1���R�X���[6v�ljmoܸnSWkSk]Ww;*�A����ngk�e��b1c����4�h��ũ�S�4�.����-<��&ϓ;k�?����6/�0
ʨ�Y�6%���NU�e!`�觏�M|Ό���7ү��ӧ��1�Z�f��J���{|/����q�W�tN�?-|rf�}W�ײ�
���-�0����g����3�Y�aS�01����d�IS�s��~#�������ڒNs�S�J&����c� �ym�_��s�q�y�t�����:P�n�z�X��7'�r�Tz��[@�@2�M͘>%m]3�2�Κ�5gf�����ӧ<�̃W�Z�PM���r�
̦���b�V�0%#mZN�)���,�����ܩt Qƌ��YS�f�$��I1��)W�#�%&,��o���������Kt�w��d�t6H� ��=���{�]����Sc�ﴘ;f��yO�_�d�17�g%�15."/�/q��|O���]즸�������+�w�1)��;b'ߩ��_Qw�M�없�_�`����tP��W'�c�j+[�����z�����Dn�[[�����[,�5�U@>�C_��K�r����������o��h�����������_�q{[KS{smw��z����!��K�s�D�&�\��3���֖��Ζ��f�_kkswצ��N���m�-���J`�c�!O�A|�ѱ£D'δ,�<�l]疎�-������N���[�Z�4�w4n�Z�^�&4
�\�S0�,>S�M�W�/Y����/�=��t����^��O8/�����T�Ѷ%-�3���Յ�H�蘄H�2&��pR�&��]�Bz��#&լ��Z���bw��ҙ�Ѐ4��Z�2(����>i���I�׿�3�SA��Q<B��N�`�����nW�ڵ+ެ�v��{K��������i��B��W;���z�#Ϫ���Or-���#�� s���LJrD������"L`�7�����,X��D+�^2��t�#���M�6o��{f͜;g�=s��;'��9y�u֬�f�.Ⱥg���{���[Q2�J�g+ζ���T�gV��,���xڢySs�,P�}���;cƼ3�!B`�}3�wߴ����>��U�ϱir̚{W,N�����������P�&��ƦD�'E%������E%����<-��%�ūJ�{Z;�I�ߞ^<��{�)�o��p�q�Cz+���t`o3!>�1	�I�w�$F)R��S�)�I�1Y�qSrԏ���4����*��&�'X�X�P�y ��i���66�-���u7�m�anmkii���k�i6��VЋ\(:�3�p�)��ݒF��������M��;1�tull�6L:Z�m��Zs�M�N�qP�IoA�ߡOgT��7��Q����s[S79͘�v��oi���X�\�=��sh��(U�	9N�����ΆM[���{z`�6wu6l����ӳ�֖���m���`�Q�k8ZyҜ��B�ڧ����1� Π$KW���a	 ��1V8ǥ�-_�a��L���l�1٣�pGT�B�<!7;�[P҇K��l�qz������a�a�ei�4"I����ix�1����������J��Aף����~uL�2Ū��6*����(M	�f9h�r�K��u�*U�M���M���r�%���Ӹ�=���M��a��	'�vab�(�w(A���nCª����g�K�Ã�(.j��	M<(jʄ0���5P��^i�ᧀ�i���t	|�-�+҈�"٩��
�5ǣ,f/ c��E��G.KM-ڜ��0�ay�
�08\����Ppc1�:�
D?G00HHfˑ`rR��}��Jm��k��RiQm�^d����%��M�0okn�ٶ������V���������~e����/�8.��<�F;S�h��zyMW=�g�Ɩ�-��[i��#߳	f���uMw�޽Hc؀��Bwk����ٶ�'[<�mi��^ײ��k{]���έm]]]k[6���b޾.�\��م$�0P!P����sO���;;7��vttu�u�45�p������ݾ	f�׵���2Ӯ�s�x�-Ƅ���Q�0�S:�B�t�υCPXc4���-�q;S���AХCҹ���rWiR�j�_?ɽ :@��AP���9�]8�r��q��+�~���4�~*��!�^t�$D���#�����F���t|Y�'�l��j��z�5�]����(��~�]�x,{GT4�H����X��Q����2ӡ���T.��^z���!)tȇ�sO�����s5����E��>٭�3/��(}���/��;��h�X����.!�M�����$"��x��w�G�^"��w��@�{�R^\{�"L?C�."�Hs��w�Dw��4�	B$~~#8�.~�p�\�<��s$ �3�aD~!�~�S�%�$��-�V��N���e�?��X�lSWgkǆ]��쩥���������V����V¶c�F������ߩOʤ���G����[���6uv�Qn�hm���w]s���-�My�&z��W D=0�X53�Kh���46o���}[]{��fL�Z��4��o~��1�a��MHUR�x�6�n�SUV�Q[���������gSw[#������ֆ�g[���L�YvZC�X�Tm�v��5�=�Ⱥ��4x|���K���+#��5�ҿ+#A��m���y�m��_�(!@�a}&���>M�הU�n����b�!��d[�2^�#D��zO�?��Y������|K���x:"[�T��0+9y�N��3��4�N��K���
U����V����'_]����^=�ot<0I)�2���55j��{�:!�(��4"��Iv�®�)���6e[�sp�^��/�1!�iI��s��bNJ~PΔWe�5�jJ��[�{t�f��,�A"$�AH�i�ø��F�D�̙�92�N��2p$ǃ	R"WQ�!c���U
G	3Ҕ m⏶bX���꡻�6���-��6o�h�Z� #P���q��[�3��t>	r�2�gڌCZeHҪʱ���W���o��I���`���4��67V����9�sYu� &H0ϵ��f���-[:��@��ww�w��ٺ�'0�Q�YE�̄e�1�b�[��-ͪ2��{�m��h�omlh��|������y��ߎ�Fs��WY(F��&�i�RX�Г[jK�J����tV���Hv�  h��e��}���r��xW1Z��N��^U�yaz��⥺����^�O,`$�H������9�}f9m�H��I�s-jq8�8jW�c@��˄Y�ǐ�"u���1�������ti�t�����o��-�{LP�kJR�K�f�p�:In���꒬�)�Z����7'���4.�,QM�W3�G��`�O�Ϛj1׈�A��z�k�"�	���#�{ ��#�8�mxF�'��@2�+�Ex)WΎxgL���:��]�DLU0��o���rj0RgzJr+���km����M�5�t7����۲qu�W_�T~}\Y�2��~�S��!�C[/�9�.kv�m�I��޸�i#����\�H�k����RG<	u�� ������)(��^��v͎��[�j[6��j��&�=��+���,^J,@FO;ɥL��l:�nu;{ꚶw�_h�l���T��ɹ�����GҬ�L	܊xg��	&��f}����NeG���f��b����~L�~���<��5Bi��'
f�cS��{�~w�$2�4�Ѕ��qS0��4�r�z4n��$�F��-�j��hE��N������G;����������s���=.�0���cL
����2�:Tׂ���Lչ����u|5��(ʼ0Ʋ(�$��緢�4'���#z���+��( g�N�q��=! G�7��&(4��'(� &ܽ���aZ��Ӽ�P���i����)�������B7 < Yu?�@���D)�[I����[]�����/�8wn|��r�c�
mz���2|�ѥD�`�Rb��������J�*ʻjkv��nk^����Q/}�kqDUal����EѠ�i\��t~��0����=���Q�y�gk�������,�7�ӭ�$I�0$�)��2�Rm���cac����*�k��6������T�}���2�]�l�$;h�V��"�C�4k��x�����+pta�/#��d�5
/&23=��4�o�98ذ�� ������������S+��C;S}��r��!�=k�chD��aS:��q����k��,t<<��R�m�g�up�I��X�>��c�������H���՘ҫM���]�H�Ϗ!~�1�ʄ0��>�]�bBFZ��+<&9��A4Јx�e����	"�	a�ɅR)�Dr ʣ���譬�S�qƨl���#���~����
H�U�H
1"�E�62J3�e�:X�yp����K�Wr*4PJLt�e0��fVMt�4���%��ǵl��a���bףs*Kr+400���&��c�E���AT��>�R�L��N����yx���E��fۖN�-ΨT'�^��!�AE��n�A0���q�>m��e.R�R�c^�r<�w?����l߃�D�-4�K��Y).�hՇ����W��gԃA��P���Ii��͜j��(�ZO�IN]�J���c}�"�abL��C��o��9�I�oy��!}��Yǖ`�_�c��j�k������Ι}���x�jY�iI�U�����A��|�0�p0cjwK0C�X''�h:x��-��Ε���O��U�GEk��^9�d�H��N���9A��8�_(F �M�0�DA��p��$�U�H��!a�)$q挜���)��(a����o��qHO��ç�EN�1f�yvCf�&�B�e������ F��@Gpg��q�HT�n���U(3�,�1ͬI��3����jme4
��-�<��HFb=K��d[��c�~�6�ޕЂe�S�u-�Q.�,&{�1kL�&��E�]�+���U��m�Ā1�ڈ��ӡŰ��LEu	J���}��y�?�	� q�����{�}7���S��h�q�9��Ks�h�V�o���a~���*�
���� & [��Y`/�1���c�|6��8���+)uNdmh,o����ܷҥ�'>�z����/~�K�['m�e����u�=�5�YLO��Tra��  '�IDAT�ajD��"֏���4@��n�J�-BSD���"G���]��x��(R8�
����KT^P%^�R���6b��p)HC�6WI:@�Z�K�)�	�ʸ��}�ާ�ub�#�*���Xk���Q��K����Iu���V����5�Y��)z�&��HK�1Q�]=���g��j8b�H��4Ƒ`�y�e�R�z�LS��6�	g�k�-�X��)�������*�H��1���PC�"���>٣�G�dӤ�M1>��� �w�-���*�X�6û8�)\�~zv=�?��	k��oO�5/�0D�o�5���f���g�c_����"&�'f�#Oe���G���,���I[ ��l��)d���.�rբ�x���_<�����ϥ3�H�m|sf���ג�+���-�̄(&��țPx�1$� ��q�H�Rb�MҊ!��=1�$���1W0�t�<8`��&!%8@w�M�,0&4Ј��d�\�� �э�k��Zx��E�댈�
�;4�U��O$�����NV��7�)ޫU@�-���$d�ma�0���>=P	��E^e�CC/��$+-�M����hj��E`>8�0x8�	�	�C���"��$���M$���H ��B�]��@�<� s�F�a�8 A�H1(K(��`��E`� �;�X�x0B�"��6<J ����ċ�  &�',$|����o�HYm9<S�2j�B���`� �}{�u����e9K����)���������.N�2b�����U��6�f*�!NlXM��[�kJ�6ìΫYr��y�an	8�5It>���5`�.!�!=qC
ON  �@��C+�� ��i �XD���ZB.�� 3�?�I�~
�Rчr��ƋĀئ�}@���dۢ��Kf~"���hR����R8�h�+-�'7����&�b!��Љ�D�
��X�
��)efu-x��r���V���8�g�C��5ƻ-��B����bwc��5fH�oFhtPx��'j��f�d���
B) H��G�q�XTq�E2����!?(D��L$��)�A��3�ֈ�oʪ1�ϰ�򜖆/���wN��Y�MwEE�s����;6t��|���fֵ�{������Å��___�ٳgN���a/K񑪥;t?J�O�93k��H��a"�mP��/Q �V��/t���=�!K��	��K�5�8^��סD9� ~�K��%S,�
�1�|K�ģ����cӰ�@)E�A�����&�K�ц����x�������;U��dش4�tk#]�yvcZ�2ƪ��R<Fx=h4��ve�sT�H	�/f��xc����2֘F`������b;M��@/�W����1Vb�
�Q�&?��
RH�I��UÕ��'b$˹B?�CNh�@Th�eQ�Q�!drb�W��5b�!�⟨/�.�┐<cjt�#mJ��|熃�g~�;���;���k{����B��O���|hp�ð��ǘ���N�<0004DK�x���7�a��2���}��A�$"�@��#�;١��!p#!�[O�妧V�N���F�� `�����l���%�p
��'ga�`1��r0���0Aיfi�O>}BuItUQR�2ϻ8�iL�*�`z����<fD�W���6�ե3=KZ�U�qGn�R ����O���T%[uI.�v�u^�ј�ztiՋ�]z��[,*L[P����/��:�
�=��xK����]_�z����M+�<붽�e���Q��g�_o������Lt-�e��}�P���&Sxk}%9K��(l蹀؄�%��U��b�*bnH&g��$L��C��.��"��@c7��T�ȱ�uq����?&]쥥����~�m7�̷�<�5٬j��������߇fz�5�4��(�f`�Q��c������]5[���'}��/���ŵ��g8��?��49��2_f��'j#�U��%�U`�� �J���7�jA�	�.zւ���s�!�� X�Ӵl�w����U�e�*�������/�r/mSC��̖�'ã����_�I�]�<w��������ݴ��nz��g�;�]�8�}��4=������wi�M_�n�^��W��!ݢ5���K��r�_��~ 3�վ���.~���҉w��v~3��T�)�W��PZ6BlP��G��Q�Mz]b>2��?Z�#	{�u�N�8��ve�XA���l�g�p�+��8,!Sx��42!�n����3���Z��E$̉��P���n���>�����4�̦�6�Aqc��<�M����4���~�zF.e���+�1���XR%}!���
�/�4{�3J����0�&��TZ?�,�B�a����)¶�I��
{��e0���E#�"j��9��}l���d������eA��IaQg��mo��(�z?ޔk�f9�:�����a�B̥Q} ���n}��^�Lu���N;w�����O|2;�v�Iڠ�w���|k�c�x���'�V�,��z���t[�E�c�,�yoS�G�>�1�\�x���w�c�{W�<��^n��B���|t���������Sl�,����_S+A}�P@�!�)�.(:��n�me�O�iD�w�*̲2��f!��H|�e<3�1H�)<�\�$DbyhHU=,`
���H	B��xu�6�f݊����OJ#�u�=�����F_�D����m�ߤ^�R3�;ь�`x��w��#Tv�j���p�=�΃���!��hA���g�E��0���(
�j�01�s�of��{H���t��1VZv�Ѫ ���wS��lB)�x6�i<����	�гb�6�J�y��t��Ѧ�&ժL��Q
F+Zq����|Tw� )��HaW�>��j����ڲu+���}���
��׽�l�tgU���_���D���Kk��ͳ�fWju���̥��ſH�e[��?K�k]O׬�UQ:׼���_8�������|�C�*�M��&W-���1������b!$�� �m�7�E_�bGX$q�9�� < %s(�$�0�"����0�{0�.@���RD�`<�Ȥ+�/��H����Y$�6X\0A�'�A2(F����<ײ�}ǂK$��痎�u>�B�7̹����M,3�ĩ-���8|�6-�>0_�2|N�T�m}���gBe�T�~>yN�/�f�Pt� �2��P�5��*���Y� s�]G��9dpG᝺i��ez5�c�?���Q$��љD�O��8%������gt]�����6�ʺ��%=6�,�R1�����RD.`�__][4X-lY��g]�ڭ_�xD��u��u����cUn�b�JĐ�(�v&��'�A�T�6æ���~�k-����ѽ}i࣭4Z`�k_�x����
Ӌ������R�b���������=�*��V���_T�c��v5������(�#��P�/,q��*S��� ��ҥo�@���6>��5�����A̨7�r5� ',3��m���h��)����N�Kf0X"��&����Bm��\[
��w-�Y69;��jx� �qPq�D��B2��)���N>�~����C����g���7Z4��7_��ҦY����pN��@�ś/�.{\���J����r�uI�������v�>��)�w���*5<I��UE�oD3[�$	�l�bM���3��ȫ29�h?"]ؾ��;=�%�<�t�����О4��pݞ]��ǥK'���ҥSt�I:��k�O/&T,�
���~�I �`��������0p����K������)�Et��թ�WVG��}��6�Q��5�r��z�ԯ���0u�vݧ;v�W����>���R߲�׎|�惭���bX���ϥ�c�ÐU��L:]��=e�������~xt��G��ߛ�ڶ��-+3=���	��������+��?�(�l�E`�/��k���xC8<�-����1r"r�D��џ��f�^�s����_����VSY]���9���.O�S����+� ��>�k��XU����A�႞mc&�/V�я[�N;%ռ�9�B�a��ڊ�C&۔�H���.�α�2*Չ�E(N<�C=�AW��p�U�e��P_&9y!m��[�����ҳ��\�!��N�jh!~xs���:���B-Z���~������W�����^?�߿�z����g84Y>#�*�����zd�� g��=ov�������ק����.|u��W� >_��Y&%�>:����h-m�����@��V)_��g_:��d���7���,���+���y�{��8�Ś�7ϴ�M�2~*���WO�ǔl�������ZҬ�閒ڏ��:�{i�u����
]�E�(�/�)نw7=��۩R ���aX$�@<�k�?h,�����hj��J5�^�����G�Z���䔆04n0�Mp)���|G���V�:�����K_��4Ӱt�8b���CW._�t�ܹ~i��@N�-Aa�a|�E��O��c#'˜��k��J'V�s+�S*����r�"�WA��+5�V��*�H�)��Rn���8{���J;f�;���jL�(Q����oI�y�2Y�*��<��66[��U�,�)�a�r�0s�e�'&,3�ϓ�E��H1g�¸��R5�r��U%�W!�@��[�=��V���][^뢹��4����ͭRx�6M�����믞ߓ�T�|�C_Jg���կ�V� ��6��N�����<g���Z���x�IV�T���a���������{�S�^n(m���殢����TqM������?����U���e^'��DX[�A���D?m8I�����*��W�O���C;���Ѫ��Y�ƕt����3�8�c�!l�E=Ӷ����[@���.�&)a�������6ô�Z]0<"	X���w����tn�ڧ�l��)�R�^[��*εk�N\�.�~�w��~��n���W�vKt��WW��G��#�;r��+?�*�-A�Ϥ����t�g��1�Җ��ʪT��)��*+��oI�8M��@!0����$y�6u�MCu��8��X��/����W�Zm���wf2�2wi3&�*en���v@�	�L[I��θ�%\�3����jz8�]Y��x��񤣑6=���[�\^�ϭ�H?�9J�V|/��-/�]Q�W��������K�%Z�ns�S�X��6¹��^rH�P��/�Z�[:Q`]�x�s�t�Rn`I�SeWe8�n��Û
;=��!3�@�s]���ڇ���i�C��ҧWj�^n:)�?#0z�0��''0�P�o5D�����L��'
f���D�&�J=�Z�Ι}�PJ�BK�GhM&���Wi��H��3?K��ۧV?i.��^��a�$˂d�:Ӭ������S� ��}�ҏR����a����,D�g������ҹ����� �}/]<(]�/]�:�v&�fSN�.�I	o�[*�)�00S�N��Tzr�=��jc�_�	�¯O��ā����i6#$�'#璘ޥ�K̟��z�_<�\!��n��j�d��n�2�F��w�W5)@�b�H����E�ݦ��/��[:����*�T�U�I�<��[�m���!����-�W���Y��8١�〉�4�~ӗ/�@�q�G�rl&�f��ү�6��(�*ާOwj>��z�=���/�	kLnv�X+�ݜ���.U����X�W�T]�`Q��K�}���t���?$_�`s�x��;D' ��w�/��cF`�>y�-&J�k�Lr�'m3b���h��K���{�W���_�D'����S�˃W�za�/^!+=tV��M�ǉoL�U���5�1:���ӤX��5�-^������������O�}zA�Qe�rM�	���OW�U�˕5O(k-�}xњGA����>VX�Ģ5O�6>s_���k�x����ϩ6������j��o̌d$��FNN�CM�l��.�ꦝ�BۧK	x��I�3�w���)���ڥy�Ŵ��M�ϝ�E>�nw��Rb�}�ؔ��8����<���=�?���|��T�6L�����^*����W�yqߪ�5+w�Y��HN�5f��n]��(æ.�?������)�-�<yz�u?���2�RT��<��g�Gʊ�9�R�(�
�~�݈�9iM��^!ԏ�z��Ϭp�/4~�G����g�P-,�,�D�-�ܳ��(��tؠU�J�i1�`��	�AM1~��,�T����ȉ_�K�pI�|I\��Hg�����Ё��/�s?�i֧��0>�L�g�^z�JOk+�1OK�h�=�8+9�INC���"e��WtE�\t~F��V�%�j�����0tZ5�n�[ם$xfi	ۋYq��,$�JM��J8�0�PtL�A��V�6�ܘ!���ƈ���f0�	��t���0US�a�7ڶ�����~$
<{t������N-��UE��\�(���	{i5���
�to��0����j]��HQY�m�O�``J�(�+�mJ�������
p�r�ݐ]E#}!C->'��f�[������u���)��i��D��hIN]r���^j�_���OO�oA_��a��j���#0�|���/R����WX��.cl�B�+�Ϡ��� �����Cʚ*v]�[�s�K�/5������^p�s�ϋ�OK��/�������JM���'��.�QX�Oq�s���Fٕ�F"��1^}B�i����K�����.�E�ca��7���!��x;� g\A��R�H� �6Sn�	De�fI�+f��,$}}�Z<�K2�C�����&���Z�*V<4��b�A#$8U ��N���*x�0(D����.-��[�.���>-YW��ʅ匵�����"�1�x��f�Jb�
1�EVk�t.ʪ5����� ���ҙD藪�@)-b�� f�ɰi�t�)������O�6(�Y�Rk��.B8�ڀ���۫j6mj�r��G;�/���/��ߤK�~�^:_�W>$�ݾ��g���Z���`��ZZ8�5T��r�`Nr��w�L���{	\A��.�j����=U�4�������T�O�v�sIv�:ӦOsQ5`�{�D��A
E�]�
�rcC�x�E�mp0$A�@"�X&B��l�ۤ�<&$���Y7��G4�x�5�_�a3�$��G������� �Bbt[�����qKN�ud8��%�`(�h5��	���x '!#F+�ȕc(�d���nB�լ��i�=|[�>�J[P�]�ZVVW�z�z���η:W=����j��l�!�J�
����<EI.:����!u� ��*�����h{�SeW�Q�6�G:>�n����^La7 �XM��J�?	'Ǆt+������O�De�$`Xb�(��B�r�}Ј��Q"yd�q^�8R�#�<
� �CmJCC�P�f΂[H���E����O�*�`��Z�,6E /7�� �B���0�>�z"�{4�~p�z~�[�	^w�E��Y����Zf:K2]�t;?�d[k�i���
0q0s�������j��c�GM{��bG��O�gK��L��o ���Q�B�
Ρ�_E�db�@���Cy�a�.xR)!�|w�ĜA`B���3r�<��J����ٯ!����q����T��JL\4H��"�s�y��W��'' Al\qW��̟�r��|������;"�U����)���9՘)�Qd�1In}�ט�#�ч�#�4(�L�5^0�[���1b� ���"���1݊	�1�E8��0)����8S5YY�1���H$��j�!��9/��af�mG��H�?o�D\E�䂘��������L���j����y�a�8�� K"���D�E#<91�o�ư� NÉ���o�d�A{��#P�Z��6:���Uɑb�n�@8SiW�;N�p �����+CA9XE���v�Rq~2�[ ����UȂx��*�v�T��F�0�l��\n��-HⰜ��+�A<��Sr�qFx�qt�<"�_�'.=�\�CxzN�A,�88f���8;����939,�Eb3���ܼr<b(}�e�@O&�/Sx�t-qs_Ȅ�fq�9���.������r�k2�D�T�6?��D��|�^�' f�bX�d+��A�W�
H���K;i�OE*�S����>�����?I�P��ź�Q�����������r�\.�cD$!94K&��9��N��X`ndAA��L}!��陭̇�|�oɑh%d�x��@��qP3<�u�2[�̿�bŉqd���nQ"荴[��Iv�� �U�(�zT\'f~�A]N!�H8?�;��G��p���.��h�����)��ӛҠ���1ӎ��  �5FPx$�G��80���~p��n�?�H@���6	��,�5��)d��x,����1��>$�"b*N&�D�GC}�Y8�l�B�3�\����.[h���0'e
��\�u	�*+-ilظ0 �'�б�n%찂ڙ�W����(4��uA��~]|]0���ּٝe��l!ɐ��z�0k3w6$�Rj���.�ً��5��Z!�pe�+~*.�V�g�
�PQ�h���u:X1n ޹�`FӰg�+ !Ua<$J��6x��N$dh�����g+Q����4,K(�(���Y�m2�g8q$'��	�hpk�9�o14�¸%�e��W����'��6���f���Q�b{/�xWq��^5�;�@r�;&���/��W�kDu��ɽ �ز=F�H@�
���,�׺
*��u:�� Z��|���g�'��B�����2�Fs�<��+��a�~T&�b����[\yN�'ܛ(g1�T)��F�*����^A�޽.��hiJyi�1���hP���'՝Z�j��ѓ�4b�%r��-Ǉߒ�i�#9 _��C&�����IV0�mgGF���O�j�$�>&rLq�$��(=�	V�&j7����C��q��>��#���6�PK��s�:֗��s��?���־�3�n�i�O����3�E��\6�c�%�%�ථ%F/ܚ7��nNr��DSP����u��ܠ5H�1슏z#�k���n !'L*��H��u���ʽ�6~�$�#KE��r��}�$�u��� �8R�V��ӑϙ6��J�?N|���������+i�I���`	0C݅?:��6���kiL���~͕������s=�,��V&��r��$��D�y萓q31�|n��z�+�+Z�F�Pe�K,@8�I0��'�����CȅQˈ1�px\נΈk0f�"ɥ˭M�7���Dy�H�	OsK���Q�f##`̏���t�n��?��	i��r����l�!�N�Ik0�k:.C�C?^JsR.\9 ���%�Va�!0���R�ۤ�i�]�1��%�j����2���9^bVȞl�������= �\�	0Dd���ژ��s�0A��gL�Ĉ���^�}�Ð��8��m}/�aʱgU�����?�&���k�3��W
*L9����y�̧��{��>�ASV�`�9�@�*m�
����
�a�ɷ&@`5�ʔ�T�,ބ)\���y�A�2C��qcVȎJ!<�F�y+5 ����6�������&Ƈ���,K8^BF������0�gb�e�u��n���rZ�@j6�T�s+!^����+����ɟ��O<����o���3||�tz�ȩ���7|��˧�9q�׽C'�K��q���W~�z�/z�|���oL�a���W�G�86y(���<�����7���W�0�@�R]7�ͯ(X����B���ߘ ���T�s?!�xN�}�����Y���@ �@$���k���*���f��y"�9����zj������<,W
|�C�ύ�zܐEna������w��r��^��=�O|=B
��ā��������]pt��    IEND�B`�PK   ]�'V�cŌ ~ �� /   images/40a6b5df-e714-4004-b865-d48720df955d.png�eP]��.
�����-�-�������݂��w�.��!�%�����{������=�V1�{�7z|�Cz-��dD�ap`@@@��ń@@@{�|� >z<�F�A@p;ݕ��]l�m��,��l��\͌A@\W�������k�u���S�+\��.�=�Xn���" C�lBC���{�Z��*v��KY(�?~J����>z�1i��9xx~U�:Q|rz؅�!ß=����~������tww7��?�=���!��M%6���wz�O����=v=���K:~���������wv��I���y��r0A��E��"����+��������E��bOj������Ъ�4�����]��ד�E��"]�o�/g't��b|���k>#�ի�������]�ޛ,�ĪE���s��&���0��\�*^�6�Hg�X|�U:��c��*5H������<U��Cx1sT�-����&vƯ���Ik��#w�Y�/��K�.M�]���5ݪo�1�m�-�rP=_Z����e���С,�ҷ.�u�K��`0~�H���$_ғ�UO�!b��a�Y�|�ܙ�	�\�!F:��INV���3�S�X�c�O�j<�/ާ�m�Dq[��4!�W1�����Ȁ}��/'MQ07+Ĥ�/J�(ml�R��m<�0kl\Ho�V��]ѼX�]c
=C�R��V`?��A�e�d����Դ\���4;IUݩq>��vW�mɩy��̮77I�wonV��y�p�ڞm��ĪY�mWt�s�wqv�|�r�#U!b�W����NDd!ra�|���iҜ�|�}�a�2���l��I��MT"�o�k�.��0�Е��*[$��i�'9P�oV�e�ܷ�Y�L��?��%���E.��jh��:vu^�~}O@LԤ�.�8Q�T18-G?��jF�>�����b;]�о9׀$ݞ]<�q�P,�>�j�&E��<*���=����Ӹ.������n?�vYJ���F �
u[s�e#�pR�}�z�I��O#����њ>=B����%��8 ~R�p+�-��Q��^������[��m�l?��w$銜�<���.͝��a����U��݄fxG�ި��|�F�A�������b n��Nt��S[��&񍣉5y1�Hk�w�U�V��]��j9�g �-[|Ԃ~��n�<}��C��a���u��jz��r�3x�ЗA?z\�~Sc��%@�������E�=��R�������@�ѹ8_#Y��W�ʁ&���U��f-ƗXJ���bv;�bi� 8��"�����(�$��a�Ndk�,��q�Nv�7[���L_�%����75?��l���wq��D�(2�;t��d+�#�|��^x�6��q9k��(�;3h�Y���82_¡�c��c��t���0��3a�ih�y��w�����"�v�Wݚ�9�.@����{L���OHgp��E�o;k8�2�Ԩ�y;�΅����S���r�i�4˃.0��mՂ����g�Z�I��rU�C2�n'n����:�_Pkk�-����H0�t�猾���KpS�� ���S�\؆s���E1���L��� ��Ær[�����&#�j�GS	K�l��}��fV�§��F��T�,2^�[�,�����������_x�h�น��N,��rm������!�H���98Q��~��&913j ]*�*NG���2V 1����?5���
���(�M"QX��?D�2�zXkS!H��%�-zl1-\��D�(M��*��i#Df[q��qK˪TRD��JA�1鏗�H��ll�!�Q�R�؁�*okC�p��-�A�98C�CQ��>	ί�0��}-k��x��Ϝ$�Yѹ��Ð<���̓�-d���+`���(��P9�o�[b���+�P��%���1F	�cEZ.��g3G9��v�Ce+����3tx��y!/`c/�;_3��B���`w
>5�%0��zj���"���9�o����Z��m4�2���/��� 0�7�R��u������I�x8�!��4K�f4D�1����<�j(s�%���05�%`IŢ
�]��%ǁ�+t�P��:������S>t�pUȼĘ&i� ��o�X����W���[	���uS��F�e�i�K��kCB��^�jZ�6�|_vl^��v�QU-�f����Dp���F���4�5(�\��POc^Ƒ0�4�����o>d��Ӡ	�C�����̩Ϛ_���&�f��|�����@�E{�*��1�N�'�#8�}&�mf�ݛ�()��0·������#��¼ U�X��$�kK��~�L�����&�h0 ��D�\ ���� �̨";/����Ӑ��bj9�-����T�}b�3%�&��~b����8G��F�P��W2ҭ�T�6B�C,Ra=�/H�8��3�t�C�����V�c�T����p�>��ف��K'<��)��#P�"hzg��ψеvO&��	9c���D��OpI��\���^>D#�oYߧ�q��_��4f.�{^�N8����
ϸH;A���z�@F�n�� G�y��� �w��!*��rU��zpgic�Kn���ᗏ>�E���x������,t��Mey�U]���B�i	N#K���K�Ks;Sc�x��1�Cy�ÖR�߳4~:'6ts
d6e��HL��5��P!�Gs�2���JгtsP��A/2�C��'�k��`��]�ځ�9[�6�\�[:t.A�$�:ظ�$�fQ.��V ��B�2�)z��L�
�:���mx� ,�]��`�'	���q)�g�qZ�2�������c����XW��/=C>foo�t�o��C�#�Z}�
r��q=�_y\l������5���po��4��8h ���4@����]�6s���T����R��>�V�K<v}ފmI�,f=�3L��1��ب@��h���]�������}\jM0��T"�)p�cuIw-y �m0��n�f�=�6�6J�C���HeQp����&[T� �.H�}5Xe��EW��9���,���>B+ș����%_�7�E�)�+/�@�� w�(1�fs��Lߎo=:#"4�=�����tv^f�M�>J��T�4��ەya�����h�0(��ӡv�8 � �.wi1H���0#=q�d66O��BȎ�Dl����W�Fo6}�!�w"��3��23�oJ}ˢ*�:<��Em�'����t��q}^(�ٹ�P~�����f"�N����q�ݘT?e]S� �e���6	�>�\H�_[&M�"r����$z�y|C��
��VA��ۿ*|�<BcGr]�R�SQD�A�E���.-����Y��!wf�}K�L�ҽE�Td�܈���(a��!��������������W��mT�$���\a�v>�PY���ˢ}p_�mv	��m�߰#!�SX�=jǣ/F��!�
Wb��g��@��D!�UNn�2�2�@�`��T3گ�)�Q��
���fn3.����}t���vcS�*א���q^9��"�#�2��J���q_fd�Jg����COz�*t��Z��T�O ��K:��ǻ�~��&D�Ƅ�ߝ��B7`)�u�"[��R�`7O�Q�~}FN0Z��S��
V�K�p��D&��+'FŠ�?��L?�7?UQ�{�[h#n"z�i�ᗞ9'�_��j����~�XTph��0|̋2��	�]ƈ��y��
;�E�#�����_Y
RJ" 3[�2��h�� 5�(u��=1���JD^�Q��!��[мQ+LLC�_�U��SY��s�,��#Bww�M�״e����<~r�0�a7�ўѥ���n�k=r_u��-+��؍oG\����+˔#2����@����M����Q7��d��0���r�O�n�tV�w�9ݠ=~堂6瘲���(o�!���V�Û�s�/�Ԉ��MG����h�8�������$yw��Q�����D�������yBU�+���
���Mh0w�1�PĿ��V��Q��at�ңp�����c��#D�axݪ�!�<r �{\�y�G}us|w�5M�k�H��(��v,�_�ʾ�R�%�̆Ɗ�Gl��
ZXhD��	 %����\/�W�P���O��HLN&Ks�R���@��̍H�������Z�S�+�Y��'�� a!l��s�CzR��'zt	o?E�FE ��iH*���s��=�RY$a+U�38-�짌>@}�8[�P�4��v�Qy����2�1yeMkT��[yױ2t�D����ρ1�`�_��|銣( pv��I�?ӆ�'T6*"��6�#�@Сq~B���V����9G��e<�:=�^��?�]����!??�|�Q�����堓n:�+k����6<�<�
hG�a�m���ՂC�&- n�q�����ɉ5�@FR�T�K�#�`���j�{�D&^?�iz����b�r�]�!� e���bY�sU���A�B�b��?194
��&�Џ�q���}eIp��H\ڗ{��!C�NK�֩j'���	a�����U�g����ΒH#/#��%�lj��H��Q�-}��$.9#绉��m3�AX�F�ݒ���S
R8P�sᯎ/e�])�/"�~�c8��5��A7���YvGz=���S"���~V*�����A�G��Zz6��fb1;{����a�J/��� ����'ɑ��J
/ٮ�0O)4*vuu��N��U���&�=���!-C�ϼ��B�+��$��������Z�_A�vZ�7�7�H����USkK���*�(�ۢ��.x糑�P�p#�*�xN���9aTu6����X2'���j�1�e��ƒ-Qx��s65�i��W�C�5(�5�/g�WW8�x��4��K��u��B�CP\�_d�`%6ֽ�M{�W�y���$��_���ʮ��)�C؛�t������]L��ۢh�Y�Qv!��W�z����A`ꡦE ���#g�48Ƶ�W��s��^O����DK��I��Q����ԟ�l'a�%A	������*Fx�����������8�G�QCm�&aQ��0���٣�����|/��sFKK�P^����XY�^��}��g�D��/d̂'	�%�Q��ZP�1�Jiu3(� !d��m�YZ�o�����xK �����,����ɭ�maE���l�q�H��3z�v'��&�t-��:Js`}bx�t	2a�G����q�L��|ھ�:ό��
ħ"u6���cw�=H��mW���Y��C�H���5��A%���%�bV�;��:�>ꁤZz٪Q�$�}�K�(|�G1{�UD����rK��L����c�����JF�a�`4�&U� `����Z5��C�у2��H,f�zQq�9�N�k��1�``�H\Asb�!L,����T�m�~U.E��|��5m'�)�R�1�w�{�:��տ0H'���gXQH��2��`j���}���]g��F-!�`@���!ވ��9g�u�O�.����{T3h=����5�7��Ie<ԿBZiu��cC��DF�2Y�54Q����h��Q?T���L$��KPG��J)�������9j_Z{��T�L�5>��^e��`��$)���ņ��[%25�:l��?Dk���$�D�f�\dT��$�hOEmB��}>��h�tn'����J8Ka"���gL|"��p�^�'�"x;b/�0~�&�7(W�[Ìh
*�aj1�U�OMܽ��?t�"t����|,����s����~��KM�Ɓ�,)�-��Y��N�q�P�B������[`�s��ؙ���DT,�;u�
�1�cx�R��N�#;�.��|�R��a@��Ť���n�NN�z�1'�cv=�o��Pv�ع��߭��('!��ǈaW�oJLU�
���8�#��(�#Qī���bo�k�bpf|,�L�%��+4W��!�R�������R>��.�ା��LƜ�A���?n�."�JmE+e�ȍ2��x�N �����
D����q�~�$ŶӠ�v^�X[/��3�Z�vKYPZ�7��
������e���*����IN�̓���	�RjM�H�?�`u{�ZE�A.6n6�,����;;��!A��-�m�h�������!�&���;� !�t�
I�Ps��3-88��y�T�=iթ)�~%�����̌������_o�������]eRw�-?��0|п�\�$uu�3j���j�K��g�琧�:�x������*�x��b%� �}�㢑[��u�`k�M"�]H�u���E�|V7h͈[E�JН/_��fe��ѥG�)ś���{��E[-ҝ4�s�һ��1��8�Q�BOY�֙-Z_�"����ɛ��?y)���a?�X/���:s"-��?�|8_i��#_�3J����[��`p4��	H�"�jޥtLv5h��m53�]պ�#�8��")>�kY�bF�C%����"H����cj�����.'�*���mD��0褵p7
�p��'�(x�֒R�y�ć]$@���:~�i9���zl}���&t��ߢ�����Ɣ8r�q	"c�(Ĳ,�j�l: --Bԁ��=�@� �a"������'�*�E�*�g��w��[J�����>���2G����A4ɡ��*ޙ!Hբܶbq��=���C@�~���Q�@9ɗ�	T���;zS�J�{�7��e�YH�/��,���؞��� ��� �}gcW@0+(+>e�Q(ge��9	ؓ�V��ψ���K�1�x�	��4F�O�i�Flݠ*���V
�16��y[�~��P?�A�I��j�� $��W��D��:Z�*C_l�Q����	Y�~ ����(
��Ŕ����k4���K�J��s�����U�S쩙BdL_ۘ���[8M���]�p�Q:���:��Z3ru�P�YFg��7�D;"���Q��b
�{�m�(�P�� ��V�C�J�+�|��:l����`�{������msJء.���=�3|2S������f��,Ӈw�;�%?$=��7�7>���};�@�o��Ŀ}��_�@@\3��x���Ђd���B�Kd0���HÅk�V`*9S�oӘI(��-zz��"���	?���n��i��n_�N�\o��N�0�<Na^gU��W������!���n�</M?�4yzxU�2�0��'���� MZ�@x�@Q�P]q\��c�x�jݹ�=���0���@ժ����̅���z�Ԏ�Eԫ��.�<���y��tʂ�Q������:]�`@(|�tG>R['�Y)W��u��K����HF��!b�3,W;G�%�8d��c�%a�\�w�p�����=ऩx�;�E�p$Vz9ɿ!Pԕ/�f4���"-E���?�N�����΃������}��3(V�}�^��'xg3%5G5i)N����������-ȟ����Vha�H``dbf�Ct��ED`f�C��"� m����L���H�]F	�n�0$���v�� �2r�'p���v�t�!����������ை�����7{#f:f:ZaW3gF"^n{CcN!�B|�x�Lm9��]\\�\��l�M���􌌴�n֎����� ��!d� �7�u4��&���7�qr�!"�'���Y�JK�7���?Y����Uߖ@�@oeE��3����3��l���l��F��F֎��
a����N���1�YY}�:|` �M����ܿQ`bfe�w����M�������?#�����l�_�q
� ��,O\���~NC��!��Wc��>�!�!;�-3�-�#- �����J���Q�h�꣇��ǀ���d�J��Чefef��ggf���g 0�22������ǩԷ��U��2��b34b�`bg�56be�e2��| 32q�0�L�����"6�V��if�obDokm�w��r�<D�t��#g��h�1��̬m\�gH���H�Q�� V6& ������������T��>��T �ߑ?�ǜ#�����N�o�F��6�J66�<D ����a��2�w��w4� e`d�d p2�)889YX��4�E�������K���p��f13��n���S�Fv�h��ii���_�����}g#C���[�}���7�� �33-�1#;-3;-�>+-;����>�ǿ�8�;���	�|����ǩ���?�����]L���A-��H`'������j-7�����K������>"!��������%�Q�%�Q�%�Q�%�W)���˔��G��qU���5�q͂0��{�y������VL����4����Q\Z� �3�U�� D\H@�u�ã�D������paw�����|�44�U"?X����Y7(�5D��494!by*3�S��(+zj��[bj�B�MM��A�0X�@i��$+��65�=3�cȩ��O6V�i{nS�Q��Q՗yo�xx� ��������DB����������K%����(0u���B+D�(��T�(H�(�3=�T)W~[���q}#OR���u)��-�O�������^�.==������S����뚻x�كЈA.UѸg�Ӯ�X�>��T�徊j�DSs�ܦ8T_�����p��eռ�8Y�Z��}������M��W�ŧ����+"LzC���F�|�ݫ��`qc�	.�H����J��o�V>�I/e%�ſ�	�ݲd׫P*}�8�T�'oJ_��*�%b��*P���Wm�54�8E�N�6t�9�%)k��ީ�}$�>S�aFW�d�m�����³;ܷ{�=1Y��8͐.,,,���J��$�u%)�>�A�H�܄��A�W�߈Յ��TO�7��n�rc�B�'b_�e��]�~/��S��l�������i��HDV�W (�'"��>�(><�b%��D��;�I��_�����x]�� @�A=��O���+�HbfuyY�[����"ʵ���i~��C���8����^ռ��$�(S��D�@��3�*����*�_K�a�o�$!B@��7 e����U�2hZ��^�ۀ�43��p��Z+��Q���H����p�zu�H*�F'���8��rZ(�������
������z�D:�M
Uw�� ]�0v�I&u�m���[�u7�AdET\���#4װ�z%ZVRޯ�|#����>�H�nur1)�U3M$�>[ �ȴr�&�{r�.�{2��!�*v�D&���q<��`k/L��${im�m������������A<ސL� �pǂ�R��v�ް�ੴgw�0�R�4�QB�@�Zti�d�0&��r\�����Y�pA�{HM�Ji
^�iX��&箼�c���D�֐�_���R�vG�z��z6�~�,����ﾓt�(�z�lVU����455=��|���^�����CHsp���,�ϗ!s��{$#�{>@���� �$����z8S��Oe����i�����>P� ˂:�7JHY�M1�����M'^/���ʍ�.;�}V�8�'-ù|�51/���%5����V���n@�y &}U]�s,&ݕf� " Y�Q�$��gI�#xĔm4ը�Ք���o�%SX;d��F�Mݱ��97B�ݚ4��x�C��x��^���.�b-��R���wa^�g�&�D��a�J��)��:\~͘ϠP��])��\����a�uvN��������]��rqq��7�W����0^���Ea���=/�!�>7�@�Vw<��Ѥ��2�����o��ڦ�t9D�u�ՠ�~�v����jG��������+��祡�΄Q�����m�i�/�#&v@�oצܴ���o�&ѠU����q_��Πf^l����g�6�(���~R~&-�Q�B�@��í�����....b�K��5��=o��x�tC��n�+��c��Q��(?hb�	~T��V4��hd�	��g�mlo�G7�,�Ud!X��Ő�� �8�&��rLZ|�~�uO�2����h�O��D���o���E���"�扃꼅=�gCL��EGJm�>Rf����.?���O�_7���<@.7mr	ѡ�>K�N������(9x*��L���z�ֻT9��e�]�������zm��A����#Kh�����9�����I*S]Eh׿�9�1;<V�.�����<�$���3��ۢs������c�M�]�DX���]��~���kR7B��!�����x��=}��)�� y2�}�`���]��VV�r�"�Y�'��VG_Ҙӑ��A�ՙtP��I��ZN��QVw�(JW��*I��Qn��,h!��n����4���;ƹ<��/,��(��.��l���A���L �}�)�9������I(ؘ]-ᾠQ����m�;��$��;�����77j٠F���t�zn6�Z.��P��a͟�*4��0��*�x�Kr|q1�x���6C�����6`g�PV�����d���@��N��E�Hy'����εo��Qj�6Iu��\�����;��%�������5�-� M�ȕ�`�wf9�x���L�T����Q)�@�~�i�����s��Q��3�)w^�k�88�ڽb-��j��0�Y�-�u8���HH�I�O��}��ӦEs�UY3D�
�a���IH��Ҏϔ]�Ϗ^���X�TӏA⳩E�:�+ŪgL���e>N;��\c���^��?�r{f���K/���(�ŋ�����奥nϯOâ���(c����l�����E�U���c�̔-ZQ��;���?�gܬ@����ʐRa��W1��3S!�H;8�X:鞯f#p�"wٱ�>� z�ۇ� X��#�:���������9s|�OF�n�e-�=G�B���0)+c�h�s7�T���HZ�U5
q�&������R̳�-M�;U����_�Lk����Xt�K�3�	����@&y|F�x<�?��,���n��A,����T�������v�P6�����j��Tx?	e_�g�D@z?�ڃ����C�׭F�<D��M�Z
C��cQ�Cǥ�G�ti
U��7y�"���Ib�@?�OU��fv�lޟ��&���{)>O)���F����g�k2��/V��NF�ej^>,&�1��FXd�Z�t�<Cc+hU�n:7]E�����W6�☄e7�Z�UI9���ݽ=�f*�7s1= (��;�`�[VTV~�t؇��{���_���~��
�KC̡��B��,E���of�����e�X�aȝ�����>ym�:]d�>���1��4���z��&�ψuZ	ߗ�R�]��^�t	ӂ*�=���1a;R����>R�k��������IS��=8]���E	�Ɂ�!	Ӆ��V����s��tA0v-B�S�:��rRx`��l�e�����m޾ڱ��\/�Q=u��9o|o� P�䘬���HO��du����%��O�����#�����}մu�U?���Ər������o�vؕ�>xr�ɶ�ze�9�R�=1��-4-�Y�VП!P�Ѽ��Y�c� ��v�����U�+�o����ޅWHۑ�	:A��Q�Q�V�-C���Ion�������r\j�_H�X䪘8)�ٸ�@�[�T���;�Ϝg0aYL90>6�[k啇6p��u���"W	��-�~��RM*^�����t^ܞ���#��#n$����������N�h�w]o���!F����(�b͍��-O���;o���9�����"X`�p0A��bB�υI{���`�H*�'P5(P{�l��M(��`*i<��:F�OEGn^�Nӿ��+�_ۺ�w%ȆS e�������V��<���X��=��a�)�e�wv��I6��o��&\�o�b�3��ż��C|��=/�ݬLUY�v׸�,��z�ɏ�������siF�i�JD�<����� a�F9hX��i	��2/��Zs&!�	)-��<&�dy��MB��ԑ�zE��ڽ31�
�
J�i�����2���%�P�6���׻��[�z5��;'w������%2|�����bZ��ܣ��R�Jw��4��@%���xI��zO��4���O0��B,�'׾�a���A�������G�����;�|C)F��`!��Ե<�hd�(dA���5�h�@~�+��'䢒A4� ZA9�U�hX�5��ޙh�#nbK�.*����D[�X�X
�^��r� ��&�� ��MJpH�6�g<��KeZZ��,����b(������L��+��0�%~T~%Є���E���1�d��Cf�;�QY�]�f�Z�ˎ�ӎy��/��̻FA�yS$CaM	�Я��kgyݫ;;;/--m=�\ b�%�T��SM�>��@�B�8�V�&!n�Iǵ/�d�*�B��@�fz:g�������p~P�d�Ί��,bh̆kP(��QG�.W��W�����d���x6��K��a}�o�Ih�;_-����rަc��f�ҡ"3�ʑ�-�0>�nk���M~]��J�vf�@�R�Q8��|@9J�{�r�ډ�f;@��hR�y�P�L�x8�|F���?���NG��7��������������6D��V;���} RQC��(��/�3#����tY$ֵH�B��,���J{��5��cq��yq��Dj�u�������o�L+��%1cO\��Ĕ[WhV�����,��(C7�Z1�0Z���M�r?�2Y�;��B�E�)�WSSU�9�R���Ԉ�V���=�ak�;M�l��7皘�h�П|�������ks����R��]y�G�M">��+��?&�X��.�
���ǥҰ2��&��k�3�Zۿ�zz�������s�q�����}�8��K�f]�h<XnF�NFT�¸��iZ�oSC�,��Z����L�<����2ѝ7"̺X�����I]�@���)�Lѵ�<w�$@�������L�Mf3�����#���ﹺ�>"J;�����3f�;� &����3q���vB{>Q�6�H`�$?2c��[�̤�Ծ�癒!*�[���ެ��b�6tC�4fB�Qi�D��8͗v�̇HE���k�?w1WنMR�9C7�4�=� �۾i7�U�]\
�R"�ʬ��;H(�؎�(Fl���Qθ۵d-<~;��{�vT��t��g�:&Lt5�,vm�/@���ml~K�E�`�z���������� M��
��61{���_\��߷�*�����fљ@Q�5�EQ��/�I�Ҍ�k����x5?o�����o}}�d1:�i�@uzm7	^�Q���r�p�|aY=������`s6F���P�q��g]��/�l3��3���F�k�b>��D����M�Ƿ!n���/�Hw�9]����5Ry���^�9��V�Qdժ��8N$��=ߝ|�؋w���A��ߦ��[���_�)���(�)�ЦMHb5�z�g=�r�q3��3
w��׻O�eW,�����Y���V�:� ���.�����_=���4	L+�����$���M����z�� }�5p�df���U�lZ�Fٜ�� m�Qz5�?%��X���GWnM�p��];<�":
���Z��^;�F05�o�e���A�ey�ғ骗r�
ٲ���e��w��L�r{��<�\ABp�oK�ic+c	�1��ܣduғ���7:����ל�ő"����IHF��k�̦��2��GR��[Peu�g�]��-��<	����hP?NO0�N�q���NMR+�J�
ɏa���u6�賨���h�\�~0ϯ�φ�g)�^<����P�����1����?C��zSڄ�*i.���[2������I�	̺���Z�4���3#j�[��]N0lOYD��,p������۲��Ĝ�#I�H�	�\�nV�)Y�a3�g��%�D��݂gh0!��H�!���Md�
]U��٣�+1�4hg����a�"��d4����cO��j��l�L+�2 K���q��в�Xe"�*3F�+N����Վ��_E6��]L�K��*И�I}��d [��_��Ebv�H�QY��(W�>��fH� y���Ջ���4|��V=f:GLhx�[M�@�HѮK���k���*�4o�J���Ob��\eb'�^	�V��S/V`����p���e�It�%J���L-=�QE� �Jײ�����^Å��нI\f,���ز���l��A4K���1Cb��T""U�?s�(����2�õ�t#�{�Ȃ`c`����*�5X�5+� 5`��X�����D�HGXՈ��k��6�*�k�j�\z��B��T�
�Jyf���	_���t�8�Y�������D۴�3o����;��b8!,��LAN��m��N���,����9ʖ%F�
7���ܶ���lE�~��X�j�x
�\�04B��U�IR9FA��;J��Qd��$r5m\(� �yb8���L)�vf&�+�n�Z��:�B!5,<�0�$*�M��c�4 �V��S����a�U�얽�fZ����#��ǻ6?�(�(O��}q8�Læڕ{���v�����ݥ�`4�v�1|��^I	���x|����#gf^j���3��qX�b�t�AY��	i��3ʉF3��K�&$�D�L�mޚ��"��@"L��+\J��Ue��0z�i�NG�T�9�@�m����y���ET�*���$�+NI_Q�������/�(bᇠ���Mr��1?��>ke��W�m�셸"9d��Y{ �)��$X�*����Eʰ\	��+�p�M|���A�@��B^�Aj%Ҋ��ѯR��_���ú˳��o���ERB	����+Y�%p��U�&[A���F�e�$�IV���E�J3@1Qv�A#b�G���u�sA�yU���Cͽ�������o0]/s<� #ǥ�W�T�t��rNK�|q+/*Q����$7#�)���m�2�&�v�e�r��0{&��-�'S"�s\� )n6���� T�)�
J~0|�T�yu ճH��g�*"Mgy.�b�W_�Ms�z��,B���F�%ع�`�G"P���E�M�^���|i�Gjgc�q%b?}��QҍS�T�h���pj��0|�����^T�&�Ð�ٌ,���'6c�"oh@U�~{��Sr��Qa�Mڕ�w Q���(�ZHiEr�%k�����dhu��SL�.�&?n�i�T�k�-%�z��2cuR����]���_�	i -���n�0���:.L�R�_dүß!�=�;ѫ�~�3�8�c=m^15oKoܧcd������_B^�p ��V4������1~����p�&�tX9c�G�ml�^�_�N1��]�khP��=?��ێ�)��߶NWu2��~���EЩ�\z\�Ќ���c�,�;ĭ5�n-PdWS��nY_a�ll��G~K�&�cЫ��V۽	z�s<o����xӐ�g�m�L����-��}"/e��+���3����Uϐ�Wꯤ��F�f�Fr����%G�(���:��Re�����,-����}�ÇfS�lĎ?E��"|�9��p���1hɁ���]ͫ�&H��&�Ky*8�]��BU�E9�$��M3���7w������Q�C�eNl�ӵK��~�(%��M�H�}(w�/f������K��kO�P��_*F�g��H($UFt��]��"��o�_|?2`��ynsi���z�<��\8������O<I���EL���3ŉ�b��[o�7bŠ��fʄX��r���������`x,��������0�����Un�{4��˙�R�r��Ap7����ps�4۴aG�ּq����}v/�9���߂��m04�J����N�C>\>0R�.��|����wu�!6�<�9?XD׼��
�+�G�һ�M���j��\�2�ǚ����y�JAN��07����m�.һK�f��~ل��\K�^�[�9��U�s[  �GO�=�-����Ц)��6udǛ��d��R�;/�R�h�0Mc��J�P)Q��	*� ��_���\��r{��Z6z�{�M�D\=���
v��,M������[@�K#L���+N *b�I�+]�`�ަ#v�e���AԞ��[����M�g��)
g���t���]�� ��.2mb��8���`�Q,��3G�o7n�F'9%e�Ie?�1,�'~oψ��T������N����swsKS�{9<�QC�b��f���|a��ʼ�NGK!oV-qP�`1�_,Ku\�L��viY��2��(w���vjJ�kg��)@l�̅���kP у<*�#fٷ�]�g��N]�����)����0,�țۤ�?�w��D$C�^Ǝ�z�<f�7>���������y�0	 ��\>/h�st�,������������qu��O�$���h��l0acO�ƶ�hb۶�4��ƞ��;������9��g�uc��Q��5�Kw��=���p<�j�W����5�\�&x�^QQ�}ve������p�]���A���M�c	��w���Ў�,!/�.��+��p�&LTJ�K�E-���<`��3�@F���ڿ�`�a5�*��#o��h���v�H
.�\�hMS?&*ϒ}��B�hX�T�<����^�}�� �.�E5�J.����q���ə�X�@�/�2$�nXF��#a�Z~$[:���Ю#_Ǵ����@�l����T;'���/珜��ʣ��8L�U�wS����O?�x��,;uE��=���DK�W
�JĬ�DBBB���;ħb~/�b��i��p4wK^�K������Fnn-:M/� ����Ƒ*r�x�ɰ����h�O;�r��`RY@z�M<�.�	������g�R?��N�E����a��K�?���8�UmR����*u�a�~�����%�xP!w}��t�\E�E�g"�6�dp���{����75!;d��T��mL6�N���ճ�D
��x�hb�!��[�i���b-�y�&�cl��딧��d
�{�h�ܟ�J��R�|և��K�n�z��&T�&3��-�4��w��	�fB����-I�����+*D�Z[��LeC/l�VVv������hx���df/�#f�����:k��e��-���~O6�6�It�Q2ohlTTD��^�4���1 I&߃�Y�l��!��c�'ss�lx�q�ݛ���˳D9%:�������Vl\bĵ[�5җ7�),M_�����TrC$�͔٢�r�A�8aO4���t(A99)�̵�j8*
%�����%Te���M8�3�V��7��𛳴P�^�Y�܆��[�N�ǻ�cW��A wO��8���Ѽ�e�޿Ƨ��^C^�����+�	b���~4�	���_��>�����?ϥ��ؖ�J�7�����vjֶ��ܱ1h��5�~:-s���F���Yg�ϻ�>^o2y�~AF�����gt rz}t���5����v��~�I#��:�UZ���S�ΪU+ރO~��R|����ƚ(��h��<*�Pmc� ���
�3a�-ؙGSD#����]���w�&�`m���=���1��,��.�����V���c����h;N��?;����-R�������Ţ �D���yuu��y>�/��b�H���=o�o��U���#��Wj�������Ii���P�y�Uv�!�1r���	���Ǒ�����r}}}��������������$�Ͱ���������t�夝o�X(�U�[g��S���b�/�����?����kk{��b��Ḡn�nҗ�?�n�b��ݺo�:���G%9	9�To�9 �A	?��o>�w�����1��+��!����	�4�B�����nW{�W2�d����u}����D[:>�,��'�^�x��c��8���c�ᑦm�������n��}�I3�i����&�OI�Z�V�e�k��O�U멉� ��@�]�5���� B�qa�Ә7.�`��K�{Qtm���66W�	;\t=@�;�>����w�]��<�QR��Ѥ��-'�7E!�<�T�ZC��?���n����9����a�����8�F�y�gc�xѲ��A�eU�J�eu����3@���\������뤚ZHqo��~K��/��]ڶ�C�B�l�B$�[PC�l\ ���uG�K��H�+����{[����B�&�}� ��d��Cm�Y�v�0�nׅ�̫�Fs^��%��]o<t���LC�8�mZ����f K��q7���+ƭ�%TI�
���49���%�'�p�;4���o����l�9o�����l��9�V|���'Ҿy�7� $��*1[��ȅ���������W���ϳt�(Ix��ֆ�lQ���9Y5��`]�_hO׸�p�!�����bkV��4@R��|��6F�7�q�I�TO~ש�k������%Sfxg �|z���6Offf������K*v=m>�n�������RD&����<;/|.��{��-���m[ƽ��!)�o�Ї�p�.�66/��帓�w!���E��P�o;�O�7߄�Gh�*z���YUˆL<��%)]��$��D���%�&H�?�����伷��wf%I�!�!��(�v3���v�A�E|���������~9߅��mÃ�m�޳�(L���TQS��C�s�3��J7��G�玮ܵd�NMb����Q����h��@&�FA��HV�+"/�2��|���ĥ�2������l�&�b|@*%��E&������|l��z�䤜�m{��ypb�-�O]�t�bx�����n������6ZJv.�Uw�ߍ�;���ɿ ^���/��vݩ��%-�C�
$A�Y��s���a/�r���7�o(����뛝�HF&&�M��Yۖ�p7�*i�}}����|��X��Jr��W�,S)yܘ���O���B��G�e��fIއ?�U���o��v��q*�txܲ3��2�Ѯ��I?�6��U^�(s�(59�k�3c���ٳ���<�?9][^���v��vF4���O�9��w��wK��ЗOܺ��F���?| �6S��9A�-(j�n�wI�5�|���p�{
�?ޒ�J����"Z╎�OT�������p��]�㐴+��Ь���B	;���WG���?�3|lj�돣<��>��lx]�k+(y�xd�T}"��FKNOOU6nX>����`��\c}Ҟ秙R�{Msw�n)��� r�6�)�Ъ8!�Tb�������ق$*��5<??���'�-��Ǹ�k$sq=>/�L�S��H��)��~9���t��d,��m4�T�\x��ᣆ�&<O(�.(8�уY�r��KH_��&�3~W��y�������>��a���g���X�{��%��!0����U:9P����cP�&w]w�s����A������C6oxmq�vF�o..�1u�k��p�h��u^M���V���1�++i#���z]� ��"aإ�=\,e����x��v^S��W	��m�&T��-=�5oϒ�_.�,�B�f,���������]f��N~�7٤�ͫv4���DZ�b�ƽV��p��N�${n�>o'�9)h���'I�}�M��_�dB-�@ځ=�?�o4ؚ�+k����Gؿ)|�SߊRQ�7��U�����5�@�n6f�����M�-������O��[f����/�rY��K��]B1]�|6�^�vH�~��8(����gx��Z:G�:������7n
.z��Ȓ��;�a���nP�� �S���㒰�T�� �'pN��	y��kReU�ͤ�Od(�/>��t���[��ϱJ�}S�~օ7͙�"��m"W��m; =���Z%q�)�/JC0'�0���C3�T�zi:��h�E�m�j,uE6F?.�ٲ}%� �M(���ꍹm��f�qĻ�+jhū����B��@� �q���Mt���o�~�n�4/)=I�ta�YCd�� 5�����)\�d{_ۍ#*oޞg70�܄�=J��t����[��_�8k��K���g���vZ%nq:����~�&������I�]--4����	#}0V�����Q�*}H-��d��m��tД��1�E��0�X�����*��:,����5���<<�������mѫ��{�2z����|��o-|_Z�2�%ޠ��UN��_\�;Gd}vn�4I+Ǫ55�;�����d!B��0PX����Y�9�7&y�F>�bVH�;�5xf����	,���9�?~�`���֑��g� OO�!����-*Y�1���f|��kq)t2�!i�jN�zIJ�2� FR~G�׍�8<�jL@�
ۯV?��4�2�xE@ȸ睧N����ܺ.�)[̩l�k7ѕ�:�2��W��ysl�(~�Pn0U�*��R`z��my:MՆ�d��ȵc��o�K�Ƽq:�o���G4��JY$d�DY9���=���ܖ74�؅�H��l��u�j!nhj�_�e��c�-vz��`�k�*����ֲ�������a%bH-k y'�ф��k��*5�rJ�G���.@)�#��ɻ��e�ʶ��3���4B���#��!�ʿ6��6J��T_2��JW N��=�F�{�7�J���@�Rf*�΄J��������D���K��df��Փ6yNC�J_�_�D�c�tA$���aȠym_�G�1�4�
/\�q���Q�q���+jP�o��u
��>޻TגKͤC�&�_��Jؼ5�3%�T�}���q���ݿK��b�����kf�bO��BxZ9�D8dc��,`	Ef�\�vD8"�	o�a{��ܿ�Bܱ���`�;�F��[q^����խ�ԢZZ�h�XrF�b9_���'1�7_0g ���<������~�T��f�0lڈ���X)�a��.��ɰ�ӕxqj���h�'Z������Z{_d_������lCvW`1��b�2_�4�`\��)�O�~��`�����7��#��'�M�aMII	WS�sg�S5	�W���vk �O"����U� D*>��I"�5���z�K���r�ku�P�d�=�~r?���<[�;�<�HḾ��k#]��>�D�C>�EA-�n��g��*���б������#؟�a�E4���DT݃WLhDW���ӣ�����9�*�qm�+GÍ�kV�R��Eḋ���F�ek�
Vm�F���5�U���^>�*�w�����Ge�	����N(�����2�6e����l[dmkƾ�#+�`@L�K�na���z��W�mv��g�ު+>+If���x�:���޶��f*_����g�9�!ꭠU�<����~0u�T#��s�_{�D��4�# �	������XE!��y(�J� a���j�躇9PŎ�ܘ�UЊ�S���i��Y�S�))�ϜQ�ϺO�ȆS"�=� \Q�|��6k E�?�N��G��H������ cXr{�[�ò�-Ċ�/1QR��\�Es��rcs�Z�|)��{=����-v�v`����g�ĕ����Rk����r*U��q���ex��g: �_-�$-a�g=�h	���ȥ��T�[�(5��15��"��M���ؗ�7�(0�Z7�+�hŵ�yG�prB��z\H
NB����ԩZ5���u-l��)�6�.���c���l�ߨ�m��Z$��+�T����Ň�bb�h�ʖ�����P�0�u?U"�Frڊ&�fe$����B�h�n�N�%��N)-	y �8eZX>��R�s��`�36��C6sB@k+T�P+U��d'�݃�m�Z$�N�"��`��!�(T1�$'�]�* �I@M��$f�Nm��[��&��|�Ă��n_���7/R

_����c����	8Ӻ����P0н�G��̼���񬿡�8YNr*R!Ɯw��Г=j�$�� ��x @����&�Y�/Bվ��������I���>b4���7��D�%���m���+�"O���L6j�X����7Ԫ����t�^!�2�$�ǎoa[�I����'L�L%o��M�X�rX���}��`Q�A�"'��u���+`:��Y%vrρ����Xr�+�2f��iG`tE��aUNG��|�U%�Ac�z+����h{�"YN�z����'y�Q�V�1���)�NU�_����ZDࠑ��;���e�j���s�a���Q �`@&NQ!㸹[���
�X%�Z����Q5� X�T��a�!�d��o���*�͚"3��#����76���WTP�����G��d�W4�7���Ц���2������6..�Y_�����j���=wf��.�5mf��)84�b��}��"������l�B�G�*��yv��͂��zo�wBv� .[GQ��QY���͵�䦽#��0#�Ot���	�ߕN��ftN�z�r�~�ID��}u\mJ�����r�}�6��2,9�a���|�e��V�l�'C�Q6�;r2=4�#���y���Tx*wUm��ٕ���\FFD�f$�tt�����0f�x>�w�0-������V�+�rw_��n��n�8e�BCc�
����o^ۻ���c�G�!Y(
��)���F9��nQ�?�3W��VǓE	K��v��H�=���$"�,P��iMBUO�o�o�qMB����Aq���2w �%N�` �tFg��b�����1�s�� ��<j�t�][�7������:��6��P�,f��ö���%�~j)�57Rh$R!�k���MY���Ed����g���
ӎ�䩠��5�3�ly��kB��Q���m������Č�d}_��O�p��]�s�7%r��&�"Ȉ�3��0����p�h�I����z6��� �p����.�6'cXU�2��e�1G�Db�Y�	UE�}e��Yd�����$�,;WV{�� %� Ǎ!�=�0�'4%�sl�2L��Ʀ�P��}���o���{�^�U6��-���g�Ѱ��.{�0&oR�R�4�8f�j�h6����d�5H�׶��B̺��6H��9�?"�*=߲e�2�.p���";�b�U�����g���#���x: �Ɔ��*���^˨��Rs�e ��ԭ�t�Y+�2��j�B�Ƃ��n�٤篹���Ks�bG ��YCJ���A��@��ˏ�ӓ�� !J�-J/MEŎK�@[�(ΐֽ�U=�����B�^o�C��~���h<�Q�#�:��h�vTg�u�M�}lDÑ�Y{��;_���K3���#�3=ޝ	�'n2���q	���N�4��`6V��CnkL�@�ɌQ��k߾��]��X�Q�
�q�Y�  �	�� 9	J  �+O=�:{�&oܒ�ڳ�SD�5�g2Y�ޙo9��^�>�ok�]z��Z������*�� �\6qQCD�y|7"�9DP�ޠoc����zD[ޮ{�_}[�)J<2���ݴ��-���2�%`�zƶ�;;I̺���h�0���܀�+ ���{�つc�O�w=����V3P>���'K�G�2��NyF���11)	Ƕm?9�us��Z�v�*�]��e��ٝ?W+����w��FA�\����u�TQ��YX�"��G��Qw�o�ńz���(19����	>K@����W�O|ƥM"�A�1�5LCDv�-��,0ԓ(�5ñ��D�cE�6�0m�B�C�4���B��[���S����匑�֧��t˘|ǵ�}��#���\��36Ә7�l&��s[���id��]Gʘ;����4X���h������SӍ���(��q�mn���^s0����jjn-�=29{���/x�T�.]8��e�/�|^���zX���\�2 �:G�n���ח~_���_�4a���G��o3+g��'�gC�?�y�Ki������'��c�3pL*�6�E�	�/>-8b�����4��֫;T��j���nPHg�^����I���D��e1Ѭ���\m��.K�d ����ŲS�P�&B�[�]�:��L�>�0�4�
�Ho�փz愘Di�?����w��|�%�}��OaHSz%|�g��R~�w���jLu��� *��y0���o�`s����c����*�H��D���P��Gw�Ƞ�u[��In��+��͹*=��P�<�$�4�HQ��+�ݸ��h��@��C�-����k�z�\�9牮��������Md86��'dRU)���z��������}37mt���~����ꦵ��S�э����F��*u�����ֲ*DrJ_�;�	�@�H�t�N�6f_�J�C'߇��� ���SP|��^��d�y�$>�TK5و�455��9e�a����<$J:F̭���,u�8��s���7Í$
`�a���J$��[���f�"մ�.���55r�M`����߷D�i>�?���w��-h��l��ځR�_s��
#���)A�{��1��R��Zqn��;e�j��屃�DM�8u\
�Ҵl�#sw�C���o�9wUr;<?9��Ifы��g��U;�z?�Ę`�S�̦I l#$�U����L|��|�:W���ۢ���4�*��+{bޮ=%�(�B�pq�ੵ4���.n�>���=��i�16RK߃J|3��FeK#$� _>���X{��C����F��)\���v ��H�Q�@�Hb�X�r2-�t�h�Ec����S�-���>,KD�?������1��]�3�=�p*�t��躆�1G�4qQa�O�xP�q|�q%�sC*A�$��!Q���"��A��+W��/	��{�_Y���a��3�{i���~���C�y(�A�d6�&I%��u��ԱŊ�)o�§M��傴���i�Q���`��X���J�8R�:��Ƴ9|�X��i%�i��[�2	�?ܦ�Z���&�޾����J�zO�l����6D2��Fw���H�Q���9zئ8EA2tf%1�C>ؓ"�]YҺ���8|�b���Ҫ���L�]E�mn�S3C�E���#��Z+�b�-�SiT
�IB�ۥà�,���`�Q����Â�s�L�j�0Q;�O�#�M�{����+���Y�M�[���Cf��y��dQ`�U%H�@��}~����1��O2j��ڱ���p�ɘjH��5��+�u�����_(��u1�M�,^��y�;�(���
!�V\�=,�<.��Q������<�B4I	C4��ӒͶ����^�rFJ��Ey_�� 5kڍ���x/��~Cox��oϽ�A�S		���9̶e���$���G��� *ܧ�%�U��N��5������M���+O˦/��T<U}j[��������Z||%I?�T�.�!�L����Z��S�I�CO�$�.ya�ԗ��v����RMG���S ���p�6��\�W\k�Arە��ޗ �B��SunΒ�����Y��#��R��R*pﻸR��!w��F��y]ck�,�l[�H��R�yE�EQ�|��T�O�}֎�tq���s4^��F ���2�Zd�B� 1��V�|�]nn]v���{p:�B��u4��6���C �y9U5�@ �Oh�Yo^�k퓚ͺ3Ĩ��6���?+�e|�Ev��]W>�b�vs�q�.j	�J*���#���Ƶ55<<�Uړ��y� �SVޜ&�"��-�6���a����KJ'[��?Tv�q�N|�r�,���apQ#}|,ۄ��x�?Ih7�W��u� G&�$7)�x�d�PC�u�n�@s��(3�F����|Pxƕ�!��P�1���]4ȏo�c��#ƾ���B�s���Mwf*9��ҺJA@���_G�[��s`�c]���H�y�ں����;@̍�h>�����*��|�����l�����t�㣺�l��*�U'8��[t�}�	�7�	X1�.�%K�K�i�ӕ��\�ur�S�8P�'iA��l�G�N9����tGd�;AJ�����{nK���J)��f��/٠?�0�|�q�plQYF]]}̾��&��T����j1�����V`�6'*
�כ�s���1��ЋKYxA���+)\g�yJ�G�V�П0�j�F;��~U�p"r[s}K�E3�`ZL��B�� �s+�khƍ�5��A����4L�m�NY$�1���)��`��c鹥��Y~�ŵ524�aƸ�8qvs��꼿�3s���\mW�)�~�9XG9�x�,9Eڞ$&c\��5���2x|��_8>���t., ��>��6�Qۜ1T,u���%g%��������n��T m��1K���bAd,G3����x���Z��ܻ�b]���R�eӠ3��Ed�O�2_��� ���M�<\����2܂_$�P.��_p���$R�2���b����M�0������~���U&ˇ'�>s-�dL��,L�X�V�<�#���K�{��"<��L�D��q��H(�_��`J�\f��E)�X��Q0��R?���~�I�3;�Ș�w�YI�LP��(�hX����>A继��0�FB#��9L�q�om7�=~����*y��`Qog��F5k��c!�y:�}�Ԛ�������U�`���q����}z�6��^��yx�M����h��D�w���E�9{���
�.�|���5�U:�e�|� �R�Wx����B�	��n��-�
�ay'�#O*�U�[�:{����85����ig]-���s�m�4�4��e�()���ꑑ�׫�+���,�F��CK~ez���u��3�َT:@�X���F�2j"(1�A���|�mr��lq����x5��I��(�y�΋j���@����D`�b�w'\�jM��<��sN�tGww��b]�$Q�)�Ά��/�����+�1�+���\e#��;J����f+ڽ��q�[~��"�����o�A<��_E�������F�A�C?ѲI��[As�m��� &������Q���
>�Ns�/���'M44�N������࿐i���T�ZY�/�Ǳ�}컽��Hz~w.äbm Q,j������K�gѵ�Q�����ݻ����?���/Mu�|�,ݡ�_��)����ڠ��g�T欔KPBD�~2��G��̙S�QRͥ�����\
���������,������`�`b9�]��=��|�y�9���mO]�L�{��`�����]��s�vmYL�A�z�0p6`Gx_�� �!~�/��o���p�e�}>����O
�%J������0�U٪MU�V�{@����͵�߹%�.����|8�K�����q���,3C���`��C0��'"3-��/���"����Ԍc�&���hRx�T������w��,�L��(G�����BT (e�Nϯ��'�#e�G�lLq��wR\�Fԛ����g*.�SI�Z�/6w�g�,�����C��g��X��S���z�<�WI�v84n�h/χ��㈠P���n�v�[V�����3g���nr]~ˇ��I���B2�k�úqls	2� �V/!Pɩ��������^W�g,d�nۇ���o�1� �x&�SY��rY_�8��� kH�T��w�¶ӱk�za|��3�>͓��w\�.s\`ܛ}x�(�,�=v:��������ՎR��jIg�HiSPk��U[O�K�܏�D쐝N���]�z��0$�w�]��Ԍ�&�NeNy�-�-�|�����`�.��0�S���Z;70��+��}��^xp��[7&�#��Z!\�,���V$^<Z )��f)B��wf\���L�����@n���Xi�U�y��ێ�`�0�z� Bj�s1(�ǡ`��V�.��(�/V�Q�s���(�����4�e-�6;����v7�hF��')�\�	��Ϛ�e0���FU[�3���x�$�t����ꪣV�e��B=ޞ�lT
��֠���V�u�o���*loW�Ĳ�N��5(�tҜ��/m�˚��|�D9�����t�����^��R��"#�5��������>�_�*	ѷ,�_]��Ɖ��1�q	'�@s�����,�Tԃ�5Mh�P0�i$���	-D0=r�@�u�"˜sſ���g�n	Y�"ou���Z�pl0�V��ʼ�:���>V����O�����0԰Z�X�B+�R�J��	�͜M6��U��*AKr��Yn����
�2�-�*�,	XH�9����Ĥɗ�A<��D����i����Z�bOy�D�BQ��.��Z\��U�o���Smٸ�N�ȥ��������Y&t�ᢡN�2OJ%3�5ʶ�_���QK<�%��u�(q�����#��1� )R�W����o�c����ɬ4aL�<�*6����@���+�v���A��M ۯz�I��pL�f��d��e��Q����8lB�gЮ�g8�ľl4o�<򲸈�"�����1�<���ji	�X7T�)b2��:��Xz����]!
9ݬ�<=V|��ǝH�?�]ps�[�J&k�_�L��*�e���D��d��4�N��7/�ȡd���M>(��`��;:����G���~�OV|t ���.����$X-l�TD�q.�$-�wL�3I��_P?e����@I�sz�@�)8��dY�F����:B�U���I�Ʉ���}O7iE���3M'9.�w�\>�W�QQ��	W�c�����P -G��\��~�nޟ�2Ƿ0���;���'e�����ː%QM�I��Lڭ��y��������N5����N�p��ے&�Ś���P0H��|��l�~|z=����O�k���Pn#�i\p	Gs���c��iB�O��%�^6g�P����w�rx�����B��|'l_/�Y�kA��p��ƃ�?"��ǡ�DIA�U�5�dp�a��_&��%����qۈH�6�!Kɜ ,��	}g�����%&H��}�lI!I71k]G^rƠ�f�#\t�&r9�������|Ʋ���.�V̪-Ǿ�͙H*��\��R���W�ל�ѐt���egBG��1���q�\�Y��y������%����!$�Ԕd�ĈQq�
L�|;�������zFdѽ��� ��ܮB���oi��j^@'�L���+0D�2��3'��{^z-� 6p;�јhX� ���e���;H�ZQp��C}�V�߫����
%��6rZZcs�0��5(2�4��V��\Y~z�A��M�?~:�UnE��}��ڈd��"��۶D�x7#T�Zwu�?�Ed�
��L�}�F�Vg�U�52ʒ{�罸R��2������zo�9��R����G�A����)�ȁ�m>���kԍ��/�*���E����I$�E��v�Ϫ�������oGͶY+�6�kQ� k�${>���M��M>O����Ң�*CES<aJ�<�r!b0�
e!TmE +am���	���GP,��4��&��#n�#s�tv!�/�*ܳ��~�o'���+e�(b�ۄ���睩�<����GC<Y���yT�!��o�k�����AdDa�p��o���MǋT�NW<]�G�������e�V�.����U�<NMR���X��k�ݑ\�o�<��*.r�m�,���BLJ��j�vb�Q\�������^K�o����Y��|��A��q�MS-�;�X��aP�w�j-����Úײ�n�p-��񽇍8{�'�1|l����roq�s����P�hE��dZ@�@��h�pG��
���B}��԰I|*����	b�Z��&�H�g���ĮՏ���$$�+��*�����2ۊ�G��LJ��(*�U	7r
o
���S+5V*�p��L�w�P�����d�UT�ڶ�bb0�c.��R�Ғ�H}]�/�#�E̓X`Bp^rn���%�{������Y��n~<�=m3��ݙm��S�&ۧ/>5qz_�5����挈~�_�����g]�gv���D�Փ��M4���=r��=N���8��/�����������ꗝ�ŧ�9�ҧ��ʿ�B�ڗrM>cΦ=��t�Rҁ΂��Op'�-��o�mSQ��'�95�%�Y��y�$�QI�Ͳ\��'����](�8����?2GD=r��K ���Fv�a�In����Q�X�DB�Ŋ�a>�\�ȒȢ��E���?�S6X���Vqf[��rHm�F��FU�e~]9)������YQ}֩�K�@� ˣFP�����Y��j��;1�D���;$pm��������b*)��N�ie;7>ƶQ�PY-4Xx x$!!���+���kXT��&��_�O"� �t�1d\�d�%�.�˧���������u�[>fƧ[;˲��H������C��(�B�9�h�d��6뼹����{:�|8_IP��{�Pâ�޷ݼq���DMs��������ǲL���J�LTz�d㒋�P�N�x�[��!/-�w2F5���r��]I��'�;�(��*���ɑ�אm�,�,���릐d��Y>��W���3қP_��oTg�g��m7sr�g}�켿�w��zH���P={��%�t�8ьɓBG`�=�̰�=~�z��]<�)R4��`�=��uZ�N)��ن'$ɰ](D��Ȼ#�D�0�aN���RM�Z2�'� <~d�H���=�=�Hi�[&��;�gQ��@��P�ƕ;�~"بw�y��*�	TZs��h� ��JL��T���'��\G�T���DF����^�tv�3������	u��"o��Zgݰ����s�R�t�;;��VSMτ��������a��s<>c�_F��������d���:�\u�d��+��׼�&�(spŁ��f�("(���y���ݺ�ݘ+�e]�_|�i�x��	��t�t���8m�eŊ�f;j-ܗ�n�
��9~����g�<�2�AC7N�W�dyςܗvߖ����n(����6u5����]��=�E�,OP�����.q������Ă*@�v�m�\� �^<!�s�Ã��>XD؈--�иY:��^y��WK>{Fc�$l𵹪�w��
�����Ǜ�y��Z%�d��)naW��̟��R	uUa��[d7d��9&��0��"@]W���;u5uߝ	�K�����b�)ѭ's�E�.^��U�f�z�z�������ѫY�H4�����C�}y���=C�ӎ���&�����l�_:��h,}�������t���(2��|39�Xp��)��~!o/���K+�Y�sr��=�ދ��~���5ˤ絻����C�`7:�9�,)X�V��{oǌ2&"�R"�]z�|:���D�M����;�c�'(�o֕��_��������Љp��t,Ӫ�r��B��(�����ZQ�(]���J]j�=De�ލ��(nvp���v�ƿ7�X�����R�{��D۲�ZMF!�Z��G�L�9���I6���1��&4��G�$�csu%=�rO�D���>�$\&�7)�dZ�LP#��ciyC/�ތ�
�w�J�^MX_-���->N$ G��W*��pk��;*a��~��V��&@;�a�:�«�hxM-PY��M�	�#�<�p�v�j��2͛=��/��Nd���~�D��hL�؆�����.>JY�����j�{��%G�o��yꉛ�a�U�W�ܯ&B+���xu����{�����[AV��d�i��/�����[ Gm���Q�m~�����/�jҧ��;�wK+;<�m�_[�>�ي����7fu�d����]zs�<�����U�����n�V������.�i��s4���D��V�����W�p>m*FJ��Ƙ�Z[q��D�tC�୙� N8�OR��'�qg��ej&�M��݋D�{.���SU�J.�I��x�(�]e�d�swN�MK��^]tM�O�Șox������������	�?�Rx��_ߦ}%�GF���/��.��AGw0�Q�L1��E����q.��z��jI
�~�XQ�\"�:�W{N�u��Bl���t+�rn�v*���/E�;�u�ZR��F�����).Z�j�WWl��n�������t��AI���6�6~~���\�ᬷ����E��4"n`��B��*K�چ��5�h�y#N�F�f�G��(p���Z4�tb���@����(�}j�]4��%�ee�	�X0"���&\�8���',����^�
�����u5�x9�0��"Jl�i��'�Ւ�Ҟ����.�S��S�hO n��^����T���(���I����!--�_��[b���v[Zx(��7U&Z���ߖФ ��p���G��JW�e�"��2�n:Yen5}
�� կΑ���<m�%(�j0E�x�
���o/l�5��F��a�'� �\(aO������3lY0əh���%9���BKN�(��9�.aPI�;�(��^7��>o�·�������#��pt >
�D��ׂH'��懕���[�~ʼ*�N�Y7�-��#�4���AK>���Q\OK}YD��{��%��ߧ�i����MmVU�T�pvq'U�e6c1��$IDqw�F*�{��N^�
�%�9��Lj���F������V�G/9��ɬ .ek�hp��O1������;�[�)�sV��\�<�.�����a[��a������W_���:�U�J�C��l��ο�I�N�*��9�r]��y���b��O�-	�.*�I�t�a^nL���P���3=A�\�E��?vSs�$�K�,�lAoW����p�ț�Ef?���G�6Q���/U��L�r���5�p�hy� ~��;��r>m!�@e#-\^�8�~�fR�����'o����mԄ��;�
�����j���0N��.���J���!�k)�R������
ww(w�/<���e֚�L��}���9s��S�Y^X���y��K�%��A���Mye��42�P+�F�9�x�_y�Ys�<����w�rt�@bXq^�#����I��AI.X {�9��셊��?Ǡ��r�b�('�ζ��U�N��x{w땱VV�屳��'9��z`ۅ]�n���$�h��^�ܼ�K<+�p��r塼i��n��t�-0/���ѵ�>`�}Sy"D*�o�i�r:/�Eͼm��0.���������g�v/���b�a�`�D���w��^�_�ŕ�	V���Ӽ1���.�U��^���S_��j�8W9eL���@/Y 2C@-�����u�c%�^z����0��4��$3�$�B
M�ܹ��XxM@�ӪP����T䔢�x�O��^�"c&���"��Z������2+no��v�}�n��hLӪ=OI�uQ&|Ji�k��HNlz������g~�s=�sj�w�lp��t���#��r�g�B���J��i�_0�+tG4����vj�Z�@�A<��R�T�ϨH�_Jٔ����Z'7��J�=�%��<��j�p����?�r���_>����v���A�}~�����*�<��#p�y�0���A%�����2����t�Ϧ�)�����?6@�d���bI��,��y�g����w�ۯI���������EKm8����+o��C�Pu+���C�HK�ྲྀ�>��T��8V��_�F��)�^��������
��P�5Yp
��Kxt����]��v~Fp"q�d)`7��^�5����ʒ�_3��r���-),�M��o��%��va�[t����4��A`�րѤ��9�	�-a|���5�.R:
������!�9��1���#���mpND�:A��t�_b{E������!����v�ͨ��V8�0a��S�#]�����*��]Obj-���!�{h�:PY[�t��H�Md%���[�f��堮��y�߉,Ք��b�Vb���\�6��`�]5�.��-��@*u�Cd��l0�j�w*�L���0��U/
�+��R�Y����×ฏ�S�1�h�m�8��,���f4���*R��n8Ӂ��s��L�z���jGMP03��f!�[	��������u{@>'�Y�Ι�-ڄ�ȧG�	�v�[2�=�5���E���)�l$!mb�[��.��->��tn�h��43U�i0�Ed�|K�/�U� ��F��7��ЙO��z�V��Sr�r1M�Xu�"dv]�ܱ��h<�\�l���R[!�ܚS�ψ>#]�&����[t���G�
��D�q��đSm��p���C�e��@=�������I	17�*�)4b����{�����\�$V�]�L���9��U�~�p.��7ĿT�2p>�I������'w��K��1=[�&e(s����D�gv��8����LP��}�H���������9{�$�V,����ݡ=�]�����.�r���y��m.�����t?��_�u������{{�p�ؖm�\h��X��D6&�� �`C����l�Wd�n�WV�)�S b��mn��]�2�y�
��#9@�9"��^?1�)���a"���S�ȥ(�綂+��@�Ƅ��vC���g|j�	���̓t�&�c��P>Y��Rk�+������+#5��B�cMnT�yI�i]��5�C��/z��Uq��XT�R;*��8��-�-9E߈��_�-3��DOG�������:�+����%X�_���D�A�R�\�G2Q5i�����p�о=5�4�_� ��61��ة�%�%�����-�r%y�h阍�O�ݫA�fޚ�˒���k���8,�77�u�\�)G�/�d��k8��<�_$1��Q�Y���żC*�8�H�#s�Pa�6�Zf���ġ���K��$\�?ϷW� 6WmK�k�d�yR��A�g��o�w�C�/�s�a��*��Elh��95?~�gw�1��$J�5��l������d$�(��a��U�~[-��Ec���c�Tp�~$눯:�(�O⿐~@�8��gr��D8$��pMe ,�
�,=���R�l{f%&g�����4�8�&�E��.WyRZ���D�̲������a�2N�����t��ȯ%�����z�ݸކ�T<�h-ˢ�-������f�����h������غ��吂VZ�]"��"�������N..��(����T�#
��_/w�@��f�O�*+�[A���E�|��_��<���B gA�!P�v����I-E�@��x�7%���؅S'�b��ܫ����gk�O|���F�D��k">A�;��?xo�f	'�'#�Ef� ,B��'���GaZ�o�E7�>�g�+L�sӃ�e�7�I��r"	.WQ9!����PH5�%]�P��r2C��y��ޏ�q��
T,�$s�;�*\3I�p���F\�b��H�qO���|=m�q	�z�僝e�`n^�Nc�$j��n�
��ڮ0r��T��9mo�&�V�j�$x�}���x	t�1�g>}kq�TvdpVRQ�m-ޮ�:��������y�K�GvP-`��HC2J�
���h�L�SW��Zb�Cv<
r߁���:6s�����ǧha����RGg!�!���W�/�>��;���A>������i褣һ�g�m{�����zk��2�#��k|v5�ol�J0o�L�:�J	�ŀ��d$M�N(�O+��t��4vRm����+������qim$�}�iFs�t*��qI�t�>��LUc�}wX6�m�p�0z�Q3��I�1��`f�D����a�Q��@?�}���_lk���CY/6���<�����B��Y���'� z�Yp�;�l|�E����v"���:��J�X
إB�}$mqX�=����C*�:�~
��.Dv� $+q�bح�������=�RHw|u	�'�"%26�s�+Q������j-�<�NSE�XS۳���H�Gng���ݷ�'��ˊ���X��zB�
"o�+���(�Ja�i	�)�z�Z<=G���餑�(Znݠ����YU�Y/|%���(��Ħ^ᒩ<b ��S��G�]1	�i�����B.@�8+5
����wY���A�B.�q�5���#�s��3A���[�
������?��_��M�m�u��+?�l����O�V��0���Tuw��np������NI�7�+� =Ã�b�3|�ݖ�ǐ�H�$�!8��FN�3%SVm,0?jp<5(��̙K��>@s��j������h�ܰ.�����ӅB�7<��PDT��<r���OY�{�1�i������q�[�㮯ۃ"�a��2���*�W"���\$w��%�[����M s���6n �F�J�q�z�R�ʷ� <�����,�IO��cJ�@#9w�N�6����|�|��0��KHk]��
kw�yw�X&�jN�R��~�.g}�A�������?������hp���4��Z�\�:]�r�Pm�E�a��)��l�a��$<\ƠG��m����#���|�B����)�.]Y��26�a����ϱ�g���o	:L�zڄ�拻0�<��Z� �"�aFڐ�X���6�!r{ɨ�,E-3�
�˶-RN�o���9��A�
LI&0D�i��]h��u�#�+8��j&��2�N������c���P�*l�m���e-ն111AkG�`ˆ1�:#v�����|��߳FS�y�j9}�+�3��M��&��o�ͲOx��/]Xv�g�,^Rb�3}�{`)�_r!��:xu����u���$��i���MA��e�	��4��+
t���?��k>��SU��n�=ھ��u�O i�Ჳ��AJU䥿�a�[O%,5��A����i��1��T�,������m��綟���&JѴ�we��h)/L������=4B,{TAQ�O�kFCdVd��K���]�[���9ڑ㣵Z���?����h3�3N��+E�\x��8�n%I�M�?���Dl44��1��B�����]݃���\� ��������+�MQ�81����AP�,%8'~�x����wM��V}W>�	lP�"�
�	ώ[���MPx�>��� ����U�����HkK`�aP�ނq���t�)��0���������y�0pQN@_9��l�(�( �c����a٫VYN�Ȟ��C�������̇ҋU;��2
�j���m�ȸf���Ɏ��i�D�ز@P����6?�L�qE���T�q�w6c���*?�s��^}��a[4��=,�$B���C��WJ�Zvʋ4g�F�,uozZYL��31+�<n{>�q�/���|�ebI�]E���h�@��J2t�M7�s�I��-�9���aƴ Ç��t�ﳩ3Ժ&�<΄�>�at@_@=`�#�.����G_�>������MM��!�wG3۬�9����2�+��?�r�^vZ6@���a�F5|J%l�g����J1E��3SZ��oƈ�U�弝��#Q��|�L,?Q4�d�tBQ$���j+��p��n��:��H�F)�ϭ��l"_yҭf[bL�AӘ�O�or��7Px�S�<*55���&����C�.��S�]�ԴM�K�<l³��^X'Ҕ�`�d�I��a-�l�ޏ/��a��l�%U?y�$aN�vx֒���ϳU0/��&qHv�n�j��^���5�>����F+X�S�&~��K�����)
F0��إ�
�5Y�~v?�jo��	��LZ6":���e2�O�i�Gl�r��NHѕ����7�4A͞��̛��2�]�
rw�+�dl
;���>Q�A(�[���i��5��i5����E?>�ꢉ�~9��D-WW������`ܝm�ݻ�>���C{��݌�y�+��W������F�_�@/I���"�����EZ0�B�d�X����Mш������K���i��쓖�L��h��i��f�3��U�ؕԞ��s9r</�� q}�Y[��5�\%	<�;�v�'V�T�����̽v��:D�b���tFe�c�Eh?�����8�����(\�7ؠSPsS����:j�/�c"
j����B|�@i�v?�M�P�]������n��Z�W2���j�wt���I�YZZ2f'�@�7몐Q5X��\5�҂�B&��{j
3r)���t6��^Z�/T^�:��cZ�l�G�!gy�W����[[7J4�'�S��A��������Z�\j	�3e��hx���cVz�G��R�����'�+�&��(ء��]Bۻ��^疇���(��crl��7Zۅ��_�8#bE��k:�bEHH;'*�6��8��Oڥ(P�L��8�C9RT�BJD ��&��-nT}e��Q/���g�vt�0I{= ,���pdo��7!�eG	�;5���{˿��9��s�	�f�-?#����t��r�̩��{���'I(QTj܅����߶����f۫�Z<�W������#��g�މ�����������H��%5m�ó�9�s�9��T�.����50��a,ޥ/"�ۥjl����9�@���5ZfE5Pb��q���0��3�߳��eGr����WC�����[�.lI�ee?�����0�y�ݰ�LW��8��q&�cB�~F����k5;������l����p��g��ɱc����:�2)�Lr�N�Ғ�����]�����,���O��a�W�KL���b�Cэ�8e���)�1;	')�6Uky�1΀MUӥ��\����(\�������bعS^�e��
�y�ߡVr��YƲ���q�2Y�m��3��I0a�A��:g�X�����~s?��S�W�_�����︓@�����2b!p��V��"���)47^��"Y �
}OY�f>�Q��Q�,���A�c1�c��
'��^�J�.,z �w�ާ�x3�z-丘����]�t�./;�/��.j��Xn�ё���s	/�W��:{���wH�Ѕ����mwH]����͘P��ϕ"~�-���Ow�����<�Og�W�o��X�4ѽ!��*�!e��ĳ�^?P�M|�N��������Nmy䋎�Y{J�7�9TIzXz(V���P�șф���U���'�$k��l,����*}�[���g"Ĭ���j��/9�{�#��tم�~��,�^�����wr�{��������o�7�	���1�wb%����B\��v�2
�0^��E��Q{�&���5*	����j/UR�� 3A�dPB�/z��u�h��%��9��!�2ס�
��GVW � Y��N�J��4K�w�Y���/Ep�f�W��;?���ȿ��`s|/��G�W]Hr����ѝ'���Ar�'mzh��}zJ������.���F)B��sD��ء�v�I�dU�ݪ��C�����|V"����깿�3V��f��o��h���/��SV��͹��^��}� �s��X��=Uh�Q��=V���F�6Vp����jr�-���0E�⺒��"��^ �>�d:wq>��������.Z�[ς;[-EǠ�o=�9��~P[E)s�}4�v�T�A~xL�](3U�q�oQ�9�鶏���x�0�2r��=�!'OK����B|��Q��ȵYO瑯�gΔ�-�^$ðnT�j����Ya�=9|/��d��_�K����������`Ff&uTf�iU2����'0zd�2h-+c�lM�wC��:�%�����KkT������>
�6��)+8��3w$�/�2?��U���eIP.m��}�,����7])$�8n!o�<�rK�XW��1*�"p�����A���QmV��������!�_�V$(NDaXAK��r�=Mqt]*�gb1d�3~�pU$���F�S.�"���XųO]xbH&E��[�� ���$���py���"ܫ�%tl�Z�1����?q|��#�2��E����x=��(iΝCfb� S)~w�lu��MV���s�>�B�����|���O|��<�)E_�*�M��+���L�kCS|�Z-�':/x
���nۛwG:h?�t�ZLΛ��r�(�1����֌7ӝ�N�(Y��y{��̫�c��©��[��뫰8�a�C!����?�%��B��q��P��۶��M{wM����˨N��n��7�L>.�6�:�
8�c��F����>E�kX8$�ŭ���/��i�o���'JL���#%�ri�����y
�����ihuϘڠٵ�,�UVD���=��Y�E�8�j����ֹ�_�s�q&SDu�-���&�z�(������T�A�ncbm��CuU��d⳧���>��I8��9cͬ�₂H0�8 ��K���b��Q�����Yq�f�k��$�D}r��B�l�i~[�=�Dי�JF��WUmw��߱<�3n�mG5��6A�tʤK>�g#��7yzQ
J�e��M)��8�Y�#�~z���@�<� 6��CU1w��7
�$^���"��5�ٜ3�|���G���q�
*Nz�N�"LD	^yn�	1�Vv��έďث���l1�j�p��aќ�>�o�
�\�صѕ�Y��f��u;��면��{]�q���lYR��1C?�j���Ӹ�=�c�Q�V4랛v,�-�}8�d�<eK�X�4�n<Q�-$�Y�Qh���������7+V��sn���m ��MQH�O���F[~4hK�{�t�C��n?~��m��1^ļ�1I��1��sW�A�/� ��1x%t{{�*އ�ݡ���V����Q�G�P�X�ђ�b<1n���J1���&���-1��?~s���{���O�cf(�+u$����l'v������*��U)��ާ*�G
���G��3�]2���O̥���{��Q`w4n��k�k����E*9T�[��к��R������%gz�9a���W
H�������|����t�]�|(`����5j� ���(�V.�b��B�D�X����W��XiK��<!t&�N����kk�m���eW��)b_v�iMM|�H;��Yc�k���cSS8�k�Aʣ�����M��B�S-ox�!\��C5ZޑpAf���ٵ�����As��k+�.�'��+)��"�Ս���-�4�U0d�4y��L?	��i��xY%��s��bPFV��x���s�1ypo��h+2@8o���D�y�?��R�?�h�z���yr(�K��<���t�@���(f�\,��#�c2�������`̯J�o��[�����>��Ixwn׸��
�;Eu����ƽ(�X�I&�L-S����X�bנp���{��F9��|�6sۉ�Ơ��
�ګ������)d<��m�P����V�����*҇�܋h����.q��3�s�Cv{�b�`���R_Vq�A�'v�1]b%�m�vd�)������ݫꕒ�y=oұ�h�����%�_���W!I���a���J��9\��3�Q�k�W��s2�K%�ȡ_U��JĄ���W�OO�#MJ��Z�TЄ��\3˘���e���Nq���_�<���������(n�Ȧ Q��B�
��亶�����Z�;�6��
x�����|+�&i<4���@���݋�1�~F1�C������#�
�)��HHL���ihR��I1��R"�k�(o���$�I��ڢ�̙!���ۚ�8�9�z�i��*��GI%���h�q�1�4���z�^jj&����=QLa
���,��!%�P�>"�ջᒓn���8��=Mg,Ͳ�I$jg�k�#iCZ��?�~�]Y�.�/��yG��}�I�G����>���l�=a�hJ�+G��Y"i)�l�V�������3���ʢ^6n���m)E�5���fse+^|[�?���&y&`n����x�����zC�VI�IE�x�҇�����2^�l������/}ǔ���_�e�o��E%��b�Y�
���TO΄蠈f�	NH�\9y��܇$�J��;w5+oM�z�|ȓ6�>y*����	8�ĉJ/t����^FO_O��+6ΰ�)��o440C��g��\ND�pWb� T6�:MU�6�^b�{��5�������3�F"`� 	"D$�$����G~��	��<%�P���n9��oE�9��������p��Z"l��1��#�8>��f�qAcK����U�`�b�b�I1�v�T� ��ו�o:��k���o�P�&zէ��T��uG�	�%>��%e�覘��7��^*b���?u�X��:Tb-ӊc�+��g�(M0� ��^��Q̲��!��$����˥�~�������p���&�6CZܓ$�i�'S";�ְ2���İK�7Ǖ�um��Q�w�|~��!�^@/�j���P'Z<Q�ߟP�R3�6[)�;�:�yt��ws�dމ�̲ S�w�%|g���[��Q�ٿ9<JK���sWpK�{�.��^��|��&��T+W*��\냾qG�5`Q`Q���I@0O��i�s;@.�OxK*�O�'�86�z�>�a�it���Ƌk\#��%���?�Ab��M��U<���?X�N��HB2:ZI��5�Bg�0'���A�c����v��]���O��T�
�gƴ#BG��m�5��]a��I�-:�.GO���ö'�Q����1n��͙:����9����]e���Hֺ���vT���f��FGʆ�3;H�9*���-c7���y���N�A�ka�9՚�3x�����D�oV���jE�K�&b��NY�s��=���OUMc��K�!��}��r2��BT&͇��Q\����v��'ܴ�����|�Aú�k���C�vvv:)�F��%k��n�|�Ai�!�J[�A Jrڴ�B#@!��C�@/�T3�R��HB���p]�{�������kବOar#tedj�K�{��M�������xL��YY��}b�ȵ�ܼc*>�r�������� �i����(n���zHf��kVF�
`3�|��x3�?D�W�g�./e�9��z���3�h�O��F>�+|��Sݪ��M[����5�3���]̀��v��a%�r�\��E͂���Y�(�g��i�B�0���.��4l}�h� я�����xz
d���rT�m�(�>�����M#U�ѱ��i���\�X�RF,��t֑������f���׳mܾ��w�9aff����7�0�ٹ&�TY�w,���8���--�3�N�4��JR)d�X�F������f���)��j���0�g�|$yk��e��U�mѪ��@H�>b�Ie�W��R~�R@OQ �4u6��#�W����=M��8�I���sr%���[OM�����0m�w�:�����g��u5W�\�J�����:�å{z��0���_�p�k�T[�	G�p�녷���Ɔ-+V�*Ga�o��]2{�e��1��2�ܔN��}suu���q�zu][i�*�)��+�g]��X�_vܣ���o�0�b෶���3}�9sA��Yi��?��T��>wO5�j���� ;�Y���}�[���	p�}y�E�ȵ�Օ��> ���Q)SJ�+�۔�ⴤ����R �`�|�o=0�%����9�,E��.�߰?�d��)��(���Grt7�QG��8�����R��o�����E=��emD���M�{���L-ط����Z,��l�� <RkZ��Ɉ��]Cܶ���p�'�\ۡY��y�9���q|�ڤq���[���\��RDu:��u��2Y�y���
�:�H��H�3��HR�ͤR!�W��2�Ψ�D͕f�d
�7���^����I����d�K%�UI��R�񈕕Ih4�"F}Zi�%�/��=2ӑ"���h��C6���R-��/�V����X���t� Pm����#|yQ0���C-Y~.U��!,�f���q��r��˪�(�v*h��R��J�`��,�hp�h�X���f&�_u��կЊ��eE�P�|@�ui(7��`g4;-���b�����uA{^`���J��pc�ܡ�8!e�(]F�.��J�hi�/��@����	��֋""mdi�����|s�����")�"\�[����]41&�[pb"�L��'N�rѽ�r>Vm1���W@P��s(D�8ED�*�`t����k�*���H��ElwT�Ŀ�߄:c�R�8��2��GP:T;�������b������ %�� �@��e&�+6�6.R攐�-�JG��@�ܴȥ�pO���+�����NR�c�0��S�,Z;;�m���q�3��
��e t��|�����-]�:9A��z�������_We��֯�����R�^;mD�@o�n�t8Wy-��� �l/I�)��Q��.����7zZ�u�'�/uy�'޲d�l��η��ZVې�K����5��2|��y�u�"�9�q�	�>�l4��]H�"�Z���C�ʫ8�x����o'3������V����B�%�A�2Ú��RĦ~m�Y��N���5�����I>MmۏTp0Y[�9���爊 �a(�5�Ղ_������4�����ʕ���šHGT����"��I�X�>\�z:�v���đU�Y�%�_3~!2Kr�@w=A������i�V������X.uqi��XT�k��0:1�V��1��"g��LFbqpu�G�����?l�,����\ʏ��-s����NJ�ʹ�����t.���a|��S���.�����\����ެw��u���^k����4ѳX��P��g3�ESt9)�����f4).I ����$�K"+��K]"��W�%��Ve�Sڣ3���fn�ԛ�[VuEN���`�s�������3�øs{:������!��H����ju�M�[��8}@%��	���C~��3`����i���Z:y����>��l����r�,m�,9��+*�?}fR�	4:���o��Pm����`go/P+�ZO]��u�#ӣ�v���^�%�m�`I,��u#K���������f+�Y�C�e��5��[d�*H�ZY���b�v�ȧI��6��:K�<+RP�#l�'�ro�L��_�s�ޅ�������V�y��s�e[��G٥]l.	��F��� �YV�l��*�HL��ԁp8>�b�sm�S�y�� qUMM��Hj�����*�9{n"_��gw0��8����/;� ���I��m�Vp�X��Ń�|T|�Y
�������-���OI�����~ooS���H�qDP���!����Ե����MZK�R���133�%�@�>bqm��&�I􍙭��	|�$� m-��`��U����-ˀIW]m"����\���f���Nd�a�msc��k��7J^�2�S�������F9�$Z��%�Q�@�����7���6��*��1ɺdʱ��y�*�b���������Ԋ:��Tc��>���L��E�'n�H߶��{e��~��Ltd@�3�n����{��t����@E��>c�
!���y���G���Ҩ�����_�v��|1X����)J5�����[�����ˉ��d�䐀�����G�?ߺIv��`�a�y]��:���+�\9<P�s�4�b�\4Wa�pڞhֺVSjґ)��1��츨�ƕ//Zъ���� 2��M��3��J��4����>`4WL(��!��Q�#��?��@A�VKK���;���ZM�a#j�D����d������5�7��~ߺ]��U��c�L���&�8g.������ѲT��)��ɽE�r.�-��{�N�Ã'/��S��7D�}ϼ�Ѕ��e�s>� �������:�<��	�{&4����e͍����������1��S��]䑑�����U����w[э�Sw�wFbǎ���щ���?;��gۧ�g{Ct��ޝ����ޣ�nͷ�[W�I�ݢ�5�s<�S�����4��Vk�<_7R�@��qOA�cL�K���N	�2]-� �E9)���cP7��o������ub����v���(��0��	���M��pQڠȅ+��;l��v�bY����U�uD��l�*��ug�S�ϣ=f�80ㆿ�+�1�����Rh���W+fwc��] e�UO^�3F��D�Q3j�HW=澩?|�-���I����W�KL?ȇ��\����wkKHz�;`�Fm_�puMv�~Z�y{�@���>�r|�s��L@z��v8�U�������)�g]�_I=�W��[[[{��tA��a�χ���<�O�I���3�v�Ž��k����G�����8���u�Y�h�����{�����!<rzK�0��r�q5���wg�r3�����������ӎ'�[77�-��L=/ �˹������S��j}W�U����:��{`����/��x��@-�LI�l�T�&ٔb�L��SԾ8ex�4qƊ�5���Xƍs���Ȱ��޳���)n-_�+M�`�Z�⨹���{��N��y��y�j�K����W�`+�:2 �C�4eį��OP��^�����/�)j[~��̣�B�~,�K���V��́��2c��MB�q��}Q�W8n"���5��U�ۺ؋w����!��_��o���?N�ݯ��oW�\�.es6�h�]2�mYR�-��H�qb?�j��\����u?(8��4`߼;2�i�l��ޭ���t\��r��*��w6��i���	_ �z_�%u�?_	=�Kz��y�f��z�E�;���/�o�o�s5���}ӗ�LLL��W>g�;/g�"�"���lf1﹁o�S�o��	�w��!t���q=-�slJ�c�vcX�Y��������(!SYY	9P��KKO�����o� ���������e��>����Xq����s뻟����i���0 zzG�	_�|V�&���6m����~<N��x���&2��.o�rg�[�hs;!�}���m�]� 8�~-�2�q���k�xa��H�F�t>�|mHSx%�<�*�ࠋ<�w��u�#C������ݪ6~�������*s�_��c)Jm���C�z�n);m�����=�0�-�g����,��~ݽ�K���.�aQgC�mMG�Ү9�㺙�u�f��@4q�ۋH��e����;/��d�_]�R��;M�[��|��S ���W������O���힬����y�x�>��4����=��i6�����o��;���}5��_I�꾊�?�Z>�������'�	ݓ��p��[��>k���|lY7��������=|ErD��n$�K�ԑ�Ә��QH2�ɟ���Y��	j7D<��N�Bǻ���7��#��$L��O��~IYu�?hs�@+?�I4��4���$*	A��k���t��L/��P G�ɉ��~�k1_��軣(�9C�bo�2W�A��U��2RF3J"���s�}�1K粆�s���߻k]m��	��R��j`���'�~]�T�J	ǧ���ˉ*`�T��.$.���l�0�^��2�|N�^����^�����	��.����B��Umg�B����G�����g!%��5�T��������Y5��|t_ ̈́�3H����3ܻ�=������� 8����}�T���ԹQ8sP[_����n*������v�*���!G*i:=:�a��Ќ��\� nO4�����:��\�
���,Ξw�Z�.Tt0�7�{Z�=��G��u��;�c�����O�B4�o� 4�^�a๋��e���y���un;�ZZ5�hc�s�9{����=��I>�v���ܝ�1b��CcG�ؑԚ���h��$��{���H��х��}�r�t�����:����=�&����T֋��c;G��m&�F��?l����Mt�]�hl��v�M���pg(t�V>�nܣ�v�����hS�u]s�H�^�}�6<��v���{��t�?	6y%J�7�D��>:���7CÇ��w�`cusg۟�\���F5kź����5o�*8���k�3d>i�]��c
�Ն�S�����wK��׉�!G�Sg�v�h��D�1ND�5��Ll��h�����g�=�?7�8o�P�����l`밐����s�HE�÷w�w�	�e�sK��hU�(�����Q�`��3u�fݲ��I9�i�~���d؃��[;��!�ÿ5��o81e$|���_ ]���H�6�;Ʒ�n���w���� 
�kcc$�ڻ ��6�#<Sꤜ��M'�s|7�xO^Ƿ[W�L��4*.-��E>�6�Vl_1�?A {؟0�٭L���d[-Ísd۽X�40�N�41j�r���7�O4�vS�>�-.���S�~[����4m��n\���s��G�}���u$[��&���~�@z��Q�7��r�o�;��.�[5Y ;A�>�����ng�@��st9���LQ(�||����)c,�>k����8��F�U�E�F�����Q���K�AU&ӭ{;0�ctl���]o?�7Sa��d� C�I���ۻ=���FG�/�:OӢ��3�����_|�R���ZFҹ,��t^>�&P��1F-�);�O��X%NgY_\�l}b�'�ǚ�p���:M��n����}��'{[x�Ҥ"��_оP<_�R��p�eh��S�jZ�Oc=�9�.�b��՝9Kg��f���h�R�w���{��O<���)S�� :�J�B#O���f4��?9�Wd�K�X�����^:�xQI��r��֦��y��=�e��e �7ƨ8�"�)�m,�d��/iQ/5���n
1p?dD���>����O-�}�B�J�:9���)�Et]"����� Z��$�d��1��.���ܪiř#��@���L)���� ���#��d���!X\_7���U�#�Dq���ײ������5Z��1я�ɵ��3���mm���X���_9 @���}n��3�~?+T#��p�md�>���� u2�OA�m��5;��+хO�<��E��⮽�"*40C�x��2!-x0��Y�}[#t�{�Vi��� �Iu�ݽ�<Ê,�t������EB�x��{`����%dH��\*�>���YU��[j��pm��=�N���,�W�4;��Lv]�?]�wSA��igqQ�2�t�I_OP����W�(!�%�����+�i�Z��#e�0���%�p4.��!��%�"�����]��:���X�f�=\�̛��h���{�M��W��sל�D
`�����Cbׯ�gЌ�W4%� 0	�MQ�qnr(sk�[}<N[z�v,�f\�������Jf�*"�׉���ޔA} �!\��^��9_7�K5=M��-��\�w���B��a��!11��>-G����@������M>HI�5�3*�� ~o��B�H(pa^���q9�íb��TVT����hJH�?��2(����n�Kp��%��www�����Np������W�?��t��K�W�)V�����yq��&Q7��b� Cm��A쫹v��2�Rs�kU�c��W+و�~n����A
�	���.�k�o���j���*�`a�e fw�A��q�hhP��0N�m�?jo=��L�ݑx]�IE�1�)U���ڐ,6��I�r���S�i`��4���柞B�DL��ؿ�JZƗ;v}}=S�S3UP+��W�M:�=����DJ|�PJ��4�K�M�qr��Tu��;��$l<��$�oPb��i�����|��S��u6.	��H���XK�M�$�~8���(Rq�ڠ;�{����9K -�b/�V<
HMMGW7�a�e�yu��J���5�a�G55��!�6�2T8�ճ�
2i�mv���?�ۚ��i�u�aw�
���B�c�l�}74+����[�b_�lEnQ�������<K�a�Z
	n-� �Z�Ml�h���{v��x=� :�sW�%�&wb���F�����LU4�_�+Ϊ����r��N��o�'?3����#��W�c\�Bݞ�P����x;��v%�M/~[���$Q
`����cMA��r"jˁe1@'B�8�l��,����2_HorƱqB=��iV�zN�6��ˇ	���d�������Ȝ��T�X��Ԧ�)��̉�&2��A���cT��_8R��� ���I�'�UU��E��c�(��{b��B?Å����yz�����vvlU�C�Х�ۋP"���#,�0���DB
H@K��>x:�T!��ǤK٫o�����{#?�߇_>�`�J*��pe���G�
��p0bzX@d}@��Z(�%g��	��d��3�A�{��T(��J���_�.�K_U~�r���y�	�qv�xЕ�֍�/��"�Vo8��>.o^cQ��,�ni_��T!��Fú�A�찑ҁF�}��cF��y%A*�q��2������(d���3҈R��H�c���x��z��ch
U՘��>�:��_0��,#���x����tR�3}��`�J����ΊEwS���\X� ��h97�<�u��V�!���Ab��Cu��T��a5�����+x�{!���Ԫd P�����Ϊ���E�A�6�ER��a�H���Z���r�"��?�}�j�>���6�Y�i��).�1J�5����e_D��$R)(L�&X�mo'�	�)zL��O��i3����
��r�� |�C�Q"H��>p�nDgc*3��3�g/���,�9�r h��6?e��ڈ~'Q$=��^�L�C�Z0��@�#��=�u��C�Ze�)@#E���9��뀈�Ė>J�L���U��� �\�)� �n�a%�d���*�~6��MX)z����-�!���a��U�io��>(��^$0�i�����^�o+��v���4ݼ�6��	O
�<�Όr�B$��KG1]�i�u�]K�R�V���d��P�$�_D�����]�@ƆGŖ�K���ff��t���r�O30�][���0�_n����i�>rR>?�P ��rk�º�"��Q�n��N���K���H�p�a/�eh%���)!���#�4�ap%H0�{�ctp-2B�����l9��r��L�Gb];�!����eY�n?;������,�A��W̩�@U��kJ� �LWCy�*kS.8i�ng�1d�g28GE�S�������2�&�O�k���7��':�\y�Q�z�H�_!u�[�т�g����g*����c��q������@vøRW��w|��[^�3���8&�,,��K�i�&�7������E=�LZ<�?z�H��%>V��9�S9��S�|�pW���خE6����JNvu䓳̻5(����o�(\4�Č��H4�8"����<R0�jc�=�����t,���z�����)��9���iC��fվA�xi�ML265�K��G7�>��i�f�'�������7�|�BN��PE�����ʊ�1��L��+�Lm�K�i����]��|̓��l�nM����Ru�fNH�/pd��Hsߌz��1Ĉ��d�%o5��A��4�ˊn)�K�(/�����K�b�>N�7sR#Ir���o��\l�V�N��}4�ph���?ɑu����y�V��a�jzq�Z��S�HxP�ȡ���kQ�\)i@�+I�·8��}�=���>�5F�^�9j��˕˞�N	>:��x��Z�boY�~��C$dT`h�#�t׺��"r��o}��Ӎg����<�(7�����{�a�,�5�N��2us;:��enǴLsy�G����|w�T���Hq�M���5[�-|�k	<2��G��U�Y���k���w��AƣZ�<D�nA�u����c�rRk5���K̓�F��
�zu]��6�|��2|t��<�1&h�TH � ���� =�9�L^4���-|!F����4w<1�{����Bp���!'&`J����gӼޓ�/㦏���K�� �.9�@��*���9��q}�vٍ�����ł�׽z�Ͷ�7��cz��.�H,r<Õ-�7j�-Ny��;�b�v���n��J��nh�PM��pJ����OUd� ��ɽ/���L�n����r�n3���+�W��P�s+�V�J���L�"~SR|X������L&*�9���c��C8AZ?�.B��ԭ���z�NWn+~�l~~��c��8�*�Q�Hڒ��2��zIqrJ�Q�zC����z��2�PY��ٵagP4�|Oz����"!�?%n���/z�ۂx;sF�6ѐ���\l6r<H���"�����%�_
TƸ�y�%�Ӡ�K�!K�����Cy�ʨ�b��2�ˡ[tT��k\���E���~�?[�grU"LrM���A��J
��U罾��]G�c,�\��T�}�I�'�V�0"��gFp~�'
ݦ����vK�ֳ���Ͼ������Φ�P�}I{쥀��v?f��|�uH��b}�&��#$�>����`].�Do壩)�K�R� �Ӏ�y�{C��6i��� ��0���{O���Z�aM���L�)��@��f�]����TM���C�c�b<(ž$��!y���&�EO����NL$d(ؠ.�86�EG��T Fʂ_�gI֭3:/#��z����i��0�ב�b�k�.}��p�����zg������E���OOW�VW��c������&x��u+ˀ�����}_���#��]ߔBzN<�U�u��Hi���#X]�٤�h�<�绺Z�8	~ػ�V�Ⱦ:`�<�Q��#��n a��卩p�wi sX��ټ�K����a���o�%c�/srS��#`�[�o��r���Eҋ==sv>���1J��Ds��#>���m������a���e.{'A��i�&u���ff7�A�x�w�ܾnZ������d=,�^[և_�e����ipAw�'v��ټ��ד�)a��i�xqV\�EJ���P���H�I��#7k-�CT����9�o�4xq��_V��C��]}�C��G�` ��hX��&# %�r<oʓ�P�4�����B�b��=����	�l��//�h�ULI"�x�gs�W~k�0��=5�-R���uN����wUk��^t�u,��BҏfǷ~�A�/�KDM���Mj}��r���*i�B�ͺ�Aq�4s�D�6R����-��Bz���N�6�u�V4�4���)�I�J�B>���3�B���0U���S�MA�9vs_	�]����2��"0��k����%e�?.�S)�E'z��.�H�;5멞^4�@9�v��OQO+��$��aS7���E=���^�`�):��F���}��L"`V}��O� �7�٭���뀺(��2]���~7w�b���i4�����ͪ�����;d��G<�p��O��iǎ�O�ݵ���|���giU8�����<zڭ3�ύ�=|�M�]��<
1�	�Dy�WML��Z3O�夨��/����w�:�-j�6�&l�j�d�+�����7�
)
X��C^2{h���x�D�ܔ����3�#���p��e�g�S�R�S�A0�K7Tӟ��]���ۢ "�0ctKp��q��exͮ��z1��L2�z�ݐu�aF!��]����ګ���eMR��d%��n�����B����~Ӎ���B��N�.��Dc+
�	���'��6H9�\�&�/�@�C.m�%^N;k�>dQ��~���U��srr2a�?=;�I��D�寞Cin��QD*�%�5a[`�/SA`�Q�ͦ��7���lB`�AԱJ��B�����oQ�G�@e�{8��?@L�s��3p[_���#��#�˅��lj!��M'�$�(oX���.����f������)xZ�@���WaJ�c�g���|'��P��j���#�+L3:q����U�V�B�B(y.�������B�/��bu��rE}G4v� �������q�R�GS'��sfj�@������G��誮;h/�K�h����$����O�@�2�(䡝s{���fe�w�����k�hpR��=�S���y4"R�X
� m�i���4��TQh��R�9R�G�������9�E��0uE�r��ͱ%s��,*�|�u|}��c+x��[�W�� 3��t���>���[����v������0�E5|��������}�sAKS�-b"�W����Y�_P����?pqyY��=-2���Ӥa���ٻ�{�)�jI<o}�eu6ge�.�?��>#lI��N��ɸ�o���a�fHB��_�P��vww���B��=gv+6.	_ ��-�A��G�����S{�y�\��`G�Uϖ���4;%0�$ns|�v��m����3��X��=���y��ƍ���~�b�8��(1_�q^��J�`e='���#��²���ŷ:(�`��'�r��Q�Jq �
���2Q��G�<��#.61��}H�:��$zDd
?q6L�p�ݦ��y&��t�3���fgA���x.F���+��]��h�Z;_[S����ɵ��Δ9�n��n��F��)��C�&���@O���yh��������4��ӞnQ�Nܚyx�5���+(Dppp����7���U���#�{z������wN� u�̧l���-�����oJD:�U�K
��GUd]�9���4�f��(n%k.���!�{��y����,-e�ώ�q��+�7W(�����_pW�5e/h�㈃K�G�t�7�S1�Z�^yWVVꛚ �-"�����p��"�*P����h��?z�����'j�8eC�;b����Q ��J��|����̜}����U�>���YY�eݡ=7Wvzz�����,V����d�$]6�q����[��J��Y i��z������G@�#���I�hrg�=^QG���
B-��zJ��kjq.uI6�W�.Ob��� t���(*�SbѪ��v�����ʪu0�l�(niii��w��������~[��'�>宎�%��S�}^kU?=[�o@�l�X������h��O\��n`F(�glJI�T�H����{Y�~;�|
��o�Q���uҝ�<�<���g^��ӊAq�� ��.��6� MC��J�Z�p�4���&猌���V�X�Ҁ�d��ĉ��Ή�e����IFL����ڸ���/���Op^U��11�����˨�[�H}���A�W 閮���};A���V���m��}?�2[�H\ �_�뛟���ȉ��C���#�O������8xM��Μ£f����j���q��hz�q��%i1��1�|f�QM���r"����R1�x�
������*�V����]����_d������KaK�ZZ�2��?ݞXTX�W-4�V�����r�*F�`K�dUc����u#�v\7mL�^��i�����ed�{N}�nl�)r<9E�td6� ��#�Ȃ�`�Qy}��A�ݻ}�yVVV����Xc��m;�de�+)��66֐>P�mR��:�����W�hnN\�W��(�߮E��b��@/�Ѷ�.h�N�!��f�����i(I�[��V���=��-���Ĵ�8(7��4���k|�6�K~�k�P�7�7�$����j����j@�������ڲd1:>UK���j%���{��7v���|�����+�C��&�.����"s�M���z�����hΤ����Ҿ��p��w~9�z�ŝ�8�#yc����������D�|�m�����@䦚v� ��R�XqryxK��|UKy%}[WC�ls�DC5��C�ʿ�׾s΀��gw�8�V���H>��'�S�z�����m�{a�6���M��8�h�t���mA�`�&�H]'	l>;����0z1U�V�����D0���%	����G����ok��!Љ;���OO���pT�´FFF�`C��0߲/�]�c��w��z��;O?N�~ȦdR���$���m~0�)��_�Rgn��o�D�f�V��_�TӅ����#c���	�9xK��L�qZ���?��	<#��������B$
�$JJN/��lY��3�*U�fO��V��D���|ʐ9H�� 欽�4P��a�wW�y�c�4a�9>���~�C)�T��ג�N���Ykkͼ�������g\T��f8����i���2h�t��oφ�ρ.m�Y[��Cr��DF�3�4����������j�G����h�����{�2��@���ނƀ��;b�U�����l2��&��p��g��R�����?l�ӻup����Q5��9�2���즥|�'��c��p�T2��l^�@O�¤���#�	��C�"��t�:�c]uu��4ҭ[�Y��O�ϳϔ߿&�6��=p�J�� �*0;%�rY
����8ԑ����FU�8����5M��#d�b9�h�<V6y��)��������N��U��޽�$��K�^�		���ʰk�4f�"11�ɔ1?�B��)/����q!䫖ն�G����s����׍��D�B��M�+�u ����!�Vy♳ �R����Jb�0�����&%����Ώ.r�&��$��֭o,;fz\3��L{���2
ď��L	����b��)'�'?�\2u`��ЦU�mU����]=�,����G*>�A��������Q�!�JK���69�9����������`#U����AA��b��^���W}�y�U(����,����%���&86A�c��ƪj����\�B��iŪQ�m �a)@'�@٠�]58�F��y#�	�P,b�+�qm�Y���F��>�oҲ����@�Yvm�f(�Dg��,��e-w�|��VJ�Z��텪z�$�����3��k,X����B���ؔ��%�!;��lY��W���1���� ==��f*�!��)�g���8����H.�C�^�S�A��S��sC�L0h��f�Y�4�C7��*�]�@|8�'��a:.f�������j��5͐E郧t�6�j2�%����H��ϰ�Z�:����H|p��hz$H���xl�����wq�W���JR�삃�?r��c�!�;?� P�@H��qZ���z8&��z�ᱺ�X�/����aln��u��^N0�^����y�|��5���6i�������މ;�΃o��Z�}1VM��o�C���&n7��ΏBnM+kV�Do\�r���&��]�1���ڈ�������R��m_f`g��UKz�K��|����y]�}����e��3k+Z���:'�#�4ҫn�R_�}�4ӭsf�	��4���Ϛ6��ަv.{&��Ih������G���:�EM5^����M�	�����z��W�o��|؉�9�/�yU��ֱ����l ���e�&>M᭯w+���ۃy�6ʖS�Wh�?�KN4Mz�C�<����~�#�ʃ�3��U��ʿ}3;�!��|/M��]�����iu��)Nt����=�ץ�����E�%t�>���z�0:N������'��o���p��ү���W��8������:2u?�`��m��?�:�"�p�[*�~�\BGW�:6��S���e2�q�����/(���� �.G��r� ��
���L:�s���ن��+^\��_5Dw>._5̸Q�DU�ٱ[�Bd�����n�������w֊Gx$PPX�/��o����r�|��~-�Hʧ���������>#n��L��`���`	�*���e�<�M4>.;��P�)jڹsf
%�k֒��C�����h���.�Q�#�%ԣZڣqM9���#T�ǵa .b0�r�/Z�e%HCc�x��������{�
[0ӎ�V��n.�~�U�2H)vlӲZU�9w?L��lK�q����7�p�9�+�g	b3��)`��Z����Ǖ�uC}}�#+�XJں�q亸��o���S�XV��=	�A�;�|$d��F�{��^���~g�X���2�3+����bH�����q{��z�	�P10����9�p�"=�[�.�|�_2��FmKヺ����]jb��5�a���u��F����Ť��� LY*���n��Z5�qN�s
>��7[���q6��Q0�N�ĸ<���f��|ΐ�nh���@�L��ѡ�健����J�UK!N#�]�������rf�b٤е�H{na�PŇ�z֡ոД��Q�ߒ�10 � J�^+�M��"��3�/��vN�vE�e�YX����� ��J��7^�$�3�I�OEC�����Ҹ�9#�2]��r&<�B��YJ4;=�j�hS~�鸺�&^g�4(���D+z}��xG�>a���.���,R��>;�0Ce�A��r�r�j��1X.Lts��7٣���hI��I��/z��su�����:�BHث���wh�'�>�酡OWj��&��w/������p@�u�����=s:��1��pCY��0ut#��i�/p�5o�W�f[�¥�Ӊ�C�Mwbcn��/̟�
%�W��~���zE��[^���K��l�ֿ�5� ��58�b�4�ڪ9p�� ����`�
P~��GA��� �!���(��+���F � C���P�Y@���FbO�lw��0����m����3?~���+��mG�2����n�h��;O�Hl]��O*"Ӌ�	H���##x���	�Ygg�Ɵ�C��3s���R�/>���2��#c�"ɐ��������VD,��o�O+�/*wP��Wӧ;� ��L[�����r�C���d����,D��F �mn��*�[��㣢���e��Y�D�YAL=�0��b�;�eܲ�[��zAl_����[[7��\�ł'�"���Ơ;�y��5�Y�1KK .Z�g�ā�J���P ��ÑUp78O�M�W�����.�$��R"���gg��M��`��q1	u���i\-n�t�/['�A+B� 'ggx3c�f���q���ꕏ�yk�H}��m~&G�g߫��|�U�cv|T���-�Om�5N4|�y��+�"{Rw���ʊ��Mq������P��B��l���I4��Ý�X�u���K��އ���2�o��|6��2�L�ih�[YE�����N&�~�����\gsrqI�;�u��рi�:-�ooaˬ�:�º�s�s�E*|ߕ{r1�\r������9� &�	�!,N�N�5J�e�C����}������8 s�F�`��|{d�kiq5m�PWח�8��n�o�SJ*�A�W��"G=���4 :��g���� C!��B�hu,B�1�"��YXay�����+g�\��06a�c����4���u�w�o�---�C���0f��]U�"���d��/����A>�Ѩw�y�������x�l��zE��Rл�GV�UZ�����Tp��< �&�X�����/��Y�+'X�*l��ک�<�։��U��)����X5��˥���$&%�"***r����*``���*��c��f�> ��;��j#B/�qΑU$�_���1�����֯�\�q<�9
&9�|L��g��3�r=:�-�'K�J��㔄���?ُ���0-i�F[b�esp�����3r��n��3�\H%�Cd��uP�(��N)`��kL�ē��S�J��vt��W�7� ��3U�љd`�@E�Ka��S�4�|�)�������&���9SN�C
�@�9f
�V��b.��	�W#�)�r{EB�5�X��q�oY1P�"�I��n@�s[��߽-����v��^#W=��ex�u���A��b�9U"�en~��z·B� ��e �k7��5���q����^��݁�]6_mL�[c�����Ѐ|�ԣ;�Ó<m�nc�v������*z��R���YK��c՟?�.XG�T&�y>n$͙%}�	|߰��$�Iٗ�L�\c���[��f���_a�1)�;;�R����)C��r�t[�g6�"��������_�NbI�G6��f����,P̙9b�Q*�Y�T�ߣ���v�9�ѥ����]���D�lL-����\=�F��_�`àK�Y<26:g;�u�����`���5��H��
GmP�P�P�Ymעe3>-C��a�}փy�p�;@��i*+����јUӉ#¡oyEEMc�~��녔_�Lĥ�9?�On�$\����^U�Z?$���T<�<��q%1�(��n�CZ1^Q9�Rq�ݘ��S�o�l /�]v	�.�+bY��j�̾���sδ�-��z����<Ҕ�?|�9r�H���'�ݜp����3/�3�����R^v��cyE��W�����y�H�@]>0�^�h���c>֐vΌ;Z��J�^u�0��%y��&�/�e�/Z�U�����T�`xt~��Z�̕��n�W�۶�qyH8�ǅi�]]��0��~����%_9sB��� �Z�*���S�f�1j�����˹L��o�: _��
z��83��}�Fн�A\�
��%c�aht~�t� ��+�R�%[l'gE	��Z�z(N���BuhjҀ�<�"0����)@Z�u$f�B����X�B� �h);�%-�ƺ0��a��v��]�r�"-/�#/ 	u�%�� �ݕ�H�X�ї���jOS�n�f782Ji%���#񳢕
�����c��;e�.�IH.�ӻ�Ÿ�h%}��D�u�N���w#�R��rrqLl�i,3�lT��FD?
?a�)��>*A+�F���F�QN|f]��pU�xurڰ~�5���`�F���}��F8�����>$""�k��B����N�.����I�,V��wjۉ�:�nn���~����}��,�ଇ�,]5.��_/�����5;�`u1r�Z�02��\�}����O�l>Ŕ���?m�=&�U:��J��tP��`�X�C�Ĭ�dxY2>w���Kf��������U�ژ�9�۪��5	ز)��O#.mb�/@��>�q}��'�q'K�h���a �E�����Qx�+x�h�)�j�eL�QǑ�=��eײ�2���-��X�EǢZ��؎���`+�(^8qk�*�='~�#��0�#����nj
����z�$�����>����F6�ߢ�錨�{��F!���!U	�Zq�8=\��#ɓ]���b)|�O@,��f������k~��6���աY{s�Y�v�An<��欜�ɪp(��&���a(e���l� ��S��'���J#a:zƚ.�A�O5R�o�U��7�R��u-FT�tc�E�XR ���"�a�D�g��<�J�Ǝ������	R�q1Z.��b�BcqmM; �WmIp0�5x��5��β��z��v��8w=ky�
����O��M��V������#�)%��h���ORW�����J���
��O)�cFB+�qKm>찀��I�هEWMsAt�P"qO|�N�`Y���5���Z�*U�`�����i �S��P� ��[�Ǐ���өZ#���w6㔜o��G�+�j�U��6e"m(����+��F���Jq�I̯tjKC}~|]~�ܺ���&띁���4.kr E�@�f�˧�{�/[�}.~BuĨ�=��}}r|y���q��ɾ�����fag(�෈��,^�i��'s̔���ܭ���H�����T(�mbb"3!�����f���G
�� E������߆%Y����ϮRmɰA�4����Q0�sb2����~������z�z~˧�c�iI��a�9���{���Yq�+�_*;:��dҁhr�p��g��.{	?7�Ѧ��篈q�RNut|���f��>��>�؅����%3�!K�)H��Ϭ�tt�J+37�cn~�d��ʩ��J��V�LI��$"���!�G{�odT� -&�y���|�4���.���EW�D��AazM ��cRH���%:�%+C��ȼ�#��ճ��o4���J<�N����VI�x�ܙ�[�se	�ΖZz�f�zN/�>��8����r�O��G�{LPZC4h�=���@��/\V"�#�g��U�r�գ}��c"���?�xg���h"xI�t���ލ|�%	�A�C��k���{p3�r��a]e��1`mVˀ�K[U�~���W��+��&�$ZQ��ؕ�Љ�(B⋲�d�`�|�<+$j�fk-�ҙ es��Jৈ��H���1�!��A\���������Q5uu�$o��GEY�<j��5$�%E��WǼ��q���3��+«+��_��"���%}�8�_�Bw�U4�?��]�E��	�����sN��~��oai���M��Ƿ	�2K5ad�^��[2�Q,���#1pV{��Oke�c��,Bмv��<WD�2�3Q�:_m��-8�����CcX�P	;�&�+�ǚI
8�Ê��HTcR�E�<0�a��b,G����? �_X�\�x����?;��O��:����[����h(��rx�������0����jZZOǩ�WF���X��hV-���]m�4a6g��JY����O�Ǒ8�=���do�ڃM���OJY��w�j���)аVU�r�8��.��׫�֍(R�J@i�>뷳�����t]�պ��e_�)n�#��������b������O�O��!����"[�<w��u���E�M���'<"�M�p i�B�w�>�+5,Z��\@`�UUPu�Õ��ˬ-w�l�]�E@������Ac!Λ9"Em�/�tC?���E׻@.i�Z[��ύ74�>b!
�&������� \�S�V@���㑕p�/����~T�O���P��&���)���(��G@2�"L�P��rfQ�(�2�ǆ0��h)�~�?��SG1��`��nn������q�o�U;�7�<=��#��QPQV��3:#�����ߧ��{�#�4���$��`|���K��A�!Ń����f�-�� ÐX�%�}���\U��-ǋ�������Ut����\�����U�,�����3�E�f��h�.��V����	e?zk(��^�SQ���
�"���]�DnۣiJ���ˌ�'�K����xWΌ
�}%l��s�{3�+��˥��ㄸ)�?im���4����,zja	)�]67e�� -��Y>C2��Y�X;� ���j{����� ������˩��'�>P(�~~Xhd�1$��?��(��e��uu�e%�`�t �qx��E�ᓵt���� (�K��Zʧ䳋��@\
a者�f�(᫑ʓVn�7�R���!(���*��*�����S&��l>Ex�,-<�[���i<��{�D{�����*m�M�&s�y��"��`��4*'֍�<`�Jӥ���L�jPS�~�sH��:&|n���$���v-�;�vw�����*��j�k#�:�2e���@1(�0�(Ʈ��>�9�º=��L�>����p�+Pjc��C�#9�R��Wp(�t�!��θ�Ȗ�r�#�<�C(���i��V����ĭ�G@3O�ų�����1�ԣ���f�#��8�ޕ��M�nM�G�L�# E�����%4ǣ$2�	��Dӻ]�'H����d��x�\*���J��ib�_����d���|!�	��35J�{?:p�������i������ΤW���G�tQ�G�'l�0\�"6��'݂����b�����������"�I�S���i"�x0ƓL�r�X�hvx�3��ㆪc��0n�V�q2S�),1�FL��c%�q�ǻ��:Hon���o�����	���sk<7_�K���z��ݙ:�
���6��#X���yE�l����X�K�$�����zE���ɢ�"��w[mtF�9��0����O��X��z��rЋRA@ŏ�Be�4�9�_�V p���sI��b��dP��T�F��S@�=Bo��<�RS-�h>�]��qo��P*�Z|��	ų�gt(<���yVo\�.� z��u_��2P����;
�� .+������m���q�1�/���d%��1�m�3Ӌ�OB>eg�����Pn����@C0S�jb1+�*�<1���Z�r�?K���aF1�����l����'`Q�6=[�eH��Eχ��ؑ��m���{�j��q�KD����F!��(K���2������W���M �O[�ݝ ,���H�� r��'�m�Xȶ�o�ZH�?"f���$��n�Ϳ���"E��ф@��D
�l�+���f���-��k��,�j
os�Y�1������x�93�(l�O����T�}2Xy[�BɅ��Ц�=�Z`�X��#��ی�)N'P�-���ܓ���v�� ���Ϲb��YT��/�(C�2!=�ԠOd0pd��G��^~mmw�,�X1���=�/�Y�oN"l�emP���63R1����R>���EXi,�N%<��m\|4z���(E?����@�o^�հ5�>N�5<���u���I����ι����B��$���E~��Dtw;��\�mkp�|m!;�m�DC]GG���}B��:���ֲ�.�4R�`��*QE�o��M1D\~yi�g}�X��x�q`��I�J�#4���D1�q��w;��/�a��k�ƈ(F2�ɺj���fX�%�������k}LE��)������{��vY�����,�h=-�4��.5�Ū�⇷n���"]+	a���|LLf�)�����5���'���Hh�rR?_�H�5cjj*%'S��.U>䖛�]�MH�7���h�%�|'S���K����d׃�S���m���E������-!�ȶ{ӭ���jzDV["g��Ȱ�yn,,}.nz��}|7r��+�d�
;��wul��;м�JXt��Y�
U��q�+ӥҖJ���X[��M�C�e�k��Ț����>I�L~:y^d�G㌏�8���f#�X����^<gVm��3a���;��h�F�. D8�ޒ��z]�mMn����\LNF 
�4���V���<�;I���������i׀��� X{*��8�k`@�K����T,��'6��W����7 T��aGE5�6C���\+c�He��Ke̲�Ir���zB���
`(�bÏ�yW���=]��|�i�����ŕ��J���������t�!3�^Sl�ӕ%0�vkƦ7�Ȫ��rE�Fu<��v��>�h-�"�޼��P��x�d�*��%�=>JY9�&[er�?��dn�,--?��c�谢��B���eUD�������1���}�%<T!4 m�$wY�b
iGa*z�+� �8R�뇑�^4��{��n�_Hm�\k��������=>̜�\ٜ�ij�x�yѺ}�j��s����u�)�pG�{��b�1b��\��D!�J�D	t��	�(��0jzzzx&N��;X�nƯ_�Y�6�k�[�F1`��{����姆-�ڋ��t'CJ2�!B
}��%X���jT��U�)�%���O��	�YC���?h��m�q�R-�q2�㭬�P�?�`>���:���a���ub����M�.�c������ ��� ��l����� �$\&ٯQ���ҖM��tK�GGv��Q��}�8D�k����tt	a�_��/��GUn�H�ܒu��~}��!�QֳXm������'O�x���yDT?�:��Z�� ��sr0��,p�'f��a���D/p7�����#C`�9_�qɤ~�~nv� >��U����CuKK(�I���|E�������4�5�o�5��FX��F��q�7g��]����l�lYߔ�&)���d�i|#��R<�j�6���Fklj���B�HEU�Z����-����I؎��*/����,��vm�=A�!�f3i{�?e�������aP��➛Aa�;D�TA."b��5S&h|l��7� ���u�t/w�[n����7�DK�2�~H6b�f�������0u��+E+}��eV?�Gcy����X�A�궶p����RB��eG�j����jq�����Q�⮭�M'"g��� ��h�ʰ(��kb��Ap�!��A@�A:��Ni����F�[@�A��ޙ��y��e�k���}�Zk��ظ���a�a��ӫ�Gt������h���?�;�?d�?���j|�{{ ��}g� �L�����>J�Y�;���RSGgng�J����F���_M��a�yl6��l���������?~-�Li<�L�{����-���8<��Y���h>�*G��Ij�H*6|"�|a����\��y��Q���A�D���U����/�����_\]{��fg�-/V�ܶ��~&����۵`�5|�s�`�������n̿~�ᠣ����J��h��B����̅�V���t=}����+��^�Xq���;B~�=�y�Swr�#5�sd�kAUL.y����~��B,�Ŋ�UT�� �K5�y�����U�Q��/$Ϥo�F@�P�nVs���
�EDD�7O޿`��Jh��aJQ$srF|��w������ׯ[k�=({���p%��]�!ja�����Ua�z"�b�qi�xzdL�"&!1�"�+`�%���=���搛5_
��UQ��"�_~����M��~���3�q�B���O�l8W��GG��sSz�;�x����̒��`&���������0-�SG:�Ҡϧ?���5�A[���l�@��O�o>z��ڕ�L��D1j;���c���m8CS��U����W��M�[:��h����ǝ܍
�)q�h������J�ھKqe�br'M�S�/[to��(p�[6iGcap��^Y��P_+����w��9��j�j�h�vF_�V���������*22�-�w����am�#��*v, �0xP',�~\�[<=K�:@x� F��:�P s�v���xrRì|/($��F,~�̴s�@��Wa��$/�����p�ˮrIH.a`1�:�}���E��/����������� )C�r�[�����F�M�Yߝh�ÿ*����>5t�����9�eN��j��Wy��DD@��-1X��j�r��RLD�Ӳ�O��-�5CS[[�h�h��Q$��%���������P�@&���e*�[1��e�dɅ����(��#�*� ���6�2�T�?�a��E��A_\�u��W/���XaSvt)�'e!�c��;�������ϙ�tʝ���>k�"ng��\��nY���U̊�[C� .B��'��璊��Bk⧝�2%Fp�������ݧQ��G�-���Y*%}P)@��4��gTġ��C&�nֻJ@릊��yG6ԚCc^��y��]+�
�%��=*d31�� �N�������}���E�t�*���]���t�45qW��~��T�l�sc���������BjԦ��o�=i%�x���\1�3��?8��̱�T��3|Ok���Z0��Z��Gnbb⺆ځ��SX@^��_�NN6H����Xf3�}u�
��B$�&�eQ�DZ��	=S�P#M$zQ� �j��!�Hn�p�\�V����(<7�Beq���i��0��/������7�U=�X"�-����{86L	v��^�]�3����n�'*�~�w�˯�����ј�,���|ԕ�J��ܑ��4��|wa������oKw4��y$?���Z3g�r�����o�пB���'}A����~%<%�j���}m�6�S�W�&뛻8�u�e����~O�i��og�>(�EI�mj�P�4D�R�>�'e��sRSr �(ӌ�7�duH�le}�" �� ?��׷/��S�����S��L��ZF�x�Rj�J���Lh>p����$RPN+�2�uUUi�eɓ	?�3�n���ꢥCJ��6�jAU�W��j�!��d42�"q���;�A���w���5œ#���E�
��
k;"�zs��s�Tr��A�~b�0QUF�����ϵ��Ͻ>W&���K
 ����M��vo��ޥ�v^�{�C�����/S'�k)�F9��P�8����l��\@h���<�O[_����£� I�b�ލІ�鴺�X�b�L�yI"��	$P��ֶO��L��#>o��j ߤ�J��Đ��-���Z?�4��I;N"/a䪤�t������h�pUZCo��b�<ʛ����@�yc����2�� �"�B|͆g��� ��=^	�����c��1�y�Wwΐ�$,�mR��o٩3�W{ЋO�+£�J��NNU���̈̆��w�������T�A���I��}/�M=�W�%[{�}w��{�q{d!�=uGC`������q홮�<�~�g�3�H���@RJ�Ĥ�1�b_m��/�|j�� Z>W�7�I���G�^�J7q(f�d�L�v��v�`|9�= ��+&
	���<�:�M�P=�S6�-�YewP�'�.�ˇ0��Y�Gcy�Z���|S��*ϩd���g��P��F��"�$d#2j�K��<6�M��PŲȒ�r���C�վ�S�ٟ�v��F$>C,wM�bG�Hw��>5��~sd�S�k��0����ť�[�6t�A�D�Fp�lmqso��!�����#x�o�x�"�D���amw���;Z��X8�I�6�M�ɢ(q��:p��?�B]SS�'.\�Xr�i�h�'�&��D>�x?��{ �p�俯gm�Wq8ҟ��6<�X��"m[Ic�N��5G�"�nX�!1G���u�vMpί�]Z����?�J�S���5s��rCv��MGH?B������j�Me+`(�Vٝ�!��:�Ok�8�^h�DJ��	�e�;ѫ\��e6��*��"L*��ϝdl�DZ%'?��vNW �ݶpᏎq��
�ψ"���]}�^�Q4X.HSН���f�B�Լop{��%1�R6@f�19xI�N����}��bl�[p��NKՑn{�_ή�Qn�٘Un����F����jO-���	����3oJ����L���Re@y��-�,Sm��>��n8�ZeX�)�k&�Ҩy���|�@��j��G��m�ܾ!۟���"K.2�ƧU�	�#�g�N_������%�[�
����*߲8Q�h�s�K#�F�;@�k���8�i�s�%��e�.�ǌ�h��g����b��+cI"�g�}4Q��"㶱?-h�{MGV�8ϒ�)��hM��W"綾|e���cD2�{�Q8��241A5x����U5,�p��p<�.6��a�@�vX݂H�a������ق�����Xs�mLf�G� �ʣg�ش��	MV�5	���{�2p�
�T��I ��&���-�f�&4�����c���A!&���L�ݵ8�F�ni�� �C�
|SW�p�\�6;^[�]]{�a�����lӯBL�	����C(�fl�D�,����:����#���>fKi�$�����K�1��!���1&��7u]]1mO��r��u/�6Yv��4#�@��>��n�9l�
8� �w�K/��]�����V�c2���քe�� M�[��N��P�3���"�G�Q�Z�튕Me�G*��H�R����+t!�6��g�qP���9BL�����D0����[ ���'�yk��!�����Z.�l�&y�&;D� Y���G�g:���+�� ��*�]T�����?�㝅A��QV��f�4jϯ�⚹�vDS*zP	[c�������|�����J�ì��I�$[�B��PIX$<��1|	���M�JC�1&U55��9���;��?��|Oo�>v���5�����#O�>�Q̩G���u��8d�����۪y ���>:��wW��j=�������]t�Yjpd��<N	#����t�sI�^/�[=��qi-�S�o�H�d� �	�r������D`P�y�K�[��H<���.>�,i��98��%�" l�}���[��hT" �'�����K�ð�q?!��U$6r\�^q���OM\r�.zAFa�ٯ�*>o�z_�m �濑����9	vL�������zA� ��t��B\�P���hʴ�
�=K
�x��X�`P&��Pi����з�˕��L[�ͽZ?��-l<���㶉	g������j�$��>�v�]h�E�J5���^�eu��w^&��U���E���{��88p���po���:})������"�m/����nsNh�#�t��&�����w�(FZ�k�7��4Ƒ�+�
?(C� 9{�	 e�|��D���O��Mث�VT�%�}�_3\��'}�c"iΌ�Q�X���o��/�
A)��fys��m��U�5�A>��bX�}�Z�S�����C�R�W%���(�o���=n��"w����#���t��K��P��m�Xe�a� �r���a�YѼ�19��]�u�ba5�{�f[[[yBS�9�,Ӽ�4���?Sc���EVI�0�7!�5EVX�iVt���%UH_����q�V7�/����5_��p���k�[fV�Oq���)��?F�$��J�K���_�{g4c Y��}]�fi�����>lF�����U*���7A^�D,PJp��.Q��S�`tm�U���.�"����O��Bu��v����?WV��.�L���f�u+�D_Ȧ�f[�$�}�-��h�DKϨ��~1�,r�:�q�.1+Ǯ��gHg���[�>�_on���d����]!�h_�q��.,.#�m�9>��׼�f�� )#�����O�X��WNo6�u��mW�N�3��+���;U�_P&�	�֡ ��<�*;���ս��g����Q'F?}ɱU�7����`�z얕�pM��a�b@�,��)���.�C�Ȕ��(��Gu��<�LMP��	Hր��vq_x�d_���b���"vz�vfI4��t5����Sq�;�Di=cJѼw�c��e����E�%����G
T�'�8�d�6Y(��
-d)`��N~����)�j�?~i�HAV�X �vnB<�[��
˲҇eͮ�J�z���!�����9���Ff�ҹ^�6��g[�SK�9�]��][ԧ���< i�\�/���o8�1��:E�Z�Φv���sP3/�J�����şU~�c!���N���F����3�e�����X��\��XC�w�n�!������`��@��n�-�,㳗[��|2�ZD����	��Q��Fm� ���
]��.m��a��v-"��5[�\d}�A�\�N�r���p� fi�3�-�=�ttt�.�-f�Z�އZ����l��/�\�Сisc��i��� ��4_��E Qb�W�Nk�I�C?7$4��&lZ:�8��,�DK��]���]�a�#��^?���FX���%��(���Pl�]zn�ؒ�<�(�)��;C49�,�!�"[v�hl,�wφ�o&q��A�1���� �=}��ɂg���Ƒ8�|-Dz#5KČ� ��w9O�W��]F��ؙJ��*OF5z{v�������%C���$)��;�*�&�|uabIU�Λ�[e��%�|9���8%�]���Ϧq�LSڏ��>l�=�����B�6\�M4��U�R�l�S�=4RȎ<�R�) �N��\pVQd����{e��B׮��/�e
Cq�*�]{�mՈ�����ܙ=��>��t��@,0(T/m�� �$��{�����I$f�D]nN���w��A�}�R �(m
9NQ�C62\�J��j���� Q�#��7�V�S-�~�-;���p�(t�i��p��^[z���ǆ��C���ѱ1�o�äI͏9W����o�����P�$žɗ-����n����t���7��a��Gc�u��S:yOo{�¥C��F�������}�G�g�뽓�['���jFjh�g�<e��RsD5�T@�l���YV�%uu��a8m�5��J�k�7�
�p����\E��G&�Ȍ���n�k�:f鑈��R�������+K�=����k���m9��X�aɟ�Ã.F�Wx�n��+5�geY��C<��/5��-�P�0S��5Ny�q�r�@$���^p0Z���7h"��z��bix�����{~Y�@���^�(X�NG˶|�ܮ�r�c̖T(��̣ٵ�km�����uT��$���v�������7=�T���S��V	���_p��;S��cT��������Q�S�>���9�D�|r"��h�	���l3*��G���l�����Ut(�x��L����W�|�O�f��M6O�AFr{��|�����fIĞ��Z�eq�ж���	��o��\DH�����YX�¶:�F��z��EO���;d8���)rA g��[c[@��:yb	�����b��+�0���zr��e��B�r�y#f"�
�0���H7B�՗7�lAWV����X�"��^��sY�}䓞-��3k:p��N��ϩG��_���"mD�M'��_�ӣ名D�2�����O�C#>��n,B�o�H@dR(�R�P遀�8�p�f\��&bJ��?ifL#jT��!?��sh����l�{3�C=j��X'$,m�+���;���!L���[tg���!c�"y�7��e��g��'��C��lG����!���D��I�l]�L���
��-Ġd �כ��0.za(N����Լ9��7���(�$q�Y��S���C�C�="q��3�6�<[��bq��4�����%��sv���s��{��^W3�̶jN�P�T��s�� ڡ����@��1�M,���Z�z�C40�g�'>0��S��~���%�c�3顖�(���.����S�_���c쵼�*P?����\���R'z�j}�9��h��p�4�k���;��e\�]݇/�ri�������\����W�̻��e����:0�a�JD���R`ځaN
ۿ����L�>�/�O�RA���MCͥ8�pB�s���?w�֏�G�HH����[ɩ#	��}��'�{"��6�.m�=�U��R*�*T��77N0*�3gi]�4�)���p��~�5I��Yƌ��?�f)�U��^�R��$#������?������G5�����Q�R���zMoTi%0ee��?���{pp�?T'Q�>�mkJ�$��"?�,X��ȶFJk
�k��V��>��8"CQ)�,�3i�%oD��c(ItK�*ȵR�.8(���*Jj�-��x���s}+}Ye2F�z�l %=~U���	~Z�A�ce1������2J~���u����-��k�15��0��#[u�/�l*>��q鮽��Ѥ3{G�%�Kz�=��'S�-'t,�u����>�T("�E�f��H��B�1��g���/�k|R���؞��py9�p3�B%�rL��Z-�����^VB�Bk�u���J��1I?���� ��i���{ޚ�hl���=r����Q�Y��|�8A�i%�"�����3�&ҍ�ih�+�v�ݭ����������֫�D�0�6��BcW�ԥR�:��S�
.:�D��͖��{N�P }��27��OV`�*f��҄����ǘ���I.x7����{�z�a!�� x������B���uR�3V�Ea�0릊�X����Λߞ`MK�?d���"�}8�Gd�;;�}�c���Y�z�]oy��ɥ��[�(�A�v�D�f�T͍�`�J���c!�ɉ�^�x��1�^��g�i`)&�����d�2�6<к�;���Z��4P�ŏfT�^�e��x�� �-/H��m��ݮ�>pCk'���zZʳva�a]evM�F\�S��QٙP��x���+�F�\����^Ȉk"�X���������?�*˥�y ��]^8�K���W4�J���/�����5�I|���+B��[m�<����H	��BjH����A�<򆫎\7B��A��h�*�s���MBfmE�Tq~9+�_xP�Z����������vȤ"���/V�I�3C���KۿnL�%��5�=A DNrp}�^����|�t���}X�џ!���>���{�n�n�X�����t�Jx]w?��^<_r�%kք*o�Q��ya��{9�UE0���DMե�"M��Kb�B�"�1[\f�ũ���K�p�
W�->a:-v��ݑpD�a@7��v����H/9�uw�jW����q�a�h����(_�C����mUAQB�G�
�ٰL��g�Xc~˪���0�׺�}g��E�r�D.A Y�h��u������"�4��kX��wh�6���g��w�t��?&���Щ��^)�
`�g2
�w!�P� 	�^��d���R��������~�c}@���ScF��l��lC�9a� ��)�t�SU������֐�����+�4>�6ˡ���'M=}�W�J���`�H�~��D���J�!���r�W��?��8�=e}X�������-�Z������T 6��T��3�

��B7EH ���$:2�����!O��x2W�5=�E�r]�N�AՑ�<�Y��w�ֿ��M�Ʊ��|���~6d�4�d��u,d�W��q�m<�c�e��7�ec���[��w>�ϷB� UPOPT����^�V�JlIt9v�9.4NgJ�^\-�Q^�2��ITM�Q�&�:��V)�����d�:�v�i/�0L�=��u�`!�8�R��"ݞ:�j��m��H��H*Y�#W~` R�i�́O�?�f������&VZ)>���Jϊ	8�`�?:��Fc�-rL�*��U�����%W�i�-���'� H_D:@�Y��i��a޲%T���	(ʃ�R�q��Z�S��_,�=O?�I�a�-@j�d˧i��7�%"���CFg�M�ଊ�/�h����t!�_=v�FH�[ʿ�L�
������s�|]�efeUL���'
nl�Yc������H$<���^�A����֚���+��_�3������X�E=ޏͲSg�Bc��j?�͞,gS+��7���2&ER�(,0���0�l^ŲZ�5�k�w�|�ѯ�յ����f�L��e$������R&������OL74�j�j��Ot�6gJ��	:�0*4Z�s�E��h���߾�z�����G���
T�,M�_LO��Y��y�zް���5Nm:��C�:�t�1A�B�v�su�Cŗw��=���^�:�J��Q�Wz�AI�_��=���c4�xh�~`�G�G==�i;���9xa�z\3���`�>����'_ K�U󾛲� ��3&t�3���X��>7$Pb�5x���a��`�tl7$�������xH[YV����������d�$� %�\�Io��������r�@��I[|L?$��ʨ��\��JLL�T�z��HB*���κ����1A��g~�~�7b����lllz�pt[�ّt	�خ�׵ t����V	���j=1��F�c�MUm�X�R��Z)J:KI����I���O��b&_y��ӓ ϻw��x�Hؑ�e�+�àl�ε�m�p�ҷ�9E�q1)�Ԩ�sJ p���� ���sI��"���A�*n&(�P��`�k�����ڋ1��P9���3��v;B�N~!"�9��7��LLu���D������>��sU�9$O�D�v%��6�,�9�*U+2�I��Md�M�x2�e�aR�O��1P�p����y����$ʠ���Mw��--";�{�X^�5����긅f�N��#Z� n�9FR&�0mK9�NF� Ȳ��NV�� Շ�����d0�J@��� tKn�:�@RBIh����9h�|��m�qn��d9��d}KK��.���RWH$�d��l�c��$�8�!A�2�P�< I�p�1��g������MK�mܟeF��#£N5�[.��:O��o���c�" �����R�Hv��N�P�N#� P[
	cVdT٠�V�!T$�_���ݚ��$n��k�Ӈ����n}B��v6vX0�b��uА�'�$�K�PK0�F< w��M�6,�����8[3`O���Z(k���/�o��/���Q��IFU�� ;����蓘(.��o��R��=��y0.A<�dX�>����D��Bz;��KG]�k�ر��:��ꍝ~8C��ŗ\���0'��vX��<��*����#1�A����<��T�B��:^�2F����Ğ墭Jݹ���Q��+TE"	{F%r>5e�eaF���i�wD��r�另4ܤ�1�eH.�H����`�R� ���|�c��̛�p��N+����+�}V�J�=��:��%�7�bi��������h��ذSYu%�Ѐ�����|/{?&0�7�5>���~�럋�� ��)�rPW�D����o۲� ��*�@�P_�u��v������
'Oq�X|���i����ŹN��A��f{�U��v�z��L�Q�k#ŵ}�G<c�겂(q���8�U۱o/.Ȓ{�F슬2@H�}h?ݟ����p$7b��~�T劥��%+����4ƧU�J7�^�l�4@*W�!�8�ǅ��]������	��R�3?��?�WGg9�W�G��@l��~��5R��sɵ�D�;��vF-�Mp���>/˝�%��r�)r���C�Y������љs]��|y1d�bdhff&��2����}�(z���n3�%|J7:Fr<;�~:�]ν���2/Q� �0�S�/�ׁ\��0��\�=�� &J���,��@9�����ӌH��Niג��_�p0�\�D1���B�ɜ�`���IW��x�;c݄ha �|�s,�!���J% �%�,R!�7��s�6}�;;*YӬCҏf��
�H$"�]�c�<�릐y%y*͘�C`���@X҂��� ��`�H�dpc�GFOǔ-��6sr��h@d�l�waOD����B�E�� �ˇ�м�;�W�
V��a(lӢ�'�.9��ڃ�F�&2����v\wܦ��B����E���! ��[�����M�P����h���z�`r�RiҽjZ_�F�F
��/
t{�(�;��O�x3�B3��H����_�ގg��#��/�}y�`�9�p$�G��N�(i�S����Z�t��t�������+�~0�����D����7y�˫8�8�"�	�A�m�E� (�,(�l�&=�y�Ɍ�<�\�cR,N`�4��5:��mȆ�_�5�|��G)�N	��ɝ�^���_�B�k�����9�0�L8Yb���sD-j��@R�� Su_�|�V�r^&^l��G[���F>F�˧�pr��Xq�:B>�Az`>0"Ic��*!V�S9v��>�����,�n0�g�_��$�ˉT����BbS~4%$Rڽk@*�j�n`\ɼ\<E���y���ś��Zr#^e�)F~O+��D6�4��.��xI�M9s��u�.T�D�"�`5��7��8Wj��������F�\Q��Ѓ�y4;ʤ�H�ֶ��{�{��z�p����h�<�5��l��ևS
��W47*T8"���/j��m��A��,{{|���g��Ɲ2��"�?����#�Dh6C����	��=���ZTF9�X�xGȊ�Ñ���l@z3$K�Ĥ�B(�j�m2N�L�����#+��jH��	胆X�*S=,[���}!�"
�����R4H�l�[�,r����,��$
�=��di>�72�������t^� ��Γ��.M�G~YBA殠�E��i�H��6:�� �6H�{yQEr�>&Ф�����(����H����֛6�b�-�K�������7�/T?t1�!�ư����ͦѡ�����,��]O-)�5�JA[m����\�O�	�E�S�'η�kwپm_(���26욅����e��Ĺ�9�����AQ�Q�r�/�O��ER��(L����$���20����Xc��и���N���pP�a3��3t�S��Gw���SwtSd�������paP0ŁiV�VIuEm��!G#!���Q-+�<�)��7�p%l`����T�|��,��!l4������T�bQiH��5�25�`ҁ�{jKZ�f�z���s�L�O� ��5�����!�����Ͽ|}�}�F�T\s��m��0S��w�������k�ш�b`�Ե�ŹdV�Z`�6���`���dܥ�A@QJ������L��7H��\�#�X�Q;de��£_l��%b�麿�0�P��a0˛����a�����!f��ؘU�p�Hg�z>C΢�e8������Ȓj�SC����dp���*�>���NّE�L�+SaLaq�x6Vp����xU�n�������gx�i����~�QF��_|�����<���sN�K�|���E�h{;7jZ��y�'9���t����D2V6	0e�U�a6tg�aJ�,��!�J�{��P�KE�4�=U��wC6�D�2�
��R�p���o8QȢJ��U�O�l�r��PYΞ8�H�J��� $B���<")�$�x�+��;:����QF���E<� -�����u��Y��4� �����=-0q������3���+���m��/[T�����(����F�M�ا�6a�������i?���D\��p���v��HJ�;D84���>�!%ped�y�Xu~mz��-��[6SCo4�a  r��#�s����n�Q����/��愵	���1�Ž�?��HX��|[	c��^�-Xb)�(_��}2�^���Sv��~������L�^�a`��2 a���+Ӵ���$fS�^�b>�i�.�WPs�3c�^��w�`�n�J��B�	{C��D�E��±�FKP^���<K�*�����$?2z��D��Ð�cR�%���Wҥr�_ p�˙�
K��^v'v\a�z���M�=%@xwJ
���/��'��Q�%��i���D��nc�楧�*�><u~�3]�ۻ��k�<�٠W�v���Ʊ�6,��5�a��_�@7�5i���,�1�	�E-�%E�7^�ɾu��N��8-��\�r��|:�y�a��Df�9<��[�-}ϳK�����#���Aր�ě�#父�����|���Ur���w�ǻ�)g?�}�Cϩ��"$DA�Vq�No�>-�:9>��rZL��|���;XR�jJ��~&՝�a:m���70�ñ˿��w�0��Jn�pnk�=�k����Q/��.�q�3�;kcG�čq�ASt[��L!3�Zߤ��d��σ�8��;[�_a����05��HieG9Q��P���2zoE��w�2�l�"$�w����7`� k�w4��s뎿c��^����'�?�,�֤A۴�IrU���G�B��M���t���V��l�m�3-�w��J���&x�˾�o����$��" А��7-mmc.���2����w'���L���>c �
l�I����;C��l8��J
>�}��t�j�E/ECcZ�e\��Dn#_�����SIzѡBDD4HG��s�!��Y�D�-q�݇������*"��7Lv������GU+�AZ����%���%đ'�?0��zfV=�&��(k���F%iU׹/�K�/����X�u�t���(afe%1rԩ]bx����S�Ūe�c��vC�gG��c[	-@MU��<�"	�5���:��
Ax�4�������f�� �V?��A7��K���绀���t4�oa�s�i9~��Ey��%_��ϡ%l��Zs�ؒxN��t�z.ݷJ	w��:7�j�f���;�屁����~Ֆ*���}F<'���0�c�mDX�$�|V�b��w/�i�,r�K��SV�}��5�C��g�[V�g,AC�[�i�:��Vj�dB}�=DU��%:�L�q	��Sr�J=5��� 5�㽖+������S�ے!�;m�ۂg)��P�v��Okv�o�������ݿe���X��,�Q��.�����GF���(�߯�1��s�nC��-�.�!��I1��V+��@v��Έ�;���_r,a!Q�j�fز�Т;�`��$�m%�}����=�\����f3�͔���cy9��\o�Z/�S��K�O����Q��P!�5{�bbh�^�qJ,`D%qV&�*�;�2o� ��x����S���#5�Pb��[��`��j��߲��Ś�m�~@���nT�%�}5�����N��(b��7ƺJ����wC"��g��}=o��2H�%�Ӓ��$�I]՛�ī ��N�ɤ%��>9��Y��$��91qLi��Q�f�Vڊ��*����5��a�&��G��yfN���tW�P��c�p�B�Y��a�իWg��l�w�Ok��"���i}�U���+���ׯ̲��Ro��[kt�0��;l3Jc6�Dҥ/��+8M�^0Ѝ�j�_$k��U�"V��/�)	˪�9�k�5��4���L	8i�t�X[���y�'����\��|/}4����h_\�\��4���}b�@���"��Z@Z�R&��F�a�Y����"YŕK�/�Ě7e��P�Zs��u���2tq�t�Aq.�I���b[�g��O�Sl�	��^Y��|u�a��GV��~�z��5�I��!���2����tk	p��n�0 i�e~��Pj��E@w�7�%����P�"*�U���y*}*o�p�����I�z�0jX�G�ߘ��5LjL�)3�DU��/���i�Iy�ы�OgBZ���Z4�{V4���F��K���K�b;Ҳ�&�})0�8�&����\b�S��L;`�,�	˳ȋ0i��I�`�Ֆ����u��5�+�������D����2u]01��Y�f��7d Ҝ��?I^���87MWxɨ#������i�4w���W([c��,�l�%��^	� �#k�E�j����
 )T��f��=��5
����z�'���Zwl[Ύ'��=���	yr���m���L��VgR�Cr����YQ�
W�o���VZ]�4S��d�l3��ڴ4M&2ט�ᾬ��!)��t�s�U��s��4�=-	WO����T���dXJ���f>���3�4������kA	Pf�b���y��Y͗���ɟ����9 ɜ�+�kV��/�K�hD�D>���j�s���ǧG�Sj�Z↫C!���F����Q���� 3�p�vQ���bۚ�ko�N�Ǵ��Z=R����~�r�z����ޯ/��ʗ�fҌ�k(,�t���8d#�����~�ɖ�y^_��tJ���{?W�g�V\�/
+���Տ�^Ta*Ǵ�1��T�4�%O�ײ3�`����5���fABй�e0�n�48qY=�-�.S�e�#s�1�\,��u���ڞE=lgٲ�V�
�Me9�X{�xx�z����?\�������p+?����g[s�|O�l����u$�&�4Q"�����|M,l���\�_�4�P��Bb�X*K~S�z%�$uH?%��җ5�wK�����u�)�3F��Ke�3��)݁b�GEC����MHݣ�tR�q�56�v���7ɗrK`�q�?��K͆qE�#	� �4�ʨoa��z��$�v�ٲonc�~h��NA5�U�l��A���
�L=M���U���32B��Ȳ�ۗ�	�'�/�K%&<⢬݈��M�דa�ZԒ]��6�=.3�*�ҧ;����2��=y$E�n��bd�������0fޡX�
G�׎a1aפ�f�f���$����|�֒�"2T���NxolAɱ�}���>5�2TAeS��'�K
&&�7�ԏ<m��N<��7����H� �F�ԏ�����{����I1�Ѝ��~�1F��%ܴ��Q�8�R&�Ǩ~Ȉ@b��ǐ>`�o*1��X:�i��\�����%��	L���7d�8H�hY5���wG�&+)�3�s�eY}�׾X-��3�#�� sVn�^2=��`\��h�a��d�A�8�ӮN�_e�,[����i�)�=�~W�t�b�&����N�GA��ϖ�sFf.�^q�n�-��笂�_g�Z
~��n�%]�q��/&K��s��(��u�FYB�m�ی�-4a�̲�w+��erϟ�·�<:}.�Ov�&��%V`п-rV:���
�^�O�Hg&���,�A�:8��U�W�55��6��`6]�����Z�φ\y��]H��4��&�a[��+WR��
r��\������'�-akC�(��9`�/�����o�W�����?o��l����垃�G����� DE��u��@	CF�����\޷32\���B���\{���a�A�OŪ̷��tQ��[���U+���@J�l��V>K�QMg�N�h��tI��H͆8����p#^���_�ֽ��E��5Dl��MD�,$(�)�wy\3�*do.�>.�=�������'\��c����hMO+�.bŻ�؇H��|z�I��y��o��'<fa��9$�:D�������Ly����C�%_c�4��^r���C��ɕ3I�����$�K����~����������fξ��+T*��
��I�'3���2r��>1��H��JtC,J��(��3���~�_ D�����S�}��n���L!�_�ޞ��Ͻ������t��$��z+���:�~U�4ޣK��np�Yt�p�~����4��Ճ�&�}��p����k
��o'���⋐@�1�ec������Qm�K��R�b�)N�R�
hq).�Hqww/^�ݡ���5���]_������ˏd嬬�s����{����T��3��t�2y.�Yi��Usz�)�(�uas�?BlU�Z v�ِ��볁2�α��Ǩˏ�M���� �U��D� �_����t�S:7��|l�6�/�M�~�cFy{�  �SF�d���'�l{ 1��f=3�7'?����	YQ��״��T��S�D�ZՋ�{��闔����N��¯����AR��HZt�Wl�]/�@$�=�^�~PI�UX]�xi�+��)�	Z�U�Fn�����=Ϋc�ȇ�\�3�j�x�hy,�2w4��uE-�$J������3m��5c&��Gx�6��&�ჶ^{:79��9G+��e[�����ݘǿ��eU+ᨀC!�����:E��`n��${�_J9VO�Ncg��"glY{.�}h.���r�(����������e�z�l���*�B��k��.b�4F|0O�������sе��:p�О:r$����_��RCx@u^/���@�A��&oO�i��Pۄ��h��k���R�쉨i�(�W�I������m�ṡ�������RVL��";~��!=a�V���M|�T�]����h����v���X}�]R&A��F�:�L�Z�q#�d�좂�����_�ydҖ�,�*����357��$�54�Ե��͑y��;9�U�S�b�౺���_w�mS��Q��%��0>�I��d��/���X:Nd4Q;T<�TLBd��L!��I��c�@bys-Y�e�6��ɗs�����ޫ�m�٘�ɢcRc���jV�'�Y�7�#f	�[ք�y)T�Ʉ�
GEz�Nw8�.�=�;���!��䪛R7�P)� U�Z����1�-nOq�H���mb2�.ծP�"Spro��~�7w;��ps^$*նT8�;�i2���IWT��������W���ձv�i��΍۩��r"ï_;��̐���8-���fAdSvtآ���y��Jx�[��_��,8m�ǆ�ɥ�r9G�#`��^��i�S�(��j�����{T~��ό!#N�7�lԥ#���������|���/7����)|�47U ���V�k���£�Vh����r��2�+TE�yS�����)W���6�x~"��X���\��.{`��L�Wb)��ڴ�JhT���|�<^���Xn�!+s�G���F������p�P�����9����q���rv���p�2/����rZKF+eH�D)��$2�ٞ��#Rr]ZA��{?\�r��^���-usa�������!����=%�q'{���z���}�� ��K��1y+��@�`���e3����9Ww��*�Ԟ�6��o0�<�����P�ޅیP����!��2*�5���i��,�j��F$���"���"�$�F�u�};��\�p��9�m��2�8���˜�r�u�	��m�ttJ������2}����`��Li����]T�jъ^��&��|���Y�e,n�֫�!4����Y���hN�� ����ԛ��ESk���D�E��_���Tשa
��%\T�@���������P�?�Y���"���3��\�g��A=�b��	p2y���w)��h)o ��ϖ(�{!����?��c2E�?p~�⤥����aM.�`F�ם�ķK�+��W���H��+��"9A��s&W�nY����w�斢gX��,l�t�H�Hğ�){��<���u�:�`z�1�2fTo�yd-5�Ť;:��]�/�c�}������rJ
�� ��v9�����+u��Zt�vu�.�~�[��9&7��Mrlr� �R2#�����t�T�,��ī������aJ1��U-�0�r�?�L��(p�����~Im��B��g>#xK
P�9��5����|���2�
�'N�3�hk������軼D}��]G��?]V�M%��y����d/��l�%�FH�_�Eo�(@W}<��3(W��
�5�E7�;g�c�sf�'�}�7>aT��38���Nc�7`hH>�'��i���KOM�O��jԟJ�{AXWғɦ�Y�Ȇ��ؙ��U���`��kyr ���A���٘ыQ��.�<)7�%АW��7����R��C\y$]:�d<b��!ʔE+7Ih��ޒ�����<{cp�1�Dq�,��s��5��t�E��_H&�6*�]1�U ?!P��.O��3Mh�KX�bD.�ݷ	�loQ;ny����i�O8����z�����$�DSnͮaS��7;oj	.�y�����D��.���!nSM>B�NacO�T����T�I?�| '��p�U`/E
�G��Sn����݉��n@��O�б��"�$���(w�*sm0IA�l��&���鴭#e�ۅ�Y��F�Ut�M�D5��1�T�`d�3C�C0#������3G��u�*�BE8��e�뷣12@H�4mv��5�Dو�o,r�����Aeb�����D�v2y~%�.��kс�{�G��p6�7����:�;<��yy�$�R*�ǂ� �[���^�zEm��t�8#���uLz�������(�n焸��<���f��U�9�D�./v]����9:	��
O�"R;�����b���y=�cm�4R����R?[����cۙ����Q�>�t/�G�c�ow��]��������9�z�Ü����4�ޢ�V��j���t��9�ϓXS&{��T� ����Y�������֡��4�ܰ���M"K`n��^��P�_�\V���R��5i�i�v��aF����_�]��ݿ�L�1�:d]����E�0�2X�Z9�@X�D�h��&Ǐ��� ���z&�A|*�_�3���C����I?���S̱��%tV�V���3+�ZΔi�=��=\���#�Q��U/��slջ������L=�9L�vn�ȓq�(3	ۀ�.,��B�_R�K<ޏ=e(q7���O�]pT76(����9,��{�<\Tz���)Z���WpA��'bm�x�8�n�3�Β7���:�����.vxn1�I<�Ā�����;�L�rD�F�*t�aƍME���{�p�qT�+0��5�����	����"�fV'G���{b�O�ﻥ�Up˚9�t�햰HF�Y6aIĕ���/�����2-����F��t�{�g�^��l@Z.�+���mX!@HΌ'0x����ws(e��n�}����# ��� �N(����z�t5��$&_�o5����i.���,�I��^(��Yr���� �:pY�:ZM��Kc:��ٺI1p��9�j����{vBf褭�k�wy���}.�-�@��+%:��W�(�y�R�(6�H��|4,�[%\P�� �z��{���{s�'Ɯ}���p�x��.5�7�+.6इ��"��-���઻������:����.=���E��y��)��������'��(�D��M~��2�P�����yt�FvMq�iC�af�	t�mm�#c�)?���6VWWo>�گ�;��r:l�S@�Pl��_�v$��Gt�<�h;{����	��TY�Y��#�!���X�eݳW-�{���C�s cw�O�����I�nd9��m��E��kwd;�:��t�7]٫����Dgɵ�Q�
Ĉ��O�SS�3ڪ��3�2��ŷtYE2�t��p��U�fP�t��#������-���=�`,�4Y-�T�g�/ϸ3�	����C]<�>.[�7��f9�Ϣs�b��{��3c,�)[�Q/�O�6�40�#��Cv�������%��i5��֞!o�^CJ�����1��L����W�
k���e�w�K�u�[�	��Bh����4l9��dv�l��&vn��(eH�{޻U��5G��.�70{K�Ns%Bnp�B����yG��&�G���{#�kQ�/F��G�����:[���
3D}��;N�~�E�nl=&R��:jy�p~��3��/�ܶ�*���T��}1�X6�f�+�H�y�ߕ������*���;�mz@����K�SˏM��5_�����X�\�
|�š~��:��u�pD�Ԅ��|CYs�ЎZ����$F�+O�J��w�ϣV�
� �ܚ6o�p��^��w�^$� 2{G�̯kyh��B��{������w�kg7c�ц�]9�2��Ug_\RN�z߷GdE[�T���u����Mļ�l�5�{IG���/ �����q#�����^�M���������ݑ����̓�K��2�|`,h]:#=�xO�j�Y�R��y;���s�;ʱs�� ��]�E���)W�zD{�H�~�|<ݹ�Hrr�YyEuA��7YW��¡A��s��8
z��TCRثkjT�����7���5�It<{N=&�*`>ΔJ���A��"�����AfN�S�����=�z*�����Ʌ­��f�n��;?�p�W�L�'��>�7��}K
�2)u��E�C�In~{��)
z���P�%��|��$z�&گ�ط�B�\���xM�y������a��Q6��l�,�t���7�*O��m���&Trj��Xr�a�$�T�0�D��jdí��?�z���GE�Ӿ�O����T	���|�i�b�?$��A��A}82�(<���J�m����
mmm$Ƴ�榦AN|P؎S۾���0�zm6:r�unڠe�55P	'��+�A@�F%<����SG5�6{�y��"�BB�?6߱�4g���sϩT"ݽP��&|ul<�5d^fԺ��l�����K2uOa�=;w�Ŧ���h� sv�3ϑs`�vt�of�oP]mgBxĮ��f@צ|��T��y��ٵ���Y�Hw��_���~	�KXI�gHK�(�23 -�bz�gR<�2@��>2�G�?����ux�i�+�ND[�N�zȕ��!S�B��)++������B\�� J��lX�"������1kv���i�I���L{�-D�u$wvv���s�b�4�y"o_�5�A�g�^m7PS�0���$F�ĞT�U� �v���VQ�v� �y�(�;��P��bW�\E���~���}6|*X^�5K^�N���Z��ɵ�A�I=z-m���8C;�ު��@r��9�����ag�;�5hWX����r`!�^/�e]�r�����,�ٯ�r-�n��`ka����>E-�E�b�5b��x�r��oS5ft8R0D*�M�l:�nT"�o�+�`{P��������|���}#?�����Km	�E(�.�`���F)�B�߿��[�����g��ʵA�
e����B}H>�޸^	�S�*z���/�����.�&���2!�T+f���_������%�����`�"e���a�\�g�ů��U�����	���燑⋓ ˬ��`z���	&h�{۽�b�i�;/�k��sJNI���2PP�'�Fl�9�G)}�)�ב�\|��g;��L���ݖ���F��/e����R{|V���GVHA}.�\���n�Z���4��i.����������q��92����Uk�0 �,(ms�H�R_����*����e�T�+�ʕ%_�����(����Efm[[�z8`�f�"��s��#a�1*	-F���e+�ꪼ�Uc��a<�4�O�`��K�}O�h��:��,4,��FP�Uy��%6_�Xq�����x�s(�����L*x3i��Cb���D�𑮢���Q�g��Kؑ����j�T��ݤ82T���WPP�m�twԙ}�q��Q�lJ�����9���o�\Й
gShMPͲC�k�-�	R�~t��20^�\��VU���������C��X�L%RL��|�9 �@܉&�3��D_�Z�m�'�=��)������\�o���e�m������`M��<���Ƚ��^���+�X	�s�n?ا��3UQc�f)�i1�K�NSЃ���s�^#��.�X�S����� -��<�6�FQ�?�{�0��wk��D ���V����g�_�2c�X��UAQ��I��M��f�Cc����y67�b���a,����b�G�ߩ���P��ll�@-m����3ϡ&O�·�N��#�ۍ���#|5�k�u|���d|�d��"j
�`���"fo-��xx�A%#��`���a��es��R���2�y�Q.c�������8��;�B-�rP��u��2���� �pc��&�� ��U�2����x�Rk9�sEH�b�i7I����J/Ў$J:2Xb�8�]�u8�FnM4:o~��B̀5\��zy��9�Wb]��\~{�1H�@��:ʇ2�ʈﴅ�:g�@��"��*"��FM�c�eH2E��K� q �ԕ�7���� E#�U���B�8A�!U��[�4�-k�KL�ЗS��i�L�'�V̅��Y�_��K�}D���\�oWDmO&�Օd0dh�F?�ɱ!"$��k:M���~���Gpg4�v Ty�R&���v��C�A ��ȹqY�.��'D���?ƛʾ'�Z�z�q����y�q��R���މk_ʒ����"T]�jf\�0
]BgHm�y��G�����msv~>wΚ�,*�k�Ry�Bg��Ik�ܨ�Β�9�o�Dor9����=.����@o_O�H��R��[�bY�0���FZ6�+2�T�8��ጎ��#�T	���.�sF	Si�[qAc���[��!Ž�"3�(>_�f���E��2j�����s��{��o s���_O�f��:uyh�xaE~l�e�$sB}�,�e#`�,�/�N$11�:%5]��1ᾂ!b��=]v�1�����=R�I�c'�r�6��C~r�w�I�A{�=�12�X�`!���=�;2\tn$P>�T$l�;��~���n��ֿ_'�K̅U�\�7���D��jFI�c��0U�(d����~�=��C��������Iw�|�(h7_w��P�%>�c�B(|2��}z��1�<�(O�:c������a?���G��p�X�e|���2���D�0�P~|\W�2-�.�D���x�u��+��Ϙ�B����y{4׆��z�N�����'�~�E��?ډd#H���i:�R*}���sٛ�#��nc�(~ʶ�2a(k��z)C)�����{�$���:6HO�s�OQj���E��� �+ݿ�|�E� �mͤQ��i�H��]I"���5�Q�5+Ѽ��u!�4Ht�Z�Nz)�h�#	ï=]�=Ⲇv��,-v7�5�g�ʪ���4N����*��`�1���>�E@��#ط��,_���<�~ё�9�I���K�b���9z�뷄rbPc�6g�Bb�r�YtsZ�O�M�3��,��c�-��(ݥc�|�" ٜ��Xۇ<f��8,d���j�Ny7ɼ��
��fVܾxwH�qTW�Hm����HV}՗�3Mf, "��B����.Q��d�ȊBZ�"I���M�*��G�A>�l�R�&�4�)�1������s��B2^�������"�UO���N��'��¥1�A�4o
����2��l;��`���t���S�I4\� v+��CpV:��xC�,��J�fDv��i91�������T�'o�x�* �L´�L�MJ+�f�]O����B%�2�
)X۠|ň>6��6g
�M[�Z5���+�M�X�-Lcj��OCh���:����d��ö��3�\�\���E]���1���W��?`KM'>���Ǝ=���#�?[|�,�x�� ����!�ʊ��� ��9��D��;�K��/� �d�>�x�]F������竹(�V9q��Z��Uy4cԠQ���A���JJ��7��
�W���x��ox(�����wд2zt?z��������{v��hEP��q�(1�B%i��䤝,�-UP��u˄?�DP���o�:�}�S���:�S�g���lW��������X��_˫5Y��)�2�����)�Sr�3S	�gK�.oy�S�������^:�xw���_0#nm��tB,�b��o���Á��=�J�ʙ��?I,�S�JdQ�v'@C��2�4U\+��Sz�w/S��Y��"C� �rF!=Ã�\
,lX���v<�-��X*�%Mɳ���dЏ!��zԀ�
4���i��ڨLK�"L�O��bD�L�i��叽(�Q�W��xz���NNS~7#XZ�ś'_!�B*M�ߧi8�T�4���F�����~��Q�MGa����gn���Ȧй�/pSm����Q���~C�&s"� �|�M��~�r-���L������!���~��hЮ'S�OdecC�nA��&�pR��ՠ�./oEv]��l�QS�l].��Wgk�	6	a�r���r���(�&��#��ɇm�R�ţ��	��4�Dv��v���%�0'��J�e/�$�m3i���pm��B�bg<�8Xn�D�p�_�N\e y ໬b�1݀/r�A�4;��8�tKċ���,�?o��u���/����	���iOT]t�?<�2 _�̈́<j��R���F�u������(�����M��,3��2XF��r�f~�N-��B��]�ת�C���x����a���{Aw��P~�.��*��76&Sd�������Dẏ�X�7�t�"%�����9��wd��[����	�?�����n�1<�ɥ�K\�ҢH(�v�l�l 
���onӜ9���\VF�E���d�s�$�~���.j k�	�+~>������	w)=�B{9��o�Y�*����w̟4u/hi����p���.�b`E�)c@H�7�j���C/��5����&Mn-S�:�02��
K�"g���y<�=SC�7����q=q����a�ԡ�v��`sv��[JQ���u�=/ܑ�t��
,��H���',�mi}*�p�6�wX������=�k���o����!��п�Z���y塩��:��܉ k�9�{�lP#���Z�{�z�T�\����Zϫ�,�!�u�*���)�#�t�_v��h�>�#V��'0�%�I"9���M����S�����KZB��}Mm��˸�w���W"@�c�����c"�t���/�C�A�T�P�����n͹"�蘁X�(c�I��4�X�Ȳ�H=��M���_�<�\4����=s�Lh�������]����KF}������;A�5:o������B"Q�<>�!�2"M�O��WɓO(9/������}	�"3��F�_a�ʺX�󪼼�a�}~	�`Iye3Z��<�},<���Z4- E�Nj��`{G��� ��D/�G
g>���@f?x�LYt��T*zq�fg����G3�*]������{����[c�uä����<�k�X�/������Uq��2��y��������u���
r�n7"�y�E�D7��I��I:�6 s�(����2��:o�3��Lʱ����_�sˤ\Jr:���$&�}{+x�	r�hz,�_��'폘2G��`�a�k��c��{H�mR�rZa��(�hoo@�3��GqZ�� ��~ސ��EW�V�e�O7����'�E�=��ڷjݶ9\��w�2)6T��k��*}���d�!׻U�V��8�+8H"Cs��r�+�_uo>���2��<����p0]< � ���=�1	"r)�
(*�ms�r�
�/��x�	���ڜN���5i-i�w0�͍mC��goI��ُtM�I΃Y����SE�n_����g:V���z��PU����Z��������/)��E��e}��$�E"k@�"n�F���T�R�1z6P�����E�]��5�=#�g�Пȟ$�[/�1���8�{D�qr�MCo����a"U3V�u��qu]�U $j/̖-&�t�[~#����|���/f`�i!$f܊mjg|���<:C/�˿��KP^YɅA��zM3Ju(� n���
+�A��R�nW1�vdk6������]q�� ߙ��J�F6��;�4�w���y�"��ѓ0e/�
^��h�"up����L%܂/�v���֠Mկy��:Hb��I��(���os��˫�л9�b�����	5�2�� �!;A]o�%��]�Z��3�p��#�t�$���6�����;����U��;)�a�+.�ٱ��/�8��f>���nQuR8��o�0���㌊#-q��!�ӟ�|#Fnn-�r�7#UA���}�A/
��t�cؚڗ<) GMC�AW��5����F�s���2�!ɤ;�X�����H���ENU����I�����%O�[Z(L����c��O0������P�<���(�����7�[7p�9K��ﻺ��+�/��PL�R��69�S�DUœs���ē5�K�'��m���b9}G�_�`x��ƒ@��o챓%	F� ������T�����������9b�빴��(�qW��5�Lz�XV������W��
m�[��0��$�\Cw�\x��"N4�Y%r�&��h,��O��e��W��ڌ#m,���������ʙ����n�ad����nb�'�7�6��qHG�����	���P7v2S+�i8u��eD������78��%����ԛ�ޏ�+�����ǐ��E�II��')��y�"�.�.�+�!���[.V=�J�Z�a!��~�WiB�+�s�y��S��M]8�����j �������FgsǗ������EKw�]h�e+����3��\��zʝ���Up:QL�ͽ-7�dʼ�w	0�!����������q�Q�[��-rj�6����.m��(����U/��Ϊ�f�"9𥡻�H�7���KԸ�|�᳜�-�Gc��qk�5��������F���il�H�H� ��@?d&,f9���O��fO�n�m�V.ṲW�iE��mvl$���)!��<4�Q������t-q�i�-2�(���G˗|�'����T�1i��>w���G>{yO+\J4�ccV���1��HLA�B�������X�T�?�uP�o����&�T�L]��F�-��ĉZFǩ�~�y�4���k�Z���U�J$u�MJ�J����̀fI�7�ߠ�gE��'B�y��uWz�ڇ���o�F�*�0+�
Q�ޒ@�{��J����{Fi�@��`25��|������ǈ;��(P(����Lb������$UЛ�d�f�YvM��w �mg��=��h���&O��!
&�������'J�1�3�v��sI�A$�M��۞��� v#�����+t�d�!��3�G������{x�&qVs�TlR��T�<�z�j�}8�\!݆�^*�ؓ�i�S����2�D|3lR��Ta� �7O���k����c�_���c�,`lS�ʛ��W����R�M ������l�@)Iɴ���s��6�d9|kp��8U7Τy��9�g�Z�� �G����'�J]C08�������̚DV����gz^�֪���o�~@��'6�)N�ߝ&�-c
��)X�p��v�m�YLG�Q��:T�J洨A$�K��"õ�?�[�͌� ���?Y�l������W�K���gE8Ѕ��"Q�&-�@����Lj����8z�U����70ҳ"��i�27�7��zL�_1IN��#i�~M$�
9f�𘤎�P�h$�E#���߰G�̗��0�N|w	�.��l Җ��*8��������Ѿ[V��+<_��'�m4C������G����C{��X:��� ��!5�||�_Ϫ	��*�]~�#+��f�����+�fY4���ٽ �������wp�Ete�;��Wb�b��.Y��*|"3aVZJ�*��o�&��4u�9���* �
�ܿ�z����4WF����6�9	Pc����v����Y.������ø������ę�#�稐$���A{`������L7O�4xR�#f�k�|2-�K h|�!ϻ�A���U�[��U�?�÷l�ly�$��bA�	� y�ɟ ��$mQt�>����L�d�XT
%�ZB�3�	����AլRq"�5N\x�3S�\~� �T�6���]ib,M-�z߲��Zy
-�f)�
}7^H函r(I��o��ՠ���#��yA	�iq��R�X��x�AKL+Ib�+��q��ꎭkLL0ǉ���D���!-���W	�H$�WuA��9LJ�L8HG>5tm�_�]�,�}��<_߾�*r��	�Fn\+�p�E!�S�g�*���/N��qz&��_j���x��.��;��-Ú��3�����?M��Et`(�լ\3a�R���zT�����LU^c��723 �Q�X.s��~�>m���!_�H��Isܽ`��LǬ���z�1��1��0�'�n	��u)oD2��A�P�RV�`�����ۺ�ޮ����u�Vfx�\��'�뗓�}��Nk۝�=���w�=ݱ�t�b  �_ۘ��i��\Vqϓ�W����+���G���2xޝE����~�����*�>k4p��?��i��ٛCOfƬT?�-��0���6�3o� �+���6�ƛ�r ?ǃ�곸�G�z�s�Ԉ־���(n���1&r��󉹴���͘�u#�﹑�ا��H~�D욝$Ith.I�*�eX���1ɽN�4��d`LR-�Q�HG�����̏(8�8v�0�����	�0X�Wr=�%:��i�ps4?��R�	�I��GZ��ʬj�d��3�vK@���@=���S�������rv�w��]Nz��8��<�L��>�?Qc�ճ�ߦ�,2�p�Ma�$�k[0��r�Є����Y�Y���$m�F1G��1Nt��w�b���9�/9��N;��Zw����������bz{�Y:8UGp s�$)�+ی^9�hDH{Ӄ����	�^rj�<��Zt��!���>��E�An4��Mo�=�=��g�0�ǜ��*�M�:Ͷ�;O+����%�_x�LK��b���2�r�������Y�J%�����QE�Y%�8��x+R�f��nG#��]=X�V5睾��7��ڛIb��G�;#N�Zc��݁x�Wcu�κ�7/l/Ƭ���k�uU4���-�)��p��p���2�^཭w��v�,$qr��5o��j�62��o�(Y���}�M��z�f՞��W����KӞ�"·��f^��(��L��
~|���g����8~� �q��D��99���4U�Vq=o��U��И�⒇��ф�Ĕ��Y���hX�Q�zo�/��I�k`���[�4����*��[k���u��!�Ɠ��������  �_e�g�z�Y@��k��3������H�1�>����4Y&'��������wC�$�έk��}ى"B5� 1�\�}yh��x�ǸG��Q��(.eV���!di<ӷ�c��f�6���}v����	h��Pg����W�Kv8��������crZj�oٽ��_夔$+ſ��PK   ��'VA/R  �     jsons/user_defined.json���n�0�_��Y"��p󭰁"@kM�KaZ蔀#����0���u��K�I�|�9�s�l��=����}᧡���ߴ�*�@p�%�]և�l�s�Y���>����قb�t��fA1쎀F������"Q�:S�4�Fb�B`�Y���QL�R��M�`�t����o�&�󵶭��!?�����Pޔӊ���G��g�bX��},����¶gߪ�7g�XW�+��$�7��	ħ��Uz�_v$HE�` R�r�Pڏe��j(}��Y��>��x�V�~���~���4���.�1����%��6x
�|E[MU�f�޷/��3��K��(w���E�\p�[Yx�c�!��L)����,���W���	n��A����".�Bu�[�܂CD.��p�,g8e˶��o�rG��Zxr.ŵt<F�������[@E&Q�=�K�z��k�C-n���R���<�� �Ts�!/��=p� V�����B���:Hw;tT	O�Fa�pcm�.���OJӂ�\$:Hn��~9wܞ<�V��_PK
   ��'Vph�(  ��                  cirkitFile.jsonPK
   u�'Vׁ��( �' /             U  images/31de6c7e-4b9d-42ac-b555-28e4a5bb4aec.pngPK
   ]�'V�cŌ ~ �� /             �C images/40a6b5df-e714-4004-b865-d48720df955d.pngPK
   ��'VA/R  �               �� jsons/user_defined.jsonPK      <  A�   