PK   `TrU���V�#  �~    cirkitFile.json�a��8r��JJ�u�B� @η\��\U.��M]>�.%QkUfG�F�ލ��=hR�0�v��Uw^���G�VM �ϋ}��pۭv���u��mw��k�����S��Us��������}�����3��8��q(���_/w�O��-׭-6��*�[QѬ**��}��t��tfq�����H�`:3HLW��
���R�Y1�T�t��A�`:'f�*�΋�
�k�Rӵb�B�Q�@)��P)��$�b�@!�b�@!�b�@!�b�@!�b�@!�b�@!�b�@!�b�0����(�q�i��~{s�@�qw�ﷇߋ���p�&�å<�%`�*�å<�%�<�%E}���/w���kˡ���zݸ�V}U,��-Lk��m������Գ�1���p�D���p�D���p�D���p�D�M��_�D���]�D���]�D� <.���Jw��B>�K
y�K
/mU5r�U��p�H~U�����K�����N���?V�s �`��)�?V�s ���D� <?��X�ρX"P���B>�K
�PZ,(�Ci���jy�K
y�K
y�K
y�K
y�K
��<v���)���)���)���)�0���N�D���N�D����H"?51��� Q;}�)"�U��(�`099��Iw"�����t�+��+�t��8�W�����O&3T��{��Y(a�Bꂵ���JGX�0t�ڮ��JGX�0����am�#,��<�vk;(a�L�`m�`m�#,��Z��Z��t���u���58+����W����LЩ	87!prB�1<���ǫ���gX>��zf�������|�l?p���#0�!��q`��ǫ���gX>��}�������|�� l?p���#0��V���h|/�r*��58}�?��\����/X>���������|��l?p���#0o���`�������/X>���)�������|��l?p���#0oY���`��Ǜ����/X>��6A���	���|��l?p���#0o���`��ǛJ��C/�B���8�������|�{O!������_�>��~<:����/8}����l?p���#0�����`�������/X>��v��,8}���/�S ��m�;�,8��?Nb~p�c�����|\Cl?p���#0W ��M�O��Xp�c��/X>�q��������|\+l?p���#0W9���`����Y���/X>�qe��jp���#0����`����|���X>�q"�������|\A	l?p���#0�~��U�W������X>�q�-�������|\)l?p���#0�8��`����ٰ�s���G`>�+�8�����+���?�|�_f�yY����z����s�N�u�Y}�Y\��K�fv��<��>/V�]j_8��HL7�.����/�����_������/t�����B獎[��/���X����,������B�����/�������B��y��	�_t�Rn�@���z����}���r��7:&'���}��dr��7:�%��t+�с'�����|��2�+G'����rt�Gn�+G'j���rt�En�+G'G���_tZCn��E'$���_t*An��9��9i/�?'�?'�?'�?/�?/�?/�?/�?/�?/�?/}�$�?/�?/��F������5B�k��פ��U��C����.,�����-ʕ5�r����g�D_�=m}Ӷe_Ҧ�X�)lk]��K*��پ!��<��u����_Q���eaW��W�¯ͺ��8����_�]���}�w�]�������ϒ�8|����gq�z!B	��$d��"����H���$dx�C2<��!	�P����Qa�@B��0D !3N��B$.j��6,n,p���8b��n�o���+AL��M� �R2�*�	�	�QJf��1��xy��!c�,aq���q����AL�8^��8JɌS� &X/��� �`q���q���'��`q���q���Q��`q����QJf\�b���
�QJf\�b���
�QJf\�b���
�QJcBИ�����}�~�2��x5F�~ �;X��8�R2�',�[XG)�q}�	�L�P�-,���̸6���6G)�q��	�-l<�R2�=��,�װ8�R2�BB,�װ8�R2�Gnv7�	��5,���̸����5,���̸(����QJf\<b��q��)%�۳��Hu�P�`�3�`U���[��@�j��
����]� �=ʷ�+�e�[`^��
�WVRay��]��0�`%�0R�뼐�����(*v�8�X@��TXM7/yW�U��TXM7/�W�U��TXM7/�W�U��TXyM�Nb��q�В-�mֱ�R֥�v��]��x�F6C:��C�k�ul��}�В-��ױ�N�BK:���_Ƕ:Y�
-�����db*��C�{1tl����В-�)ѱ�NF�BK:��7FǶ:Y�
-������s�`fA'/;K0�N^V��e*��C�{�tl����В-�ӱ�N^�BK:��NǶ:y�
-���^>���e*��C�{ul����В-�Ա�N^�BK:��GTǶ:y�
-���^W���e*��C�{vu&�̗�В-�=ֱ�N^�BK:���ZǶ:y�
-���^p�*�VTZ����U:yY����В-��ױ�LG��Q��������U:y�
-��r����e*��C�5tl����В-׮б�N^�BK:�\�CŶV'/S�%Z�%�"6�Y���-Zi[�����e*��C˵]tl����В-רѱ��N2��d:y���ˬ�|�
-��r� ���e*��C˵�tl����В-�pұ�N^�BK:�\�JǶ:y�
-��rM-��:y�
-��rm0���e*��C�5�tl����В-�jӱ�N^�BK:�\sNǶ:y�
-��r�<�*U�P*󡓗�:yY����В-�2Ա�N^�BK:�\�QǶ:y�
-��rmI���e*��C�52Ul�t�2Zҡ�Z�:����ThI��k���V'/S���h3O�NT��TIԦ�TIT��TI���T�移3U��3Uխ3U��sO��T�g�d�$j>�z�y1ޛ:�5W㿩�Use0�:�4W�écBse0^�:�3W�1^�:�2W�ũ� se0^�:q1W�ũssu1^�:=0W4��x�t�^|�i�ƋS����`�8uD\�ƋS���`�8u�Y�hD��ũs�re�^<�`�+����Y�2/NC�+����aO�2/N��+�����E�2/N�+����!<�2/Nu�+��b��bz>��b��b��b��b��b��b��b��b��b��bz̆�b��b�����Ƌ�7/n0^ܼ�Ů�}��5ua��E�WmQ��i��]ݾ�<�"��i۲/iSl�����h�%v�lߐw�m^f�H�e��m���)���®<�T�¯ͺ��8���9.Q��<u�/�Lw�uw��0,�??���ǟ�v�?����|�'����h1HȌև���8c!	�q�B2�L�$d�Y9HȌ3|"��g!D !3�<B�@Bf��ĄH\�ƅmX�&X�F)�i�����(%3M#c�`�`�d�	n,�,����4��a����QJfZ�a�qpX/aq�d��&X/aq�d�U&X/aq�d��"&X/aq�d��,�t�+XG)�i��	�$�(�+XG)�i)�	�+XG)�i��	�+XG)�i��	�-,���̴0����QJfZ��a�=�=��q��(%3���0�⸅�q����b�`q���8J�L�1S?�8^��8J�L�,1L�8^��8J�L+@1L��M��&,�װ8�R2�BW,�װ8�R2�\,�;XG)�iq0�	�,������GuЪ�vv�*���
��hU�]5XI��tQ��*Ю���j��&ZhWVRay��]�rxh��
k��5*���+���1��]�2xh��
��xhU�]5XI��tQ�;�*Ю���j���ZhWVRa�5�:��NƥBK:���YǶJY�Rڥ�w�N�E:��
-���Zs��d_*��C�k�ul����В-��ױ�N�BK:���AǶ:��
-���^��dc*��C�{Jtl����В-�ѱ�NV�BK:���GgbA'/S�%Zޫ�c[��L��thyϕ�m�fĔ��t�R'/+u�2Zҡ�=p:����ThI������V'/S�%Zޓ�c[��L��thyo��mu�2Zҡ�=�:����ThI������V'/S�%Z޳��0I'/S�%Z�{�c[��L��thy��mu�2Zҡ��:�UZ���\Q'/�t�J'/S�%Zޛ�c[��L��th�ƀ�mu�2Zҡ�Z	:����ThI��k>��V'/S�%Z�]�c[��L��th���m�N^�BK:�\KDǶ:y�
-��rM���e*��C˵]tl����В-רѱ��N2��d:y���ˬN^�BK:�\3HǶ:y�
-��r�#���e*��C�5�tl����В-עұ�N^�BK:�\SKŶ�N^�BK:�\LǶ:y�
-��r�3���e*��C˵�tl����В-לӱ�N^�BK:�\;OǶJU>��|��e�N^V��e*��C˵ul����В-�dԱ�N^�BK:�\[RǶ:y�
-��r�L�:��L��th�֧�mu�2Zҡ嚥:����Th�2��S��n3U�i3U�d3Uu�3U��3U��3Uխ3U��sO���$j>�z�y1ޛ:�5W㿩�Use0�:�4W�écBse0^�:�3W�1^�:�2W�ũ� se0^�:q1W�ũssu1^�:=0W4��xq�X�\���˕�xqꈸ\��b˕�xq긳\Ј�ũs�re0^�:m+W�ũ3�r���N�ʕ�xq�|�\Pb�����E�2/N�+����!<�2/Nu�+��b��bz>��b��b��b��b��b��b��b��b��b��bz̆�b��b�����Ƌ�7/n0^ܼ�Ů�}��5ua��E�WmQ��i��]ݾ�<�"��i۲/iSl�����h�%v�lߐw�m^f�H�e��m���)���®<�T�¯ͺ��8���9.Q��<u�/W�?;t���n�m׿-�����v?�uo�հ�n����o%� � �X֋�WoE
F�}~w�<�l��E�&"�g�����D��.�~��F)��������
��S�8T
��|�g^�#�����u�߾�2k̋��?�ie8��R�F�<������~�e�k����sC���34��������m��
���G�o���������*�o�wFw��������M�as�o|�Rn�Mo�<���6�p�[a� I�7�|���'���:QW������O�)<��)黶��
��C%}�!w����ETa��W�����]ww�����w����a��o׋��^���$i6�%�8�'�K�q�PH!�0��*!�X{��b	3��R�%̸7LH!�0��2!�X{ӄb	3�mR�%̴7N��>� T�a��}R@%@�k�i���G	H�f��(� �RS���6YJ9 �tܥiN�T�� ����*�0ӶQ) ����*�0��U) ��;_gnk�X�h[��\�L[q��h[��\�L����h[F�r3mG�r �k�r3m��r �k�r3mɖr �i��r3m
���8! ����gX�m�M�3,/�_�r3�r ��_�����K9�_�_����\�L����k�Y����!H9 ���r3�c�� �i��r3��r �i��r3���r &�3Z�xZ�\�LU5��xZ�\�Lu=��x� �T�a��"R@<u�xk�WG��p	`T�Y�K1.N�w�����^,��NC�_��7�>>�b\�Ǐ����A��G`������u#��X>���~�y6�ϋ�#0_%���Y#��X>�.:������|������A��#0��cfpz�a��/��
b��Lȋ9�6�'%����w�A16D�"`B^D��!:�� �m��H���&���h��0!�	y�5چ��LHhB^4��!:;����m��P���&���h��0!�	OKN`�[GY�s�^�����R�Ӗ���		M�<�6D�-`BB����i��Є��mCt�&$4!o
B����		M�;��6D�-`BB��+��i��Є�smCt�&$4!�zC����		M�;���C��+`BB�nC��y
��Є�SmCt�&$4!��D�������T�<�B�)`BB��,��0��۫�
�ӖXjt�R��0!�	y�3چ�LHhBޑ��!:m�����m�N[���&��`Zt�&$4a\����2}�I�Y��K���ŀ		M���6Dg1`BBr����V��V�Y�Eg1=�&$4!��@����		M��A�6D�-`BBri��i��Є\�mCt�&$4!��۰F�-`BBr9��y
��Є\�mCt�&$4!�!B����		M�%��6D�)`BBr�'��[��{��yJ��Sjt�&$4!��B����		M�%��6D�)`BBr�3��y
��Є\�lC��S���&�2sh��0!�	�Dچ�<LH/f���K���9���'�=�R��Ƴ���4�*����ꦙ����ه�>_O?S.*
��]b���g|4\���C���r�N�+ u����\�'�gz�
�#����r���0�+ ���L�\�'Ƨ(���I=1>�(W@��-����϶��I3>c'W@��5�Rǌ����:f|K��x8)��%�.�j�DO���Rǌ����:f|�E���1�s$r���ܐ+ �����\�'Ƨ�
H=1> W@�N�N�dK=�I=�I=�I=�K=�K=�K=�K=�K=�K=ы��H=�K=�K=��zb#��Fꉍ��'6�x��j_��EiM]Xr}��U[�+k��@kW��=���3���mٗ�)6�m
�ZW4��
�v�o�;�6Ͻ�E�����+���z�,��s�j]��YW�gz��s�K�K�r�/W��~�uw�uA�nq�yq�,��.8��>?��p6������_���fl�-���%nLܚ�9q{��=J�Q��ܣ�%�(�G�=J�Qr��{Tܣ�Ո�=*�Qq��{Tܣ�����r�=��	����{X�a���5���G�=j�Q��{�ܣ�5������{8�ḇ�n��p��q�=<����s�=<���Ï���{x��p��{4ܣ��_����/�of�p�w��%Nw�.���O>w;��Ѐ�{��%t<�y�yձ�1Q)!:ʟ/��2�p$��[��6���W�#4/:!a%ܤ8ߩz)a+#��z�	)�d�yY�o��_7`�Ȳ����w�S�W|�TƗ�x��K��R_r�K.�䏗||�9^j�������r{��u7ۻ�"ú*|A�}?����f��߽v�qnY8*�OC;�E�6e���Wժt~�E�����n�ڼ91���������h��O�+w��� �y|�����?l�q����[���'X�����>�m����^-~�o��_?�6���6�-��}�}���?����?v�x7�����.o�����������0�-�����p���<m��d����� $%|3���.��mAƽ)m���^5�Ss2�B�Ekۍ�JW��Pm]R���}��5Q۴vI}�	��C�:��d�x����~��"xF�����f8���EY�o꫶1��?���}�@m���S=\��M��R=hփ�4���/�T��Q�zмGy�z�{�>�ɕ���M�����D�v���Nd|�B��Q�z���i�g�\[���B;��������׫D��&L�����+�/�Ns����B���+?`�T�3ߋ�+�f_���K\�M�Gi=JJ��R=��9��Gs7�zKfobn��s��l��[U�%�ʋ��y��5�_���.��&�W���hoη�����'�׉�6ѾL����w��BϹ;�:wg�V��l�ʜ'9���u�h��m�}�hO���|�㝍_���u��M�/��|{����1�n?����_���4\�7�Ƅ�t�������ʏ����@��]�?�߅�%�c���R�lK����騳)׾�uk�zSr��k6�fc���+W��OF�=̺d�YG�����=	�_`����׸��d�7�6��Ѯ�ʼ��������B��\[[���uS�a�.�����.�e�lCZ����i��b����ͮ�rf�����K��f��p��>��^�&�ݧ�G�~��ѻ��%���I�8ߤ镇+�y�o�Y����yj�*d���W͛����W��5o�2m�*���E�Y�E]�ˢ�{S���E��%�T/��q;�q<�������/�?~)$۪�c;��^��� `w���aL�����`��z����>mׇ�����>۟?pKט�/�6����:Ol�����_�@������>�G���[|~\�f���~��C�9�ϻ�ջG��������%��Qp�]���~�=j��O?��W��/����=����n{{��?|�>�{�n������/�4�^���o��9�>�䮶OGM���L���=k��˻ŗ��7��^����˟���g�/��W�&�.�6�f�I:ݵ�9{�g�B.����,��v�<���^hv����{�����$�����������Ƌ�����fU�_��\�.p��L�a=�d���W)��?���\���v��EߏT��iJ=��K|��>�NT���V��.u�=��B�:�lFYљZ�3���u&w�3�Z�<�zlվ���c���l����R�F�w��~�^Ś�*uy�/Ϭ��϶*�+Z%G��e���f�r<~t��������a�o�.d|�n�����������揻_�t~�c�����?PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   `TrU!T��-  R     jsons/user_defined.json��AO�0��
ʹ��6eko�]vBNhBM�K]R������qVƄ�Ip��ޗg����V�ށ}SP���	֡�Ԉ�8�Tq��RǊ����P�w5��%������a/�Y|7CE�$�R	��<V�P�T���4!e��\���8>��Zt�����*�m7e;�z�����[򵨗�6�80���ڦ�MC�1�3�R�[k��-��,�M�i�Ə��z�,���ơϹ*�q��|�,�D�=ݝ�ލ%�i̦���l.��u�������bo�����ҚG*Yӂ��xc����u܌_PK
   `TrU���V�#  �~                  cirkitFile.jsonPK
   1�_U���R�$  �/  /             �#  images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   `TrU!T��-  R               �H  jsons/user_defined.jsonPK      �   6J    