PK   �IgU����  �    cirkitFile.json�]]o�ƒ�+��4��I���� y�� Yd<A�TF��+˙d�߷���Xb��T��b$�]����bW�>-v���^nw}�G�{\o7����]��y�)�Z<�7�~[��k�/n>����_}����k�Φ�ge׉�U�*��hx[�ʾ����fU��-nn��G�dVs2*���Ւ́��j���/���~��u+V��]��7�Z��hc�z�ESI^���UȖ�������N��]Q��Q���p�ԵPڵ+�k����6�K��5���|��*�K2*�+2*����± ���N9�!���XP�,�C8�PM�p,�!��!z�$C8��I�p,術�����I�p,豓�X :���)豓�|�̂;=v�!z�$C8��I�p,豓�X�c��a����f}�<Q?l��z��3~D�m�߉pˎcٹ��w�;(;�e�ԏ����ʎcٱZb}'�����Xv�VX�)���8��5�w�;(;�e�j�����ʎcٱ�b}g�����Xv�.��+�����Xv����������Xv~<�9gX~�Ϗă���.��8�����3,?��g?���=K�8*׃3,??��.8I���`~~�
�I*p�� H�_\�U�4���,?������:X~��ϊ���w��8�������`�q0??�g=X~��ϡ���z��8�����=���Xg=<�"�����+.���.X~�ϯ�<ǂ�����*��������s���X~�ϯ,��`�q0?�&*e�1i�"�:�Ijp6C��z�7�k3/�x��L���sw��̏ט���KU��N�r�Bt�DqW�%E�r��s����̙��+*�ʙ�8��ɾ����'b��d�=QǓ�s��쩘kO��d�\{j<&�o����֗������k����D�OV�ϵ'j��}�˜�}IԾ�vF�ڗ��+��W�'���D�I��Q��?Eԟ�����SD�)��Q��?Eԟ&�O�����D�i��4Q��?Mԟ&�O�g��3D���Q��?C���3D���Q��?Kԟ%���g���D�Y��,Q��?K�_I�_I�_I�_I�_I�_�gKf;�FY�f�M_�BT�.�n�Usb$:�<���-��.LcE��]z���M�y���R'Ξd?{������hӆ��T�*�2�X�+�hNbm�<YI'��σ�/|���ow�����j�Y�@CD#�P�4�H�0?��t���B1�(��������R4F�Ȣ|
b���2�F ��(!(D�6.l��6�n�X��	�9(�r�X��	�9(�r�X��	�9,���ƒ� N�8.`q�4�Kq���qpX�8�B+�8�⸀�q�Xt�	�,���Ƃ� N�8.`q<�D/�GV#P���0��B�pT�_sp�Vw�x�x���\��18�G�5�iUH��w�Q�~��uZ1��]�pT�_sp�V��x�x7!��\��&18�eG�5�iJ��w�Q�~��uZ�����pT�_sp�V����$\�Z��>|��+�@�K<,ҷ�Ү<yפ�$��<�W���~���m��+�@�K<,ҷyR�,lU1�_�ZMvB�4,���<�ؤ�$�	yR�,l%1�H��Iǲ�����"}�'%��6PJ��m��,�@�M<,rf!O^��m�'��<yY���xX�o3M����&�1�H���˲�����"}�'/��6P���m��,�@9P<,ҷy�,l�B�H���˲����"}�'/��6Pb3~;������6%/�_�Y�=�,( %�^z~�А����p1a]ί�	�Y�;�^'Bu �b��vF-OLd���=0���g��D�`D��sF�O(cT۵rFa�о�3*|��V�Q�qQ�6M�Q���ŨXbT,A]	��%&KL,�K��%F��b�Q�¨XaT�@=b��F�
�b�Q�¨XaT�1*�k��5F��b�Q�ƨXcT�1*���F��b�Q���؀�'0*6��F��b�Q�Ũ�bTl1*�[��-F��b�Qq�Qq�Qq�Qq�Qq�Qq���S˩P^�O��U(�rI-�
@��
�K==��Z����Vj���l��G�z�[��}��H7��~�ܿ�w^R �X��4 �0�H!�@@cR#�X��4 �0�H!�@@cR#�X���\�"qQ�aq��7
� )�,vsX�F!= �p��o�(���N��aA��\��	�,�����b8��߸8,�XG!= �p��q��(���N�8.`q��\��	�,�ǐ HѨ�bd j� )�5P��
�k���Lv0�Q�~��5P����E4*Я9�
�B<0ٹ�F�5�@R�&�Ѩ@���(@
��d�"��\H!��VD����k� )����hT�_sp �x`�K�
�k����|��kZ�Ӈϓrea*@
�E�6Sڕ'��"}�'���6T���m��+�PR8,ҷyR�,lCH�H��Iò� ��"}�'��6T���m�t,�PR8,ҷyR�,lCH�H��I˲� ��"g��eY؆
��a��͓�ea*@
�E�6ӔX��lZ���m��,�PR8,ҷy�,lCH�H���˲� ��"}�'/��6T���m��,�PR8,ҷy�,lCH�H���˒؞Q���Y�}FR:Jd��H�(�5�g ��D���Q���Y[{NR F��M`� �`�uNR FñmC� D=��c�i�)@
���8���� ��c;0�)@
���XbT,1*���F��b�Q�ĨXbT,1*�+��F�
�b�cT�0*V+��F�
�b�Q�ƨXcT�1*֠��b�Q�ƨXcT�1*6��F��b�Q��O`Tl0*6��-F��b�Q�Ũ�bTl1*��a6��-F��������������U' ���z����Q^�\������|���Q^or�/(���?�t7w{��������W���]�X?�7˾�כz�������6t�^�U�6]єͪP�RE�UQv������U�n��/
|Tm׉e�,*gX(�ˢU��y[�f��J�������- �$�=�������_�ޅ�m�TU_��ˢQL��ꪶi�:<��$�B$&���0!���U	�O$��ԇ��t��]Ů\T�G�M�[�9k'�VV�X.;Q�ʶ+���ۼ�$��''�"���%O�b�K\�@Z�r*��^�br"$��1)#� �	����Ğ�d�U!o� k���7D��2[�o%0Rd8�QH�bA�I�E��{�-E!D'%�����Omeɖf�*n�	�I'�%��݇U�|=甴��KG�z����hg״��_{��Y׊���K:T�rR\�~![-��-�`���'�?��<��$kb09�sA�B|���P��8ʙ9��с���=
�����ș��ι���G�|�x��s�=����;.��>���G��<Fj������Ů������fӅ&2n�K�f���r��� � �pٙ:!��G��e�=��O �K��������1�Z�dB����Ր|�7�ߗ������N�]��-M���8�/z�(���j�4�8d�������F\�F��T����{����	��
Ļ�a��e9<D"D��;e�ڊ�����mJ�r��L ��j�};l���"�7�/��x�m�D��@����D�;��Nvs��V/͡�p���b:5n��~���pg���������o���� -�͚��!�G��](1h�s)����y���������R[ 	��[�[�������͸�2\:#�j\:#�\:��\�=��D,��+u����ug3�{C��c7�"����,�+Z���ޘ�ʮ�������k��2 -Y��)��Z�D"��}�<zd��G�(x3�of�k��![TM��v�x�z���y����c�p�{Zo��������oW���o�u���D�Y��AV"
�Y�!�P(�Ȃ��BkDd6jc�?�FJ�Ii�k�l�~�#�Ķb$�2tR��2���Ȃ����!� C��남A[�]9 ��1���GT����0���KT����Q�0���OT�X������� �S��t6~������� �S:����O ��1���aT�x* ���/0�� �S��S��o��X�d�1�Ͻ���`�a�q0?���'�����`~��`�I����8���
�?,?��j���ˏ��,���π������Xm���`�a�q0?V�`��`�a�q0?VW`�U`�a�q0??>��@�30C�f����>�g!�4��pt"�љ�!G3�.ӜL�RW����)a  ƥ����0C�fx�f��Ip�sR�
�&���@�-���r4C?È�!:w3�h�~v�Ct�f����.ڇ�̐��Yi�06:�3�h�~F�Ctf���j ���)�	t#�S*���r4C�
�Ct�f���
��s+`��Я~A����r4C�r�Ct�f����#��y
�!G3�n����w��[���6�� ��Og13��M��δ��e���h?Y;:{K�iA�.�G��^�%�7Y99�N �~�Rq�����s��d. U��ms���n��@��t+�\ �����#%U��u��7j��:���͔s�:��4�@��tm���!U���SI~�Su*�SR#��*QR�(�J�T%*�U���DE�]R���JTT%*�U���DMU��*QS���J�T%j�5U���DMU��*�P�h�J4T%�U���dS�h�J4T%�-U���DKU��*�R�h�J�T%Z�-U���Ē�Ē�Ē�Ē�Ē���9[2۱�0Z�B5��h���j��m�����8p���{���ԅi�(��K��M�y���R�Οd��I"O�?����eϳ�U�^]:��k�@KbY��q�$�Q�����֝�p� }���G`qs��#�~�ܓ����w���g���(*�fh�[rߔ���7�5�͹oϽ��[��[o1��j�o!����[Ho!���x�-����Bz�-��P�By�-�p�By�-��P�By�-����B{=\����B{�-��0��x�-��0��~��[��d����[Xoa����[�����z�-JoQz��[�ޢ�.H�y�N��Lg�����..�;'ħQ�~��W��v����&��N/F/�V^�4�<�up1�Y>a�)��u�'�x��EJO�1
;t��oqb������V�8���~�/��M��ᐜRχ���~>�����!>=Ğ1��m����z�����ǽwo�\
�J���t�cEū�XV�r�,[މ�6���z�K���j�_�)��͒36�����m)�b�Zg���d�?�1J���FQ���?��{]�e���I�P�/gvW���c��<�]�3س|U��7{���4|��n�����~��|x��_^���=�w����M����^-�h��_�:�¿��6kGx����~���Ϳ9����;�|�w����}���]�?O�]�-n���ȇf��n��i��Nx����\1���➵�~�u~��R^[}Ua�U��Ο��O�n�Է2R�E�;i�'\'��*+���r}�}�Y�6I=̫�v�v7��,�-׻�}�|o��v�Ju]���wW�RĎ�����بM��,j�E�J��8`���V�G��-�R�@����Ǫ��+���L���x2O%�D<��W%��+Mu�Иȅ�<npu�a����nhS27%>6>)�c�X�Xy�Μ��'��	;����RF����[ɸ��[ō
?$x����)6U��E����TD��hS�DD�OE���*��ؑ�ŎT1��Q��GWk���Ʊ�C�25�0�0(�PàC�24�0�0(�PàC�25e:2�0t���<�0tDDmT�&$�P���~�?��_�O�z�[�{����_�6�+�
���RV��\����4�I�_&l�����]�j�B�L�e�V���R�-�0�{�0$�1&$����M��G��˃����Au�R-���n�r�F�M��G(F�2%٨���U�vJɂ��9�o����,zնB�U�U��^$�(ߋ�������о���	b�c�m�3�y�a&
����	��6|̓~�f�������)�
��06�>��\���[>���{!Xu-�?|��s�P��r�yl��!���j����o_ǌ~����_��������z��������������ћn�z��z�p�`��e���Qf�~��fOX��㯯�+���}�^'�+� �>lכ�/��� ��ݻw?h�����a���zs������^}}��`;Ń�9�������w��NeoF0i�Q9�"R�2��l��D��+�����i9��z?�.,,i;�XX�t>et$ҘH$·X0{V;Ŏc���Y�R#���6�SW؈%1+"��v.I�D��ӑk�.,��������"O��&���F���;Wj�[�÷\kqV;!"��k��b�j��VB�k4�z%8a�%�Vھ�<��":zYN�$��r*���4���(�ݙ�Gw2ܡ>j,������+e�Ĭ7���4q�ɦH�Q$��i�ET�G����?�����ݺ��a���?���wo6O��߶~�����}^|�?PK   tFgU!�+�� �� /   images/0fc7fbbe-b47a-4373-9472-5e3944978531.png /@п�PNG

   IHDR  �  .   �TV   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��Wtk�y�������z܇�_�����}�mY��%˖JRU�#�f� 	f �9g�9��9��$�s�i��RU�T�v�'�U���sd�g�m�o�1��\3�9�ε �����%�w⑭pd?��b������>w�S�a��4̳9so�;a��fN�gO/���V�W����.7�.ח�6�q�t9�7?Z�9^�=Y�GX�|�/͜�Ξ�-^n.\l-\l�`h7;\�9^�=YK�͟n,�m-�o/�o/]l�������������n������������:��,#�������E�8��K�G�k��R�R"Cr��rl	�_����������������������z��u�t����.L�ǅ��ŝ��l�/�������_����_������7f���+'��G������s�-�SY����"G������B�p	���*�8i����&z݅�h��^bzo޳��_��$�;s0��l�p�����VW�o"=��!�"7�@hw~jg����ID�WB��mjwnjo�M�/��������ZԽw��|�	����.�'�B��yt/B��Klka�jȵŅ�� �B<�z��<��8w��t�=w�6{���;\AVe%81�5/O#�j��[��Tҽ=�ٙ��&|{s��Y�֌g+j] [�Jȴ4e��Y���S�9q�E�+a�Jdjc&�=�[��;W�HC�B�0�-��A�߱r�Ő�ok&���;�JxVC���g5��<1Ӝo,n��s�J.�K��� �j*`\�B�������R`b�7�pO.��"�Zg�潰�y/.4/L�8T��\[q�BΖ%��cl΅�c����}9�8�a0��@��B����E�h�9������	�@�24k��-�'W���aup#����W�#��9�Ȝi�gm�q�54��q�/�̫A�jи0,���ް�?f��i#mĨ�[�f��1so���3N�g"u�ĝ�Q2�ĭ��E5��mH��Q�`tr 2a���]����V(����[!C���ơ�itΪ�L�C��И>>���#�wN.:�V$���c&}d�/<��W�Gԁ!m`X��M��M��&��~��HopB�Є��m��F"����������x�0S��j/L��U��zC�*���������q0<>2�v�k b�zz%>�§�t
�\�+��r�J9��OX�=�svu�իW?����ͽ��~ȶb�̏��Es�D�xn@�����g���A�=1'�E����i����G���!�D{yq��쐚�#��;�VH���]���PoG|�ѳb����T3CVX�6����fFXA=;��M��c��>v��#��3;�Fe����������=�bN�[}JfP�ֳ��� ��� �����}��~o?��8��� /6ĉt%��s�CL���zU3��붱K���0�ϞF)vPK�嬀��gx�)uǴ�ï�zt%:��������?,�_5�W��!75��U�՝!����ѯj
�뽊��Vl �|�z��o���ɏڎȠb�*_2uF�[��z��-��qK�]���!���*���)#����Ժeuy�[Z뒠 d[�6���.�S�z�H�#�>e�[Q�%�|���~�%EԡΧB�*���#G*�VIsɩQ�C��k����>��z�U*��Kl<"e6a�STi��Uv�ֻ�!�]�Q��xOx��d�P=��a�]��+m���-�;ދSA�SP��.@�J;���Sa��R� 
����,�r�b�8e�Ny�G�dO��}ZA�
���)�ڄ)���q��-"��|DU�~MW����)ir˚<r�S\aᖚ{J��M�Z��9%.�C��NI����Abɮ@'P\�R;���-�p�L�E��UbRs���S`�.4� e��M(�r󍝹�N$��B\�`%V�-��%��4�$C��Na�CP�R�2Vd�9�8X`�ɷt���]�����)�v����E���iU%.�q���b'��#*s�=����ꕖ��I�*�b�GL��A�J�8�6N����K\�5G�Pܠ�d�r�]���Kw���g��[a�Uw��UEnU	�ɯq����f���փQ'���H��R��%D�-q=>�Y�[,��Ud�)w�J�{��=ٞ7�.���S�cd�P+ċ��B?�pC�{j喙zj�j�f�W[{(�ΊɎr��L�4i%�X��]icS�l$c���X�jaL47��%֎"k{���~JXag�9X��dW�z���)׭q'�	�?��xm/�8����:b��YysBњP��0DZf�)k�7�J�����..iLH��ژ�&¯�iabU�<��4�|��<����S��� �l�W�0(*
`���⠰p�+���{�|����"?V�V�dK�2���+*�r
}�</���ww�;:Kܼꐼ��éOW�������p���o��h�n��S���8�r�����-= ���(nN��;�����.r��]]od�gX��S��B[����v�9��g�g'챃Kwu�ۺ2��䈻뱫'����q3�݈�2�=YNN��_��e�;�8XO�i�\���|��<rt��2����N�M�w<�w�Ҭ�G�v������A>������l$Ns���7'��A䑣;��A>O=��i��t�s7g:�8:��;Z;��Ck�#+���0�2��\T殕C2���0��!C4�	k�ΰ�d��ԂeX;���]�*��j�;��o�xb�L� �~�ʸc�ߵ2�Y��m�Hp�B�A��g�@��M���6T>����ڕe�ɲtg��P"zy>�0ah�"y������<��A��eZ:2��O�m�Ṁ���F�mC2�kiC�w,mw̌;&&>�>�
%>�wݷ�3�<R7�"C��ɞ�co�emC	XX��9 ��-�LtD`w̭�M-(↙~�Ƽia��M� ���qt$���M'�]�����w��GN�]랻%�q��n�[���:�u�@�o�?�39����GN�O�'����u�b?ru��{zzy90D��]ș��1hS�{����{n6�&�:I�����x�n�	N![Tv�Ձ�8��сLR-�\ #��~�~�c u�$K%~����8�>�egް��t0�[�7,-�ۖV��[6�1y��Ї��t z�}s+�\h%�q�0�i�6�eX���o�P��23�M�l3=�D�1�!�ef���O,�t+������lmHS8I/1"�Ȱ���G.�3���p�ez��>f��Y��,�wUz�Z]"�| �åmdת�H�b�Ƅ�iNk�W�"�	�n^NK�kfE�d�s5Ƨ���1uF@�	��"J�W�*r��=�!^q�_��%AA����
B��0� (��a9Ӝܩ�lW��'#Ѓ0e�ޞ'��?7��I�w?�u��ُ����^�
7�MF�Q�϶log��X�����R�E�b?'�ە��Og��{��?�2�]�� 5�ޞ���q��[�j�x��Нw����Q��L���\ cЃ48�Jv�Ɇ�qu�rt���`�c���;�6Y"��lDn��nX7l����o����}WW�\���9uӆĬ6b�`>��-r���5��ߴ0o�ۮ(V�����L@�8�m{� |���:p�Re��(�#[T>	2&��GA6�us3&��\/[�!�:�Q7�@LW�v�ݵv��.�C�����MV/U���zLT�y���&6���Vpv��
K����嚹嚱�#kAUɅ�l��%�ե�H�O�33�O�{��wM���P��{�H������$U)����צ\r݆���^DR��T�с>�ݹ�`�oo{��@�����b��`�`T��v��:�i
�`�}q�;��꺓��j��f�v����uw�q�a�H���q��u��q���@���%XL�oj�� �U%��!R���0�#�#U�V�OE�	�l-�;��Z��s�]�����[߳4�om�nk}�JG���v��o�B�~e��Ԉ��--7���~���6�˳�s���&f��YbcQ�l����A"���6V���e��6�{k�����屹)��{bg<v�=r�=r3�܌Ǟ6X����m�� �"0�ê��^�,l�C{fET�7�˚UM��y�aQ	4ׂ�s��y	5!��	�f���A匨<&���&,��Kcܒ(�(����$�#��?'��q���T���sBܬ鞬inF��x�'-�MB?����-������˾�c����v �:�<�&���?����C$o������� ��e�l��3��~���A�B�@�@t@ �<?ț�m�dt�	[���	�[�N��ޞ{�nL�[�ND��:��\ru�"�9�SV� Cd��I���.��������m[ۯ��w�k�v���x\x�w�I�FP�q�5;)ߵ��߱�^���ka ��q*y��B>���D̓w�-�����y�#!��8���B��Z��\�I2�@@'����R�J5�T/Ue�mjFx�D�ݰ�î��V�Ms;,��.����!�$4Iрr���NR���16��|{�E�~ml�!B.�_;'b��Į[�%�`����������pi8*cf %Bp���@�!tN�+`p1�v��� :
�%yw�]~}�X���������ĭ:7��=H�.���a�=����w}]�]��\���p3oy�!
b&�%0M�Se���-]b�w��7=��C�=�'!b�ɾ��F�Dyx;����b��ɹ�J�dp��,����:��k��wm-o�[~mkE31���n+�]1!��� ��3	�-��67�'���h����o���Nv��U`j����:�L������r�v;Z9.B����je����{3��Zhk�0ӞX��G��G��GA���!�����nM:��@�إ� z"�J�At��;�43!m\R5,ʡ����m^R5'�̉*B�8�fA��bVT>#L�qQI�_��A��0�p~T����ؓi,+$�
�eX�4�Ag����=�Fgx8"?�w��u=�w�8Oo��?�2|�)Ki�7��ϰ4W�cWV��=(���H%��J)²��Ɛ}\;�	)V"��pӝם��#�IP�.��@�#����c��@0(@�;�w,m�4�mg��h��$�&3���8�4Sq��m31Bg+I�K�������W`���.��f=�dnm�)$Ce޶�ej�G��Z�-��I��͊R��b�%�UC��)��1�8�Cdaa�U|��Ȅ@69�a ����n�fµI�0��(�@-2a��a(�]K[�8�Kj���&��w'���������W��Ik&�2}_�Ԃ��__�����/'��~��
��5Q�&�E���'��B��N���07����KJD�]��A{1B���X�7�dT`�`H��l����6 �f�����btJ�&I���������Gl�1��y�p�; ��-Ej0���S��}�l����[�.p���!,U��.���I��{I�L�$`�S��G[Py��љ4�Nv�@����7� �a� �T�7J�}�<0�,Hij�>Ⳮ�):��X�kS�;ƺk��Ʀ;���M�RGg����l�7�,4��Zo�qV\U�.�	��L���.��AUX)=��V�j���ҭ���\�w]-�ܭ����4/=�C�v�b��b�{X���z'�5���~0r`�G��z��`,H!�9��Q:�
A��0zV #gE	1��q�(.,�	�#��(77̅pΏ�������9؝ᦃ���!AF�{<�sS�9-���(L4�� :/,N��	��p��n����{H�z^��ߓ7��$�a���6��b�"������&�&<r���7�H���Թ�e� ;��B�<	t�a f��tR�I�ޑ���1N�B�A2�H��P8�[
�8��R9#������嚓�@!8A�@�PH��$+��df@�)Ij�%8�`���=�������,iQ�h�k�'�Ւ���K�GH�%q
D��f�V��Ե��w@RCs�w�e����@-�l�/�Ϳ04"���i(D���	��@G���IYFd�zm��c�͠> �{�vBg#���w�)ʃ���=�7���@�
��BO�#�]I��ȻV���!�����x���@m
�dt9���.��X���@�k.&_s������u|D�h&n ar��Lij!]�p�aH��R�75�QV�� :�^'5>ư�E�|RX��UH����;��&��B5C;�At�Lg�
﹈@I��Hw��ޱ4�L� d������ޝl ��[�-m՞n���ig�l-:[㈵�h���j=�:���o����~;��q۫�*��:�Һk8��{�єki|b'���h�x�tDyZ�LW;}��4�)�v �4[��'��q���ڙP� hQ휬nAQ�@�5�-H!�V�K���	�g�eγ����rNR<# ��)��.��H��(�t�X�LN��Ί�2��'Ӽ�)>�{����>%x�c�N���d��O�\⏧�����q@p�������C{�`?�N�C;4��ɽ�$�S��pLx8)j�����a�<=8����l��d�Hc��$L�$�v\�w�R�9���=;)eyDr�wL�%��g�C*�w��!9�)���fH�9�D}��0���o^Db�#8�4�t�}o�K����u;�Ad�R�2I\yI�KT|j���|��4?t��8:���P�$�SZ��p	D�d&&�m#q	�)���VJ8��E'�m $}k`^���h&2����>���_OBw�S�}�Ќ�)�P�"�ߚh�AX������2g��S�������w�����T�)d�SI��E�-nz8e4]G"�;�Q�I@���
��+p\N*k�������?�p	1��,��d4���ԭ����!o���{:��;��Հh@q8�VT�P��D��r����Js���۞n�t�g��P ���l�!Cᯅ�j/
"��=�q�������\m�5�[��!���Ɇ{�m����,���-�1k����9Ѡjavh{ͺ��:=�:��o��'Q]8 �8X.G��^mvV��*�ܴ.Ci����ђak}hk}�hI�=r��܌G����j��xY�ގ"�f�X~����˿5&�� ��;΋����d���N��	eN@�΄ԯ�3�,*�à��f��QAAL��g�9YQ�2t��e���g>,������ 5��>�}_�=7;h0 ~����Ay&��&i�ꁏ{��M_0��[yR���G����������{ȣ�'v�C������"� |`g���]����'nnv@������\<P	�Sw��,��y� v��u����Ņ�wrp
�~��JUu�nۻ`7l�k&&P��uK�K�m+��'�׍��災���<�"��`�s�]����}S;�hc#��f�M+vǁ��eJ�%LL �"<J*eP	쀓�)�o���1�Ӝ��֞Fv�Kx�ԅ��I���P���n�:�4�
�Bõ8����u�N�q!�����Q:ѧ&X�vݷ�]�[��[�-#.a]7�u�׌,�E.1 =8�DY�5�=�P��0�	%'��;Ng�b�׾5N �kSGޙ��g�#%�w�[vq|��~�6���8�M�C�O4�(Ǒ�	Ưƛ~5�x}���H�{�M�&�M(Y�^��lTr�KV�Kq#pqS`p`���Dr;��߯� n�g$H-� ���y�:��O"5�|S�B^O7B��67�'�B1و K��F��#��K��זڹJ�%�&��j�������+�z�*�A�m�׺��b�V�!J��D�$���H>�@X�=7[�/�����nlx��KA9�������ߝl�1����Z��n�r�,�
KØ���b��j/O�_}��껧�^}��է�^��ի�%����ի��~q��2��4	p��f���f�w���vWS���mmN����)��sB3�ݞ�m����:;Ͼ|�=���l��¼�(��Ӓ"t�����Йlq��d`t�,?��A�<#��67���G��a�gNF�l:�E��InH��%eq���87(̞��IF{{�|�t/��{�{m�ĸ��̩�|*��� ���8:���ߠ��Ѭ�%(v
�{O��;�������B���/.�
�\|򪙃�����n%��	�*��%>I锬|JY��y��A�[��z%8X1�*t�˼
괶2�.p��\Bd���zD����GV�CK�CK�}���}�������ԝf�d��H�i�ɳ
*�*�P��8���D�Gfn�C���e��\\K24u���Ol����i6.�A�������G |�c�ݷ�ܝd�۹O�=OL=96A�GQ`f���&^��瑹E �{�N��А'�#cw�K��$-��X�M�Hs���=�D}��N�o��ߜ`�7ue8�7�.���.y�U����xh�<0q��o��I�=c�E���י���a��o���c�?چS�ǘ�?�|g���D�{H6�D!rC�wƙw'��X�=�2�ݞ`��P7.�����6R�h���{�1:�m���`Í�#�8�x���d�S^�	.����;��ƅ�"G৓n�쾽�k�ڻ�n�=4>��&>	~�����°RAH���1Iޭ����=��&��$Y�9{p0��M�|�Kn��I�	y-I�lM7��c��g�t��
��غP%�{8Z|$ͱt�5��hH�����}��;��in�;�:��X�Uւ��Z9��s*������f���d�/'��16]74?23)����gi�&�s���d�ի�$��ūW_�z��o�{�ͫW_�z�X�m2��_|�-����;9=���f�18��nZ������sП�dK�єz��΄��
|��Ms>�~s���nOC\(h�.]B���2jBBl^�2ʜ$��!Jm=�͉!����b��9yj�0M�
�E���Y��!�\���*+��҈�((.I���� �//�/�I�������su�u����ᰤ���Y��9��<H
j�l0=cJ����CC���8��%_&y� ��}��H�߱���ֵLk�=�T���iM㔺5ܛ�����9�����g��b��!Vt�#6L��3��0	��1D��X����+:��1����0IV����5~Mʹ���*k�tT���)���"����ؑ�#6^�ѵEGi>Msx�֯��j���і�P�WW��E&rh�5���}�r���&ʳ��m�
���-G)�b���%�!Rd���H�ZU���+b�,���!fh�έ��5^5ͧ��J�97��*79��8�evI�$��)+tHK�J�5�z���ŭ���k���X�륹5unm�����k����.G�VY�M�J�2�����QV8eT�g�̢R�4�$,���|X�Q�c����ϝ�g�w��u#��<�5�P��	N�I��_��&A�M\j�"C\���a�U�k���0\�̋��=�͜��4tfzr&�,<��Fr$k��Te�,�?�"�c+��ae.Y�M��ENQ�S���a�KX���$y^�K
\���ы�8(�!}�GZ��Q�[V����C
���nq�OA�RU5���6����TTY�O^�&/���J���%!�8�J|�J�
<�B�V����%�Nq�C�k��� ��+q��D�<�r�FƒKR�"\�[���.ɲp )��ݙVBX�����qA�`�	�c�D�ߚl��d��-����6Խ?єfl�tt��;�����w@��Y"�fp~�駟���Cq��i2؜6����o?��՗�~���w�}G�^���_��lX|.��^;�
�r=-�.F��剳�~줃��Π����w�͋I@����m`gR����j�Pfũp\9GYar�Y :#^�$����taTX#R��G!�E�1QNT�&�&������C����"�.�*��E~~`Z���N��=p���;����߿��$k|�򣻋��}�����Ý>�cwu�Q#N���7��~o���i��9Oa{����Q���i�Eؠ���1���46��5��c��gZ�5����9�"n��L���A1kV��tKv͂U�`W-�`�9B��]��T&,H�P��͚�F���)͒ݒS5gW�#�J�f�I�E�jޡ��*���M�����E�vɣ[B�Fd���ػ�%Ⴋo�ӿ��[��.�1�*��Z	��.���vͼK=�Dq(9�8JGG�	�)��y�z��*+U�"U�s�*Cr���g�}�Ӟ���]����z�ޣM�����.{t�T��[�8*��Q���V��K�w`98�Z��W�e�~�˾�?�X���ʸ9�W�(�"s$���P�y'
J]2��C�$�ճ6t�-�[��$1:!���?ڎ�͚D�	��	&�!T�M�Y��ͻ�JW�Xa��v�.��R�� ����Q�,b��[t	+�B�cF��&1��r��	3F"�Y/2"������aټI�`�/�E���i�h�(�3+m0ټE�d�]u�F7��}�eO�w`czp'ܿ5�������p�$[�n�7|x��M�!�O� �ȏ��c��IŬQ�0!�~ͣYu�W��u�b��]��ۊ�W��YO�jhh+2�Ҭx	�D2l�%+��5�rщ���l*�(N5�>wK�i|�'���ĳF�̤0n@��L�	&^|�qJ�a�~�����j�gC�?�����4�|�����;Z�`�Iqv����}F����o�����o�������J��n��'noe�W7�R����&�c�x��w����|��ǯ����w�/_}��g�����btU�{j:���V0t~⤧��nf��-'�G��E ����ʇ�,�Ny7Ҙ�1#�k��5��]9C��(��&D�`q\�$��<LI�9	hIAD�凅��aA�47g�@�� �հ��2�^���=O���)I�O���e�9yA�c�Y��eD��w���k���>v�q��d��ܥE����%�S�C���P�0>g�M�͘�bƱy�q�1�KX����a}dbd�<1o�!�Pl�$�[��y'l|�a^�M.y�-��K��9�aэ�3��Y3�L%C8��ć㖡�� ���Ȭ���s4a�q|D&����ŀu����iً<a�	�q�g^L̹�f|���s�|c�Α�}tƁ��^�8K����(rN�q��4"���9#Q��̹mK�q�#�.x'���i��P̬L�D\�����������Qd{�4�5&ܸ||�65��H�}S\�l�ƒ��XFc���ǜ1�x�o[J�6V-sqì2�����v�PԊp8fK}��OO��Q�p�2�6�8P
�!l bđ�Y�X�6w�qDl�	�D�b�����9f�H`�q��-H�!�I�P�;>5<�����c�!#�$n���1Z�汘i$jT���a���	�F"�����?a�hhb4jDbӬm<�<5����1�:��Q2�H<8�Sxt��Ab�A�AEe���ߧ��cH��8�p04I�u�E�}�P�1r��Z�I�6h�}С�#�q l
YC���q04�����1��e�M� ��V1s�4��N��f��X��{	C":���z�U�6�OYG"��٢�#���d_xR��N���z��q���Ѩc4�H�h��3�vL���C�Xҷ᱑����(���a�>��bF�ؿ�l��D�����q����_M��|��õ���o.sv5�]c��&��^ ���@���K�ծT�y<�����t0X�-e��Yiy�2K3�2
ٴ����������ӫ˓����o���ի�}�xTk��T���p�d��N�s�;�����9S�>Z��7&�1I댴nNY�P���Y Z���T�H���y�3��8�D&F��D� tQXT!V����!A�� (*
�ˢ򊨪<�̛��AI�����ex�����I~��<��98�A��O���zh�zl�Nwr�a����Nv�@j�����</z���&O�@3���϶ز3��D]rDV���Ԃ#��Z�{��E�3��/��s�?y�?o�^rp�+��E����48���#�%���gjѝ�܉��Zq�����5ou-:�K.ς�=�0c�G��.�g�8��ۼN�H
]�x=�9�c��Yp�<�y7�@J�sxV� W�8�2rՂݑ0�P��͕��<��θ�v�Q��Egh�Mz �
��;*��ֳ���O���O.�,m.�g<S�\;�`s�'zf�Θע�9;z�9k��&=�o��w����ŀw>��X?:���,�=s^4�=�B���p�eK؝	�3a��X:�,��c֊S�"ל���gͦ�>g��`�d�M�<	�kƀ���tb	*曳!�=Nj��ML��⣖�'ap��|�q��,��f&}�Fgt�����������C=��Y㓸e��-<a����C��;6b�"∎�ã��#6�S����ؘ%:j�##���5<�wƆq	��w���(�4�o
������>�B�=npD'���@"��D���u+{���v��k�;+����͕����B�s�#fTՀ�P[E�8b����a��OML��0���䳸��rt�~z�yz�~|�vt�rp��b�������#�D��ϸpbz�05h���B#��0:"��R48�,�Ɩ㞨��p�F��!Ot��Y��\�Aolh*6�7�GY^M����������?o ��i��#uo���j����s{���>Z��h?<��z�	��_|���j�fä�hr9lf���� ��.�D���똜�W(�ҳ��+�?9}���G`�׿�����/?��/>;���6{㸃"��4Xj�mM�NF�����ȷ�I�A/v���i#�G�mx<��⨴%.���kfd5	9��t��rV�t���k:ϊ�o�I�f��Q��Q����!��e�e(hp9�_���sqHR��D�>~~H��<q����iq�O���e��9^~����ړ�x��vN��<(�s��1�#�v����,�������}?�T���en�ci��|��F�A��\�Kueʲ�[��~�Ges�-N�ݣv�����R�ڤ�.����+Ɯ�!�rȦ��F\�A�rܭq*G]�����7���^��)'��q����69�:�F� �3�F�՛D� �[7d��vB����"�Y2�dհS��}_�]5����y�U�g��԰S3`S�Z��Do��Ze:���*G���v��o�ZUcm�Q1`R�Uf�ޠ4kt12����N�H�vR��Q�t��&2lV�[����o\:lR��	a�Q�㈇����gY���?�8�z~zv�����MLH������ӏ�2ݸD;&֍�T�͸P3.�7�t�j��L�!����<{�z:5�L(d��8_:&��Gxj�Le�*��O2�QL��C=�a�p�[:����X]�,�=��}L�po��?����IFY��|�S>ܥ�QsT�<�P�l�K:�V�tˆ�DLAC4�҉�*����n�����A�j���T1�#�ʑ�@�t�C4����x�S��F���n$V0���Z\;L�+�YJ��`�P�d���k����!�|�M1H��*�0D`�A�t��A� ]9�R���BT[9��W�,���O../���|���g/O���=}q��C>"�����"\��nT��&��������ˇْA�x�K=*�F}+[{'''��Γ�\����ˏ�}�����/�/�OO�w6�g�Ö>� W<Ёn���QE}h��_�Z989� �?܋��'���c���A[3�TѵC��Ѷ��v�G>��m6p2�wƚ1����?������F�l|g���$��袏7�F�6�����_��G�I�J������1F�+s����g����A��O%��s��}-ՕY����!�@8=�=y����?�����}��o�V�9+�,�z{C��!��:9��]����;�f�
��
�%t��6.�H���긴j��\'_,��Ĉ�}���4!!��I:�(`���y�¨87��J~C� (�������{�{8�=D%��@g�9�.n��[��z��)E�_V5��U�%.qU@E��hAuuPU���ڹ����F���{`�obݳw�����ϲ�Y��vOW?n�����쾉�~c�����R�ub�F��N�x��n���F��C�]���f>�s�X �|�OP2ʓ�H�:E�L�0�7H���GX±.�A ��:�g��bp�D��I!�"�v��``
2g��tл�Z�&zc=�ԡC0�-6p8#�dM�`�m���6}k�Wh�l�l����y�q��P6"���LzŰ�����3P������;�q�p�	���eC"K���L�}xТ�񄃝����&T�{�7r.���]�\<=<:������~�t�!k�K�y�IՀ���<0`Ԍ�%� nWO?�4�X�`�o�Mo��g'��tO�s��5��d�&�m�L�������Go�mA�g��{���f�m��&MM����K��� l�n�i�մ���:I��:Q�|L��)FD�A ޡkB'0�5���v}-K_��G���4��ă���.b�#�E0�"��0��&��������١e�����ټ�t���=	�V����[߃~�6q�ڸ�,A'����׊>g�ľ��^[_׍B��;��ݚj��N8Ј�=��8�rG[��Tz�@3�eLY����/^~��ً��Ƚ8��?9�;>C����Ջ�H�<M���r���*��5�6u4��������L�$��>9<��Bΰ��/Ⴡc�����/>x��G}��~x�����Abs��m�ј�4Գ��������r��[{���g��-�/�{�dCM|=��[����i��:�`�b���Ȗ[��!f����і!t�������P��us�����`��o�N�|��c����#�L=68��`��UK���QMwg���N���-�o�D�.�'�~��j�ak3ګ{��n;��V��lɲ6d�sl-0 ���6�&�����> ��4��115*��%qqqT��rA��=��g�Ku tɌ�0&+�+c�¨4����rQDP������!�E�S r�7yF���$/�_D�we:z�<�
��fZUT75uS�Ɛ��S�����/����~I��Our+���_�Q��r����+t� �R���+�u�9���z����S캎��P�2�í��6�8��RO��
�;�[2��3D�:��`7��=�2�#�F[�[�k�{�lq[`�o�YZ�D7g���W����`tt�'Ľ��$��o�@R��7�*�����D`d�50�ԫ����v�m��9���O=C�W0���t}}soC[_[�0WeW+m���6�@c������Է���}4�`=���;[�Q�q���l/,�cź�N8�&	�R_K�@���U_C��#ʚNWbk��;���'�[';�Ǜ�ȠS�i}K� ��� ���ζ/���10�{Z{�;��}(q�d{�h{�xg�`ݿ0=�����YhN�0�5D��Ńk'�G�Owώ�!�����Z�kj��C�q���N�X�[k�gt�p���^W�`�O�m��Ъ�UڊJ]%���H�������U��u��&]#n�Ʈ�D-3�sK�3����U6.��e�jk���ު&}5����A�R�� Ě�5���z8cn?^���3u�p]������>�Ω�NZ�fs�8�������~�B1���1��C�����7��ŭr���h�|K/)���f��{����}�W��V����[s_M��
�ӢoD�9g��.�e����������������������6"��{x��srz	R�>}�� 9@ƿ�����ii�:j���}�������m�m�qq�N����ήH�'�;���;GG��G(��v~yy���^~x����Ɂc�ӡg��ju���3�o�\���]П^^-n�C%��6u�;�U���5,�W_ե�
���c�BSe��x��W�-?j��H�?���H ���w��������u���Ͼ8{��+TC���[�}�~�P�����~����mwc��/��x�^}��n�4׏�+e��zG}D��!��)@��Z�-��Q�� �o�"�+�#Bj\T9#)���Y���|mD. �c��("��4e�	,/,�G�%ab������.�J�f�+H��G^�(@3,�G��ӝ�7H-�JhS�=�� �����2�*VTɎ*:#� �5���aLW�T3��>��BN\�5�cFt�HoӴ�!���� �e�ן�����n!,�Ï��V�P3<6�^8�?��L�m/�m�j'E��Fo#8�W�����o1 1��z�-��f=�=";������K{[kG{ӛ�ۑ� �.s��I�Ԣg�L�����ӽ���!w?�nkoC���3*r/���Ov7�w����-p��$l�kj�7���m�����z·��� �V]S���="5��3�zoo���JC��R�k����P���i�e�z��������Ӄ�3�Ǘ�Ǘ���+{˶��7ԃY���3{;��������������+LԳg�ؗG'��+����om�c0�<�l�{@��.onzb�vu�	|z��v�v�Nɣ�+�P���f6��F5]�
n6�53���Dx����9=��M35]�ZF=*r��67�C�ZM3E[_����1�����::6��4�n�4W��%��buy���HU�H����������64���B�����ë��WgϮ�/�g�ֈ���դ�G������il��D`~gy�tw��p��h�|y�?��:t��2FBSoK��s,dA��gG�'�Fҟ⒝�ݥ�e{��xbk�͓����ë����eǌ���Q��䯮�U�k)���f�QS֠.mP��i�k5����M%EUN�������-:��&�3�|xz�����\Xp�c�P`b�k	��8H0}p�M}v���'D�b�%x���z�PC��F�m���1���;����s�d�Ww�g��C����յ���������ӳ���gg��}�A����LtwP__�?=�?;
����giSa�R�%�j����Qz�����IV��.�����Ɵ����ڟ��t����A_��Ps��A���m�~����>�L���Wղ�Z����f����3�ϾI���}v��Mj����^Sj��0�=�6�ۚ2�M�VF��k0���x��(h Z�6F����4*,����� � /�ˋ�a@s�幢)yU#&΋����iA^HT>C�qNYqHR��rw�u2o���gPl̻6y���.R�*����4�h�؀rP���5;�M--ƆVc�XK��b��&�`�qj*l�������Vf�����tOK�#��������_d����e��}���;�ecMg?Y���{�f9��ˇ�[���?�ݪ����������݋�����F�g맬���ã�����ftm}y�h��p�xM��mT��i��t���������g��3��Av����횈8v�/w�/��N��NwN�6���&)$a3���w}q��t������y�\Voo\�X�����n��lZ���BSU���LWS�TЊ��cr̉������S-�y��Ow�N1K!�.�=�>�����-�z��ZU=��]�[?:�>>�8:�88�<<�9<Œ����l�`El�7�Z���l=�s�TX�'K�[�)G���{�k�{�w�/�\��TVǻ���t�J�(DG5�v� �~�sz�[���TUcT�^]\>"Ϧ����eM���X���\=C�3�N���@S��.��T�����jJ�����X�ۮ�g�I}/�����ί�..V�6'�F �JM��Զ���}��ݕ�s��t���F���b����e�;Үc��k]���������W/�%?8�z~|�����ۿ8'v~	K?�|��u~���4�Z�t�XTk)�:J��<eU����{��tU���Ue���Z�����f�OA�g 4(	a;��>�vti%�JN��M���:ɘ�Y]]��_�?���6��F]��į�W#l�k@5z��s�����O��2��������{6��fiDZ�x��p���p	�> NT�����~`=��W��*Օ�:uwH]_��fTǅ}�Q���Y[�ʠAK�.����ҡ��4��\u��!�������o�h����Cu �?���j*��(�p���C`q&6ˢ��[A�ke~6p���?ώ�/R_i������-�Z�趱�3-�H{diH���@k<#������L�kC��$���¨8h��#�5y+#��t���0?=�͘�C;�ԄaIT.ֹ��'ޞ���������l6�!W;�����ζsʽ�����7�h�[��������h1{��3^̛(OV�'*$��P�4����U��*�E:^��	F�9cE�B�h}���\�p���?dq�*� ��fwt�$����a�Ӱ�c�i-�f��̹<�xxȂA��VU��o�;�߃@x�����6�k�5*�Q�kea��de�pfm���O��s;���ۦ����XC*�����f)&�����s����i�+K�����������B������4]ɔ:��Ӯ��C0�<�yvp~��;S�	8d�qt�XT:te-�m���PM-PU���P���1�wei��r��s	���Fbcku��	�W���=ל�E�\����2���] ���܎.��Vp����!V����';��d��Ѩ�ѥ�C��g�66'��6g�k����#�y}g�knc�h ���R�g�_�hj�M���<>�-�Z~���6j�[k'�ǧ��U�ES&�+S4�&dӛk[��] z|sIhP��h���Uy��4[K�RS���
Z�����[�����OQ����gik���X;:m�qG����
E��1�t��BӐf����m�EX�`�c�����:]n��l�]�wpJ��(L� ����)��'8��:�����Ydc�5��@�T�k�+�dg�����V����і��U�u=�XU��,/Q�P4-"�>����D��O���9�����:q��^�j�**���
Yc��]�2O//�o�-l�'�w|Kb��FۈUE�� }�Iی�`t��EC SKt���R$M�j:E�X%G����b,��"���?^����$z�
�5G�!yt}�(��0���ݽ>�X���FUASWҴ�ae���YW��[�1T��g�jn�7�?�������������ڟ���6��7�(+�S߼��|$�J��,��e{yq!~��o<�����UO����/���淟�<]�*�xi��2w�汥ት>�ڐki��{�c��_,�MYVG��y�A!�܈�R��I�Lv6 h����{��B���D�rIX�7%ș&/�exi�G.����em���|��<q�����>ae@�V��J֔��ƨ�n��U�	��Zk'h���A3}���	K�3��&�N�4����X�=;s��2h�׌W����c%��J� M8X۪�������Gō���dF�\Q�q��a�4�׶����Mt���V֏vaOw�ҵ8�y~q��%�ѳ�O/�qo����3���A�-l�zfc�5C#���Ŷ���1����VM��fJ�cJ�)�e������������Θ �啩ŕ����������ފ|L��+�s3d���*���ӓ�����Z�tzi�5�+�U���T�Ќ�ڪ"�HYU��sM}ӛ�'(�tew'��q[�=����:@y|v|�e���n���vԁ�(V`+Y%�H�tldrz:���vp`��K�]���4V��� ���ך�kK['g�ݻ�ӥ���¼-<�ﰌ|Xml���\��z����V�M�\����!YI����Za��U���lo�\l�-���ҦRY�ڇ��gW�p�'�s[j�H��&SEISU<T�=R�?��?�Uf�kkt������3@茮,��|�������Vlsӻ:��7�wV����0=�<�
�¥y��eS��[;���z�����2���ٝ��h�����͍��R|u}e� ,>B�S(ܓ��������.9����Y�d���r-�XYLC,�*˱**US�t��:Z��"WY�+�,��+<�s{�)/{qu��ً�ӓ��u�F�HQҰ�(SW��iŊ�bYc��-�N�q��s!1�u�I�U�Rm%���BS��M����������Txw�=?Ӧ���\uM���\S[�n����M�0��\_��q7�d5�
$�ѵ�F�3[�gg)@�ca�����\M��\Y
τ�Y�.�1+�9��[�-�M[�������qo��j�~��zK[�3ь̅���|vy	E��.��`}kwc����vL�g�<��f3oo�'E��Ͽx��<n05ت{��b-	�F(��Ǣ6�/h��pw�_��D�����sBɟ%o4��ȏHr��5���#�c���t��q���ũ�L�p���l�Y~!���ޝ���EuAQ����\�2^�2���Surs�!�8����O���ٗO������ۈ���"����߼��w_^~��Ʌ�ug �3غ�����CP������g2�����J/�e��m�hF����Q�Ҭ��l����0bnc�
����_^�?{����_���^�^�<��eh�Ճ#,��4�V�ֹ]����������{&8�����(����gO���.������@4�����E��-���u����KH�̜�aZB�����c�jYs�����d�(�j* ����Y�Ʒ� �̮/��}�RV��k�����b��.�7$mTs��~8���s�g�\���S+��*X��`ha��E���%�Aߨ���P� 4&3 =��*-���yt�ts�hfuEk��S�mu�n�����k��V��Lk��QϷ��,�n�W��܋�F%�H�&�"�;�����g(5K�2�1���sz���I|sMb��פ�����ez�}]����4�Ev��p�7:>���zk�u2��m6'�D\峂�%r:}H�uz~xvU���kM14�ziXGS�x��ķc(x�^�q�`|n�+��i������(���DWV�,�1��x;"<�q{
� �;�W��(�T)J��eX�JJ����<eI��$GQ��,͑WH�%��ٝM�LF��ųgϞ>�}r�O�
�T�Tu}���HQ�'��+j
e�e�֦>۠n���
$���"eE���B�:���C�'�3��ե�Qe��>_^���櫪
���*���T�岦��yv�=���&���1��S�AH�o���9����&:����������A�d-ĸ�Z���h(�F��2����.��R�j�G�+��RU����#]��h�?�P�VE����kmU�����:#�/���믿�I�*�xe�d� �~���B�`��ߑ�����}�B��*-�OL-�֖kK�����9��3���h�4��of󓿵O,�aQ)]��0��eM�I���"�e���s����,�+�pr`i���v��M	�\Uƺ��*��7A�L��YY���������}��g��o��H3��|O�������1?�����{@���U?���DF��,�=����
���㠱��A_[�o�i�=����Gd��H�M#�jy���Y��˻;��)��M��Q�-�o}2,�X;���1o����ã�{�>�.���ζ%�o�u�H����"���������~du����>$Kȝ��z��J�@V{G��[k���Rq&a���1OW����5u�
��=9���uz�yxY�e�:j%-URg�?���A���$R1tJ��<�3(훋0T�&���Fթu9���v�Z�^�h����Xh�lq@7�{�;���Z�W�.!�7�z���Lڌ�����)����C�|�5��*�#����1|����s>ޤ��"�$ �vx���x�;���[ nՔ��>��;>�<<�m�
'{s$���2����! �@II��i����c�O���;[*�H��Q"e�H����^Q���%l,���]c�����K�S�i���5WK��d-5b��ϳvp���������|�ZfcqBn�)��_������D�V�ȑ�As�9�g\�G�\�Z�^X�����g�7���rY#=��b-h&��VjJ�U�9�lyQ����+���J,S6��(p���/���`��xvwY�m��T�JEs���HV[$o��Η��ks$��ҚC��d��XYS)cL�Lm�^��Wv���NxD$�z��+sT�d���.�PU�5���ϙj��k��bF��*CJ�V+TU�������:|	 ���O��P-��TQ+Օ���2MettoUmm�h�5�-u5��7j
 ��G��++��k�G*E�_}����H {�/�Ώ�������o����G����}����9�櫯���7�<�3Ef)�B>�Z�	�s,Я���򃣕��uu��ϩ�o���)K��,+$Ή�3����럦�%_�gO�����$�����2=�,7/�+̰wg;z
��</�F�+��I�5ԍ��*y���e����/?=��;d�6���)�c���ԫW�[Xw�1��o������F�B[�O��w�9�j
V��>�BM/��R�1�X�;��<�|F�\^���ˋ��s֒�#ٺ��_w6!k����"���j����!V�W�6�H��sc�`}{ok�p���{�bl��E��V}��^"������D ���:�o����涶���o�&�:�N��bk�aY���Ɇ������Vcb�i�T�M�.��;8@� ���2g�G��Pd���X+l����֚�<�=8���Z%�P���bRU�j-�7VȘC�S�G��I9���5�5*��Q �(�3������j Р3Rb6���{ƨ�rYK���]Z �1]���+�r�X1V �&����_><��h���ˣs�X� ҙg}|z���yh8R��I|cClꃂ~��x�,��(�#-��)+3d���X�E�R01��ƙPKr��Y��i,[Q�)�-Q0ua���. ��\��R$�2IM��5�l���i'��G��9�V�ͮ�������1����Z%n�����mxG��2S�W-ho�J����z�l%@������e��a�U檊r�%�ʲl�\�./�'.�5���CS���J<>9;?���z�E޳^=�X�[��/Xb�a�y<��y'�z��ͅ��|��6	�,U�����KZu�I ��7��ĨpB_ ��V��|��\-��Ud�_Q���#��E��s�ْ�L-]F�BzY�°,�7�{d�Z�,%���P�E��}�2�DM)�P+�U��2Myu/���R��j~���P^�C��R��P^�c%�NC�@}�������_~u�ry��`g������믢�gr>9�xz����׿���g���������X��'��ͭ��2���8�v�-+#���jZP�n��qrO�RhND
@�F% tƴ��d&�9��;-.����y~aᴄD�Bp�8 .�K<�27�t�tP'�[&�=F�t���\-}����������?��D⯾��u$e�����}��'����y�ڏ�G���K����^G����碼����r-��[M�Qt�mC��}8�l�m�Wϯ^���z��ttr�|tx�v�B������Ƽ¢��Ұ�,U7V�9#��
>#O��>>���ѥ免m�������t�pfmAc�Rҡk��8�����s�L5���ˋ���I��QУ�[�.q
��0P������XY������TP0%
��х�
U�v��7���Ѯa�� ���;%��ٝ :���pqw�0NR�N�t��hvg���Ҕ��a�ouy���P�k�;#nk�T`HĖ��ӇXϭ�ė7���$����Z;ܵ��jE N�\>>�?'��_0�[*j�Wgi4�л��� �f��\(h~����gkG��a���*������Q ���戨�eeOT����ir�YE�������48���tp���c�	V��yb�����z�@Z��/o(S��#^ w��W�v���*I}���E���»��꿼�70T�� �����ΦȤ-7�J��C�bbe���Z�TaE�y�����`��5���HV_��+�d�y��$�K�Y��9�t�s����Q��-�[">���up�W������O���6�Q����ճ=�z\��ѷ�id���|"/�R2SI�M�U4۳2��X�A�����na]�'��PR���Lua���X^�DQ����t�����8���K�%�jj���P^KS�-���Ã��p��$��D���ɪ��bUe���HC)�Ua�PJ���D�o�-.�G9�oUU?�T�5����C-��:���هW_��T ����ˏ.�/..����?�@�Ϟ?����_~�������?��7M�����ZkC���a!�m��#��G�-�)��h��[5M��v�4�vN���O6����gC_Gɻ�O\ :3 �v��������L7��'ε��9ηw�{xu��:[}���}��;�4�Vm�-}I��!{����~��o�@�������R42��L�!�/��Cq�������O��W_}��W�|��]V\����&��/<�?f4������BU��0�:�RK�쭩��V��:z�����&���%H�sp����������2�����tZÎU[��V����h��m�=�����
:C�.mo9��!���Kll�!��ã����is�6OB%KBy=���/4����$�i�'��˂Ae�������$�t��5����k�ՙ��Lym���DՀ�j���%�*�4���{�{��I{u�z�1���i�sk��h���@�XU'�#��5��8��΀!0ڟk���8�JO>�:��Ao���	'f�-��'���Y-m,�@1�NP᫫���a���Z8�?�"������b���!�fȩY��j-߻�����T�"��"tLĶ�7���99��^��U�
�we)�" �Q<���qrE5�e�O���*tE�����*]J˓��B������k.ڪ��r$Յ�F�sн��T8Z��E���4����c�}|ꙍ4+ص�v����>�ݚ�\Z��,4�h�qtBlk�{B��}���P\��L,$�2V����j	�L��y�����OV������IE��w��L����ʢ'��4I�.��b���Jn���9��̆c����{X��@%_v>��k��={v��W�8xz�|��و5���*��Dg��1�s���}P:���q�|~~@�l��}9�呢"MU�H^�X^�t.G}�����8��@VFLZr_R�#�*�4ɬ�K{[d7����|��U,��)ʒ+�v
0M^]W�U��蚡�'j�O%���u�UT؏U�?U���o���q�O?�����ᡉ_~����]�Ç����|����}��������	Uk-��6f�Z3LMY��|sk��k,�E�����~����ϡN�B��� :k��X�9qFH :��=М��y��N2:Z�� �9>a��a��[��zE�s�����E��i�율��C���|��$������6��%�w_|qzx�9MF���$�d�k�z	_�as=BW,�`���N�}ivnok{g�����f���e�����������k�ߒܖ���t��
at���L���'�,/.�ס6w�f_7���A{4�����		�s�;��`�KDU�
j��"WQ](��]�����C��������4\'���'w��-$����� +� ��܏e����|A�����l�h�9ڋ�δ�:J���^P�sF����d�BAM��*CQ��nj�}#���$)��櫪��Ò�������/�>v|~�����G����} J֞��ʚ�2�|bv�`e������|��s���<d;�:���3�������! ��k{��Ս!�Gg��W�v�S�����/�>}Y��Y�݁�,�7=�T<�Uf�h5:�osm��d��d~o[�5���( @�an��ά���7�� ��ٍ,�s���ՏpE�a}�&��td�i�FZ������8��V���F�Y"{+[�g{WgK�ێ�p�����8"�X�}�o����#��������}��l���Q�#�{�!�]8�Z��4L�,��J���ѳ;�c1W��Q$j�M;gvw1��w��1����K�>�����0@� ��d� 4"�j�g3�5�ʺqc��]n����K��E��}��PI4�0�)dO_~p�����.oR]*o�S�$�ODq6���kL�� }v~	<���7�q0[JKSR�+���y1��,#:Z]{��U<VV>$�ޗ�ޕ�ޑ�ܑߓ����qC/X��::#�j�=;N�HJ ����(��.Ԕ�jS�.��P�uu�T5�(�����꪿�T�����Ҋ�WT=h�P׉�{�^^|��e�a���ǿ��8[^��^��S�`�ŋ���' 4�狗������G��D&UKy��	�9��FД�v�� ����j3��J�-�L	
"�� /#�͎�"��A��� ;*NҦ������Q��$��*{ZF'���>vq98�N~�OB�(~]�]3Y�:Q�3ޢw�v/ֿ~��w�Kf������K,(�?}����������d�	�LF�������ޥW��Y��Z!����*c��%�Q�X�限+�\ހ\�sx��������1����~���[*�~L����S=���T��%�{� Xg�k��c
Mu���\��7�n�-l��m���eO��F��Z�_�#�.�n��v���PF�UP��yʪ\Y#}L�X^�oA������|װ�2qGۀ&��1��\Mԩ��U�2�x$KHYM���V/�m�.�Ce;�|aC���n@��^?"�����S�.5SR�PJI��5L�<{�g�s����8U]���(P� ^F���ӧ'�d�sR���K�
�lnl��g8��2�Bک	8�76�v�� ��=��p>:
0�3m'�n��VKۋ��iwx{oi��]�ݟ^^V�BN��oz}+���#dB��#�WP�h������kP�	ͫ�> ���u}�����������1(�;���F��~)�G���-������:����
k|nz��p�����c#\"mN��I[��S�����j�Z�wMFv���ρ-h���#�|%��	�k+�wQd@�����9�#\����76�C���F�e������8:^;؟����Bi�n���@Z/sL��$vw��F����bi�2`�nma,�67%��|1���j(
��,.���e�@3hR�#e9�,��9GV��+e�Da�r����Zbc���~�_�^^]<{	�N-�����>f��5�VS����Z\�^�9=C�B7O���z']Z�PUyOY~WQvWF��PV&�7/�ѥ�:/�(�-*�#.�-)�)*�-+�#O>���`AS$m�u+�[��@?���DN˕�g�J�/�窊
5�%��
m9 ]�[[J���򯕔�TT����Cy����,�@Aɫ����. ��!������/��O�^����� ���?����~yv����>���~�ы����D��\QcnȘlN�lα���c#��kvO�f7=�MS���<@��>M���#WZ��H��L��x��u��}���p�R��U���ָoe?���]�7��ϣy�)�x%��d
?��
��4�w����㓍�͕���xbH?(K�|!������ ����{wo?�x����A+.m�V5���rsYjSA~kA����qON�lP���������jk_��G�NI����x��������������(�������=��(PU�i�*�UXd����&�D�mqaju���&5�b��;_�$�Oz���[[��%�]W.�B>�*���<u}���g��/�7w �綶,� ME/�ց�qMtogq� 
�>7U�h��"C�7e%8�X^�%j��]��]@*�1'�i
ŵ�2��Ӿ����;��	q�������H�$	;"��g�d`k���IޠRV��n���%�"�����H�:/��F�W���a]���H��2�FgBޕ���Vl}cfs�X�%�A ߼8�_�����t��ry�lqK��϶��ؙ�܉nlXf�t��X���ѱ�{a.��
�-��@�#�m�y�g՞�a�ciu�������j�o��BAÁ%�����ǵ�����!���݃��=\�����j��7�Lj�����̳��L��剸ꉤ�yX��\�?>\8�_��{��"��� ��֦�g�6��X@yhs̅.^�?\I������BK�M��:Uw��V�f�Ƨ���~bgӽ�J��BJ��*G]�/��:'C���M�Do��A�+k�8�<kˑ�m�1��/GR�� ��0"��8�,����"�9MUvWRp_V ����e��ك��X�\,��Ղ>�Cm7������=�������ӽ����RK_O����h%pU���B´&Bɝb�z�:9ֻLE���
�3���-}�,���S�D<�`��@s2qE
�X�K)\#�M��8	�/�E���lyY��8SQ@穋�5%e��2Me���'r�k@+*�ZV���ҿ�V���ʫz��_�����s��P�Ϟ]MO���m�gG��������ߞ�?{���O>�������'�$��*S����F�0��Zi�|��CB � M61`4���F��o�7�L�Ո����t��oB~;�����J�u�:�)�n���z��u��7�ᜱ���߼��5��������h�0���)O@�7�6v����մK�k�h-M�LF[���΂ɹ<YwwWcC[U�i��{:o}r�/~���?`���ԛ���_��_��C�I?�'���U�\U�sA�ey>�sou��|�a���DƔ�M!Wۀ|̑R�>���/bH����X�S�j-�S�ՀK�f����,a#M#�$Sk����L��g�k�i-�j0s5�6Mjg()�����
p*MY�XR[$���ؗ�\�&���T�.��H�t!�g}#���X�6��3�d�ﾼ������ww�vf��}k�\�*_QQ_(k�����{����p�0@ap}y<�V�
u�2j��:OV�0(h���]��Dh�5�]ݞ]ߝY���`�����d�j�UL��f\X�/,L�FĎ�BIs��.K^�!���QM:��e�N�f-32�8U݅�y��>MM{�����"��4�tm�&�AF�F�Do6��T�6��Z�X��[�&F�X��9���[�Z\	������q�D_.��>.s�,�����;����>�Ca�I�cA}�mȾ8��G�{���3�������?E�~(���i�}�Xн�\ۈ�m����:"(�=7'4����3�L8TY��1�X\�K��ꧬ���,)%G[qZ� g��ˮ�Ů	u��*MZ�XZS����\˫Εe�e(MX?��3������Ӕ����в"�����W	�H��hhX�,eu��6W^���/i�6�r��Q�|�x������|e��r�h�87�cՖhZ@g0:OQ[&aN���ΐ�6�L�K�R��-+�!�����e~)�E�`4�AF#IYrK�4i�-qa���X�"���\\�����k�*6V�P6
2}0������uI����\u�m9�G����PU�_�%))��������յ��v_��󳃽C��wi~�믿}�������������?"П�卓��yq<��0���%��4c�#c�csS���b�=��]?x�tq{ڻa���˼�5�c��@OҺ��"���)@��t�t�o8;ȿ�u��?ɷ�!��:�=>��\9^�4TrǛ���O������[�W_~�ч/W��6�i�(HZ�+��;�l�����TW/�b�����_������������@�0���y]l��-�]{����������w:���h����Q����X��כ~o���"Us� �~����H>��d�+t�mӀ�H��Y�XZ�K�bJ�hKk
m"�Q?��Y�k2e����5Ž,ŔE7e�{K%Mي׏_�|K��{��ҪG�IU���JW>�{"�Ս�9�	�y�Ӥ�W=���/e�(ō,ǈq)�\^��@+�t0"KN =��n.���V	���0τq�M���ق*��Ieeda.���Aޖ�ۊ���cz�c$��;y=UށE�)���#qU���1���k����z,��u�(�K�OD�O��G=���bIG���ơ=�ܗT�ST�QT�V�ޒ�ݓUeI[��v���e�U�l{�/��`�)�=g,Z��.-N��8��}�qa�Ba��Y�C.�s��d�
j�ۚ�յ��X�/�]X_�ߖ�S��-4_㱏����~����7hx%"z�����⮔��_�/e2G�r�Y�q�ã�oDj���<z��-] �T�HAy$���;�'f�#�)Ƅ4S\�XZ
��������1\�b>Uܗ�ޓT<T5��5!�:�n�<����I�%w9dEQ�E0�p�nJ
o� �;R �<SW��$7"]�z�Q=K�V��O�ds�"�w.��w�wtz��Ք��m�y��`���ש���bI��>8<����b;k�Q9�
�@ߒ<��a�Z���%P$P���� ��e(j�Ko�K��
n�oI�PB�}�>M~]k��dj}�Z�,Rץ�K�!��M��U�E�b �@W{SN�����+U�_H�����$�|[Y]>�֬f��CA�'�o��o_}���Bop�϶gO/�ɧ�~��'�~���{zr��ųgώ�A�$�k��p���D�S�}#��J�D��8 ���4' �xY�΁n燾�i"����R����㦋4��d]���j~3��o�S���rr+���&u��h��vW���W_ ���o_}���/�m�,Ǣa��>>4&K�[������Hk����|brI2�ÿo��d֓����o����O���d"���������?�����ϖ�?:���5���������t�28T�Ŧ<U9�´��#�dJ�3d�ry��2�,9+2U�O$���j��:③�<��Zi&�c,� E�-E��	`T�z��HQ�&�I�bnc��irHf��S{|)��H(wE�{B�]a�!�쾜�X^}�
�@|Bv̜�[��LE3���e��؏�i��2x�bݶ�X8:�/�i��bAm���P�D�s�z;�ĵY�*,�A��)+|"+!�HJ�!�x"�H�S�u9|Z��[�&�<�$��+�Q��P\/�)�&,K�z���ʃ�J
��["R�[���b�	���ꖤ���t�����,��%+�#�(дu��mE��.�_�X��#)(Wֈk�5�Q��ҧ�Tst����Z+,����*�+$�nA��$]PR"oa5j�E�3T�;�p�o�oʊnJJ _�{��Ǽ�,a}���r�[~�[r�_|CPrCRr[^�����ϣ�	��hxU���R�^(k�V?B�k��r��'�x �dH(zN���[�S��XFƃ������YQ���[vWZ�@P��ddH�$�7y�$�����U��D8�^(��|�oI�Њb(S��yW^4�Ȑ� &�5�yX�I+��ԛ��e���'�n�׾�w M�3u|����9(+7Bn�P��l��I�7/���}v���g��țp��n��B�+K)!���*���&���ˠ�2�zr�5(-�-)�))�Q�\Ml�_?�;>!��cI��A�`r�<& �t���|]�{�r �/��E��e���HQ�O�ʼ��^�������K�q���W_=��8:�j�����E飓�����?�aϟ>��o����|���VV�.Ο=}v~r�jtH����*�Ps�P��������Z<�Nmq\],n��Ʈ ��ۓ��J�	��z���� @��t����f��d���9�me���������{6v��W�V�����q*��X�|������I���o��">�q|L)�hJ�D!�pU��y��'�����'�}����n�x�ѿ���p��4o0�G?��?���k�w�T�DU�q��i��l$ y�)�e���2�̴��2��ROf�f���?9��H�� F����䁼�}(����M�C�;t����<�]�*
X��o�y�}U�e�}i�yHf݄rQ#�Z�d��D���KR�ꆸ�����s�r_�z	�mq�{my��Ŀ���K)O���.���
�փF�
 u�Ț@���&.���Z����@9)^�U�@^��$�##s8u���䎲LA�ޓ��+)�&)�����({_^zSQ~S����gߗA���>PrJ��EY��\YV�<��,hP��e�mbJ���U��+8ʒNU>S�ߤ(�SU��
%YY��,i��#�ĩ��)~O���8�]qλ�<J�������즨�]A�5a�u�@"��� ����Gϧ ƥ��i���S��X��n��DTJ��g�쾴���P�4���衢�>����.�W�c݁CE�q�p�E�7�� 5��uq�I�=Y�}i.��IՌ;��E97D��%�d�cMx(�*׳���I<]�G&��������E����'<�hrxa{��D�7�֏V���\�Z���RVc��e��6<���z�0���G�
�p��R�ۚ��d�k�� g)�L�>1?�t�7��b]�VxF�������=���h̗�E�'����[���rIk����bh/�]��|C�DU
���zWX�W܂�*+�S�����G���W<�k�T�b�HX-Q膾��(��~�������;��?������g�?}������x�o��oj�3ўL�ޞ��cl�glz8�T0�6�Y?���Yܞ��:|�2_On����&��y|�{��[��n�uW�5�]gۻ6:�3�=;�]+�};놕y��|b���LU���Q���鷿}M�o����O6�Q�w��_-��&�E<>���Ngxݞ׺���p���d��u��R���~���~CG�1���������������)K~*/�^V��*��i:1���z���E�n�1�=)�L!�&.y���,�l|@'�EJ?PU�SPY�(df��E�6Y�d'C���l�WQ��=Y�;��w% �uY�{�B��	��,K��!C�eI&�u��𠛴�4� =�a�PN�7L��N�#;��u�J�ei�i	��&�jKrq]F�
d�YE��4>���v�YZ0�М�JRyT���fɋS�yߗ�+�G�ޖ�ޕ��#-MZ10���P�^W� ��$D�"x�G��LY^�<�D�AU�7k�غ|��P�[��[��-�����4�<ioO�ۮ�iTeQ���Ҍiv��������䎀��p��wD٨R�v �d偾�����]������$��e��KIO�����䥱;b�	��;���w,��Ȯ+0�;rKV �+/�-ͻ�(��,DwaT�h$�7�!-La�}� E$��8��4��<L�@� K���8羲�=a6���&_Ʃ��:6�f�WOw�����}�2-E��S)��=�\T�D@����������������p�e^�Ȃ�Y�*x ,������탭䏈�\�_���.��q�%�dX��%O4��ee��V#g{W�O��^>;|v�qq;�QLOb��ހЅ��Ѩ{�%_��/N���2AS��<����G-#ߙ$/۩+�u�d�CZ�#a	 �W���T��9TԿSW�XVqMS��i��	�f%<Q��d����W/��k��q��� zksg���峋��ŅI�xs��Qbl|����� ����t�5��~pv�5���NХ��� '3�{��<L����纫t��q0޶ӯٓ���:_�-�&�CkG��[am������>���t~�����lgk%5h��@����l�KD�����7�/�e�7 ������g0��k?�7���ﳟ(��AQ�3q �X]��*~� �J�i��T����ጢ��Dy�ȿ�9�Q�J)jCQ�	���(&$Z��|�N��B$���R� ��Ia �L '+���8{+)���42�o�r1o�����W���.G��se��չ���s5X*�>���.��hᲜ�����a���ȪSYR2\G��I�fI�R��ǽ�h,���|'+��7ń�҂_K�ߕ� ʰ_�ߖ�\���//��*�hp�=2x��4yn�"/G�](ϬQg�j3�u�쑡B�`�k��7V+��;F�����y��<�>�I�IU��rr�i��tM�mi:\�&ɽ&�~G���,�����3 7EV�(�=Q ���A�'5~)��PS�|ge���0|�%�������Q��TA��J��������1�� -�^�n(�}q>�р�4����Í �H�W :�g�t������@*{,��r�O�l�^<;F�q>~v9��:��T6�ɫ3��4��<�_��������'�_C=>]�?��\3-��u���+�<q��>]'�F���\]�\�8�BTU[��:]VE����(k�5������9�z�Ջ�/����GB*�	�+lP�&V�!��w|y�\���
%�l�q~��౴8S^���(%��@��ԕ�6ޑV�D\�ײ��QS h(��*��k%����RTe�1*��+1�PĨ�O�������Ͽ�8>x���^C{���+@����Օ��}�5͓�u��+�h���w��o�軓��ME#m�q`������u�}��{����O�;v�I ��-oWj[�;	!�_��¸fm�i�x��v���uu��X��궱&�K����Ѻ�߷��������	�<144�)�b�9��N�o+�?��Oa4�SCߋ��{�������8����Ҳ�Ք����L5Ysa����@�..!�Vuy�.%hK�9!R�5Z2Mr�+�(�kF�%mҰ8��sLi�RP�F�0�++���ބ���a�B1Ag�l|8rGYJ&�� �뙏�қJR
�����2�5L�f(��;49�2L�״��A�ʨ<K�p��ݲ�b�ɕy��r��'�J4������^����[C6��vN�E�t@U>�\~K��+I�/�y��##F��)WD�&G��:�Ȳ�T9m�@��7�k-
MR�5�Ɔ]s��x��p��ez��1T4ڟ�(���m��(�
�����G@�8��� ���=q�5Q�k�%���K��	�n�S�Ûrr��+ ���"�y�d��T�!l�]�Ǒ	�XO(Ic�w� e� �C�ݒ�ݐ� �uy�])R���Pɛ�۲�;�\�&K���׼��?�EUSn�Y�qUӘԻ��qL~���?��G/���m�fy=WS�DL)7H�C����m�+�L~K�`zuU���qsd��%�XT���v�l,��C~���R�ٳg�����J�Z�l��K�MT�I�5�3-�n�>}z��9����������*sL�&�J.)��Ĵ�^��� }I�Q�ӕ�-��K���+�$%���ByU��V�i��6�jk4�Z�#9��R���(?����31 �od�+)��������qFC���:�%"o���kO�>��w���_�����������hy=�m��JLM�'�n�oN�ޝl��.k�N������8���3=��{�Λ.vJ;� M����`]���gg�gc�gfܰ�߱��ݔ ��T�<F�uo^m}�m���~:�.$��*��46G��]ݸ$��3��F������.���E��B���~�_�P@�g*K���s����K��"�h�]
�ݗ�?��� ��:St�R�N*�R��OU~O]�4\R�#P#�\h:"눊, �IMZ�=Xr���HRw$����� QsI4���Y��u.���Z��6[X�DX��B��z�A�l��P�� �T��"KE0��cy�Ei�������+�!h)�W�HM���I�������uq��wąI�\����]y��YQ��O )��yA�"?_�]�W����s�r�#E1C��(mq�nJ\��Es���������h��X��P�D��PeRE��UN�2��<�oJA�<���e��㸺|�yݿ�~��{Ϝ�p�Ď�Y��j���(5U�����Y���bF�1�N��ڻ����<gfΙ3S��ru������?{���E������楚J8�C�m(Vi3��B�s0<`m�jIY�r����-Ռ+�#āL��w�ޟNC�o�qb\�ӯFљ���C1`
�g"��>#�w�X�%��Fe�9�q��^_�{�:g��-,=���m#}�N�%U�yXlLȨ̾?��?�Ǝ�d������u.��D�!�zrI[�(�ѹ���Ym�mnʤ8<9I����'�k�\<Ud:벟���ܩ����==
�Ҁ[��~�wd�no���+̐�g�f�|,�zUJ^:�<Ic�<Y����z�T޹8{J�=�\�`iȵ5��/�;.�e6�j��M����c���_ص��ۮZmS����f����#3%��h8z�ı�gr�J_�d!d�QF���-A;�|�k����G&F�'FG��F������*��eڝ��*��V%��'@��|�����}��P�Y���p���;�a~g���4p��7�l���;�cu���۫��V9X�v�>-�Dy�(����^�s�-���:ZK

�����P]�e�t؜Oz����¹�	[��������������������hn���Lu�]d����|P�4�WK .�Z"P�$]c�b:�ܡ� 0����7*�b�����J fa�P�����pH��'��l�����m��/|��R@J��[��y���τ�A�!�^�Ä��X���&q�Ef�6�����Z>}�2?���G�׀�U,l@�6Qd*���1�Av9E�X(MABThN|Pf��Iv�Ba��I}�.)�c�Nΐ� H��)-�&D���hh�c# R�]�P�X�íaJgDbf��순����;%����&��o�;�El]+ڲ&�wc����������ke��Qzfh�=X��C���� ���}f�
p�r�9
Pe��ᆇ�TB�T�IXAH�~�Yps�)p��:Us8�
-�94� m��N:�cK�&CS��e���N\Ɨz��j^� 	�u_�����o��>�SB��H
z���T��7.u�!�`=��8�0�������z�����?p�И�SScSӣc�����Vwkb�ِ�����g< �i���!�Dۅ�;,c���R����������w{Z{Ƈg&&�g����ppJ�8�����
:�=�S�7�c�낂Щl�����T��(��0?17�1�}��z���]��ٱ���Q���	W��Pﭡ�:wgB}��B�z�
"z�M���Z�����d�EdI:�'\�}����c�5�+o^y�����&&..A;�}K�/^��M�t���t�o�2��$W&�Whw�j�W��t��������'��_Ď���Z�j)L�x:�%t�w���Ǡ���!���=���( �c-`}l[-�8vT�y՝��9��zJV�M-�ϺhYx��5�-������yWy�#[�a�\Aw�l�5��SO@ſ"@{��ӛ7o8�9�ߏ������w���#|͡`4stD��И�#�c���l
���1`���E"5��y�"W�0,0zJ��%�d	'�&Q�4 ������̤+��� �=5h�+���8��#�������B�L2o��G����T��n׆X��fER͙P�&@PFd���<Ȩ9(��(M��*�By�E&HCM�=�,J�M��*7-��t�n����`c4��F[z22;֟����s����,J/��_/�K>((���D�2}4I���Cb��LQAfI�E*�Kc��c�rk���L}�\ۘ��cQ�	ْ��w����ꠃ�?~���.�Q��+Ml��=_�p�Dw��:B��Ps���c!�����B�h�p�q��r�5�;�݀�
��~ ������A����q@����&�2���D�݃��JB��u���͏��|}�	G�"?%4�������	��`|��h��Q�`іV��c��1.��|����0J!��䝇�]�\�3�C�$��(��$����|~�[�*��2/=���q��� ,(ÑA��ȅ���w���YB�J�:��ყ�)��,�h�=v�������g_�	�%ʐ��h\ t�^m�R�9>��P��IrE/>\��,Pv����=�a6��xjnqdf�=3�2>V�ݴݖ��L��#��c3�:��SA�E�ϑ 2�FKT��qڤs�,`4������ߖ�&GGF��4��c��3Ϟ<}��/\P>z�So���wp``������v�����X�+ai����]1?�kwT�����*�$��]�`�?M�u��<�j+J�tZ����}(�y��{.�zG��5���5i���1�m�H��J�Wq4��I����b������O~N��ۛ7O7ݾ�cwf۳�˫2�N�zi����Į���8����|��������������]L[�$m"_;��̙�BA�=��,]g
ʌ������ 4��8դ+�-K!tP�l䢥�361�=��e��j�0��*מ*3a�>�����Z�[2+6��BSQ��h���/��/��F
��	���K���v�I��(!+�
��뒳Ϟ(�O�9��bGT��Xg���)Q-$��4��J�:u4�h�+,�^Sq�b���9W*
o��_�:QdN�9�L��Q��#Ԏ4�%��厣"!9ʜ�p�0Ƈ	I��xT��M�"!Q�u,�#���dSْ�m)�δ{���$cAjNq���M����S�O��6����/��۽m��������Z}V�ә|��dge�͊���.;2����EXB"2E�P�� `��g��a�2o�%DI��f����o�j��\>�����R�L>e���q'� ��Cq��5E�Z��cR�V�S�E� �>+yB��rRS���l�K�gB�͛�!K�^c9�M����`	�T��B�	��/��������2�`���Q�R�74�=@�L^no�6TR�:�F
��F�S�r>z	bo�"P�Vl�on��;���.�C,������ё�������������z.M�n��B}+Ш9[��<�78>�=2���'�� �����������Lm��k�+<�^P�1�?��AD����,����#���ڔ��K�CfiQ���O+����O�<^\�C��>��)�y�_>Eȅ3f���-��]���w��nn��Wc:Q��)�z�hv�k�TD����?�4;\��P� t�}��k��^[�V�|�t腓 ����8��롚�`���P�P�[�R�@���>�'���U�����+�/��|��ݯ��{����<��a����,[v�#wtx�]��O�l����S ��i0������惏,��h�a��+2z�Y��?w��Y�k-��RW A�z+���|֑����M�Q�7�F}I��v�.��S(o5��,��ΐ�+>h �/0�z���{�X�L�b��~c��;Ӑy�%$ddެp\)2T�*�ϼZ�^j�li���V>���{�y���Fu�Xw��`��@�x�mw����bۭ�Mu-�.�]����t��V�XW�Hg�hO��`�Ԩ{j64=14;����3�z���|A�����[����K�5w���7^�9�~k��������Ł����M�.�7�n�\(>�u����F_���;�7��_�����;����w�[+2�\����xiDpp���OO?��=��p��0�\j{�q���Uu�VERY�Ɣ+>��͌YCCmaަ �P��������A��/l��{ma;�|	�"�F%!Fn(�2`x3{Ȋ� ��Kʗ�ΎC�lh~L�m���6����f�t2TIZF3�y�"��;d%:C�C��,��hN��F��&��A%5ξ\w���Nw����ƞ�VT��X�����v7����w���|�}�|�Ȕ�oR��ܡ�Щ�A��ޡ0P��5)���E���7.�����j�hu��a�;�C����}]��o�)�
:���I��X�$V3�
��J��I�P�q���mp�gd�d�	�P�)R�Ơ���'l<�����ᡒ�&���u&�ǂ��
����9j���U�cOИ����i��{Me�å���`�-�i��_�x��W�^�~�˯o~����ݰX�v���5?h�w�����e�y���񚲸�R͎b%���B�L�}�"!��x�M�Qe|��V{}y[Irù�'6��a�It�	Fפ�?�L��i?�R ��V�lЩΟ��Δ�uO����7�P��wUAN��aԛ�zk�#��^3?iL��ٵ�����o6|�������b�´o!l�@.� +�a�ߊ=*�!%�̪�x?
@3���a����t�jD��!s��P�_�'���=�G���L���c��ehdh�� ,@g
�2R���������2 G����L���41������#Cs�C���#|~��>9g'�f'���#��X��_��\��X��6:7=2;56?7�0�����),�O�-��3K�8O/Rm��1��.Q����3�0=<710=�;=�6:�`��mxx`v�o�R���3S|�?5�79:8;͖'�L링��������a��@Oσ���k�;]���������ŅV��������J��V��]��^m�]}��"�Z�:�%��#Ķ�K��-��B-{���!`�N!h�)�;d�@��)�q9��Cp���u��wG�lAY�D�]
㷃AG�D؋Ko��� �^c�>S $<�A��Lv�|���� ^ ���G�����!�
��d��H����~��$Au�Qj�M��-��*��]��woA&_m�[��u4���?h.�s�z�*�����)��(�[���!2�9Hv��9")F^'�MWG	���8�kJnߨ{����
���|�����n��ӥv�1����� ���Q�p[p+�c��EiMv\����|���NW�W[[.6ޭ�{�V[[sok�@KO_��`{��e��x��?P�ەq���̣�,��6ՇVFg@d�Ze�1F|'H}�qZ牤�iqqq�	�ϝ6��NB��|\�Ȧ_�mjr����n��+]���h>c*8���,��)�l-T�X��|��\�}9�z�+�����+�s����T���˕��Ԇ����\:Et�H��AJo�M��X���Gv��Y}�P�q��srWrrqBޕ���^�����^�l�֐iԟ<z,����u����߯�]��r��7��3ڙ����}F���3�{Y��l�C�-��Qg� �(�F��G
Y�3�:Pu��5�L�*(n����>��D�!3�"�w��a	�xa�Lx��I7лM4g4_�t怆���I>����9���E飏�_��7<88C�Dg��>�[z����������lvni~�la���å�G���G?=z��K�`��i����ESǡ�ٟ��s=~��O�{&�ßh���ŉY�{|f���=�lnbf���g��2�7G�M~ns�S3�c�ζ��{�����|��j�/]�r�|]aA���d|���j��#��/j?�{ť�rr�i��Ci�����A�S���A����=B�V�7-��w�h�m�s���F�'n;�X���p F��������4s�	��;ĸ1�y��x jWh��]F��� �.�=�g�b{9�c��s�	�LAӓ�4����a��b:IPG_�:HR���Q[N�*�>Q�Lp�Rs���θL}xFJ�i�`�#�ɏA٥���ߍ9�RH��Xs%����:pN�sV�&��̧Sr��<�F8�1������:���)qԜ��Fp����\��!8U�$cTG��g��O�Ζ85��ҳ��ӉG���+n\)��P}������7.;n6�\y(�̧�*��c��#�b�M�Ω�"7�c���}l��Dm4I�mb�iKq�A?�D�?k�w�J���j�����/�@��}K8ߠ��={���466���~����W�_�^Y��0�Ӣu1	�q��"Ŗ"�R���24�zk�f_M�u@�ܽ .�	ʣ��Z}w������'��?��Sm0K�\��&����IG���W��.��^H�E�mm{���/�߼������꒢��O�;��e=hl���������w�M�� ���`4������O���{���N�g�����
�=,�52��k&q�����	f��k�l����΁9��X�G�1���ch�W��F�W��B����;HiO��	�C�G�Cp���������@�4J��	λW��FGh@,��Ç�_;>���HU<� ���ѣG�������"p����!�>���'�g6�ؒ>_XjQ*����3��8����'f&�ha�%�J�qyq�
 |#�xl�蠻���מ�ܵs{^E�;w�^�RZZ|��邬�+��J��.V4_,�P%�\'��1���a	 z���,,�B�
Eb���u>��N#7y�q�q�q�(�/F�z�*�/�7ܤ�Fc>���D}����rh�F};���Ί}� Й"@���~@�.!`�1�s��f��P�e
����
nB�R�;�易�6D�ҳ�2E�y*R4����d~:�_����Px��|�J/�4�BAuP����X�
�g$l�>������ƨ�&10��{�d�z�o�,����,m ����\B��N�n��	��G��I�s�a��� �,(]�.ё���j�>FfJ��2S�����S�ͩ�u�q���G6�����l��xs�R��C��!r�U���Ѭ�'DG����#'O�I>f8���*.)�v��_�v�޽��Ǝ�w[��k�s���+7�����/��^��/<u�DXEJ�"C��O+��S��\��T���T�]�Ft�$O��
큺�U��=;=��{������3�uG�R�Й����)��7�&�PG�|>�}E��ʔU��k���c�ct.���ŧ/_���ͻWO�7�t��S%��wo7vw������_���ia~~%��}Foz_D�������t��l�C�>���}�g��4S :�`#w3�`�x�9��X�,`#
[�Y�����j�Й�N]�1�kdAU���<r���&]��R���+���&�n#��A� <$ȃ)��w�'&F�fA���E�d������3E�N���́Θ89���d�?��|����P++h����!�q>SӴ��@���[Ok8����N}iq~�F�[�����w��_��Y�عycBRbÕ��n\�(/՝9)�>y����ʅ������8]5�����Ln�[	Ш�3�t�o#���>[�~`�O���	�G�@���	I���c�ڢbu���{�0,�� ��� ��{�ߋZX_D_�/p� ��m
�i�Ǚ���a
D���a��"��f���P@��l	pD���P*�u�MA :�t��iS�l�����EXFf��������6�!�Kw�ڙ����@id��juF�]\~��S	�2�OO2=��$M�؝?̨&�7��w������C�� �	��)���"��s���(
�(B�2.D��)^H$P�_o!�۳���*����C�b�CLs@�V�d�İ���v���S��}�v�2��:0.<(�G)	O��;�|85�J��p��	�Ng����r����Krr��r�َ㺓�üB�"�F��0֯P��@��P��D��L��L�u���2Ֆ�Xj$���wT��*��-����4�N��ݬ�r�\<\t%�H&�\�
��6s��c�I�3��֊���c�2eb��b���/�����??�)�u��fٲk]u=��K�������"����Xц�hM^�~��}�)���O�s��e*�:$�:e�s4��
_�2�&a
�� �YB<�x�I ��n�P�̂珔5�Go�Y�����%6"CY��Koᛴj��p���xX#94�d���O9x���%QP�d��z�d��0m~�(3u�5u���@������3MMQ�]� ��}��2�#��xN����A�&�m��vY�.�3��=�z���,�Xf�����a�M�4���� M���J�9M3<B�;�5S�Cí�zn\�˱�Q�i��3�	1���$m�EW��C�Z�מ�+������-����XB���<�\a	�k�@U���[��H�	r%낶�`�t;t��y�i�	�d�/���G Β���S���e憦�m��u�P��7������&�}B :;��LA(��,~�E}�6ǳ�kenŁ# �(! hl��z �
�IyGYD&4�F�4�.����B`�9b�!��\��'��:{t�#��E�/�g��GXs�����HyB�Z�;��P]�����;���r�MO>:�-�;�A8/c�!c�%����"}���8Ȫ�el�P�4�&��ad��V册ȵFهV�G%��ed��F}��9�@�:��m��d��7k�Ω�����ܴc�H)G�d�"�V�|���S�����ΞMO�e�&��F���E�d�3�Bsc}cw櫶��rH�oJ_�ʿ*S��-W�6��7Uh~� ��{�*�w@ON��ߪ�H�;Pw�k���$_�"s:o�L��2�[W���	[*���%m-K9BQ�9\��33���ի�?���U��ق�܉3���o5������>��{e�������+":�@�өx��k��ߗ3�kVx�䐯�T�u�W��k��/,�mV�vL�]JC�["X��SAݾy�As$K�
�o���D4� �)r��`�b��rڱ�Z�H���+��V��x��;X]��:xG���"0����,�R�> Zb?W���5N��iDb0P�`$&�g�h�	x%9i�M�Jʒ��=]	+���lG�d��သ����6�˴����q��h�Pv����wGX�v*B��|~��k����}�ZύKWk������뮢�{W��^���okP�P�S�~� >>K@�Z#��^M���I~������ �y����c�a)3�*��J�,\<��	���Yr%��6CSX�p�q@�>�w����P`�����hJ��s���m��1���^� �C ����U���M}dB� ��9�@^��7�3�Wȋ��X�{M�T*��@�P0R,iid��bׇP�Q#-㉅�Ɯ/������L��K٣L[u!X�J\#]�.h�6T��Y@�PoS(�k5���" �i8s�%A����av�A�쫳�k�RHf ��L5 ���v韭4���W����ʡ ���%��$_[�?�U^��(K�ܐy8�d��$lG���H��"�E�fLҟ�LV҄��F���a���T�rds��
�d%
�/Jd��Ⱦ.Wnp������B�����:n�+)��XO7:6���{���<��)�ڴ]��I�\ɛk�h�ySu↊�M���qߖ�n*��Sy,����8�P�1�t�����'���rLg�O���v��@w���4��N�����͛F߽q˳���梸e����~j_f�C�I�z�C�>K�6K�&S�:S�����S���!C�s�d�]��l�Ҙ�,��T����Î����y����icah>@��Đ��
Sf
��ѵx��15MO9�o�~"�.{�@��т������ë���/9

�S_���9F����1����c�#A���q"%P�m�18r��������3ގ2�OO�0��r2��8"����G'� vXY���<E^ih�WL�
��]1$���zth������`���;#-wݍ7�o��t����uu�߬7��Ju�c3�b[T�@�Sr4�F��e�	��� @3�X��o����A���sFgU�b>`&o2t4��o�BAH�Dj�?3b(�a���� �$��o���������ȑ��
�|H��CG�~�-״�MڜE�aN"�<0'm˟L�W�
�B;�jf�����L�'�:�"�	HZ�R��\Ha� +��M�^��Q��&�ǝ�1|'�-q2��@3o>�q��۾����t�0�c	��HW�BD�Ejc@[#E6QEOɿI_klW�;Uej�j��O����Q�K����A��Sû��	�E/�'�g�6�W��;�d���m����4�xq��c>:�4�x�=�W��4^Θ=�����LņL��9�o����@�o�Agŗ%���U��+Ԙ��|W��7W�l����*��J���UFƺ�.tU�xֿ:uGm�֚ zk�㞍�U	�Ϡ�w�ߕ��X�t�����dLa���b������߽y�0>T��c8�϶��w�G�#o~~��VAcZqt\����=L�����d�"� �[��h
� ���ɡA�^�� �� 4�
�6�������}sB25�����{oSn4��0�;��Dc%PNIfEȁ�T�$F�m���a}L��-,�2^�8h�F��/�#�y� X����˨�:tu]4���$ 
@O���:>62�l��,�8(	Fs4����L�d��u||ttd���G&ƇAj�yjz�mI�G���i�_V*�z:
4g4X9As�B�ya��gR���"Iihz�
�g�{&��`S�]��bgtlb`x�Awׅ;��s�9119�H[jЄ6�*�pr�	^��S �Ͳs �0���!�CЏư�Ji�%?��r8�f�= P���)yK(�LA�� љ��b�!��f+��ӴHm�����ǟH#���&�CA1�D���԰̟�7$-���G ������t�������$t���w�+ ,`��� ��Y�����k<��Z�eOl��hTɌ���̭A"��ϖ�@�h	�n�B��)�O4���a��!66�S�E#}����B
t� �Ί��C�O6�_3�dN�GY�3�+��Os�k�����!����.��.��e���$�Z/ڐ�&=�}�W��/M_XE_8%_dI?�U���H��󷥪��� 4��,��r ��+��T�Q~����j}�u���������i;k�D��4n��V$|�J�X���<a�+yGej`�1I���#-KO�z�����MYv���n\�3=9=��5�(��i���'h�h�g�_��:�Ϙ�b-��E��C53:��S���F�$���r��2UZ�@�j'4�fmV�:�f�U�S�';�';>,[�9�~���칧�~��������l�Q���z�dм+6#;��M��aN-�$�#�p��u7�`{1F���L/'�K��-I�0э�[��������.�h� ����C�CcC��21�D$��	�&D��o��=9�&�0
����#C�cC�#�S�$��پ(hK�1�kovVdlp�����	�󓙛��q���P�s�cs��s3���cS���#zz�߻r2�DbN��&a�����2�]fO:`Hes�� �� �΍�NF�����!����-E�����w;�M�͙��(�*���8��A>��krqP��1��`���c������³�9>zjfIB�w0�D�����Da9,੓Qe�E-�( ps����q@�<c=r�ᩦ�D+�F��4DT���;IQ|���L������ 4K��+2����R�`�������X����C,a6Q���[$ -ʤ�-ve�|� ��G��9�fi>�R�5S�g��>����2�h�غLt�*[�z�5�y��L�H��E��%�!|���.^o��,K�y6���\���/�%��˾.V��)QU����9vC����2�
���n���銃��N�=��ib����JusaJݱ��#�j��զ�P���cm�&W"�����]I?�'m/K�?*)MM+H\�Xz�ӛ�/��������, >@���-��gpfjڇ �ϧ���}#+^�;W�{Vaz�ra�1��o:U�٦��F���x�U�YF���īX�/I�Lͺl�'��k��k�56�gV���טּp �*�7G�Ʊ��{�J���y�����R?G>NmlF�����Ļt����̥�oHS���^6,`.��P�W�q�e8c� ���R�8 
��noog}|ɕ� ����������r@��BFN� ���'���He=���F�c�������i��h~4Ng:�e���虰Nl���`>L�ŒR4��<�����쪹})ٞ��GGX��,�n/n �e����5fsR���q�h9j���� %:S02�e��3�Ǡ��`������=��B�}����mQdV����ᛣܣ.)���Au��H>:Y� ���A�!{Z(��� ��5AhR�X�A�<�,�5I�M4ޕhm����������#����1��Q��8̢<=K�EdR�X8��פ�5�}	9@�8Cr^�g�g�k�������nS�o'E�3GE��7�$"�Ɉ,
���P!R�K2e�Vj6���D6��)�pHY��Dk�*��ov��_�2U��˔��gi�����쐱V%)ôj��,�'���>S�Y�b�C���63j}�d}�l�S�I����y -��H�Dt)���Y��"�[W��G ���@sYv��ѓͮ���ZMkij���c�k�l�I��]���:qcUѹ2������S ���#�3��'�>y��嫷?-��eٲ�˧��g��z����_��m��Ϟ���Pg�w�4u�_<{��C����y����f1*8�[�e	T3~����5v$�'YZ �>3k��U�ZT۲���LM�]!l�����BVx�d�6J�:��i�B<�x�y Mq71�� �ta��T�$�Z ���Gl��A��xc��H����2{x�5b[����uxlp���f���?�����=|�fB-g4��Е	�f�@LN��1��������AWoKOW�`�����(˕����ݗ��X����c�ML1@S��e��G�n��e���@fЙ�_cz��y�������xSwO����9ǔY1���ԃ2u�ɓm�u#��XC1��0�n3ö!��Ԙ��DX֯o�)`������4�~��J���Y�:(C�W����q�d������䤦�AJ�d�.-�BN k��)���G�Bxq�~y ~wK��z�|������>7�q4��L�9.ج�7+}�
���b6�L�ϛ�C�Gt���b+�G��8��O&�9^lH�I?[n3��(2�,��.c}l�1�9&�,�N�û��$�� ō'�H�^���͂��B@���7�n�BX�%2�%��dV�®�Ph�ġT�j"m�pK$ e��:$�N��k]�jA�&7���]L��X�>��u2gt&-��)�$O�&K�6K�ک\��\�)�-���lպL��Lɧ� �t^�%��џ�H?ɑ���,W��P�e���h���)��ƥ�?-�^���B��Z��K�ce�*Jk�ߕ @{�zOO�ܮm+K�?V{����=���z� ӛk�)�
�N�R�
@o*K�U�Y��(N�]*�z�t�g ����B�U0�.^��0�851I�V���� Я^�Z�_�ƫ��n�]Z���w�^��()T���Ė&���,��V�:�t�EFs74wk�sF�X����%3�++������@�D4��T3 �Й�vmYV{4V�]���-����xF	��(_;/�,���b�\�x*���ʔ�"ym�іˑ�TZ�H���VR��FW����,61C��'&���,��E@{���z���6����]�ϭ���}�jk˽���~w��r�@S��q�7v�Cc	����ݿc'��f"��&_�̋�'l@3G�GG��O�<�����9�����Ԫl�aV���B}q��#^�c�m	�f��n���G�u0��3��:
��Y8��x/6���x4�^#�B�I���Vv�-�b�����7S��!p�����zp��w<
�
rO{z����`_sw���U�b�ȁ�g���P�Z�H=Qi��}���sr�wv�cz�z��K=wWKU�Uf�"���A�m���F�!{���9�#hSDXcS�u���Lչ5���~0��<��>��9�n��p���n)k>/���d��(
_�s��W���b��<���� sCR]�H����S��u�wʭ�r�r��-�(;΄Ɗ���L��.���r(�ԅ��M��9�`����cfk	�X�7���L٪L�D�Vg�@jf22�l}�|u�dU�h�#���a��)��� �<_�Y��͗���Π�W�.�?+S��qix! ��2nOe�AW2)hޓp|���}
��R�^��=xGm�*�h
��T��}e�Ɗ8��,qOy��6AU���n�ɳ��?�z�t���<;�n�ij�^Zx�����F����£�ǳ�3x;'�gF�'= �_N^�N=��_���aS|e��5K�Y�0 �#K�F�UժLb4-8T٨Z���(՟;��w��LωAN"��`���d�9uEaRX�n��B���XM`(x��J(^	0X��^	�����
&c���F�Ҳp=<���`M@x�qL���_1��{��O��TYs# =:II`zj[X|Ⱥ�LS,c.װ|��'b���1t���z��z�k�\�3�8��R��[s�\���v�g��=�785�]<G����}��O8nDd�Qv4n�R:.���e@�Dq�_��73�S�\]=Y��%BL0��f�h��\怆�fR:d�"�b0�ˡ�tf�XLAl���@���ܣ���0���ؘA6�?K��� �{����{~X�2{Ai���
zФ��7�O��Ѵ�;8`��Z@ge�%��Px���u|p`nzt~nla����L���ն{W{�UfJ��r[�4+���B���rИ��`�"��x���53�;124;9�4?�D�U��g.�,-aY�����>}�S.$���f�۔x)HMS�U�X8����(xgEz���͢p�<9�ĭ��Ή��鑮���75�d�Ei��`�6��)U9eQJ��Uz�*A�W��/�?�d\D��
(菲�g{|P� 4lM�zm�f]�z]�
�I�ڙ�ǎ�UN1WЫ2#�d��|V��$_����j ��"՗ej���Gql��~_�CU����j��U�������e=	�����oU�����>|��06�^���:���T��\PЉ�\�ߕ�o,��ѕ��"1�&N]�Pv��̓����I��+Ev�Ӗ@�&'�������O?=����᣹�����/����/�<��O��ٓ��ƪ�"S��Zc���II&;Ԟ���&4;�+��_��������P��D!�� [$9:�8���x[`�4�5I���+�`����7�u
��S{ȁ���f�0G3���Ѓ�` ~�����m����b�o��Q���q͎B�G/�2�(��ex��mfy�9jh2Fa���t��mL� �� �r�b;�rp�b$��{:�TJ���сzu�9�H�|4?��Ν[�=-�C���Q��(�<�î���� �1@���qŰ?a��Y�Ş]�f�ִ�9���A��ȝ�n[]Y�Q�:;u�c�OЙ��J5�Z�v��% �{��:ck�ŏ\�Dd���wDdE%��9,`�xB�O��;��~�ޟ�1������1��<���f��D��j��I,���,a��F�t4}�9��C��p!�r��q��=336����ON��Ȼ5<1=63C��ַz����{�ٯ����A6��n@**п!��d���`��������]1�w������<�κT��u*J������3NN9�
��	�m��G�ũ�Gm6BT� S;�oգ0�ZX�Y|�K�Z?]n[��t���J�,:[)�R�u��"=��ˡ�ad�h�P��f*V娡��e��չ�5�ʵ9���J(h x�C[儉a벤��;�1_�-�4G�>W�>O@Z@���(��\��lʯȹ��ƥ�X��+fse�κ�]թ{�R����+Nܩ��44���y��˕\w"��Ⱦ��;kR��w����x���H�v��"�M剻*�«b�E��ק?[z���OK׫]%�,����1@�OO� ����R���充% zq~�^��r�>}����_~1u��1��~u��@VܷV�gv�g���6�W��.[mS��L8�|�Sd��tT백=z�#n�36<?>*S� ��|�`�g����(�����x���%�뉨�.l`y�EBX&�UZ#0?��2_�!�͂�V M�8v��RPr@������ߤ	�K�h�`=z�<	���}Z������fД�����f��颃Mr?�$�$�ˀ�h�ټ׮��6�2w�v!OŲ�|X��� N��I��Q?�2���;�#?V�:~�i�;�H��]���PC45d-G��4Q�mE�U�w���X�aؒ�hf=	��3�0tX!���U��Q�r:�5Q�B�H�{��f�����>h�}�	��t&�N�l/���Yb��h�����fy�I{��~��50==1�013O�G�Q4�����ܔztthb�czl~n`z�kb�r�=�5%HP��x�(�%k��"MFy�A��$%HA��ndl��<6
[�o�m��_����q�l�-ʢ���R����Y�7�O<`��^��x�T��D��3����q�K������+іd�E.�E�2�Xa��)t�kC��f	�ٮ�(S�Щ�@(h�f"��rT\AC;��R�Ζ��Usм:S�̱~]�\&_GV��	�1�?�� ��"��LD��_��p@s�:o����*����-�	۪wצ�I�=�{O�����꺪R�O���w�R��5���63�7��~W�]i��I;�B\���$WӍ��O�->{�p���<;�U~������O��3��`^� �;��9��K� ���dwg��(�Q�Ջ���B��}�����o����`�:+�L�怆v�?�B;�(gLVk>�(�XU�;���cwص!91���H;��X���xm��Y
�P�\,�"6Sk;8KDf�kb4���B/�`��x倆8�ۇƳ 6��s`w��Wr�`/&ҩҍo�)�T�#MǊIACF�hL�1r�_�fe"ڱmV����,)�(����s��l9Wf7(���fe���3�U���K�Z�����A#���YD���J:36ѩ�.�˲�s����������;59<>��k�w7��eT4����v��x�1�C�c�f=��psy�@8��Y����GX��Ӎ2�2%�ǜ�|���F�"���MS������Di��ǢFEHc�/S܄i@ �4*���4��A�c4�m�6$p|�����'�Ʀ�P�Q���x�������[�s�ܿ�������^���)�=9R|�B�%>��ஶ@�,�&�������!<6��Cã�����m=]�ݝ���nw���>�
�papf�F��=%¢�H��b������P��z��7A��B�ʄ��W{��O�N��/,-������}��Y#�K�h�C@K2���+}�j��z�@T�U<�����W'�X��.anh��,)0M��r����ȱ����ȕИ�+�<_�i���B0ZFU���.�|UJ
�t�P��*懪�����I{��T��i��v��Z�T:��( �����#�[��~�L�Z� Rc
���4�����'ִܞ���K/-^()�.(*,�j����3�p��l��`��<y�p�J���ƶ�1�ճ>~�d��=k���ܘ}Θ���N��v�jA��{��P��1�34�l@AdSb= M
��ݢ����F9$ t0c4���?�V;ً�I��F��\a�i3=����9��Klڑ���L
�1\&G��[(���Y�E���D�x��z��&eD���n�Q>h ����a���eNN��#��'r0�����{AR��4���|���Wx� �q�M>&����v�T_U��z�g��=�?<�ſ�w���҄�f�%��Y�tǙa�vf��	{��Z6�+��5v�V߿�Zd����.!r�>h�.x�>x�.�L���!�GqpՌ9_��Fq��ެ���ܰ% M�e�>����	��v��z�AY2 \���cҲ��	�lG�]/K0�4���� P�0j��/K�����!l��-Sà%Zj;\~�Z���yu������v�`Ã�c�&���\��|,�<�u�����N�~��i�c��ԝ��U�`3�)���|�Q�6y�c�)jvbˁᑖޞ�Mw/ܹZr��u�R���_y��F[{cWOW� �A��o����w�Y!:�,��%s:C[�.T`4^��_!*̤һ��F�񛲑	1-..B�LN4�ݎs�J�
�]@k��,��]��$]o�,�+a8�������?ۣ���.弆�^�����МM˘C23��2G�k>���8+�tt���J)����B��E��˴�_�k`���W4�F�ce���4 zWe��������lvc#�]���+8����|I�ɰ-�8������,a{i|XU��0����
�k��ٕ�#Oz����4��h.�ߛ�~�{���ƾޡ���ٙ�'�' ��seY�=Θ��2��k�44�A+?f#����h�h�bU�ό�ЪXeU�s�?���]�Q~�4':�
	@S� �R��1��z�����,���yD4l�W4�Q� N�u|����W,�X���`:Ȏ��-]4�Am�l=�`�D��ݿ�44�?F�Ǒ��hc��Dgn�(�q���Ms�d��	k�yJ��� *��!:��IM��]
�HA��D���W��?hn��&M_G��S�_�At�YB%�yN;�g^������~bt��P��@F�����6��Z�儷��$�.D@8���]��wz���/eG�ndI��ef㮏@�������z�'�d�y���2�����r�Ȼ����t�h�ohw���B�����������)�a��dW���7{�{Q������G:��ښ�gE�ǅc�pSLDz�,=%�0�FG;���gx�kt���@�� ���)Yy�Ya��(�z00 @C&7ܻ{���l��d��l�<#Uk:�h��L��wo����sFMO\ﾟ�&ԈG�r��g�n�.�l�������B�j�1�����a���7=�s㳳M��j�LЊ��C��R(s4����M���T��ة��ߙ���8�,x�y�s�g�x��Ng4�:�簔 �$���3%��$ ����k3%<��&]� ��(V�\������+������\��2���wW%@A�����ct��^�������gBj)zgM�����ƼI,�#��2+~ki4 �j�:I#b,��i�����U#sZۇ�?}�0��±<��L�3N�_�~?>q@/--=y��p����7��z���S��h��ճ�g��r��m�/*~�Zd��O e���8V9T�yP�D4�J�h2 ��b�;�� -Hb�?� [�3�aЈS�,��a����
��V���U����=�Yn�'}q�Ic���n�W����p��O,{�.����A#%�H.��z��ο
���=a㓿g� ds� �8/��ab��^��L�)���[�-'KMA:�����o��D�f��QfH�Ք]l�h���ߋ�����`���E�9:x���)�K��ԫ��2�΍o�'~-��Z9x��熊<�c
��y�ی?þ7m���p�N�Q�:�`��A�����%��ޛu>?�{�dߧ���#AM��M�YfM!|�@M��2r����4�� �w�(�(7�B�-����z?`��7������G|�g\p��l� ��Py� M��|��!�v�u���G�N�����i�/��� �<�,0JB��HA+1$�.����7���[4��W�;MJ|3Xd�����j]Yv;+����nw�uf�2�����/]�S��S����jo���l�o���Ѽ�
[B� ;�	̒�!�y�%����A����+2��uwQ�:���A>x�������;�ƸHA&���ȎwM�ˡْ��un<^U�#	
��^0zu���tU��c��;�y�˷C��G��#��C̍���� ��fFA5�sCs����/JW9 �U*4��J��}e�[��[�-*?���X�������Nq����-�	�����W�	*b7�j�)��RR�(/J.�s�����O�WVX�׮4MN?y������g@sO����ӧ�>|���Sww���wQ��f��-��?{f��0�G��S�t^c���_f�~�Kav��
7�N�����(?T۳�����Cf�X��-��Z!�31�B� �	�9�E:$S2Fg�h3'2��tj�c	K=�&�t?!'�)/$�ہ��ٜ��x�,��~�Hz��zAf>�s�ڃ�����6:@�C�x���Ï�����l�31�B��2G�Ѣ� ��G��Bp� 4�t�<�[�ё�öK��;�;�Œ�;	�����>���2Me���,eߘ�0��4�y#'��h�m�;a)�����Pj�d;-�La�����`�f�N����o΀^��H 4x�)�0�U��a�%N�Q�����-��eZ�"m�+��F�Y�f��/�85<n׳��,���l����G�� ;��y��2���-�s��	���t�7��D���Fq�Nk�Z�8��;2>8���(y���H�A��6Q跟Y�I����ؐb�PYu��������%�7bs3�u�}��u�,�dQ����W��ݓ���A{}1��/H�̔��� ����&Uȹ�3���zz�0��S~��ٶ�^�Ղ���@���71��QD�	���%H�L׃�C=����k�MuW�u�����yV����٘�}ZfU�,"�S&vJ�-��f�w��/�b��`4 �a��lrF��P��J�h�R��v�6�v�G�(��0-��;Ͷ(����֐�u��g�?ˑA>�+�>h�ʯ�5_���X���j�oʣ7V�}W	�&l�J���Q���:ɷ���u���E0�O��HXҔ_s"���8v��V{xKU��Ce2l�+qCy<�LV�C�&�2^Z��}�f�!�p���sws�+�p�o����~y�fif�_�N���L��4X�_z����Ǐ_�x9>4�t�\�P��3�*\i�s�E��͊u�t� YoS�����U�����R0��B�>[���?�J�fd�G�:���f�3�3!��0!�&���m����VP�%3-P=4�x�@+�H�Ϝ���,=?��wԒV��>zR��y������@5�7��R2/���}�P�ǲo_�P!�ű�!�we���f�v��'{�|Kdp�T�ն{I�'�uQ �^�'���S�@#�x�d>:��z,�ƕ۽�]��Z��bb%��{ ��94�g��?+|?����N�_^i�!������|p98]�WE�}o����h���2�uP2h���s��|����`#]1���b��(�)c6���Nu6�i�z������ève���i��B���ƒ�1gK�O�<ڑZ�-��vrQ=I���7�;��Fh\;Tg��p���b�6̮��J�4�� 3���)"��1YgO�r3Η�d��������!A��4�H���bj�|b�cx0�Je�^�c��#��h`
�2������r��=8�����|��pލ�H���D� �.=��SCa�kP�d�����7>�7>�:0�_W{�f���	Ѓ�t-�)'&�{�592�Zj�3�R���,��t�'&��z������N+��
�/6	�5�;�O�H,|� � ��.^�r[�m���R�;�V;�>ɒ|����)�,S�y��͗��/���%�`����Dq�G3���������:�@mZإ��3E7���?�Ot7�^-��@�՟�����c?֦m�!�cxCA��ߖ��6��o)��q%JK��/��--�?|���������~���oo~y�����S�����_��ׯ.>��<y������C͝���ёɅ�饅���X��70�Z资]%�3�g� �?�H>����D0 z��)��Fo��CA��Re��0�4�B�@3�ACѠ��Z�8�Y4�I��)/�cp4ˈ�ӊ���%�`4v�e��,��G�7r��(��X 熅��0���[�A���!�����C�Q�,@qE��3@�||Za1�'�W =�>����Ƒ`4��]NOj��B����%�-�Z�̨l����y��Iѳ��L�����C0'F�s��`�Ɯ��L����|��,G�`���ij�����m�|N�+=bsF�ܠvB��&9:�@i�XG�픔#��Eo�8����a���C�|f�����	�෠����hH�=4�����3d�v�H;rn��,�Z s�o��|�"s�� �� ��ʚ<'%���x�7P�}*u橚� * ������B��X]�8[�ܪ�a�<�(�(aAFY�^��d��ehQp�
*hR ��
�@����~���u��X��P��(�@�7����El�	3�e5T����ZQt��͎�6_�	�(��D�}K�o��m�ܯ��7*�ǆ��}�M��֪R��DQ��ƞ�ޡ!���ɩ���5��X�S��Td���o�#>1+)�ʡ��A�����M�'��XD��@�xJh���V��1���.��N���ϝ�Ol��2���3��s�tC��+���L�7y�y��5�U_�+7*�.��&φǨ�P��B�X��*~[u��(h��4��# ���16���{��Aqʅ���G��ax��(�X���\�MI�w�q4��#J����Z��]\z���㩉ku�W���߽}���G�+.����M&�O�Þ={@t�����M�M.LO���
�9�7'�k�z�� ���C��S��B��b:�C0�$�9�WAn[U0 zgV���ZS�lR�`��8$G�P�V�WA�z=�����W�2��e�,�d51��T�`�(2�X�w�D�c��c��/6V�@�s�,�X#P�s�k�:Ȧ��v�l�70�w �O���&�qA���I2P�p����;<�I@���g�q(��M�]�]"�*Py�)�0%���P^Qq»J��%�ۥ���ޡ�����"P��K�4����01�
�P��� �4�=�����;��u��zxf��ޥ�s��-�����-�P�f}�&} 4o��j�)��;M����[u�v �i�@*D��l� ,�� 2 ��~[��-d���q�����Τ����nr��=��|�����I�Sv!
��C��&@�Yji|�},��g��s�G�Y�JR�>F_]r��e6lzz���M���n�i�丐g;|�(]aIT:�#L�H�:�$�3�}MJ+����*�5˂mj��ZWG'��~��P�%W�QC��� J�qX�X��AFm\fFU����>�ѹ��C��'��/�<)�(e�Qt� 	ɵ�{���S=��׻�g%�I�擥W/���˓,NN�O^i���LS�U�L��cS|���ҦY�^��|ĆS��U�?�H�V9��f�#��N+�fpy��ҥ}jW~nW}��֩ݔ�9;fKn�ּ��yq���?��|��ޘ�ޔ�1W�!W�m�jC�"��R͆R�7%��ʵ�ΜδP�bQ�[+c�U�ޮi��
f71���{�N>&������۫�'!��c-���
%��P��7���s���K-���M��>{������K�zGп�{���B�������Ϟ� �_�z��_��OR�ˇ3c�#Mi���l�n��s�b�E����8h��c3�f0���Wۨ��ٮYoS��O�7'5 ;I]�"s(D�(j$��٢�BD�"H!�>f.�.ċ���e>�
�eh��;0���L�Y%��-�[��@hv��#��2S,6œ�C��a�?k��`!@g߽�h<�$Z�16q4{ͦ��L���5���GFem�}���D��P��O�<��	�(��ˬd���

v(��pc��|Ņ��;�}����~w��`�{��������}}<���������O%�y �'~ͳ@3���h�݋�g��ҭ�0
և�h���l�v�j�4�.&�Ԯ ����n�?�&3O�M�;�~��'C��bYjo��y�X�!�x)��e�`}��	�� /�/	��Ե��ƟH_�G��9�d�@o3м,�),:� �|H!������;�}���h����������ѹ���[�M7z�.w�=Q�;^�K->iR�(ŝ� c=�%�.��C,j���UW��B1�c>�^,	3i|�.{�N{�u�119K��0411;����w��7DY� ��@����[
�Ff<\�|�o|���k�-5&Fc$qe�{]}�#�529�<Щ�0�����)�7ğ
��9��;Y߅L
���ULc�8����L��W;i�5ŗ��ϝ�/������;��J�]ia�ia����䰲���D�+9�")ҕZ��_�H�=W��@�}�zsA�Ƣ�%��ʢ��I5s:[�-�wE�Ft� л]��G���x������;�M�)��Ck��;��&�:V����M��&]��4����m�I!�Ӛ����Z�g�/.�YZ�{	��gl�����y�0���Lo#[� ��_={�t��v�S�������tkG��d�*_�զ\o��$��f��*�H�4���>k �uv�Z[4�k��Ol�����ڽ��ܔآ�]i��āV�%I,���S S������x`�E!w�����R>�@6�>)�5*�|�pj��Ѩ�!�b<H�����9��n���M=-,{/��a�2T8�u�ʽ��^�9{��3��K�'b�G3%�þd��7��1�[�Ԡ�ņ�$����~��:4 �>��S`	m �M�pC��ʼ�;7j�.��]nm���	���y�����^������v��zz�������D��=g�<����H>c�� ���jdz�� g�����m�P�i�)��y;��}9���V:�g�ї��g��Eb�b�@J�9����5<�`�m$o�)<y������h��vF��<;VR�!s��D%���R#2���T�������*�1�P/9Zbohkm���b�3�NN�O�@MO/��&�F槻F[G�n��X��T& 1:�H��-��C��p}�PQ�>8�?<�54x���H�1ب�f�c�������0����yyx�-*ܓ#�7�E�&�q\��>`4���щ������ӽ#cw{{�.W����ԵJ���\zp�659N�*�zǇ]w.$�R�V�ܩ������ �@�_-��݈�4�Y`�}dS|�`���?�H>�+�95�T�!�����f'*N�CKbB���9�a6�ˡH�������M��dH#e�*IMB�+y_Q�|�E1?��n.���e�b��w@�zc��:v[e��ʸ}���'5U����?�u���*k*J���9���0 ��2�S��5)LD'��+'G�K�~(M��<%�9R�rixf|af
�����ꫳ����������'?-q������9�	����9��_<{���Ͽ����OO�G'f���z�c���S5̲��₸�̒O!�M�U&�!j�9
��r@3Ѡ�' �E�ڢ�ak��O-�M�ؽ����Ը�ճ��vI���s�CFsh���Y��D�d1<���T�e)�F*��9od�(t��*���ʎ�h<-	k!���w�5�� ��c��+BɎ���X������T�g��8�D]��G�b[��;��N�xo����_/�5!V��)�/�Cp�9�6!4[��l�Gb?�"0(�u�(c��z65�z��q�4�ty���|��2��N���
n\��w�z{[cO�{�wh��i���_&B3��p��206N1 ׻�+�	���z���i�,;L��i�� �!�%K2�C�f@���f���h&:CV�1��5����̣ܰ2��ɡ�#7��B5[B}a|c\��@=VX*%���\Z���	�` `{l�9wt�^�m�@ƌ��ڦ{���Z��Aw��
6�?��0M}�g�-=�YZ����ŝ)�]�Rt&R� �����o����κ�����3:Rq�A��jV�8��ρ��00�ǄrW&�$�ܻJ���������{��с�� �s�Ht��&Ut��k��SӣS�=�c���2����<¢�������n�?��MO��8W"�Y�ʬ� G�w" �\pt�ЪX������Dg��#;�D���^����6�'V�Wv���Z�Ҕ����Sp��W&�k��_��/��w�x���q��a�_��?�����DJ�����W⾢�=e�?�h7C���l�ˢ�fؖ�8��G������j���OWp@���M���>:������ݵ)�jS�פPB;f;k��P��X��,acq��d/�qI�aKC����O�f������5p
��˫���X���1�2-,,�� ���y��[Pe������������=Vj��g�l0K?�ȡ�a_g�~f�|�R�)z�MIf���(W���T��k�����-	҂�1IJ�
���p�C��u��9���e
:h�z+5(�<s<�t��MF
Z�F?�im=��0�l���t6���( �k�G�y��0��X�i��qp4rq�����$�}�c��-��[�8�	�l{������z��P7�==�n&e�ѓ�d��|�X@�"���b=db�q@<��F�$F��^�.?�!?xV�J�y�^�C:��.:T����g(�s����rk��.Jd��^�<�b�N�X�U\������m������#���y{�V�K�6r�LM|����YL#�b�5�a�MkL����L��f���z�Yoo@y7�Q�gZ϶�k���&����\���Ҙ��7(&�J;(h��}�`�@��TF�'�������XM�9{CMŽ[@ޕ����޶�)����ih��ٹ��� tf�gj�q�S_㌴D�<���j�_�t����t��h�݋b}|���Jm�4_~�)�˾�$�,�X�2k�����瘞rO��]*�c��R?�<(+�צ�a�X�r�ss��}�c�Q��H�*�.�t��M��Z{�Z����3sc33�#���%q�8�3:(3��3a��h����L�j��$�?�BS˰���*�Z��s��[�fW~\@q\`v���+R�?���f�?爲�D��T֞;�`�|=VI(�<�]�(�*uY�3Y��sBR�´ya���*.�2io�v[I̖Ҹ�K��/Uo*Uo,Q}_���P��+
��>��,�=���FU[�ыg#��v�N�V�H��+9��V�l.K��4��ҸM%� ���]%ɑ��N����O�ǆ:�j+�6\j���>����/iqy�W0�����_~���Ç/^��y��󟞴6=��������`_���դ�!�v�]�I��,[g��6J?�j>����������DtX�`Q��We�����쉊���yq2�
:�!qH�|�GA!rՌ��vJ��4p�e0�����䌦��{�4F[HrR�ˌ&�	�����Bgk(m�{�gt�Q�<�m2d�dI�E�)� =@
�w�ƛC��C`��`1}d	�qJ@
�<0<.w���4�t�������p4_�W�hp~p�����>�8U�V�)�1��q�,B]�WP�����M��GZ$�Q���PE蓢�SU��:���֖r���  ��IDAT���QO�T~����B��׾��+w��^:�*',gy6Qw��������&�]Fjʣ���@�d���Y?�l�k�#�k��fҼF_�]�_&G3봍] twOs?2���я3t��߃�@� �a����z��ʽMA�lD(,��t��D��_�&8#!J�&:o>)TTܺ 0@Ͽ|��޽���(��[��I�Q.c�s����{��#f
��C�J�-�Vo������j�,��b}��P�5���n��ԇ�K��Y�Ac*���b��}#��"��!�Ys�<XЪ��Zn�����k�xp9ʪ��x0kT�gu ���L��LN\h��`MTg��c6�	_���˫���R,m��`@�C�5�W�>$���^N�W�wH��Rw�9�r�::r��Ӿw�L�{�����w�0��ݯ�/^ON�il)*�=i+T�%��"S"b
D�eTU�wiܮ`:zs�P��e��6W쎊X �PErTىR�nth����F]��xCzd��uGwV��yKU��*b4��lv����oKb�)҂�ۊ�˓e��/��Gvfdh���څ�5�3�O%,�߯�.�/�����ⴰ���ً��_����/����ݽyڹ�A���wݽ-׮;�'�D���e��d�ZT���N��� ��%l��SCM�d�j���Ҥٛ���Lі��/HT��l�٥�Vq 4W�������4Q+�i�'7t4uia>e̙7�І�W���� 17(SlF(���?�K�b�2Ǵ9,���j�~&i�!�z��zl�F�C�� ���U`�F��������C#=����]�7��j��ȽR�Tq��.1ą��f��˚FY�T,�,��Z�1L9d$�ؐ�8=�%�)��PD�!��Q$8�Գr������m�Bk�� ���܆�V�~����LW��'4O�L@6��^n�u.�`F���kSh3~p��a�)h?�BG�lp:��iM �����'�U�N��=D^���7(�(�>X��k �3���Aj�ƚlp��d���эr7�=<A@���gb�0ȓ��a 4�!p�|��@�&�jT��!骈�h�p�x��R��y�~w7����!LOθ������eꕾF*7�:!�d�`��]�|����ɉ�"s�f�g̽-Ȳ@�"�mq��cS�����ڼ��_��</�(Ъ��&��s:�'f��g��Ɗ�cM�js���q�G[�㍩�5EC#,�����<D�����٧��� k�7��>�U���,�Ъ�����oF�F�CS�����[����b���}�푦<"��N����|(?{���w�ސ������_`�r�c����={�ۣ����7�E	�<���ം�آpeuB`�m����J���?�kI8פ�v��,��W�U�$.?Y������W�Vq�r�����c�kҶ�P�3��N�������~]��m(��>_{�4ATx�T���=>��y�V�՛�ye��v�^n��f"���_�7o~}���˗??��ן_�z��������K�.T�_���k�Նpo��+�|=�YIQ�:���
$3X��iX0,��䏶i?4-q^Y�C�R\�
���*	��h�A6	u0��:Kh�=�3���@ZN�~Q��B�h�f����J�1�c����⺘c�7��E��5�a~�	@s���7�C�)��u���hjVbP���.���aT���{z���䜯Իrc�'D�"}\�QiU�X���c,8C�*�'+��y�D���"���A�:ࠦ�����������rR���g���~N��C���c�@M�ΥݸJa�<�<1�O ������P�@��K�U �N=��Y3 i������L���`4���h�������d5g4��� M�[�� ����9Ё~_���c"2k$<d���Y�J5��X��ޥ�D���R���W�e�qq'��DgTA�D�I�Eņ5��%~�� #��0�#24�t�"#�RQx��?+UAX����閑��U!:5��#��bC�p?�aR���*��f
�j��'�x����P��[�Ƅ�ڲAVh��5t�I7)p&TU�G�Ա٧ot�M���-�a��[�r��m���ZǹR���Yp����mbv��a��[������9_�<l�۔�w�c�R� �1I�l��>�fD�E��"]m��2��%?dj|�Py�?w@����jz.�{;���sp��_�����}�nCÕ��W�ܼ~�V��A����O�����pXz65�\}���Pa�=QW�t��W��,��X�c�vK����λ�b���,��(>���`wkϭ��5G/��;@都�����)0�zc�����Л��v'���lr�����ު��Yw���{l	"�Moz����:���DZ޳8?�����W�޼��r�ҍ+W�W�Օ�_�Xs�N��D�ܩ�aUaV���®�
z�Y�]�Y�� ��$��q�̗�Y4_��;)>�Te�����*�Fb��:��w��R��HY�2����q#�,7j(�D�.	 �~�'q�/�@��\h�М�
(���gh�Z0'��@3SmR�7��Ǌ�:��F���ATW'����4Ou�T'4�˔}���Asw������w,��E��zU�I��4��,��7����OƆ	[q�8g\�]�D5w� �p�%1�����}F�$��@�h��_�W��S�bHi :��N㔺�G���#���h��
�q!��ƞ��˕�4�z�^c�&�M���}	�_���,�~X^w�}�hl�������+��X��PEد�ۣ��q���k[�FC���<,7���4�f��Ñ͝Ӭ�j�3A���D�
Bm{��^�ܖ �BeO9^�;����H�*�,�7�,QA��4�,7��9�ۚ���yI]Q�{s�U��MR�@O�9�>�;:Iъ�S����E� ���,���}��A�S:��@�*�~�V�����G&'F/�ܔfĄ�h,�����PC����clxbf��|&������������������lu�1������������8h�ݘ.^��%C����J��.s0�C���ZA���[��(�́x}Xi��g#�o^�~==5_W{�bv�;�KM>���Q��D�O;i����7�Ɔg�?y������������8S^ę����YU̡��=%1^5i��bՏ%�me���ݥ1 tTɑJ�zh����. }��j$�=���0����]�՛E�Qt}X����P��8�����㒬���e=�mC-�s�k��l��Ξ�7�"��o�>y�_hR�ˀ~���G?�ߠz�뻟_ܹ��p���5%兙��{�9'�:yx��&�,Pc. ͺRK ~H(h��65м2ǚ����s�ؓJN��Qe��6��.%:�����J~d�J��� �Ʌ9��`�>���Ml�M͌�2�����W�>x��2Gy�3�A�7��O���65T2X���k�	�PcZ�����N��\;{p@OLg����a���ᶁ���ݗ��ݹ��*N�1�e���Q�*�R�Ij�$���8���sX!��.�	���Ih.<�;l�U0�;d��w)j���$�a�YbA$(Ì��Վ��[�C�,�%s�����@������uuT7^K�?{H�Ol���U�5@�Ԡ!/�3���Y 3���B�Ӄ�r���7��`�4�N\ Jڙ�P��ؒ���It��b�U�p4�x��O^#���{)�������B*�,�[�ߗ��fO�`���q���H[�d��������P�h0���# #�̑��(D�G
��hݝ� � k9ļy�?�FM�^$ȃ��Stjnz�h?�0� �r��!>DP�[d�P͂��f��|I�E���Ե\�w�LM��	:��*�^��k�嫯I�t��i��?1�îT��ۡVG��a����ig��:�����ř��iI�5��S7�e��E�5F�0,c�W���x� �ʪ:P���T��:��z��_��_�uxx������t��f1�'��drqD$,�����W.��kbS�Rm�U�(�*�l�~��x��'W�*��E�`��(J�����[��X��P��T�Q��,�`i������18���w�ROuJݱК#{kR@�m4h,�w��"n�+����"���Xn_�|U��X���$-�8-�����Cݝ�K*mV�!��ݞ��g�&F�{���/o~&F���2E��M��m՟W�^��3�ֽ�������˗��/՟/�/.�q�o�UW��c��� ��Fj���Pc�'læ\mU�������c��"�>�-q��G�3S��O$���l�5��7�����ՎH��P	]���߫��L2���������:�7��PX�!4sA
~A>�� �h�g8p���}M�CjὛ-h�����B8A
�b��Ђ���ͽ����.��^�tƕ%�;��I��%>&�i�����!�B֡�N��',�x�p����A�V�=$��=	O���;C����2P
r8a0����hRD	���W�nt�NL�V>>=35=ˣ�E-O�����HSO_]ӝ#�&�w���P�� ��Ɍ��pd���!��U��Ay�5�;� �&�c3\����&��`�
ى�F�t:G<�"r1i{��/o-�>h�ʾ�<���nj!�#��*W�!CD�Q�Px�R��Ή��ٙ��鞩Ⴋ�tE`Fml�������Fd�M�<w���gx�yp�2t?p��ܨ�0�0@+��Ǌ���Y���w���pAdWX�4J����@P�F%��G���]P����ۑ^�D���Da(e}*������A�b,���t������'����1�+)�)�b���Ɏ���KU��#�2d���s���DsHi	���kL�O����	>�
��^1�¯�/�����c��UQ�70��?���p����eyvk�B.=�|�|"�r�T[qj�I�_޽{16�TX�"�G�(�.
+��U��V(�Z��]��T���@I���D%O���{�|�+��xHMھZ�@�p�J�RC�z�.*ߔ����*��a_��X��[�*�Iͽ���j�y�ܘQ�Y촖������
s���\��������Ɵ�g�˗���}Kt~��E��۷�^������4���֖��O*t���M@�A��D��U&)JWO��M	.Èєq���� �/�7��#���f�%�۞"�M;Zv,6SI�
[Ea6�s�-�;4H�,7���<>h0o�= z�.t�m��d R�܏�h�V֥�r�����+J:�����ynl���Xf>A�Rv�A0�E֓�-��GFY��Yg�16��������b��⛗3�
"3�Btq��4������N��U��b��>�Q�(Q2��R��v�0�'#��p�=:?��@\�%�g��p��e�&�ؖh�Zx�����ή�Q7T��<��
2uWc�\1.�L����}����֚^�㧗��pJ 4�+����!��P��g���DNg����u~�Ht�O��h��� �QV�P����ޥ������ ̅�"��ahB�~�vǝ�Æ�]�S�/$@S�	�ED���x<xU�
rS���2.5���ꛘ��]�Yx817���8�}ZtVa��	�0s�Ȣ	�)%ﲫ}������C#����W]�y~R�Ea�M���G���2O-���o�1�IMq��6R�DZ�C�JX�I-7'+���C�08:㘭n7*.C�=��Jn� ��X���� 8��-{���}]7Z�]}p�fG�ζ����[P~`��־^l����p�l�R�U�$���������������3��fG�O^��%g�.�*z��������T�j(�����6��p�zCy��Ą��d����Ƣ�ʙɥ�<���7��Qv�0XQ��-U�.T�I�S:�f���ʓ��Ǫy��pO[����5)�4&!��դR�����U4\���	��$��	�_��}S��4������1;�CJ�%䞽�z��|�Ң���gU_��M=���{D���i��@g��:c��7��{�n_�p���$�n7e���P,?��O�iWn��5I�[�����z�z�#�;10�Q"�ɛb'Md(�י��T{�R},	1%'O��G�e�8�j�d_��u%�
��!0��<E�Zh�xĒұ�?rL]i��(V�Ё��=��#�\�bK���#�`oBU=� �3��qB3K��>�}�2u����
���������	Cã����[[�/PlF�)�?C	�|H/	�))�	��3���:Uܗ���y�Su�ҕ�d@@R��I��Rr	�~�2C39�Ӗ%	�|w��C�|�X\�!��$	�����9W��v�OM�L���N��(�|�ey�X���m&' hh��~���6]u>@��m�1p'��AL@�8" �)��[�b��=��i�6�۰-9�y���ɒ�qh?"JR��@g���
��<X@�>�/�4�QP���W��;�A�t@3�	�{�(��'أ�'�W�
2��uW:�zG�F'f���g�f���Z��dǱhKr�5UmIR�I��e�k[�]��c�?Cc�5��=x��9��d����,j�����
��?>dʵ�/+�U�s��QWx�Ė^j/�Ry��~���������Ρ��}]鮬SL�E�C1v�`"�«�=�#�,��dn��ʪ+S����%�Y���N�ZO��N�;Ϥ��昊/_�����v��IԚ=>u��{��`�)�S�?�G�Y'��s��;�N�?'�@Fx�1߼*����Ώ=++�:wZ?42�>���uuw޹�P_V���	�>�|�0�jlx�q�^�u�9e���E�
��b��� t�U���� -)9^~���탂�kw�a�G��u�wԦ����.�;W"
�Y<��8��� ��|���	^%G�9��u�m�W�׹2��t9�s2����z��W��󷿼�h��_Ҽ�@�ۧ��E���Y�n�wf��}2?�x�FUyEEqyAV�1���2�!!ʨ�ϊ��(!:�e�XUkJ~�c��XU ����|����|`���P����-q�y�ó�R*Τ%�mQQV��.�ép@�P0&j<�q�]�[�7����X>{4��Q��뉴cF�h���FZ��QyY$|�����VO�Ĺp_ I��8<�L�H���70�10�*?���ހ�4��?4���S�P�8����7�|MRo�R�A;��.Q��b�RjИ T��<�T)^�ӒIݚiXk�.`Mg$)��Z��2�
�5자7@f�qC�h��F��5��P����:284./�/,�-R�?_ef��V�t��+����������<�tJ�ғ ��^�3����"�J��]�e`ڇkm�X���pE�~jK����҅�J���3G
~�<J&�#i9~�p|w�����h��0:�d`��x{,J}|��(جR9��77���L��O�x����=c�C�7zo�[:n_h�~��:4;>17>º�����޽&��,�`�&��h��[\�Y��2rrpfb`r�b��ort՗�������гh���Yp�^bH
6�|����"�}���<�38E}�)C�{���YFb�16ܨ��ī2�E�8�=$C�OT��kJo��t@HS�ZT[���o_�}6~�i�_2���K�hع���	��t�f��]�u���Q���w�޼z�K�������������P߈i��kf�2������ΙD��#��$�e���cw�0�Fy���x��䨢��Y��p׃���Ҵ����0�@�P��=�2iceg4%�.�'R��|U��@�!/zk~\P�aU�a���{��K3��i'��fkqg�ܳ���l���� �W����!����i������2�������Egss��6�5Ǒm��ϝ�g��8����j�^�ά��B�
~jӰ�:2�z�a�~&�Q�7�x�Q�9zw���#ʂcǪ���F��b :�f�9�~�0��)
`mh�fh�X7�s3hr'@�c�N}� dY��^Fz�!Q�꩚LM�,��V���X����4x�l�)��5V�.Z9��'?�R��(km���{���n[w��(���-�4�t����-%YjcB�A`�Q����NncT�#FVv�Z��'��R�&�rОO\)���t�B$"�l '�/<�:q]؀�-*8mr����إ>�(az��J������	H���I�M�2�C5���O���z��M� �-Õ�W�(�X�t45�$s����q��tb�:_�\j�3�^���4g&�&�D �DR ;V�OfbͶf��v9a��_��
�u,*s�v���i,C)
����N�0��n }�@Y����[=}]��|�>53F�.R���9���攔c~R�� ��pS����c���z��Y�oU@AGcϔ��Gݐ�8����p���G�����3KK���%�:Sӳ�3ig�Э�v�r�5-¤6˽��(�Q�$��t7�N��LBhO�����>Qd	�)�͔B�fф[1���!�<DP�5
cJѕM=}�C䤆����Z�[N�;%�[�B�/�ȿ�G|�}�.�?�If�<~< 0|���/o��2�1�ʴ�GN����3�;��h��g����ƬBrt-��b���)��1�_�]'+>Zv���ip�z�7��]8T����%K��a	�h�.���Z�煚/�5_jar4;��B�SSsN�YK�}\����&�W�ܙ����[�����o�>��ѿ�f��4�+��Upn��Ͽ���̳���׮�����fY�Ź�9v�!��-�(=%u��vh?��L��Z��fj�y�E�I�ϣ8X�5v�R�ʬX#��Y�_Y��N9SJN.9��R�х�1ye�	ԯ�&m��X�Q
o��
h ���Ɵ瀀Z�g&�B�Y�.��@2����%�^$]͔��B��Bi� �	nL��۞7�=@��&Y�������E�.�K+{�z�힆j�#���v��Vf_��X�(�Y&��Q!�/�����I��8���c��� ��1ǫ�=�)P�dY���<e��dF�� �٩��`^�YbO�_��=��?556MQX,Z�MX��x� �8�g0{o�.N ����z�,������ĭ��7�������-���� 7�ׇ��m�4Y&��#���b��ryIcu�ݠ]X�
�#[����P��R�����#���Tx���m����R�m
���g�*��[���twQb)\;0��
�CSC�#����wE�����r{��Z��|$@P�R�l��7Ŝ,5��C炼8��q�I��Y1����$:�*�%	�s�Ud��q��*}M�-5�f�Kۇ�j[���EQ�Y���_��!VI K	�9fP��.47��DA!�:4|��][d��ꃳ��@�t⿝�\���:�ɤ�q�H9����kҹ���O�;{�#�x��a���;�e-�ls�ػ�o�����*�+
��P�j�kwk����+��ǩ�OV�c.����ƞk�ֲĺS!�G�'@�Δʮ:�Ь��+6*-�/K�1�K���~Q�eA�7�����,L�̊O4'd93��N�'�6f��7ܸ���%��e��}��	��� ���Mϟ?�駟�6��Y������7oC>�9�ق�� ����Sԍ�';�K��"��Z.� �5f9WаO@d��:�]g׮�F�6)כ�7�|s��;R���J-LT�e
�T�D� hq�5*�l�lv$��=Ѥ��p_SuW�V#��>�H�
��
п`h�]B�R&Na3�ޥ7�D17�V���v������^W|���г� ��Xo��3Ħ�9]��3k��+�����{�F)��;/�=�}�W\i�SֺC�%ڜ�L�1"s�� ����RBJ�<f���p�80��)AD�������P?���rYָF\Nj
.��LQ�[��α�!��eh�:σ�|� J�:���X���+hh������\��\1̛�\@�T��N�dT��DˑC��z���)��e��!.E��Fd>\ۑ������m9�)e��Ϭ��@?%�P�
���f|/�/���?7�`�	i��,@����\�����:0�;820<��w�����N�T��Hʡ��~����ڦ��˵R�1?��O�lv� S�2T�9Rj�;��18������>w{oo��&�Ǿ�ю�����+�ٗkd��P�"�����}"� h�P�g�݅��x��h�@��zu�9��A�g�Q/ k(����BWy��9<�$����/�67��7���;t5�j?>-����/�#1������8/�44%�A��_�����o�2�guU%���Cm@��J�*ꪯ��<f�ef�3�@i,�H,����^E����{�4�Jb�J%�ꛯa�?�����\��J�;@SG�'4S�q*�_��|S��T�Ey�Weq�/J���!��*�~��)':�$)�}T8,�O�59�k��ͪ��o��6�����"�ѣ�_~y�Y�/L�n@��<�E:��|=&���5�{p�����|��J]�áO=qJ���ɢ��lp@S�AFgZcU�Θ�@g�V��Q�Q��n���ܤ�_p"8��*��	���L��.�ۥ2��٥aV)�0�D�vJ	͟3T<�(+u��E2SR7�jA"Ҽ�O��,W2ጀKA �ދ����/��S��#4W�؆�,3�`ʝ4u�� �7�$Z ���%�{�n��)��%M���������ww���N4��ln�q��mOH.>&w�B\+�(�����)�)�oĉ�5�a�gK��+6�EH�p���\�m1��\d;�w�ꭾޞ���F��9��K#����@z�3p�<�iQi¥qY��?p��\AF~|����ց�Tg�a�WF�e\2t�gّ�v&�{vY�Q����	��؝_�:B*Eڐ3���45ZLbs��a���-��j��2�ɬaP�X �	�S�ӏ�_ـ}C!�}��E�>%�UX�����}},�vOSo7�!?�z{���<*����_<R`>�.�2DA��'P�Fyt���7Z�.77^n�W�Z���W����j�[���{�����,��[�n5@�t	!E��6d�?<�^��ߤɨ+���y�w����~}[�6紟Q�cC�p"��=�,SwS\)�@F�Ș`9_~��%Е�������꒾�i?5E��=#�0�`��Nꗟ��hh�>�񓩷�~��ʲd��vt��v����a�}�NEQ��[�o�^�^<1�Z(=V,֔)|��{���E,�����nb�?�����z����ӡ���פ�I�Q���*��TM-�+������J��"���,����/Jb>+Ґ��@�y^��9��b�R�&-�w*5�Bu<�p����*����?���M�ߗ/������_��?��}�b���	�$�/^��#M����׷��ڮ]l(�˯�˹\S�q�H�������Vrn�g)��� �d���ɧR�T@3�� �W[���� �'��{[��Ɉ�IegNW���R�3�2�D���tF.�*\��B��һ�:��Y�@ �"ڲF?�LC �!�����j�xo��o�>$K�c�Jo+���n 2e�q��\",_t�(3�:�^���V{���U�>2::��M�1G`�ycr
U�)������������������`�4�\z�D-h�K���H�_�3	OVx0?)�F"�	������0d�6�)�]Ċ����/��7�i`Y���P��Ky�=#�����L����4�]k��jkK�++�(�"ý��$P��֬�8+�Yp�'~��6�9��;Xg��,������Y\�(�^�gMZ���^��8��Υ�wnXɔ;���P,������IA��w�e����g�5Dz�>z���D8��-λy�����*Sea������o_9[�s�����K�Ӊ-�~gd�:
� C)e��Uьa>�� �*.���qJ�O��Dg5��Z����<s�պ⛗�n4�4��.�L���K,bcBp�"�$�t�L��G�W�b��1*��97�U65V=h�xp/�|��N���A�A�ܸ�����E(_%�T]}I���e������܌������q<�ó��HV��m0(�4{}�.�z���o�*]uE9�9 q�G���m�o��������$yQ^��SWw��@u�H�X&	,R�+�(�9T�W�)>~��zp����J][���j�M��V���2��� zSU29�+�.��a��%1_��~^@���<O�i�����$3h�Ӕ'�i����'s3+��>���O�u,Oo߽��Ջ�O�<���S߽?a������ޡZ���ӗ/_�?�����������7�4���*..�˹q�&-E}$=90)""+e�5�+A��U�)�k��g0"�<�(5��?͌��I���h���mT~n���=���;v�Z����T9e�ϰH�$�N��:�����B�O�D&�$�C��ɜ�|4/Kl�MIG�bL4������݃թ��^�P�a�c�QU�R t��FE����m�EZ��7ݺ=����H�ٹ�i,��d̓8:9��[�]\��_\\z�����å���Ʌ�������,	
kt� �[��9�8�ٷs?8��	~B(�å"�@� 5��B�^N���cxot�~=4Ȳ��/�G=:59ʕ2�2���2�����&��ƚ{���4�-w���3�S��y�!�3��>�g��/�K����p� ���!��[wh��v@�D ����Fܧ���hj@�r���G�?+�/�� s 0�qp��Ѝ\��+\F�i��B�<7�eFă����	��52Gx	oT2�iu��8�!5"=A�O�<� 1�Ff$���	M��S����d��P�E�G�w^��Qx~ � ��3j#��0��[�Q�S��p���s��������� ��N
�@�Z"a<� wV �t�~Z�p\iKW;trۙ@]�A=�
P�	��}�:%)������p@�c��!��)Mn=j<rP���\��S�?�`���b0��l�z��>�]#�~��ś�b��7�3���M��4�k���|�v����~����|GfA��Hr�RV���.��/�K�<w���E��M�W.t�N^J�=z���޺#;�9�x;!1��ME,������b`�k>+�BDZ��$O�>K�I��s�|s�&07E��ѦȢ�Bc"��3f�)�����orr��/��d�$������Ϟ<����U�M���9���_�z����s��W�q���������xӝƺ�z �������si�g��"C	;�گ-J��O-*��U�֢`g�Y���3����*;��`;�?��Q�Τ���T|N�{<��쉊���ڸ��!瀎rЀ��v6��%�3�c�����xF��FI'��O�Wy �=i��C�["�ë�G��$z]����l����tf��3���z�M�K�#���49��&.��5("-'
��6���g�g(m#��ܹ1��@�\POM��/,--=z����i�����d�����Rp�TfՄ��K��'I���4�ӳ�P����~r\[�/z���ywf����t0�˲�-VI�b��J�,I%'D$3���$3��$�������*�{��}s_�g9���ʈ�ݿ���k���I�-��Ph���6���8��K��rK����3l�eV~��x��������p4c����������FW�]		�J_��cUs��;��[��,B��B8x���,�(^�B{��7R}L.u��/�́K�+�o��_l��G�7aU8;�*�X���/�>��m&�*5J�Q!6j��+�{�f���?]��J�W)B�p�"ʦ��am
��E5����R�m\Aj�E�_d�]rJ��&$Rߣ(�skݔ��8֑#J#m�(�,�.���"���#'�ےY��?�9E7���a��!	��Yh�*̢�iq�����K,�7C��,�4>^bsS�֡P"Z���S ϓ){�&Ԧ��r���d*��˱���*O;�!�ɪ��w��ßVW�vw�^�[z�k�?����s�ٛ��?������jsg��Vv�Y��H!�iP��w0���7Ǻ hI_~H��8�G�Ч(�]��/:!��G����F���A:j0����h���oʍ	UYZ!=;�(�I��ntݹs�Ek����'���yP�Jxe�����|���w �ov�(c�����}�˟�i78��fύֆ�j_Ukc���.��4Ő�����8��(_չ�W���sih��W�:�wb��'( �E�����������keyu��J�ګLq�H])7�N�*�f0�h6�5���uF���~B@��5�̒+ u�*�lHhH!T��Q�T�h���Lald
�" ���@.��<�����\��.yH�<ޖ���� i�m>��� ͤ'ж�� M��߽�p����� ˛��ɕ����rA��R$����8�A��!$:�<!�C�_.-ɉ���P��"��0�a=�82R�'Xӊ����/����F�`�.��vw �Kg,؍����"�˯&���_�b,) ��e2!�����w�L�%�L�}�)�a���E���Z �� Z��N��m&l���.���MB�}/�+�+���A9���MSdQ ��m͓1��@U�q!�����P����s���5A�V�z�C[<��2�N�sQ���:v�KdD�O���O)\H��5�Y�6δ0y����U	R�N�bG�o�b6H�SBT�~���&٥�K6I�]����>��xZ��	����'�e�g���4�'�6��h���/G�+J�VD���T��D��X~�i�����~���?�ᯃ���ͽo����i/�;K�5<4u��ә�ep췿}���W\o�H[�A��� ��F^Mܿ5ٓ�4�;?�������}ӕ	@�Οu��0~��l�:������ر��H��>U���������x1ה�X��T���5uv?Z^����������_�]p��,���O�q#�����B�������w5?G��N�WJ*sN;tG�!���w	B>C)�����) 2K������8�?�˰��!t��\_��d���[
ڊ��S��U�L;�e�s�'%���`o0�lė+���i��ՄE��������Dg'�o �,�1E��#�%����Hb�@f������C:&@���笱 5��g�I�8^b�N�{��(�%!Vu�=�}���������ED|��;6
�� ��c���wP͜�o����@m zlq��q���"UX�Z�@�E�N2 ��Ǳª���#Џ�o�X45 �d&)����`E!������޳ə��E>���:�ղs󫤛��x zrn���D�������P��&�¬��W-��K��9��A�aFU ���&M���U?̊�Q�����C���yh3�Ť7����fy &��XW0�B^����.��"�� ��s?;~U����,���8m�(����t�J��s�^��U�)��4+�;��%��jY..5"���0\��S e�?[�o&x/Y�WP.'���ώ�n ��S.�p��\��xY @��CHWf���������g�C�+9ޙ��V͏�s-�ɠ�{E��e{�d����E㥌h{}ٷ�z��?����W�w���7ow&G����Օ��oW�7�?��Y�����_�����S+�V� o5�BM!���tC�վl�X ��䃛ݹ}4'!%���9ӝ@����2鋎��;�@�#�d�·���[L������\G�T����t_�3uyy֬�O�;q*!2�$���[g�T54�������W���_w���{�\���?���ˋ+O=�w����������u��*�ҍ�W2MRI�)֝�]u�*�gS�T��r7�I;s�Lf���s*wF��$f죚f�u�:S#K�����׺,ٵ��
�YYAtN���RT�3KM΍���#�0Ģ)�׉W
,����-�Hި�AÀT��J�F#ȆX�IR�c h
����h8�e M�k�fa	��(K�@@�W��42wq����ڛ5���ݻm�g>
�<ѻ��7뛻D&(���X( *@տ�b����M��i�c�~@��B�+ 24�|Ě0���?�&QbPzJ�úv4���$��J�x��J��xxhv~z�������/���Ú/�4��������aߝ.�ms\���%�Ӗ�Q�.wn@�N��(�EiH�8���v:��;X?!%����F��FӣP_"x�Ǆ�u��,�Ku��X�!K�o��:HN�{��:)��+6�z�vM�:K��:��OB۬����H��m���A;��tޚt��ZS�3��<�߅G��Ȅf��n��x`=@�7�;F�TT�%q�j�ֱ��������`M�`EeLڅh;��4�ЌBc�9	��Q��ubIG�:
�����Z�O�'��PL�W ��d_�4�i4GU�T����_��w���]]�~������>���͵�w����������Z��~��﷟tz�e�u��f �`���6����8� ��ܾ����K��;U2��L�|>ޞ@�>kO=�n�Q[������������9�x[6��J��Bs�B���Q{9��,˝}���!g�%G&^�-,�&TW���|
L�|=���?��7��_IS�O��7�_���_��7ۛo�=hnlkjh���s�+yWmkQA�F��U�d��${F�7��z�Uv`'�!���碁�ܡA�Լ/*�7㣝y̰���كc����!��+oFB�EZ}=���rk~j�Q�Q(�
�Y��)��)��:��"����z��b�c�v��Ǻ�`� ��uÁ��7���42�J/�0Ic(���x��VAjrwP��g6�xץ @�p�aӗ�0�V[n�995��I����6���v��f
���
KݹN�?�D���a`9������̄��Fb�ǹ���M�Ӓ(fA&�b�a����6�]A3��E7�I>�^(,�&�M����a'@%*%�����s˳K4��{�y(}`@��v� h��2�����<ϫ�G[��6��5A�%̥t�̰M�Q��mi�M�B���eC��x:�K��u�y�N�@kS�52L��bѺ�E���Y1xF�Y58y��梛�R[q"����i�;�}�:�p��D���"v^-�w���,��Y'���tb�\5S�{u�Sr �,�4��uP�#7y?hH'%/$b����'~!@��/8�
&���+P��S�]�,5��H�dO	`������"N���`�٭"])�������E4�'(�ߡ�煉{�$ �?\O�����]Kx??������K�Ɦ��߮�n:�-=������e뿋������������c3(8����u��FQؘ,ka�n���ƴ��{C�A��cqn��j��םؓs����� 폴�L�?�0;bt{�Vӡ3���&R7>iL=Zo>PCRz��@��@���pޛ����Rh�>�u��q��Q��F]����n����wdp�������g�6!���6��w�ˏƄ����?�������7C���߾y���C���eBI�%3=�dJ5��J�*�����+��ē}�i>b�dK�+�H;;(ؙy�u�?�|�?J%ʇ��R�3�����c������'-��(����Tr��(�ڬr��9|&K����x7�tP����X/�@~^k�;�c�2�M�O�f)C�,/���™H��ɅvߏRG&&�x>h�[H�	�� f�+�Ng/}�S!�����&�i��ۭwo78�aX��l��9rrl��R��`�m@|fi���`a�E�P�:��%������%DK*�)��� k�Ҕ`��4WI�9��0k��RD��ZL�����ϟ<���XX�k���慄��.���Z��YX~=1����̞mW���7X�:�v L_dӝ@A�l�c<�3j:X�f�4���&Az��ޔ���ˑ����.� ���*�jP{�Y6- �i����(�7N's���O�'@�7��S�#�?������7�&���Z*h|���84M!�� ��N%�˂a&u������P��,<c"P��\m���X�р��g���}\�5��/��L�i�lD��V��":��Ag���4��@X��N�dQ����.E��Gb��S�EA��Dhgb����\����� ��3<���o�67��׵L����w��/���̿��Y^"@��CCS�#SP��+/^�y�5כ��&}`��k2J;���E7^0������������+ 4���l�����Y:���3�.20�Xg���40�`31�`�q�a��@��`��@��`�a5 Mv�R�ߧ=��|�1�Vd'���}�Y�9�T݅�_�O���]��j+���}������N{{mmk_߃G�^>y�������?�����&���Ǧ_�|=z���ڊ�U��i�T�����$I�3������D̊�e#�Yd�l
���KwЩ;�^A�n��C���dCE���5�|T7�|��n��ʼ��"EmAn�5�1��S+�r��ig�,�-������!����Zpxwɜ��!�^5��aE�܈T�ؘ@�.�E��S��E'^t�,�㤠W&B��2�4:����b�L�Ӂ<b��%�iL����s3 �1�����l�Epp�I��k��`����a�/qe����읡G&13�.E-�{ah��KQ�$�hP�QWE���0AF7��t�z�P�;�3J$oO�N����L����('ep�H/�"�b�o��1844�8�@�C�h�e�/$;�4-��=5��rb��VW��)�qM�&�O����Z#��(����;��N���6�h�@3�r`�t0�����S折�β|�ΧmQg� :���Jt�H:X����@��*v�B��\�lF.��YEH��N�N�����SAJ�a����In((	�݇�|����f"�������KB2=�3��풅�H�"֫��W���64��������/%8���J��)c=4n��:XϦL�Il`�:�n�FN�PeG�Y}��/���RP
N��[�[���	>çy�]K����{I?ˏ��@r�f˓���w�߾�����ߣE��_�r���w��7k���?��?���[����Q^���v7�4��4P���d�i��7^����$��~5y�:?��rP_^@/t����lp�hl ͤ��5����������};��W���
�A���K{֛��˽���v\	�8������K�̌N�x�������]Qnq�
J�6woG����n���k<����{7z�o�4w��j�gi�]�9��\QJR�cC/]�x1&!>Z��Y|5C�O*6$����c���@9��d�(:b4�B��������=�|�K�RmP���> ͡js@��W�qWZlcIJ]Qzs���RC��YU��{�r��G��9�d�n�����5�$7��a���l��Px���K.9H���v�!4Pc��;� hZC�5HMR��O-��@��t��0�*������4MaA�pل�+����	Pܚ��Î���{�d��hyܩ���J���AGR��	.(_I��"��&�"�?���^]0�X�[��vMU�/�\�X�2�Gh�)1N��)��Q��DA��*��|6931�:�L��9�)5ď ���'��(� �bb���5٦�vBR�Ѹ�����dl�1U�=�Q�$�,�_D�@��8�e	:��`a�UB��q
���:�b�%յ���X^:�Ϋp���!���PE�Q��׾x7�L)���wz��>s�p���F��b��,̞)�ĉr�S��̩Kq��Ee����1��
�J�+n�"+Ez��(QY�T���E*ue��<-�.�p9��k�5� g4.b�(�R���b��b
uER'!�@�F�(D
2Aa�ň�XA�����)��D�KK��H�rMdyʒ*Lǯ'~|=�'����kIP� ���I�1�T�㺾��������7ߢ�����o���K��b������?��w��_Xy�n{cc��V��јը�o66�^j6���E5gi����͍��z�>ܔ�w-�/?�?�b��A�0��9܎wf}ٕ}���i��6ӡf=��â胍ƽ����Zn�j4{��Wj�V���kV�xU�ܪϜ��޴Hwf���#?v���G����Sm~^sQAcQaSqQuAA���������,��k+��%�����˹��1�B����	q��&󩯿R�Hs�25FU����Rn�.I���}���+�4� ��a�4���P~����GJ���C��G{��L0N�=���
�_�|�N����Pbl*���4䪽j��Y�N�|N��9��ƀ)�����P�4��.�aD�����h� eꁁ�|����+NǠ���JBa9�9�Qh��
���̄(��n�����2��|'�G��i5���4�7^)R��a��}KKK+++,.��}�tt��w�Ї7��+/���ו���I�S�l20�7⏅�%ׄ�kW(+�ՙ�.`���G�J.O-�]�x�n�,���)Dm����.U�[瑑9�q�2�f*h��]X�[$i��$F�$�������o��YXy@?wv�%ٵx"��'O.�b|��	�qQ	��d�a#ԕ��6�K
��AD�Δ����9�"ƹxX� 6K7�mp�M��{�g�t�a?9�]��I��ɥ�kq|���EF�J�p4�0֦5m�hL�,� M2H�pA#(�X#u�)�ⲣ����y{*�7{nTj�$�<�.�%���}G���y��ث�⟀Hmu��"���5:���X�ތx���b�`!��hj�W����h�<�����2Q�t�eN=hf'!|�����ᶔ$Q�p�5���N.�j�(l:�`4��0�Ө�
Q'����Λ�p���%�$�4�C.�ϯ��-�|P$��(��B�{���'}T�rܢ�ӓ�fז�g��>��X�������o߾�������_���������y z{{see���S�`07k�i�B�.6�5=�%[�\x��=?�&�w�4g�_��J��|��&��O�]>ٓKIG�X����Yo��4޵�]a�h z_�t�_������6|T�=Pm<D��_����t��94g�0ܩ������Cb�A{�Do�aWɶ4���a�ʱ_+h��k���5�.�;q���/��c�������w���Sr�R�tVw��<��Α���u�eW���
�Hx=9��)5(�3E4;��C��u�*����|z����^�{������4-!D�g.sDC���L�Xr��Q�]f�2�<4 ��9E�S&{��h9��QsM#�!���?�u�LcUX;J�;�D���W�(!������E1F�Nb�(B�������.o'�g�� ������d�x�� k,��6U:���9|�Q����e�3�ʔ�s0Gt�d��蜵����'/s+����<�GyHx �5�\e��jrt�Y�M�e����т$\��B+^����K�DA���o�ߚx�la�����~�םU}%S�6�\�K��L�8Trgzn�����������ܱ�5�}�.�>�.a9F�������9�j�5n?o^�/�y�!������t�h|��?D�-��=�z�Q|NB6pn��&S�,#�In��a��x���4�F.0�O�;R��9�9��C�;:���t�c�X�z��#�ˎ|kʈ�`U�5;oW	=�ڇM����O���m,������v��v��ۋ���L���}B���Y�W�_W6u�A�[�쩼3�����'�/{Go�}9h�����`p�'(�5��D��j���EkQ��{�f�pFK~��21��!N�ZE�I�|��p�����U�zo������g������#w�O=��������5~���Cߝsy�ҥ�{��<ʥ��0��kR ��R��650FT,��T��͒������}p�����D�\����w���?����o��əE�o�+����ڜ���YZ���d
l2AAG4fh�v\S3�/�ݘ�|нW�z�\��;�Mq� �7]��
�To0M�2��ΌϺ2?������:hTa�:�ЕzӁZÁZ��#���p�F�R��C>�'>�Q�����F�{�c�Yƪ�F{�<[w!2�4)2��a�OD^���U��s=;�≯���Ï�D$&|p:4!*�Rr�ܕ�)5�+�����g�A��E��]sHP�Y_u�4S��r%ܠ�G����¢�������j?�~BJ�L>~G�	��O���Y�]�b��i/�e�e�<*�G�&�(qZU�ͧ"d9���f�	"o�@0��S�>ME��9�Ƴ�d�EA��h&ax(���K���r��	Ls����4�};iT!xVzQty ����Y�jvuF���������*��`���lt^ZZ�������G�[^�@�YY���{0�,՛h�_@���SӨ���&�'M����k}8�����͡����pp���G:`FG9�\Z��S�����)��jcy~si�����Ƚ���w=��Wk�i]:��f�U<�ǟ ]�;����o���MB�ӝ҂�8 ����Q���  ���L1�N�!�K0�	@�CBᡎH�MQό��b4e�`�FC��v3�0$�4p̆k�A� g,��{��\�S�5n�Fc���|�T1أ)\�NϗCy��-G�	D k�H�b�j�+�w�q`qljsafc?�ڷ��nm���|Gi���}����o�ۚ�Z|8�4�y�����I[A�-ɦ�^&�L�hj\�]L�+�g_�,�̼Y�__�z|m�w�֓+j�� ��A��4��.i�S�,��w�Ǉ��'�,<�nV&;��E�S"�c��N���������7[���kK[d+o�qϰ�w��h����%�a�k��Ɵ5Z�ns�K��Q(�ˆw�_�|�D�^�����
���!W�m�z&''o�߿u��/��'��?����}��ǐ�l`�_��׿����V7Wh ���쳁k�9�ќ�LA���m
kN�nJ�5_�=�� =198<���l_N_>��Σ�нyPЧ{r@g�����������>kO?��W��M�)&��`��p��`�t���hNg�GWU��^�A�����Uu®�������Ժ.�U���d�f_�^�(��.ɱVZR��%�g�J���0-�$K"\�w��RO[�_Z5����"?�)k��HP��4��	�\5�<����}fq�8����0B�����P o�-�˝��>1�!O��H2T�I4� "��)�(>W�3%�%T�LF	����df}4�VF�g�cqB�h��7��}ll+y��A卋#~���D�fy�"�=Cj����Iv�d�AbR��5T�}c�c���4����O��@�Bpi��PG!M2�.�,���t?��s�&�_ ��@{"��D�Z��*�(��lv|beijeyx~���#��g��@ �+*���ځ��ggg�(���[��v�������䋹����Q �����Ɩ(3*�c�3q�jN�]@��v  =�� @�	6%գ.	y���`����C��l!b�|I :s#����.���y�}���q���]شfh������6r�7�X|^,��t3�!� q4�X-�ta8�?e�)9�va�4�G!����#����[�M��vms���*Mَ��*��J�9~�nac������ɉ��G�/l=^��^Ys��|&�U��K��yy}��ֻ�mʢ5�:W�S"��J��Z�$�Y�x�C�td�>�3�7k������YύF����PD8�2wv��3\W���f��~K�y�m�]���ze}߸����nmӴ �Z��sCb�K�J����'}t]ʆ�P.��d ��	{�'~Q���3��ף�wn?li�|5���R����TX?F��3�������7���[[]��k��6��o)��i[R�L��F�N�iN�6�����������=y��ɽW�{���rq0�����/�h�X�َ�ܞ;֑y�͟��p��PSꑖTl���v;�Vi�Vj���F0��t��0}ȣ?F;�V�kʧe)��)�����tm�`�)�j��"ŴGf�++ĕuѕqޙzZ4}e�}n����	��\��.=p.q�����b1�.���ip��g��,�潂X(�x*��.�g���U�%mvm�-��Q���R���.��E-) �����\>CS�l�,Ҁ�L%��u@���3LC2s��âݔ>���M��q�$��ÿMZB���	by<x�z��mrﺨT�ˤ�v���RR�bR��U��:���؜��K�.���l �!�Q��^��	x;�t~yipj���X	�?�%9�RQ�Zy�k�ѫ�������7K��4���������� �HAG2)M��vy�=��ɍssSP��!���?J����o�V�ޠU>�<=�<;�����[�Π���MY���v�=TZ��L,,=��W$	*|/ G?&�̓��� ��b%��|LS�!~^Fg�&�c[�Y�f2�숾d�����"���֜�|`Q �Ě�羔�S�����k�gq��b!��5x�VP]K>+J���J��E��Y\yr��"s�o�-�.mmr4����[x=5�lt���(���:ZQ���߾]�=���ln�Z�:7ڡ�t�����-�[X�?�o������퍧�#�5e�v5^� �?�nol�C�[k{094���]�U�Ù��&+o�G�u�ue�������ڦi77p?s�k���KcK���sKC���3�S�˨Wެo�Q�,n�>�z]��3��.�T0Р�O��(%tA��EI{�%�J����\y����w�״ww=���G>���������]��o��o����	b���祥ͅ��Mh��������mb�)�^��x��ؒܜޔ�l���@��ܙ�
ݕw�;���ꢑ����FՓ�uo�W]�l�7y6HDw���Дz�%��CM���_� z��P���"�@�;Pn8PN��C>��f�G�ϭ���P|,�?�)��IZe���6�Q���Muت<���9(ҬT��N��^�'�&�D��'^2�d�g�sDJ٣�n@�,kIM{� �!�)��V3�љ�>3qm<�1}�I?��Mn��[lY��>wQG���W��r�2�KNg�O�����	��A
�Z��8����aAI�K&y� ����{�9�y��74?����rS��.�I2���;Ƃ"��fa|���9���L�Uī�ϟ�
�斈�0 zy�d&�F���ʏ�C�N���_Y��]��HIr�%.��&3��zq������եŭm�  rEn�����t˳V��NtPX^�۟�,�!��J�kMMp@�) 3ͪ��w4��O?��;\�
Da�1����w��� ��bWu�]��'��4Ļ��a{g`��6~m@�����l�M�>#��(W���b� h`�N���D�;�fuq�����DĬ���j�#7�N�Åڎ9�cDi�������Y�B�aKko�^MN�y����oWs��4M((�/�~����~����Hh���m����ņ'�R��PБE�K�"�8������(h�;���@�1�H�Ɉ�Q�5�\r��[)jͮ�{��sh�ll�f�V��y��hQg7^o���������v�./?���y��ǝO�=zPw离�������k��&��=��Q���~��|}Mq�H�a�

�g���J��K`K?.��h"��t���{w�:o65�=z4���Ѱ�����_�����o@�w�������қ����ũ��uWjM�f]h��L��l M3BDG���?V�/�Lu_�וs�+�|��;ӕ:���=ѕ{�;�k.����_���HM9H���V��>mM���|��t����e0��W�BDSPt�	��W���� 5$-�z�Dj��h�K�'*��G\�a7t�n?�����ML�������@�Dg1�`p��X̼�{���T��`QϼW���4ӈA��k_��ákw���J�=��S��k�/��$��!ٚ�zE9�@0�c�6��Y�pz��C(	�B�&.s>���`#�m�m�5?�!�`͇�QDW���#FSC���R�wP�i�D�_�GAg����63y2�b�ȡLNglp���4/	�s$͔)v,�.N-N5�l�	�W��4�8tf�ժ{/�'g7ެ���[�\I!y@��幾W����$QFq���L��(b���������*����&�=��4c4l��4���o��h��ã86h _�#-�MN�Ņ���bgM�]FYH�r�!�i��\Z;��1�2�?;�N��g,���Q0��T3wn��f��ȲE�_�`1�~�L�폶�qYL�v����C��$x]b�Xx|I� /Y�C���%�Ţ�sS�xQ�U]poj mp?;� j�gc#b[��,[ZlN.3$���4�AaI+k��;25M�'RO�,�a(�
����q^u�� �
�=�)u���g�\�,�߽]��ݮO��"��6̭D2ڍ��hr]{49���= ���тf %��fkwͫ�ihz�VVg�Ŷ:iA��(Mf�H.1'��&��p��U�#�h�0�u�Np���3bK`��H�zO��gE�m���JS�/�~X��cQ����|M�G�W�ִTU4?y4L��ę��~Go���q��W �w����X��^�[�}>t��&�ؘߨ?_�9ݠ;�`<�d>�ln�0;}K�W�����ܞ�	ݗi�7���\����gz����9Ցs�=�Lg����Y_�����!�R��|N=ܜv���3�]7bt�h�z_�������
����&�T0v���O8����C����&�tҨ�qv<S�,S((m��?��F~g��#4s:��>�?�39䢙��2"ꊕ���V���Y�Qb�L�!�^��t��9�yh ����uN,���p��l0!� [�+;�:�ڃ�A�cY��B$���H*�� +e��c�2(��(�('ph�Qd�i�O�>�4� m���PЏ8�g���D��k��=�(x� �~�1.����gx3���z�����������[R��~��t{{�qa�sPY�I��y7&�HQ���<^\��J�XJ��vga0��p��Ú�/���e��? ���S@�{ў`?�ߏ̻��;�HM{�l���fH�"�\��
j��U \�e�?dcĹ˂�0��LAS��ܱp��K�,H,*k�g�';���e�C��:7�4�g��q� {�*$'�Uh�.�-�S.o<�������޶�s|�>���t�"��扂^j�̮*�{���/.O.�L,,����5�:��!� h���N�ԑz�A䀦��7�l�Qk�Y/l�=�z�Q�O��J�eE�hȫ����Y�`�h���c���V :ҮJ��l ��,:;�&�}69f�,�	6C��/��%����OG�Q�p� @O��ݛ��^�U�~_��C���Ȯ�a{�UEV��U�L����_�ٝ�ږ���/��($���W����nP� �o~����Q�������KO�5�&U֒y��Yw��x���L#M|@k���=;714��o�#��J\gnP�+g��``4��._��[�W�u-�=�lG0�M��-�O[S�d��4�)F���F�a�m �`��p]*ww�1�2퇠���+t{}���҆�^�g����G*�~3�ctp������ )�]��5%�c��Ody�@^ ��K��p&�.�gc���8��9��ݦ�]�g}y��6�����.����Y�!w�y�F�[.�dvRI�E9�(��OQM�,��F��Ú�a�I�����9@\�.�\�iC��vR�p�k��q��g
��`�_D��$t`�w��s�?RPh�K�_�x>;;6���2�����c��+��X�X��.���]�\[�����6���U��D�h�$ݤ��T>�f�Rf��&�
��ς�Uo�"A4�<���U��4�fs}{���渢�%�/�; ��U,����_�66��iL�����>/Ği��9ʕALd���ہvrh���"$-���|
pFgD�g��xʚD�d0:��N\?c	?e	;e?m��'���]]dC�fI�ɯ��P�����d�E�?ĳ5^K�#s�۞ޞ\�T��3�@�s�-o)K�cK5Q6���H<�� �6Ml�AR�Q~����������x�󇆪�p;��,ƭNpiS�i%� ��*k㰅םo�g�,w��#��l�,(h��TO_���/��倾3>�VYQ����	�=�иa zzy�ƫ�)��C�Z	n����� �]+/K���|59=���+�6]^����|b1�)S�ܪx�L������gI�#(������í�P�亵����;��՝���W��h,���_�~�O�9��?��/~����ف�ї�F^�~��n}_uzu����`�O��O4N4�N6��6 ��tE����p��cqa
��3�;���}�q�LW.�\w^Pw~�1�iu�梁z���ȶ���S�_�����іThj�Ҁusg4�|�5�H#�j�p�	"��k
�#M^��,;�Y��ˍ�V�~^�@��PZ�������a�+r�g�6EY��,�HM�4 �t�� ���\A�݇
��a8���C��M�қTs]��L��䴻����j�*��f\v���<2Й��<�Q��L�t��:��W`���c&�)�h&4� e�t\AsFckh�Up�a@�H�-�ʦ��ˤ�I<����Żh�k�E�w�Yt����ᡥ�9����� ����.�Q�9���F�"ɼ�<��`�u��o�}������+��[[�o�{�'�&:C>�{�
2]�����q��J�� M�;��������۽��3�&�2��7,C�\����+u�����{v�-W�O�ƅ��x'�g	�B�91��=g��4�
7��c��Dg!��kcm�8ڲ�I0�m�<�5�Fx�(|d�:��̌��$#5@�{�s�̈́�0J<>r���H���n�D����ҷ��hQ'3eM���#��XQ���=���c]�	
ȹ19v�N�+�G	�P����p�Fi�W�29�D�r��n��?�����F���Q��ы�T���v��:��8;=��Սͱ�9�݆D�.JT�Α �`jzx�b:���;0��xs��[m�E��x��\���[~���J��;�}�SM	��nKK����!�U��������MX���1�����\�͖���6�{6%�g��v��,)?/����d�ˤgE]���*טL��׊��5�ϟ����?�9������_��?����W���o~�����7������?��r�����[�=y>�����g�>z���V����e*����tg�����i �u�P�盌�ͩ�+���@����W=�-ٽW����LA_>ӕ�u%��5�~��I[�����;5��齥Q���m��;���ϙǃf�mK?�l��)�|���s�'� M�v��P�06z�x�����XN��KCZ �aDpp������1�5�Jrح����^v0X�b3�|,׿�Ra�@���i�1�:���G<�/���E�v1��w��S��nx�K���%Or+�To��4��/��{��i`k�hV� 1��IuQ�.�������r��
$���L�?B"�xPb:�DSd.
|��z��O8�Og��tƕip���WX7�7x�0��O�R.}F��������қ͵7[����Ӱ�������sH
�9Q$9��2��ˢ,����z
h&:�x����4@=ͪ(H��n<�c�,~cS�u5>���Z!��9K�3\�\%��?�t�"i$��v���AO�;k%�mvT�Tϱ�
Fg���9"(o�-�e�;/�c�
��a��َ@�(��f��8/���@d2Ho+����36B9�b�>e�ĚEt�Fl�]4q����H�3s-�������ۂ�_/�-I,ǻ��TYuE�f�hT�h���<I.3ŀ��JsaGc��Lk�q�E�QjnH�xK��uU"���Ա8��0 ZfOu��������Y�gG��9���jy��Wk�F��*�#��ѭ���9����@��T�NS�Ck5�uV��^�7rxje����`��hyp��9��Pcl
IY������(j ����[[X^({��uq�Q����}�&��U�_[R޷�>���Xd�K$ST�1H>$,1^��QXW�������_���,eێ��������?/,���ݾ���篛[�<�n�ƚ^��iH�3����AYPͧ���皍ͦ��yS�_A��/��=�m�|��|�=�/�^�r�����+�]�Rn��]��Vu�ӎG��n�ݨhκe�k��y�Lg��L0����O[IG�5�C5Ҙ
Fh0A;��à��1@�5�O;Tk��.�0�4���az׸�8p��T���GZW��Q<�  �Nⵗ ���|h�q W�X�?V�Dg��SO�qO���|U�3�ӝ�]n�Ye����]Q9���B5<�8����t�~0�����r�2�)�(&���EGJ�S(�`�@�$ȕ�+��eꔇ�e;�����|�,Z��	�a�̭,PT7�;�9��i
��hY�1/ޤ�E������N�D�Ֆ���sS�o y�<�-���8�8�w{!jPl����Y��B�]2�G\`ͼ��&f	���/��\��gW%�l<�W�C	���p{
޵���3\~�N��_΂�TG�����՝��X���p��������D�&��2Ӌ$��J��t�"shrY��b�9�h�c�Z��H���3Z�"��@�� O4w��D\����<�LAG�Nmi�
ψ��O��U<%7��/R��;U�vt���H�u�ma�s`nb�EIN/,?+k��)Հ����'� ��5�{a�F�
X�������!���,��C�/��q���Zϫ�#�8^�5��"��(�rbe����1-V� �Iv������ZE 4^-����d[V�UjS�X�eݵ�g�v���Z����)Ʃ��_l`4*$���V��q���cs��+o��k����ڍ���D����t���*��*?\&t�b�瑁���IP9���:�x6>?���_�����?���Ksh��E:����}����g/oܼ��zJ�e�եFw*�sD��d���Zm@s�Z��Y�κS�z �B��Ni��=���y3;8��k�)��O���Dt@_~@��K]W�{K��E�����疯�~��W�C=��݉�y�-��۲����2`���kI��t�@�]���u��ju�� �}u& �p]:�P-0�F��jwz�2�6�4��C"5EO��W��hp��x}�:�|�6��w�xe�W��>&vС�I�3wIf���{t>����܍�����������̪�U�uDg��s*�v)�vF9�؀�$�Y\�g1%�Ã����I�]/9h#�U�[��`4>�Ρl�	�
A�y3 b苔E�&Ua&�������`h��$)�P`7 (C�����A�1�p��D�7m�t4<�_�^7����t4�Lt^���\���_.�4*�������n}Z�n�̈́fNghL�sv��T��AM��׈�|;c�DA�^-�YZ�_��o"�K���s�Xf��?_p"�p@?)i�&��(�u��]ɬ׎�����1�e5""��gm�@- �m.�q<�s�Y+�L��AkS�!�>g	9K�gg�����A���`��� G\��|\TgS�N�CKY�!�Y'!茇�SƳf�8��qNY�ӘYQ003@�w�{;�<P[s"-�ч���Jh���<�Y�K�P��i�����;�}�H�2�a�Խ324����.���� ���L5�����+��D�9֩��(惤�l�'0�jn���c1��� 4�lIg���a@�K2�����N���PB/��E�	K��a��M���<�;<�0��򛑕��*�1�	M��.�GN��"t���K��&�Ȯ �?*K9b�����o4���c%
�� '@ؿ]�k��5��tvu޿ug`bjmnns~��K+��-�{�r�ޣ��]���?y��Ym]SFn�*U�ZfVy͒���Z����j�Wu�3��o*�gk�k����	����l���3���L��~�9ڒ�K��4�^!�F����kҾm�[�������rucQC����ޮ�^��zeGAXk����o(U�-�00�h�v��t�^@�7�k��;ؘ����П4db^����֤� ��}MVe�qeM�1 �X=f�fh�(&��Uc? �|Τ��W�1��wF�����������g*�Z,�wN����B�U:�Uf*�*�G��Vr��V�1nu�[M�:o���R˰�i�*%" �������WЙ :��@���XF	�N�K���q�q@C/����Y�W�(��W���I��S�9�`9�YH5_ø��.�jz��@oln���gWV7v44>�� ޿B�3qp��;@8���zks�\��5Fg?"Q�^O���i���	N�=H?V�Di�O���Hr�j���W��K$���s�֙��Wǻ�3���/���x,��p@����(2�,&����>��`��t҈`"�0g2j�2�̿A�(��'�f�Yx�!�g�!�;4��ѹT%���$��6�@�B��p^ :S�Qe�S�5.��?��:�����U?�8��Js0N�,�|��ช���v���oTE�(Kr������
ҫr�L�+�T��Yw5��j���j�t�"�j���n|����ȫ�9��YX�]\��_��]���{ �ŵ������)BF�]g�)J3[���@A��g�4�+�m���c��E�/�'8��r�XZ������گ��Ԗ�&_�1�M�NM��T}��T�KkËK}S�f�Q��#A�s��CQ�s�� mQ|
2��4靠��	�CV�6m���\�uI��lЙ��^�\��Wz����k�--7n�z^����u���n}s_W����(���[�$�J�5��<-��t�Fu�V�e��X���z�W�Qu�Ny�A}�Q{�Y�� ֜�i)�=��/,���|�6֖�{=�'/��
4�oP���}�e{GQUknU��[�Q�|��������vՋ��������Y��s�i�<ޚ�ys}�-���T0��hH�Tp��s}:��A�nH��a��"uK�Qa<Te��ȇ*�P��]@��󚣙��S��!�F��CU���Ә^&}�L;+�|���?dS�0:k�8)}h`�ey�����[n�Qm�//鲙�ӕ.-�,q)i� ���Gn%\�MV.���&q��",ʫ�vf� Mt�pv���	
Dg �m���qiC�&@�_���+��f���!'�!0aE9��"<x��A����9���,�e�����"%��c���]M4sF��s�c���X�;ʩ�4׹X��v�\%���t�gcC�O�](G8hx�hA��~���G�Ȉ�dXn�>���ZZEk_����#_�o k\�9c���_�?؏ �tb��^A�@���-���=�,Kz�}N�t%S��&�~[J�o%�E �r^gr8��cpE�c����t��s�hk���y} d�sI�i
�@91P% �DR���0bu]�l���6��E �Y?!Ȍd2Gz㋛#�4~umsi}}da��Vk��*�]jT����D��i�v{n�>^��~�0�p���W���:^ݹ��Ltb\�hQ��P���y���{�c�������Ff�^�M�|��)�!���[�W�n�y�8�WkK��P�B��<��t��bv��͏�i�EU�UY��m�N��J�2@�ili��F��n��� ��܊ʉ(�t��)�2ީ�+ow����nh`zpq�y襬�y�T�]�s�t&@
|�#(���
�G���æ�Ԣ:o3i��\7Z��������2�F"QK�:�&�lλr�4=��+Ţ��z�%;'����Eu�^r]#u��R/UN�ˏW�?��V���^;^���A�U���&�D��tkjDk����&�ű�8�t�^ë�����^��+�{.��|�'�=��]״uٖ��-ٕ�&O��Y�����}�yc�v�p��[NEwqhs^`[���l��/�3h��`��fa��4�?��|633�ғ��ưШ�J��uP��� ��ؿrq�m7C36``1Y��w����"�8����E:v>s/T_In��z|9}��֛U�[�%V�Ǭr�9���.�!����2jr���I;3����4�09�\��J9�)�(P�E��tF�9���nh��I��נ3m�t�(Nl�9�3�
�r�5�(�(�����L�Ν�I	c�֬�˓9P+��%��1������aa��zl47�x�-��޻"���/�9��L�cp:�W�h�8憋/��N���~�� f&�-�dzl!:�kPTd�ٍq���z����$*�5B0��|;�2�Fb�Ej�H�F���#@c'����_��E�9��O��4�EqPD��`8�L�lHK��B�@R�� @�9�j����W���V�I�3�����МΌ�8�.{���2_3� uO�;u!rd�΀�g����A�0G\$˸�&�;R!���͡�UА�W�o=R��h�K{���rI�z'����-�צЎz���۷�o�Q�R�ܻխ��幮�{
Of�K�0i+�U?��p��������������������ӭ�=��F���gW��ߌ�.yz��T����*x6=���nl��o�^��i(��Be�]i3|��ǆh(�ʛ�����W%�sk��J�2r!2@�����Pp�Z�g&��h؋�������V��h�ȭ��*	�P�n�A�CE��c��";dQ�����B���WV�
��'u�Mpb�:+Kf2I:�ɠ�NK-�b�u�[���2��x�9ħ;�S~V4+���j������ת�7�a_��i5|�@���f��
�x�ѩ� �u�4 }��2�3�峝y���&vj�sK;
��s<�z�Zg�1�k3�Wj������_�l{��|Ҙ�e��myg[��j���9�F�������(�7�3R�;�94�����8T��g�Ѻ�#�f�e|���a$�+(*���
Ho"2��xm�;a��@3D���b��]�c�_fBs��ۛ�_S|�����}����ͫ�b*7�J�K��Vp:�b�噉e�&^�S�ȍ]Ռf#v2'u�04�ɲ 2B�����o���ѐ�|"	Rл�̀`j��f��'��ApV��c��-
9p&���F���t�M}��������X�{�<���������U*?��?�
�O"c�������Օ����=2�
!���h�?5�NDڭIδ�&ǭO���	h��
5�Y]�!��w����²�A�=�Z'�ڴxp�;���1�������ȏ��1&l�	ͺ�r$q!|��ɝ�D����B�
��P7�Z*G��"�c�#�<$~��0�}dɦ��OlP�&;+���~lð��L	��c<�Q΄wR�3)�-KD�_�����P�x�`4t���!S�e6�U� :�����FWW����4�����bcqs�f��8�!ўZ��`oo��󾘚�XZ�|�bG��$��.�|�����so�^L�x��3ū���ɕ�7[|�������VGh��U����EƇ���k�QP��;km�X�Q�ȗț�,� ���K���
�k��ŕgs���OZs�M:�����"͝����f����/*>|(���#�|�]~Ħ8n�\t��.S�+�D��b-�B~�7��yR��L�Du�E1bj�h��2�q�q��9S��)?�$�Ƨ��c`t���z�:��u:�����fZ��δ��ep@��ޓ3�S��&�3z����c�TNRt^`畄�e]Na�5Gc��Vg��[j��4{}��6��Sl�Q{�Ս��[�=%��SZ��7�o�<Ր~�!������f���XI;\�J��ԙ���	Ӭ���������C3	j���'V���HMڡJ�6j�{3`������a�@>Xn����3|�OH"�EL���O�c8�6~�N�h(���snT^ﯶ�n�>h�ݫz�k�x��f����w=Σ`�R��]�0�*�AB��2���rΑ+�e��=LsF�{;>ev:4w�0�E��̠s�{�j���I3F�y��.���A���P�ӧ�g\23�\hg?�!WygK�]��P�`n~j��ڂh0 jt���f?�8�a\�r2�P�-�	�8h���Df���z��f&��)�����8E��(����	�!��zctp��4�3�܃�;�_�����~�]i��kCD��8�]�`4�4U
��|R.��,#��%�����ְ�B��I{4!�g�gs�s�ave��qYޅH=����Ɏ���P��؀���1�Vv�����7͜ZQ��H4�4kj�[��T&;�!���0w,���[^{6=��PkWF�Y��#	�w�G�r�< �9�H3�ů���E=[�������ɂ6G�h�she�l[oS��>ok��&�����F_��]fʬv��x�%���$��������3��[2��"�Ϊ+��i!��U�͠���X`U ��VE���
4c7zI\��s�R�To�:0����Lɣ�_��� ���4�?�?�?w(~*�~fK��8U�J�zɡ��P�����l�V��2��W%�S���E�3Ūs��3Ŋ�e�3�	���U���r�!��B�i�:V�9V��hBs���|�~�d<ٖ�M���t�9�%-�-K�|��������ԓ�� :�;�B� �tg�)Z�^�ȋ鸢��)��h�k�����*��JCaUjaUZIUNYM��]h}�~k�A������E�*���M��i_֛?�3i0i0���8������P�O�z\ ~�w���W�T�C���L�o��P�zk�_q��`��X�n@�n/�{x�#�ɡ�5�,ϾT}U���譸~�hvߩ���+��B8k��W�,����ze@s���3�N0�@m���S����4�����"�t�9�<��k挦�C`�D�Ay����)�Y(���є�Xg'w!��L8S�4Qh��و2��,&o>r����ى�>��1}Z�������
��1@�h����Q�\����#�a���ޑ���>r��FƼ��#�u�[�j�R<�8'�A��bs�3g4��Kt����}ï�V� ��j�ˍ5�ә+w~X���
;��y����66?wk�y�����|AH��%ϳɶY��/HA3�CO�N �9d�|&@���3v���p
����2����PR�6`=g�.=e���-�7���T ��e���q��;љ |��p{Y���/ڹS+.�C"ڕ�a�';�:G�ñ��]@"�}6=�S�1�ѻ���*=��[�]�^<��|��s�oH�JC����ⴥ�"�F�N����/�'�VV6������/��\ע��0�&�,5����r`dv	ߋ+l�{�My�h��w��[�>��VU-��!�C�z����WS,T�\\(n���i�~E;5T �L�Y����<�!�x�
���~���<���҃��k�>)6}dӂ��	��
�3Q#:���}ħ���?v� �?t(��=���E�^A~HP�+Y�-I�K�>s�?��)�#0���[�) ]�=R���\u�J}�F}��֟��ԩ>�W�W�L��/��_5�i6�Z�C[�U-��;ɒF^N?�'�u� ݙ{�3�l7�8�������mW��L[���R�_��\��\a�Ve�^�VX�UP�[R[��p�=����:�W�+�O�o��|�RK��ƌ�Ӡ��7e�>���5��� ���߇��9��g��
!���Zg k��c
���t1�y<�v&��2�3� +7�0��G|�##�|�<#����]0����V�׊��<w�7˯7��Z����+E�Q�|*�9�'�pS W�?(b�^��u��g�b�Nji��8PH�k|�y� wC_R�E�%�b3�,������)����j�����^J�o$����� �,�kh.��ـ���?q@�R�u�E��J��&��
�����s�4��(܍�r���
�ǀ�q������0@O�<�R��d��%h���1��t�q.�ʓ@���S��<��7�廀���5�a8\`�b�1��G���h��)��@5�"A̳V�y �R_6hx�-"��J��J c�_B��%��X�hj�� �R�448�vi0�@3?� �мk4�����@6�w��rw�g�O��X@�hn��cGy���c��4Ѩ���vw���V ���ڒ8A�Vp�hQ��$��rG��Y\\_���ŋ�	`n~�f;�y�B�����$��0$����}���iZx{ru��Vg|Ij�M*�����4kG���i����$�lL��߲̱�C�S����6}�M~�t�Q�vlh��
l �Ë�P�qVM�HMF���מk&�	qn�ĥ5�rn�z<��<��F��/ޝ�ʺ�r�ĸ����]	FS�� 4�b���M���x��"��#����J���(����d��b�1�{�Q��S��!������=�C^�Zñ�!��x���Z��j���Q�U���Ǜ_4�K�D��t{������Le����^N>�mO�՞s�+�\g�ٮ\�+!�����)y�ۯ�5g�ΐ�y>U�W�Wa�Re��ryڵ����|G���yW�轎�{U/�����,q-W.�g���<ِ�uC���c�����Pө`.y�k���\c"��F���e��p(���+Mt ]A�~|T!��4wt)O;Z���7�DE������k�v1�f͵5%7ꄛ��;���Ue]�Ԋ�9�)����2��|�.E�Gɵ3����a���܉ڂ�@3�N�T�� &~%�(�)�'�EG�E����4VE$(К���f�u��AyЙ�8����$t�/�S8�9�!v��j��ɭMv��q��0��2PJw�0�ȌHcS�E:��w��p��Xa�;=3���8�A���zW�D�т��C��v�(9%q ���n�-�3�Oo*�8�%�r��J?���C�)Ͽ1:8���̢�w� ���[b"������������s�n�V ���O�+�v9~+�CHq����,+K��'\��I8���1�8�(=I����,l�$9w�E��}N ���f&����*xGX�E��ϡ΄0y�8�w�y6\�ә�,���c%@��0�Oh5v=�?��0*0 z`f<��$Ѧ��(n�ॊq�(ū]�h�I,�JKݭSӋ���p���I�F}��'�@�����5��SkKU�:b�u�VY��CR�U�J:^�,��,�
Ќ���B�@g�["l� ��UnѧV�>���˶����a��k��&�9�4�y�0���;�AW�d�]X[�[^��f��&G�m�J�4�Щb�Y�:� �a?w��~ϡa��Z���N3���#Q�� ����8e�S��e�>vJ�{�+�G*Շ+}�CU�CUʃ��#��O�TΠ��z�F�gM:��	�m��29�o�0���������Wc:��ݔk�LW޹������uH�sӛr�R����+5�>Un�6ӧ��j�*����r�>�g�,7�AM7�����_�v�n�]7r��q���,��Zx����+s�5fU��em�g5��VCP�s'�.�ɿQM��.i.�9��k۷��vȣ?�3�y�xI/�K=Y�s�2/��$��zRSI��;�;��[�޻���e�֜�\�Ϥrk�f�[�R���(�.��H�Z�Sj:�Y��c �\���!c"�>������x�{@d>Q&>��%��� G��₠Li�,�Ɏ�Q��-^T�b�E��S�h@�à�	�b=����)I�.�6��Q}��ڒ.۵�Ҍ�|��#�2�A����e��D^��o�aH��Դ�fQ�*hSb+�0��o�z�@;,;�&p:s#�x�ξ�@��n{ԧ�q�A��3E �5�2�?����ͱ! �z��_�_py�I'!�L�����b�߾�Љ��2�����Y��Z�M���O�b��|������&A����@-�ʳj�|8���s����g����18�E��8oRӌ�\A3�5K:*��T(�p�s}�HD���%��ԑH.��*L��X�ƈ2�+����ṥ��s�[Z]�u���l�A#�̰�@'�C���4Iņ4���W��%aж� :�aL����Q���
-<��X}�#��jW@����Z�!E��MU���@L\a}}h�S�`��9�3jJ�,j :Ȧ�����U�������+�ou$X�av��K\���I�6�&)nX+d�=�Z�G-���>��203�88�v���Ц��q���Gl�i�SEy����D���������~_��>���{��]R0�c���G��+�_�8P��_.;X	�9\��Vˡ��hW����_��N���k�lɔ7_��	���F����n��-��B.����g:(�]t�դ����+��S�W��T����t�*�\�����^���ә}�4_jzyF^���Ng�ӎ��;]��^�����>���si:Jb�j��U���N��&�c�XM:HM�f�O�����5E�U��O0��t�9\N3��`�zLǼ��ԯ<��Y�u�d�ִ>_������[u��u�Z��Tݫ�ݪ̭�3x�Z�^�RR��[I9��!��]��&���TD� h�k�a�A
��)�� P1�,27�S�mp9�!='$ð@��'���M[��m�ެn7Z�*��ņgmM�rA)�q͋.Dw�S�/�Q7���0�J_^�����S�k�#���^:o՚��X	��o����� �^]O��S.�bL��B,O:
��Z�73;A��?���俌����Y8������EG�jg0h@ё���--MO5��L*S�F �9p{4���@"I#��w�������%��Ҽ���"cP�ߋ#9S�6�-�j������ZXx8��J�5NP�@e
�ѐk!��3��0 ��툪�@d�Hs����\>Q�wV�p<�<)qF���pn�f�f�1���]��}�-R�`g"�|�y��F�0��<�t)�6�a!BLb�u[(������F%ٍ�８������ެ<�,�����D���Jp$��dTX�C�$�R�z���́g3KK�=�K�w�hKwU�Հ�g7V����_\۠�,[�sˍ���L@m�(?/����M�5-�Rh}�plaie�k��L_/N�U�[5�6E�]U�*�l\��|�e��g߬�>��h3D��P;IG�����qP<v]VE~׳[c�ӫ[�� ��������޶�K���G���P�F�cڡyߥ��S�SuBG��?)�s��;d0��N�X{�!}ߑ�����(����PV�+WͰ<ҏ�)�}
��J(h�}�Fq�Vq�Ns�A�e��X���F�g��/ZǛ'�S	���)��o�N����'#w�_6�}��W��\>Ey�sw�X�@5e�Wir+��>�ɫ2z��r���OÆ֫�a۫5�M��􊜼�²6G�ö���=�w��﵏�)�ny\�s�e�[��ꯜ��:]�u�&�tm����/�Ra����M��&�����O+��|��+L_��/7}]n>Y�P�P�Z-��L�Zf��^�[g{��~�^����aW��Ά�mU7뽽�e�e����N��c�0g�J�R'{4����lĺ��=j6"�H�]`4�?�d�QJ�'LPv$�x;%X�%@3�d@�����glIg���)�W��^���ى���wo�]\~n�V�%p��2~}|W���E���8[��A����o���N���h�����X0,�� �ԣ0K	��l���^F1��R��X0ME��\E��Ӏ,# +:>��`��OA4.K��\��B%�1FG� �
#[8�q$J�����ɉ�ކ�2e�@I��"P���6�"�� Af�pjdz��K�a���ҀF�_�'@c���I�C�Q��&Ʀ�O���Rp Ч-4VFj����1p�� ,�06�SrhX¾)9^�uI(��]8��3�&?	;�lY(љugm'������m��ſBn�Q4ۖ-:�� m��~0/9�9�a8G���n ��(�4ަ-h��=<2<;?��F�g��X���S�S}E-��Z����KE8՝W\�x<6�G���E�hfq�����vo�E.hbl������~�- z~s��Ԁ{ɪ:琟�Kϊ��6�%QQ�fp�<��ز�Wci}�6�_-Us@G��z�t�,��>q����;�UbF��œ�s������f�߮y1�race����w����7C����Ţo��Y�GE�!Q�߭������ڟ����20�|N���C�s�F3}-Ş��r�3�=���A�>0��'�}��}���'�T��U�T) ���}� ��p��H��X�t>Ҩ��I�e��Dk�ٖ�K-9����#�9��&�����v^�r�+�lW�3my��!������/Wh�+�f�\�z�c�ڭ�x�d>L�Uk<j��64��g�3k._m,v�U�=no}�{�^�؃���u/����/���w�]��ב�Z]w5��rpuNpMn`u�����Ui����M�}��Y!�W"��4�6���)ڬ�NGzy��ʼ[���Jo7��W>�nx������I_����[;:�������Wa��%-��믙�f��(wk%n94���$�.e�[�xxn���ɭ�:����YvB��8�/8S��U3('�������IA��gm�s�Ȋ�:ТWU��]���~���_~��w�k���W�l�`��<��p�Ank�u��6}~����������;h��Ņ��/r���,ԍ	
���f4.hvQ�~rC3�$�(�<�;>R(��4��g�v�P̯���f�: ��h�4���{
y��"�A3�|&��3�b��]\z99�訊�E
�Qe;�t6rݖ)�sZ�Gg�vo���6�t��a�����;���0e�?
���Ą��!���]�X�~�E|�:c��gh7y�/�o9�@N�-�_��|YĴs�yGτGS2t ˿A<a�k|p���ř/��Ph6	Kd�%R�E��XBq)�'a=�l�"�D�=
�"�z��GLc����kV탛O''��(6cimcess�-�tpq��Ѓ�g��/o�>�n��p��y<���$u.��Z�IU�VV��L�d4��m�Aa�I-Y�/�̬���o�6�ן-��׃���v�!� =ec�Ģ�)Im�skbaO�?�^\|pa��[U���qbTIj�þ��yz�뛛���W3�W+��L����*���r���=_�Z{���-�)����N-�<����w+�z��ڢn(��t�?u���{���9E�1��O�iQ�g���H��w�~�J�����K��gN���=W
���У�Ы����Ag��)��+e{�����*Ձ��j��Z-Y��P��P�t>Ҭ=����lkFpK������� ����ܝ�q��|�-�DK& ؙ�q� ݒ�[mέЦy�&�ح�8VyT*�B�+<*�WM�in%�0m��`�ҫ��̆��˹���JŮ���/o����G�7ݩ{�_����������A}ѣ�˷+3���>��˪��]�����W��=l*y�j}�&>i�y_��^��?��=�|�U����i7$s����-���w��z�x����g�ƞ>�����,��Yu���Ú^��ti�N5�	n�P��r�(1.K��� '�`��@�
 5wh8�������Χ,Ph�h4�8Ӊ�vM�=���Ñ7[o��}�����Bۃ&�U-���d)M��lP�0t�k��E7�_�ln��xqg�V��P	�X��6���J��I��1X��up��Je��
e���T��Uл\CB9��\`�}s����y�|agЂmGNL��N�`~$>c/w/�����b-�?���&����C�v!�h85JSG3��� ����4�]@󏄆��ɥ�g����2~�4+
�2H�2���fh���?�E���o�a0h�s ��L���P���� m��HP3�"
�`�����a\A_����<�:�̲��d�dTm0?8�p@���x��!�K�䐺��O�-J��Hݹ��4?�w ���������֫�޾y�[z���j�bݖVA�ssm��H\9�%��!ђ��6��2�oa�ͳ�I�+��E}VT��KNؒhH���*ʞZ����9J�BU>��rvy���t���2C������=���������ֶ�_���o��k}��`�������*	�o�Π9p�?4;�����*ϭ��k�O֦�g^�vy<��D�>A�NQr)M�v�a?q�b�G��[����{�X��R ��n%`M�����K^؇>	.�TМΐ��0 v�A}�Q�Y���O؜F�n-�?9@�^X� �[^5�v�G��]�Ч�sN�e���s��.'�fg���Ԧg�� hs�V���J�h����«P�4��5>��B�.�*|Z�G���U^0������*��j�����+�ַ�����?t�o�.����w�_�i����V���M�7�n�j��5�hyu�[��{���v`�խ��=�O:k6�<l�ޮz<�-�����#�xo��y���ns�ۭ��aۿx���[��w�KoW��̾�}�󼧴���4��'sk��X�&�M�ISǻ��� s*�\r���'�Ĥ 1��$��4��%��&��|�h�AP�w2L��P��\�~��<K����~3�8\\]b���R.ة_vɥ�1������7+�45*4�̓�WW�-��(�-0:����N�.�2+9)_���T�'G��$����$����1�FI��a+��P���d������b�������/6��5ft>.5�0�xl�z�kW�����e4�q��� jA��`�p�)�����;h�]�7b����6 �����{�5��a�\���Jf%���u��L9/F�c�	���1'�d ,��In3�S�����n�E8�YG"G��Q�~G���9q⌡9gwK0�"������٢)�M8�����OHF���x :ܞe��Yt�����gOǧFgX��
e�苷���ېի[[+� #�YZ�XXb1�4������Ɛ2u�-%ԣ�c�鶞�	
�$��̛�3#21��������x���_rj�l�+��wF� P�l!����NV>��cI�[fgp�}�+��ݷ�߽{��۵o�W��Zz�����:����ķs'�0�<4X�T��{bpv{c�۷S[�O����o�:s��4JJ:*(�w�?�h�w��_��gN���rq8�-�Aj�ئc\
?��������{�a�k������5 4�P��h��y��@�
G4�6j?k4|ݚ�MK����l ���☛{<t�c�=�� ���y��=ٞ}�3�tgn@G^d�Մ�L :�.=�B�V�3z��r�g%�,s˒2�m�v)��,��Y-w��8�W'��S<k�G����FC��\��V��Y��_S$v�<]�꾪��M�۞v�?�i�G*�5Y���A��yu�g�F��>Ԝ�[��46�m��U���X[m���r*��}�Fw�ٓW�Yswf|lmmaso�����w��q�hpe�|���wh�y�fbe��ă�'��U9RQ/�b��
c���7���`�:̫t*��N%(�2:'��h�(H@�@����=�%�>mO>#H�>� �%�*X�E�e׾x�bfE�~���z�iY[I�Ud��é�biλݯV���߮mn�esʍV�hN*���)�t��` �}X�qh@9h*)Q��p7K[J�ui�U�(��*�0�u��D��.�ÿ�"�/�����>����/�SP��)������A	@���Q�P���E���`�i������Ԉ?%���)_ؿ�x�7 �����
��t|�s�%ަ�S���[�����3c���&`�2�
p@M���*t&#�2�m ��y@����h�q�eC.i��c�1w}�3�h� K(tt�-"�r�t�FC]H,S6e�(5T?���a��L�d�4�$a�i�ŔM޲��7����c�v�-ӄ����L����-L�<��z8>��j�}�G�)-4\(S�m���Ƌ��WK8qjiehq��q?��Ey�.=#ȁih��.��m�i�9�����`:0=w{t���.�j4a�2�b�i���/��x'A�%+�[�ŵ͹����7��%���T�뙙�_����m�j]��^/nnl����_y�vdk�f�^�7�3Q�_�p4�� ϩ���T`��?�K~"J� ���d�?9$?�~*&�F��
���c���7�c�lo�|��@��H��`��p���A�`��v����hM;՚~�5#�9[�t��zvv��������(���|�#��\�Ϸ]�h��T���|5�.5�Jg.ט+u���P� ��)����(uJiۣ��Ur�6ŭ�h��y��S�UМ��J���,�ܔ^n���e�2��3���+W.��7������Y�����rv;,-e%��Wk��V�\��ˮ�Ȭ�H-O��Ɗt]y��<3����كGs�xcV�FE=�Ǝ�⩳l�4���
���߾}��������72��*�^U��VCA���2ġ
u*�k���pH�)�g2G
�p���v��uHNI@3䀎�6Dt�Wl�+==C�����o���ޮ>�~b�#�Ɂ6�A�l.2�YnM�NoPe>m#�S��o�mi	vM"'��UN���I��_r�\-��$��7�=`Al��Qج�N��kL���ɩ���ڞ���솁���y6��!Uv!�x����� ��T�?���k̭��Nw�7�/ǊJTܹ��>����`��\_�`zt�M�E7�5>ss����Y@p�����yY%�Wɷ�"�dl��]oW�ټ���4�:���>b��#��~�o�TXm	�6�9g�?Q\��w�%9��J�.&��=C���	�H�8���Դ՟���+".	��5��bt�~�|�N.�5.��4�e,�
5��h�X1&Ɲ튏F}L2���hJ�i��X�R[Nqkm����������1��3�/'g!����>���;:���i�۶�myqx��R���E�P� �!M�`�jo�?��8>�7��rGyP�:����~^��C��,�j	�u\�9�����~߫���Ǻ_�+4�e�0{J�]n�'��5�<�FE2<;76����zd�����Ł����3���g`/�f��6?{x�ΝbIW
�i�ӫko������{hc���?X�:&��;�{6J�����{�?�K~nK��-��~.$�#ְ��t�-����W��4+y,��9��#5Z�����TШ�:����cM�ϛ�\>s@���(���~�W�/'����;�AA����O���'�rε�q@�5]Ϊ5eVh��=H�YU��{�2ct
,�%K%	N�ī�y52�:ť�:Ր��4�s���5C��9����X�!��t>=ح���fCy��"5�"-͗�U���IK��3���^�ѣO�0�H��D�ƫS��5�fR�^����^��ē���3��Q_MO���x11�lb������)��|15�����_\F�<�������v���sW���I�:u16PΤ�"X��Y��3w=���� 7	g��S�����B�1�ӎ���!H �!����X��U�����в�1�>��s&[ea�D����gs�so�I�,-���>�R]�X���K��Ia"�b�fcR�Dg6@ܟ��ڟ����
���A
�V[a�Y�z���y��Ќ�? ��������_�Џ �:`�f���j�
����r:�@g
,C#H�E�������T^��"-�?�	[�#�G��{�p�����2��223�xx��V�`�E����P(\�T��'��0�� ����?�-�4���He!п8���Хhp6 ���2�҉��th�	�������A	F����Ab��0G ,@ӿ ,��ÂDre�>C]T�Rܤ��P��'A�(g\��0�50)f�aSPy� ����K�R=e���Χ���~8:�x|뛯_V�w^�������z/ו��D���5@�%���v��A���Up��2�gO�䅖�c��ńzk�7H������J��i�JsM��ZS�/Ζ�@q�(�\i|�%��5)�L��n��<}���q�g7^��|���Yͭ~��E�j-m��^]^}�F��3Vq��j�/Œ_fN���4�粫�a`z���nn����������ڂ�I�W�QѰWTCG��R޳K���=��=;p̑���(�G�{�w$��|�b�U\r��,���ҽ^��r�H%���*��*�:�Z�gu0����):�%#�5G�Rx�5SУc/_L<hl6u\	o#�.��_�fݒu�93�5/�6�Ψ6d�����SPU壑�ˉ��$�$�%e)	.�x�4�-Kv* h�hhj�vS�{r��T|�w)vz����F �q�[�ҿz5 ���7z��ƀ�W�v��njB<�-W)���ߕ�F�`��3�j��7[���x���n��gw������ ��8z;\7:���}wz���l{����؃��G3ϧ�痦�֖�nL��t=�ڄt_f�����CDYt��wBC>S؆S�⃿�An�S�_Y/"pNH��ˠ3c:E���%�-ʢ����4���糳<�lek��n�EC�04������e4� �Gfg�:���4qh:�|<U���[������<�442i�h�;���/0��ʻ	�I��Iv��?2�H�!Ѫ�h�5���6�u�G0��>b��O��^{�V�d���iNmI�U.�.3�9��`.6BGP(+�������
X�yUA_��$�o�/~Gʿ�pp�m� ���`q�Kb�ǹ�80$=�dT��8e	&�L�
���\�筡�,Agm��a'�a�/8i�8t4�72���B؈�rkX�`���w�N�|�N!�� t0��
h�d�G�
�"a�0:�It�=S��(�Q��%�E�>�#F5,��Ib"��Rbe�U_��;/gWZ
�}e�u������2C\	詋*ӆ��#�KVU@Y�9��=ƃ��&���#�Ü�0�*�DT��k.���x��|���yVN����?�Ҟ������?$�"���ҋ�M����W͉����g��{�����U��B]LYzRY�R��s]�:�U�˱E��b]t�.�ZjH��ɝW-�QE��RM���qha�n�n�����s�k��h(/ooMn��]��r��մߦ���HT~�P}$�?�I����E����=���S���a�����e�l�@O�ȑ��#�ϝr�\�I��X������ڣ��c5��j�_������_5��i2�jJ?ߘޜ�m-�g��r�Q�P �~�t{���gZ�@������T ��SiYߠ�\���;�a`�ĝ(s4���!�1 jЙm(�h�W���:WJ{�k2�[)���^@\)u�!�
��x����Z� 2hN5�GAP�Q_��-Ñ8"]��@��h�)ŕ%/�E:�ʚ+/�T�eɭ�h��a'�f$����b�P������u�>'���LL/.-ln-l��m��V=����(Qꠖ�/�o��\5�# 4^Y`uLcU΋I��	d,,{�ؒ�	��r;��#�8T��9њ��r`d��i�m��Zq��U��2�����É5������i�� /�MA��%�`1v~��B3���? &Y*�L�	(�$Q�hQ�(\�{^/,�,����D��.�WVi�B�,}(b,\2c���&�o���K��W [!�&'��vs�b�m�s����9�%;�Ze!�2ɕ�94�r�z�PKͰ`^Hi����gZ(�yw�ߋ����zu��e��}4���V�Z�1�i.A��8U�0>���`���W�*d�8`�� 4�L~a����� �F��+�/��%�h��Y,`�Ǝ�
#���l���a'�L"Z$v����㠚�:Ƒ @�HA��Ć�RJ `ZH���x�:ޢ�/3Ɩ豎�P�F� ��рq�X�s6��m���ݍ��I�&��jl��"�/9iO<-$a��%���y���x��������A��Ҝ��������w��0���!�?�.��ߥ��/�S���������N�r47��u����)�E�H�&�"��)�m2X�]n�E���M*j'�*�e���u�/_�ΣQtm���d�� ���6��|�]��*?(���GZ��ە���e���vPT��'*>�K?�I���t�(��H9�Vv�>����k>��~Q���1~Y���x��x����֌�/����a���V7�fU �WSO;G� hH�����_���`>ِҔ_}%�6-�\��P+���B�A)�9�<��1�)h	�D��81%ѥ�%{4�r�C�+���Q@6��ie�5$�G-q�A`
;a�:��JX��8�v�Z�aMGzI��ʉ.���ѡ�%ٵQK�X�Ø ����fah�ǉ�xќ �)1���QP�jse���ә�������������D�<�A�x?!9��Pl�� ��#8��tpB;P�!��M�(ꃩi4��"���u4=�]�\^]���vcby���.���~�dr}u~��������%M��m�]A�SHb�Ô���3��C>�=���&� �Y���H��#P�]�hQ#.W?���5b1�{�ͤXY@G`fh�����A	�p8�0~�E��������ٹ#����x�6L��'���llz�;�MJ@�f��ٔ�ʂ�����fG�+�Q���2�__ª���lRr$�&'���r��Lnh���
X��bl��Y�\(�)���G���!bX�B=r�z���9;A����`�A�7(��b��jY'�K�� (�?U)~yT�Dg@ygNn��\"� �vF�|��ZC �\A��Q�!����=�	�S��#����� �b��X|dC4��P;�P���iF!%�&C\�vPk��S�r>���*8�>e�?i�Ú"	�o���^r�}qR�G��%��kK�'�#�d_�靈�Q���Ku���;�������K�YN��91�g���K� ;�ü��/G��������������_�/������}=�bIBPYB�5	7&�B�4�x��s�ahi�4��07M��PD8��.�B�.l��|�j`zn|auta��̬���O�7�ԯ��o|i_{�Nx�N�g���>�K�ڛ�����������|�m��s��Cw̡�̩�TT�9UG�q��K��G��W�g<Si:]a>S�z�*�35���3�֦��K�3��1b}�>�T��t��d�� ݔz�)=�9W�t��k�1=3�b�q�dwjW~hK���, ��T�.�krR��dԤ�)xX
�I��(e����I,i2�M�=1br���1�s]���b ��U;� 4(��K�vɈ��p*�(��� ��������k"���'a|��D���!K���O\
�5�Bp�j(k�0��ƺ�qnm�C�RE:�Q.5,ƥ�I�Ee�C-c��zO�������糳c��#�3M[S}I�&\$e�B2 ����Att%�e=k��[�_b쁁�,̃��l�-���	x��6C�	�(Ѩp�=y4����f����nkm{iu{��[�%�]^~9=Ry�9�T:j$�w�3�3��cԉ��s��|��]�M� 4J)ڃ�b��+ z���.�I~e��h�젙����i�h�D��]\���E���ybvahf���d��_Ax���\NS)�)���o@J�i>'rq��W|�o���>�~>1�zz~dn�ƕ�&�r�@�ئ��쀵uJ�ʃ�ۛ]\���zv;���B^XPid�-"T��Ћ�`��bH�R:���g6Z�����]F�P��ȶ��4�
�JZ���Ɵy�Ĵ6�7�XJ��F��P֡� hR�"��p���v��0�fX��:�h��\	���XWl�#&�!��B>�� ���a��b��Y��CD)��`O��wUL���-��5�a:���ĳ����sJ�dƿ&|Us�0bO�ſ3�����������?���9���]�=Z$�ڦ9�4]�ANC��*�� ��U�iI��q��G��ܐ�����3���oe_8Qy�,>КdO�)Av)J�%���Q�k#��OҩN
{FqcEϋ��&�N϶�0W�	��q�y��y�-9��|Ew���@�z&i�,m���~&i͓�\Il�NlΉkȌoʀ%4g&�f��3$�Y��lIsvrm�[s��y0U�eE[��='�-Cі���T�����R�ӒZL1Mư&�F�|��|�!5�)G�T����8�fG���onӷ�AA�j��_A�Ϛ�?kH��6#��Jlu��鲹:�X�Q�Ni��!��L��cD`�8&Y�r�ь�9M�Mk̓@�$�1`:�ԙB`uHi-�E7]GL!!�;S8�9��X�*;I���+��ӝ�x�����;d#a��w�j�� r�9�E:�	r�H�:�� �+�y0930??���d�EVe�D��`9��"�%����hc�́s�/���sw'�k�iK��2�,�.	5�4]yكɩ������w������򻍷�Kk���7_>P�ӣ�J4�P~x�<�� kl�-�t��&!�B���ؙ���H;���@H"�ʊh�31Ʃ6�m�_��_���;
|b���jA�8CGI�ҿ��wƀ@/��/N���#3�ӳ<B���x���WZ�Qe�Py��=]l$z�+>̝ XS��fN@{%�a���-�{�>��58�tlfpj~rn	臎� L��e�������%+l�>��YƭB�А�C3��/�F]�8�y!�d�3L�/؂�b�q>/���w��s�a��glԑH�fø/�X� ?������|�g��hV���8g�������m�$������p�sD���l����`��+���䳘 ��L�w%�9�㜱ю�(1
d�~@��9�씬����������Zx�x��36ܲ�Xc۞��7B����SB�YG�i<#''��]�Y}�z��0����������!���r�g%�s����0�!�*�{�r�󹨴�� �982�R��H�*��|ʩ��T��z�O�"�>'��/�7�ٟg���0�5����y 56�Ra��n�k�K�':)�E�̞z��U�~۳��n\muD�&\**�\Z|1�80��Bd���c��b�.a#�$$�(���.D��*<�P�q'H��qE*1BeS
��`�=����Ś����TWDnUB�/"�<*�<<�""�:*�.6�6��$S�Cͧ�M�����LMS�_AONAA�4h���ڲ 蓭Y��>Q��r5�*Sߐk�2k<�a �
���@!�ޛ@���	���"E4@�#�nB��G��4Y?���y�"љ�DpAX����!���~q� 
so��C�\�S
:�+����Ǻy6g�0��Rĸ�i�/��>��0�i(
˻���܁��ň���+Λ=���/ffFWf۟tfx3Ru���jړ��\���tg2%'b3�2b�kè�	�4��5�K��S�4!۞(*�m�%�u�w`aelل,�A������C��BL�2̞B��& ��a&|8�Q�y�C e�!G��e��ڙ冦�B,y9�
�����# _MA�[��F�o��t�i.�����	d�z�� ���q@yrz`r���轡�[�_w<{\���ۚ^c��P�@��[����X�ʋ
l��3�DB�y��B�>�$]�.�i���v�>}zodl`bfln�B�U&�I(�:�ĸL(�����7�ko��6�(��B�w�xz1O��ٿK9�3�W'��!A��{�%[p�� �71�#h�O[�ϖs7�6�{���|��G��ar��ğ�Gs�K���E��<z��7�`	e=�� 4�FcL��N�`{L�%��� ,�4�����#�#�H��ax�hWѠS{L�-���x�5�[妖Y�)FJ��~Q�%���دl	ǭ�_�	Ѐ5sz���Kc�.���0b��`��3��|����>;rߵ$��n���/է�˾<�8�;�;�`8�ԝJӞ5*O����h�	4���\�(��*�'��}E	����_������'����b�f~�$����=���ڦؾ(B_S޻QBmhQ#R�j��f����M���KB4�`m�%�%H��`N�������-!��`SQ������ @[x^_pf�`*�h.��Q�]�Wz��o/Ë��(�;�≂Y�����"V���c�ژ�갂��ܺ8S�*���|���h��ͅ;
zz�����׭����̓-_7�o���)�ˆL :�!�64��*t*�C��%U�P%�!�I���i�Y�)�>BL���|�U�Hl��1ɻ~�x��DIl@$e91��D��#kr_8�_/�,�ܮ�dT��|vW�E���V�Tܸ�HRd��� hsZQ���J���)�"�\)�b-YF�������������H�����+q6�>�dK
vP�}�Ҫ�$���ΡCb�NPF�$p�9��<�=-�C<%̮���G��Xd>닣f���T��2c���Ԣ� ��@��)�Y �I��̆wøvt��J�&X���h��q4S�@p���R���������w��[��m��9��6s�B�f��Kg��]X\��[��}6:~�ի�w�]�-��V��Jl�>�X^&�v�Q7&~�sː��/R$r,����3vbu��S��e��bMX�Q�+������`�]ٞ'�_�o���t���in�̽����v�]�d�`13�������̨K����t���|k�����̻��V�[>V*��#������-������zo���ze9<�2���v ��3�|x!H���K	���7�^�?����'�A���`}JYz�8���P`(��p8�����bq�Z����g��MМ����A�����P#�(�b�FL�`��$�u�p?܀Ѡ|n`+L�%�8�h��]ϱz�6t&��!Z����Ąkb1�� ��m����r��L�y�:����r:�S �`����Z����AS�A2_P�� �An�+ɡ�J��Iv����҈�̊P-����Y�Ἇ)�s<�UYrH~1K�V��+��
טM.ȌLK�%I��I�LH��t)(#EF�+�j��咞K�~*)���龜\V��Tc~<��t��j��b�e5�Q!jõ�C&XQ�3��G��%eYiU�C�����~cKG~skfk{6XS{vKgnggaw7�����������Ĳr1��³��J��e��riu���F�\��ڐ�֜�ْ�Ӟ�ә�ە�՞�ם�ߓ6ԛ?؛�Ց�֦�i�j����f^L��j��J��F�$�>�W�݇7�u�l��S-�M����:���������	g�N�*�V%צ�5��2!��&�i%��=(�X#-&�:ꡅ&���
�t D�Ԩ�*����{�%6�Ԇ�-A	6�ݘ���>�D-�|���I�9�1Ɍ�v ;�AÀ�dx9�vH�p'UvF���c0��F���@j'��B~d�bZ+ɯg |�x1A�ڸ���۳�졒��y�\ZmQK���Y!~�#��R�b�	�P�~Ԩ_�W(o�c�)$f�=�4��̦��3b�n����l.$X�b�8�Zhv�x������NP�[zr�	�L�0 �>0�3�x_|���
D= ��1�������;�Qe�� b� 6h���pFN���..�����K�#}�Ffqj|�<�P[,�Q�u�0-� �����P�y�0��#��_��c/k���0��sj5�gi�Ԭ�"Y�V�V߻�8�pnx�N����a�~h��J�v}�~�y��Ǉ����ݾ%� }%���(�Ii��ɽ�w�??)���Gp�-0��:O�@�� 4�r��AG�/b��.G ga�G�(jBOY����������C���XQ���B��(�%m#�@��F��b60�s\���!Fk(1Zj��J�R���*��B4�����x<�.���Z�;�	jx�Yr=㇇J�k)`���5d� ^� ؝W��L��t�
Z�:��&A�8�����A�K�?�}B�	g�e�4T'��~�s1\x���. uw��V[�������O�~���_��:^��4�[����q��f����[a9q1%қ%ҷ��/fŽ��|�͗�W������p�x��%��5 ��
"+ Pzf���0K�֔���o�;yp����yp���/G��v����΃��	�?�������������`���U?#�����{���c;Ķ?<���|���;~�?����]C��zr+��j��V�,�!Y�T0��%����sk�K-���І��ӵ��k��)>�I�P�ѐJ�T
k��"��5s�W���J@g���%�gI�?��2���
~5@ʱ�@[�81�-|R�5�5pbLHD��_��D�ɿm�a����*�����;�2���n`�i��;���"҄�z��&6�-��L��s�Rq���E���#��峺��]g�R��  �8�ǧb��4K�6>D��Fqܥ���B�K��IFĥ�ث�7
����P�6��Z�uᖚ����wl9w�y�;~�g�m���ϋԢ.Ypl����p��I���jR#=� �`H����Zh��@g���saaX4p3��~������wn�����p�!��� _|��I{��%}`7P��H����f�촺�����q�4�=�e �a��±I~�J�ո2���HD	@�+��kڸ��	�2�%-�� ��s�N`���U�ܖ��������MGo�kG�<��mß�N�k�����Z[�\[ۀ���}��۰5��^O�-�)!��(����I���
ӆ���n����CrS
��`��;T!�R!�%l{]����T��N�1�Z6�,�Y�*�Ef[/ k�q*
p�6�h,��=pa�{�}6b�v(�� �9VG��L=WZ��p*��l��A5�0��D��F�k]L����=�H!�":�d�ڏj*1)�T��4�-��{	��"�V�?Q�>Q�Ψ	��2�(Wuq�ԱΉ|J|�1�#�L���^>��\���8�UyJLyU��z��? �z���~|�ˏ?����_����=����D>����������!�F�N̉���
O���o��#-���s鑏+���x�BQ,Z���['	�����k*�-%��D�� ���|�%��nY\[����_~�����K�����:������������s:�������v���Gw?���w�|�Ŏ^���o��w������?����JU5+�����^�߬��U˘��#�����d�r��5 }�1�\C ��Z9 �b�2�>�P� �K͵ ��W�� >�=0���f3�&*�[kT:t(�����=�؉q��ɬ����>�* =o,Bx�X"��.¨�E.�Ǒ�^P@��Ŋ
���O�ȁ-`�ʂ��is���(��M"�Q�4I��
�Q��&���5p��\�]���t4��Śp��C"�;X�j���P9=3��^rm��G���YP5PuL���虐�v�֓.���-����ķ�D|珔�@�󣔏�|���W�g�U\;�u��j\�kha*!˘5f�9��} ˆk=�� ����u�¸��|Ӏ��408lkj8�>4�Ƨ�p���
d,�X�Ek�ھ�yo��=>��
�@=/���O���H�?��b��׻�pN����$��$-��� �A���o��pTH/���o$��;���z�n�����i���h��5�O�U�|] ����(�^�Xr���HD���}`�f����q�l�������ّљᑙ�������)x`lj���36��gq�k��ǥ���zDr�Q·��CB5a�ڰ�T����u]�`��;�Q44���0�ݑ:*A��[��]�����bC��cxڻ���2����ͨ�e�D-3RE��8R��>ׁ�4 ��LaC�`��f�8O�r��s�ZF㓮�!�P�H�(�P~/�D%)0�Ki`4�4�������oD�sdUI�=���u���1l(���P5�qAE�������g�D�߀�\G��#�Os�0�y��GW��<��|.)��N�Ey+�|�}��^ې{�`�� ���z_|���w�i��̯�̬MO��o���{�����30�>z�/�����ӣ�.�p3£RC"�i!%�T����O��>!��FZL�`侪�\ɯ�^��Qv59��w	"�+���g��R}Gi���N���o��~�����������~��,�z:{'��;Gk�����l�7�k�z��M5u�C�}�KK�{���G��������?|�ͷ���ڊ+�),B� }�V� ]+g�d�a��y�[3]��4\A#G-��tu�嚤��Tre��!]T)�]�lb,Ƚ���`\BC���· p�F�Ml _�b3l��WP�/Hi}���5cf��:��B�v1O1<���!
�d�KL����.��Rd	�\�c���V1�(K�+PXs�f��<����s�%��yu��d���
A�Y�[�=����,���h��5��"1�RX:26��]��}[ێ����O�I:� � ^ύzK|�1�������ga^|�}�􋏰�<ƾ�8��#�O�~���K��g�cAM�����eD����y�ǹ}�칷=�9�F�A�[�Pk�x�jW�"��P8�(��1X����<��"�p4*�X����P��6js8 �+&#y���xN,7U/����y���ln���9��V1���%���D- k|��Dn�Q8m�Q	@Ӱ�K��P;,F�n Q��(�O�o�b$�IzYR��ajrlþ�t�F�^?�����^���X[Y]����j������~�q��t��szph�����������4�EģҐGe���?�Z�ЭQ��p}8xvK�ҡЎ��!����X��6&C0���E���!���˶�r��G������� �s8�wl�n��W�]V�Q�SÍ�h3���H�h��T=?�Y=�5k����w�o�{���բ&5��F3�L��F3Q�F2�HB�֓�t���t�@;t�Qj�.�p.n칖�[Σ��ή��7�\��h��E��]V�ϫq4S����u�Z�i�^M~Dx��Q���?,�EX/ʃo�/JR�s]~���?߹��������{���C��ff+d����Ey�Rk]c}�ڊk�Ώ���c/��i՚�Ҭȸ����2)0��\����&���@�/F���h����#�8���@zp���F}uk�Ғ��o¹������{��݉_Ym���dm���$%�TU6&&�K�J_"�'�DJ�$)3����%7W�є��t���.����}���8��o������&f�Օ��&�^� ]'�Y+�S�j3&��=�E�d�J��95��v��S���%��V^�I��ˤT�H3 �3�1A!�X�5�� �3��cL4�с.Ew��F��f^$k� �^���UM�A��3�1p�	���@gT>��Ѐ� (�qd��G4'y`t3hd!�"Z�S�
릺�l���������Q�������P�ix&	�̆"78pi�� ��ENj�	!�FsBu�H�\^Uֱ�9�F����e�JY�����!\L}�w�Y�'�W��xF��֓ܠ��7���3��gAO�?���8�ʣ���/}�qK���"u�8uB����Av�\3�I�V��&��[դ�ɇ���:(�F.i��0Q���WlN�\՘�Ƽ�(��O��щқ�F���m��Y`(��F��nߊûl��:Q�Ȧ���@���< �g66�K[��$���fZ�F�ZK9�D�a&
 ��#�h2
LDK���ū� ��X�"��zM�Fu���C��]�N��
ɄV�jK������9�.զӳ�pnn���������vZt�dQ23N�@���j���֩�Ƒ��������ȗ�O+#���Q|�	�ٛE1��h]D�!2\�X�"��!�W됂*���䖆��,�����7w��s\CU������{�;�����'���֮shs<�.D7H�h-����Z��Dg-������s������m���������wv��;����)�m�0���F7����CMx�O3R��ɷ(�绖|[��]��!�m�**@z��}��_�jTu� ����3���x���ߝJ���D7�L�z-��q?̔x1!��ZR>{ۿ D*�ܾ71����[V֐�Q��H�#�]�u�����߸|�敠�X!K�$�M����A�+�`��?��YZ�$ω�OE�2�{*�K����t���PU2,(���jP��(�Z8��% ">5L�aL������=��������dl��3��6�Z�0j*�Ҙ���8����Y<�P��LT��yY�r�D��lr���)�	9i������ή��O`��g_��շ?�����_~���/�ίh�E hr��Z��!!�6 =�>O@� �m˭�����K����gk��%��I@G�f �QG��ea10@S�0i�|�pmc��%&��pn��,�6=r��
O�	�!u����L�i ������`�6^�gt�ij�/5�;Z9��G�
b@��p6���L�\V�"7���k&������;G{w�޽{x���]�>=9�{�{wkg��OfV00��H ��U?r�c�x�Q@^�ND�fZ&�F�%`�Ƿ��^�O+U��(�7_`_|�y�x�Op�����煿�	y��/�e~���藥�/C�O���^}�y0`4P��I��@��9��̠��r���B����(ڐ5 L��#F�8�6�����8
�Ct�Js�A��ٟ�Ǳ�7..L9<KϢݹ�p��;36�ĺ�i�g~up�6�ᚶyf�9�kv�9ks�m�������jt$�4V�K4Zc�_Q�5�\P�����G��f@3��5<QI
 o����t�|#庁tEO��Z���|6�jAѠMT���Pɳ��f�{�����k�񵭙ŕ������Zc�9?_ʊ���3o>���y���"��P<]o��*\���v2�oI#�Q��A����H�]�'���XCT�>,L�� F�h�TC���ҵ��\��B�pݬw��;@8�u�ۅ)^OF>x$�����A49v��k��$���C�͑�Lg���&ca����y
kV�ڌ�qp�*���ֽ�u,7h�f�@��( h���&�a?�x#9Z��r`+��A`���ڝ��t����moxp����{�3�U�Hc�^xSϸ�&�ϫ�v��"~���ʟD7�G<�J� �jN����ɿ��ȹ}�����?~����JIiU^nq�2M!K�	��	���\2�K���DD�B�������-�$���Y�%m�=�O>������U�����SoE�97��S���3bQ�z6������sű�Ԩ��um
�С��i
?cD�c��۷{��{���Wv�׏f�}���ι�Qkeg��4+�8)!͠6�WVW�-f�:I$L�qr�ڼLcQ�:7� -%��Q''���r�tQf������zljm}k���շ~����0���O?���g�.��i��I�lR�0�^�p�6!�&�]�3�����zm�"! :�9�rs�$�R@A_�J�I!U$����eb���.A�5HF�����s�B�j�-#+Ή����Krz �5�m"; �@G�Dyd�Y�%͏6"�0�1�{�	d��piP�1XP�}O�SM2�5�v�{�;?�:��@�w���]��^:ֻ��lg.���Cρ�i�>�2�o����D��c������3 ��L�(�"���cuy��^pz�]���IM�:X�&���O�A&�>'
��"'�-n���s��+2�5%��$�$�uQ�K��g�!O����x�w����P;^�,Xr{�P���߂}NiJ��p`̃�@�f-B3�A�13�d���GAu�dX#�k�3�R�&6��31C�	!������R?7�<3QP]Z���:3f�jѷ5{�S+,�����ld�j|�q�6�4=^9�o�mM�6���qEE�A#��6�� uq�8 X�~�w6�P5d�6;�jV�r���C��ߒ8��` ���#�& :ʄ�NM�	.9Ix
��W�5�v�h:������Z�b�a֚Y�@���������������������?��'��O���R/Wem�f�g�&| ~A�Xb�#��g��e���!�dDFG£�Q��#(�"5=�FiQtD��.���ߚ��;�#���7�z7L5��E�c�a��N���S(���p3ઞh��D�A��x hg�)7'���Da�eҾ��C-fv�O��Upݪj��l�e�2��d��Ǐ�L�x�8&Y�M��ޘ���]�����m��]��36ۆׇ�����iߚ�67X˺�V��+Ч�/'�|L|��Ĩg��Oe�o��g3�q�e�������������77G��H�kM�=e&KV��D]�YS����R�talL:�o*P��R�s���_}�=&D��]ci/3""#�P!?k��Oy:;���[�d�c1��U1p�2�r�: �e�`�	�ֱXza�P���q[�DS����n�{��m��u���K��Ԩ�]�=����ѱ����������C��ou,�����	<nܭ���D�
{�k���_�_t����{w>����}�齓��>U)?��K����V���W�þ>o�j]�֘r� �r�!�t��L��b���!MZ!�cy�4��,�x3b4��h:���5h1�'|0�F߅�adF�X�2�F�7 ���`���h�v���QL�{���Q6�igP�f�`1�ֱFvy����iF�(��v�ά�����������)�mhqe�昷{]��������������6ڠ4���4B����`\���w��vE�d}����kyc��\�r�n���wG���b\yIp�bNЋ�зQ��"	��4m����Z�6�hJ�i�J�i̻��W��ω#��� 	{A|�B=�Pa�Yp�q@{w|K��D�2N�n��,�D���������� �����o�ɡ�n#-܄ZIឍPT�����01TC
W3"�|�1�iL!��*1Ӑ@,R5R�FL�P�3���O"'0��S]�_,�,�D�#5LTa�q�㋁&EH �����Ȼ����KO�F!�Ŭ��eBz��:�W�2�%����ě��˪h̿�ڰ��Q��y?"a�o"z`.O���J�^cE�#�|,��3"�\�1s���є�Y����x��_�����[�?�������_=��_�����Tg�}횵����lME�Ei�+	aO(ßL�~^z:5�je�%�ctQ��(mD�>%^PpE�:�Vq8��f�w�O8�6��j�  ��IDAT��A)��]��-���r��T��`Ygy_G������ݹ�F�n�^��o�>���"j� uA,c��L ��h�O1Q�zAY_����o#%���/ٷڦ��&9���X�LM6�� �H�A���z&� ���^�8��-�����:5�/L�RIY�����5��*[QYZ̺TD��E�6/�(�����|L��2��t�bQ�Q�	�*;��d�����|��?�՘R�3�G{�;�9�m5���R\jx���b���)�]Ç�b:����[�5#,</2�R����\.�ɴ��n�Q.�I��A�_ԢL�kpu��XcO�WP��
�r��wtXR�\R�W�9]Z;d��ї��L %@ڿ5z}������d����d�IR����ШWN_�q)���&癍UmmCC3SSks�;޽�?����U	+��J��]��]�]���V������67��������KM)g���%~R�8]!�\���V$�k�E�B��9�e�~��~�6"7ř�P�0��SE�:dt�P�!��.��@��0�"�8e��x䣀���Fr:����|�40$�Q�J%�l|���Eγf��L������ͳ�_�X�nk��Wd��y��M�Ʈ֊����)]kcNuY���̖&t������c"���m�-Bb�8�Tc�"O6ހ�Mc����@��ݿ�>��Z�٧6W�m%��C_�<�~��>7$BA�1%uv熪�*����{K�F�GFj,Ŝ<�yܻ�7�q���_Vľ ]����m[����;��mۼ�E5�0�21g|��׌��� ���0��$�Ew`��ܨKz�v��Wи�����E�
y�X=?��#��)Q�f-����|=;�����bt�8*5����0  �a��Z�2�����!X.\>#4��b����m@u��I �� h�#�k�C��6j"ϼ��@�G�ak�g��T=�}A���7�7��w��	���������쭪��/�������߼��������sO���_��_�����?����pBж����Tc�������2��/$F|�B/e�M$�&2N��@���c��1a�� u^4TC���&�f�N��v*<2��Y�ߛdT�Shy
R���#���3+���ӛhas��[v�7����jf�U;�ԡ4�x���5�@��sB����p�`a+`n�6 z��Z�J-���9l�n���d���/nm M�x)Յ�s�>�͋�N-9�գ=Ԃ��Bat����X=1�f��q����w2���Tїդs*�IaOH��RF?�B|#�jN����M��=��/��bxd��H����8�P_YiVo.L��h����"x���_^R���շ��,tJ���RnF��猢��Oe�=��Nn0Ϭ��l��CY`���⍆��1����Z�N����T�^�2j(mW�����B��H���%�IS�Jmn���7��B~Z��O_!FRR2uZkC}{_�x_�������޻s85׮)a�WQ��⫕��U�U��*)�*mdSж͕����EkF$��:Z$����V\�K�V�Y�B)W����x
ܱ ���y8L1���
�\Q��zf����:�ψ�1F�L�l �/ҿ�^F)�(�����:x��F}㱢�x<�o�PA߁�D��_�U?7������98t�����B9�X��H�ZY%��%T��eH!�I*9C��nk�qz�ǨE����%ߢ�]%��-(b�*|d��,<%�($�bkQ���Ԧ{��k��@���� �u^ȇ�`n����;Q�3l��R�[���+�I���������)��k���$�o&^K$���{^v>����<�t���Ȼ�_�,&W��h=4b4U�n�#ӡ-��1�4��:��,?˛��4�V����3Ct(�� 44�d�P�z��
�b�9�0�2TN*j
��gB}=�4b������ο�U,Av9����kzT*��<!f�7��,��{S���A8�B��Um�6�x�X��̤��CO��^��_���F� Yݐ�В�(تJ����//�o��G���g�m�K���������������m��n�q�.i�Ai*�\\@?��tr�K�Q�'Qai"2��d=0:�-��E�����ib���)�m~r�	P�ٽ��{hnJT�D��81���B��C*	�yU#�ë�붹M�ĺ�un:�R]�	UC�(�>L���T�Fi⢵�����rj�����$���h����sx��N��ꢱ��U	i<?VK���t�(R�����k*��Y�`��� 4cJ?��t��yҠ|��|fP�(���cv�{=�n[�x{D>�r�t>��'eAO& ��+4��a*�e�UME�?}��w�8��ܢ�����������;��73�t��e6�cѕU�7�}�����pGgU0RC#sIe�S��g��O�D<��aa,����t�3K#�ɥ����AA/۷ʫ���f���\ޮ�U����-}�X��ͫT�w0��f(,��ѹ��!��Ԍ�쬂ꪦ�ꦱ��c��ݓ���F���ZF"Ԉ�WK�UInր����]�	�=�:WZ��u�Ku	��3���������UI��I hQMJ�63� c��X�o�5!��|ut���Qp�K�IQ4*s�Ө��ƱF�RA0�F�F�z��atF
p��
S��eG`�:��	#��e|l�O6I�d�pǼ��>8�9<�?8��ȷ�\L�+�:!\�T#��L@4
AtR�ANפH����{�:��y������#�\�GY�hB ��ӌ��x�G�6����o�W��U�cdeJP��� � ����6�O��[rz3�����y�x�Z�Z�<Y�8թ�L6&��~O�Z�e%�9�=	#��z���v=�=��.��z�5݆�"T� �m��DEquFz��� (�U�PZ
���-^��3�w��� ͋�V�vFb�q`�z��F*aF��FPT��;GP3��;����a�� �Ӏa�p$(�oP؆�t�k��B��(��6h�<p �B~j���U�O}]s���|�F
�Xk��G��@yMF~��&?<TS֐��Q�۫�|�$��G�<�����{���1������]{����ӣ����4��rw[�h�Rc��_z-1�����Ӊ��ƞI�d��2�E1D�18���ap0������|�#Exb�~hc�0�g ��3��(.P\��0?'�~Zt�C��Ӳ�
�>����eX���;Wg����ي��ao���&�����k�soΞ�{[x�-ޅ���#�(-S��.ǖۇ�#���q�� k�-�w�a\K+˹,�7z_z�-��S⋯
��_\��}-!�v�o��:��;��߾0�%zW��"��R"���;������F�l.�����>/���֣Ґ�"_H#�ʤ��������߻���֮�C����bzx�/���kGD�*x2��dfz��;�?x��;#Ɉ�J��>���!=��D".��ρ|60P7}=�%	���H���TM./5�J��emE�
�2K����yJ��@��QV����R�.�z(%����%�$&*�R�2[+��m��G�cS��d\A�o�J�1@?LTq��g�F�V�dM���q����g*�g++�+�K���DA��m���F�*f�s�X��^��F#�X�?naz&Zdê�a�y�A>���yq@���hL}v��!��$��MXc5��ql0@�p%���X��jJ�h(q�P���T��w��߱{�,j�^�6p(l\�w7��U �i�������Y������o'�lo��Z�Z�:1�(�C��a� ጜ]&.<���O0�u��;�\�u�kre!�\t���whNf�l5i͊٭��_�>�\������������j�d�r�-���$�%�I ��@|5��rJDV�l:�<;�k��-6�X-h���ʊ�0"��W�bD������X����p.�$��!5m������ ��ka?��pT)U�AAr$���J����x�R�]��@ģ⮫QHpwh�Ԡ����/��ͨR���`넔+�8�h�ݾ��#���}��FVj��+�a�W�7�"� h��-,��f��Ǿ$�yQ�
;�0��<y���`���VWeb�G��_�]y�ш7�K�����u������O�����8�sz��u���2�/��N'\ˎW�2�O�Fк�*�q� ���৥�(8����������}��Cn�v��s�M��$�xgY�>��z�q�᭗�מ��x�Cԩ��;2::EU�s���?J��ڹ�����?����r����t�)��W�7sJ�[�K87��n��	R}ˍ�V�������/�=�����c��O/?ɻ�
?4^�:��l�`�
����Gl�C�)I����1��Ă���-ז>Z��:�#m�c��<����"��
8z�^��Z{��7{{}�C-������i~tĽ��;~�w�`{[AbJ�")'=���m}e���?޿���2��YD�V"{���t��ЗR�+�t�Fe��@j����EQ亞������!cyXN�A�S�˒$�.5}���w��/��.��"0lQJJ�Je���[�n�O�‎�]��\�b 4�:㡋��ޘY�lɊ�U^F��.W%�����+K�L$U -�s0=,��c�\DL�"��4�n`E|��(/��'Qs&�I@2�}��`���@����E4�a��� ��V����!�F�#HZx�T&�#|�I&�(�]_A�a�
j������o������%
���@��d�0�(���^6���:8�����v�{�.{�hgvuANs��21J�¢��@F���h�2���5�U��[�5Z���X�jodK���a��)��+3�t&;8KA�ˈ`�t^��bY�fM�b�b�V��^��ι$�SFx%���������oZ\���,;Q��y��weJV��Z}cMX��p� hF�p��:"�3^��Z 2�E�Q4u�&D�Ph�gV�ЌǇ��W�Q>o����54��I�����X%�@���n0�Kѡ�<0leu�F��F�P��ǿ�������Ѫ B�zG�6Z:|�(=fH7U���3��u�MhF_*��������}�U	��E�XTKY��T+�&�>�R�e	O�#?��U���b��������Z��s7o��֭�����S�_x���.��fI�a��hȴڑ�ޠddF�/���2��R2��\zx!UZ� �2ƒu��(mT�*�L^�K	�����州PD>/&�jK;�ח@����C��@(l���3Υ�ᖂ֒�<ɭt�Y�}Q�[��������y̗Y�g��O�#�>�	z��(?�q^У��b]�|JB��.k[�G�}1�ksy� r'7���5��Nf����i�x���4�9E���'��&E?��>� �ʴ#�g U*A��;��7��r�����wt�Ոҗ�w};���޲�k��PN{U	\����x9��j�b��F)Dns�<��ǁ�Q��"3!��Ra[X�qn��\�ln6��&$jƆ����+��[c�������r��,�OgD?��q1�rst �Q�f=H}E��2E��tYKʫ�-U�CURB�*=�@(iR{�~���b�-�1q������B}~�zn|��퓹�]+��F��^���%��60�ǳ��>�:נh�@��Q��Fe�?��\� ��U�$��E5JI��i ��3ق���B���"��l Ǳ��0�IF	U/������1�|��W>��M1�(L7�:��(f�T=tk,�jA1v@C����o�Fx���3� ���������k+��&h�+v�˳����;�#��g�ڭ��l#�f��
Yi~�����ko-�8���&Z�f6l�3m=�[c9�9$zkl~�"�M��M�:�������u�2���^�ot���j�t�a��z�:���Y���������Ͽ�ԥ��uj�������:�`KZUKn����,�u%�%锜v='1���qn�wus`u�kyA��U�Q���Pjuia�c噐Os& �T0���0��Q�_�P� rFc}cq)��B)��S�-#V˕���U�e�h�MSM��r��o�JED� a��X!i�Q,�Z��V�0h�@f �,j����)z�Hc-=Z#Jo7�k$e�X(���U6JaǴ?�l����5�U������v�gu �$�c�������Y���k��ķEa���jӧ�5��m�x'���i�g�h�B.�t�9j�{#eY?ڇ>�mv��F듴f��S��c^L'��N9�ϊU35�����|VE�/Ay����o ���}L��$�T�fhh�֋�	����ܹ}t����C��}�;�\k��/���S��@���,���^�^��<ɍ|��(;�I^�ܰ���#`Z𮐢�.�v�Qw��]�w{��j��.jn/j�h�����ۆ?yww�v�����d�+����^L����4�+��w�X�rݸcˍ���0���uo��uyo*�/��^I���̦�
�l6�
����}����)�?g���彝�y;��N��	A	q���~vrt\b)�N�i(�Z���޲��Y�b�*�5�Eu�^O�����}{�XH�I	1��Ws��!>��rZ����j�T�Z�\֡D�kh�H�
ZURRXl5�4�el�&)�Y��N��W�f�^[Z�ilaZZ^FF�I_�0�x��`t�Im��UR�����AM��
f�X�_k_h�֧F�&]�U�t��B�a��L��F��P&�*�%|��ۍ�7PeQ &�퍕�D��P	�H���=�3�A��k򻭕S��A��}r�6ڶԩ�P+˓d�	\�XlI����fZږ���cm�m�l�$6B��K(��2��^�fR	JĜ!@
V�A²淭-c�y輰��;3Y���=;;a���|0;��u�п�_���'�&����kl��;��>�Q��ǖg���������G{�Cw�TG�%`>̩�B�Lt��F3�YzaB��{ic茺���έ����^�~c)��JKig�!QJ=�����Ϳ�7/�ݿ{�?����ɴ���JgS�R�|�AQQ����$����J���\�&GRf�j��n�L�1�ea*��� -��a bDalE.U�Dav�|Ƴ�)��1��C����m��h<~Ѡ�AD�i�Q^~o����ڮ}c���wz܎������Ҕ�li��e�����[��*J�~�p�V�X��Xt0��׀r,�k���fw�u�f�}�c�)퀑�c���'�rQX�	l�B�7��1�o�4 ���×A�èm$�L�Y�8ٹ��Z�:Z�Fi��3I�7đo��q��-�E��w��&�'�^�>���b���c�m����p�\[A]������ˉ ��K�?�߶����+�l}�C6Ą�#��?���饿W\$1���#�RF�$�{WA'6�.�9�6�6�{��GGX����>�s��ѝ�;���H�:3�Z���Q\Id,��'��)!�ʏ{]Hx]�� ������������zM)������vQ��w{ƶ�a�\��K�켢��U 4r���������+�S��2�I���J�s:�\�PQ[2�rz��p��Ǘ=ކ���t��J�۩��2X���غ�	�ӽ�s����㯟���O>�-9W(�$��I�\.'ޠ�Ev�4���wN���{���q}n�o����~Ǭ�y7m��M�5�M�_~y�󃯭uYĴ�p-����~.�p*�pN˺d`��: �/���n/WQ�1J��]�nL-�OO/��ը����i������'��߽�_c�>���haNQvVQQ���Z���{r�;2֨��3*Q��U�7k$��T �����E����zq}jXM�%���ꄏ���+�X%�����*h��E6��Aq�p��j�@�� h@�DH+SRMi9]5c~����d����G{w��>=ؾ�W���ڬsnhyx޵�>��Ov�o���������*�ʙ�hTf��*r�f'XP5;t��l`�����A�gc� .�u��sbPa�a'�LE����Uۢ{����;����m[v�m�:�G/ xoD���3��^���.J�i2��+�|~�����ުg�إ�x@%���[��F�BgZ�<�Tfյ.�.���4lnmL֯�X��M%�[+U�%!��G����Ǐ�����߽��z�iҕ���k�;��ǚd�M���1�ƜR�^Q��Ja��dG�):Yl!/����iP&��[�� �Ő�.��4(-�aM��`!X���h��Z��1vh�P�;:µL�9�csn�0�{����;'�n������b|ͽ��]\H�(a�S�o����	�	 F`���u�H !�GG��l�CEw4�[�tZij�����k��Y�q�lM��䄩�2N���U����!@�	W�@���K�X���	��� �<�ȑ�g��=G��G+~�i��J
�m�Ua���K	:IS�js��ds�k�����o����?_�3߶=V�ңi�I�ĿM��Eɍg���K�{%�p� āBQ����q�cL�6�jA�s���(� t��Ġ?%�?�19��4��,^D�����h1��//:��K`�kvx�) �}�ٽ�O���>��pm�=��h�J���䡩°Tap'8���M�g��2�����xt���G���{�N_`bm]Z�� �T�HI�-c[�;��G�ӝ�#[�_5����G�JCs��yҰlq\NrQkâ���{h����֖��1:E�#˗E%��%��[������co�o}��͏.L�P+��EA9��������ۃ_~<�;�������@���Z�z}Ws]���Ə�����_N712�C��WL|���C|9+��Ŵs�9-�v9:Po 4(h 4H��MjanZz2eJINn�V�����w���xoku�����H���-���T6��֖��jY�Z�
ѵ*Qp�4�6�W��0��a__X� @+�r�kq���Ry�"�l� _��W'�Jl��eZ��q�c�$�g��ђR�%�x��a)�Y�[�����;�sx�����ާ�>��w�ݹ����'p��C��g_|~�/N�����c�2%�*��D���G#e��6c�fA'��l� Ѐ�Eۺ���U,'i$dM"M���h��g������wo߃��c��n�\��k��B]2E#'i�S��a�;��|8�͸�JT#���n�����+K`�%V��sn�:��1@7���|9Y� #����/}��*ԙ3���^����=��k�����U�ۋl��㍲���e���7�_M��J���bFi�T�(F�&+h�U��M�u<D:�<)l�"!V��c)�h	�r�Y�ۢ�,�D�Ѱ�|�2�	������S~���i��;GG'{���P��O���gS�Ns^��kQF�Q���u
����b9؄%v�h?�i !�&N���l1�m��m�;v��y纩�2\E��&����71���klE��РRv���k��H��I��0��0�o���?���	��O�g��UR^���̺�6圸�[�T0;\�o�Y�ٟ�:\�ٛmu�W�uk�*yď8g^�_z1)�,�������L�5)�1Ib�p��$}������$��ʠ?$��O�x>1�&�&?���4�bi3��T��tLMMnn,�P���@�xw��~�pQ����h`:�:_;�S9�Q7�U:�d쫳�4����zj�C�#uC��.���x�*�������l��蜜�!��?<8����럛��*��,��(�ꨜ��_t���G��#������93U��U2�U2�e��4N�G;�=c�M8+�9��㭝���ܦ�֒�6̄r�J
;,��������~����������|�Q0��֎�v?��Yc]{g[��?>�����\S�tJx.1�*|9��d���T��z�E-��t�I�tTLA���B��]�m��n��-*.Җ,��y3�m�ۿ{ǿ���x<�3�y��\uZJ~c]��ý��&���^E����V
oU�#���̡�I���������Ԏ��+����J��t��\�Eq�)yU����J	 �B8,�,���EF�O$i��
�ѱ	Ӣ�_ZY��w�Ϗ��܁�� k6
��]��ݻ��g����O?�G�{��[si�t$�QM;l`�|@�}$��>�, �4}]�ޝM?r@/l�蛬L��l��"P�L]����}k޹�o���*>�����[�ot��M94��d�uI)���m?\��=Ϯ{�>!/I"�g$�����Ѭ<�U .I}Ѿ�
��o$< zr�i����L�P������^�Pk-n��\8��[o�l�M9�l�r�.Э�h�o�W�J��p@��~3�~&���|�hI�	%�`�� �1��p��=��0���ǋ"au�P��S�q�1&r�U/��x`�<F'(쬟��v*��**���-�' ����#��w6wlUCU,5/R�@$5��� u�c}a@��#@g90َ��ľ�A�	�PAb�ip˶?����ڪm�Us�L���P�ԛX��X�>x��H�ƈ�O��S �f�������d��{w�wy�\��q*�U%�eI��Ko�N�(#,I�E�%kå�֕A�HK��*$$}�:����+IQ/�ſ�C/�nMfZSsZR*b���)�xV����?����#��Og�?��rj��.�� ���t��|��:Roj��7;k��e�m=��k�h����l�P"0�����g`~�c��f��r��q��a���_Y=��0��4��>>R �� h���92�==�9;�13�5=�1>��p����/o1<3�O��mi������X}��
ӛ��ѡ�����n�d�u�+��:��D��ڱ����vm��y��zb�2ڧm5M��'Z�';���<'ޟQ����y�����/��t���8��2��g�~��=��7v���o��j����I��!�Z�RAA��M�@� @_�Pq4�v� "Z���ВC5�ő۬�n����m[�[l��[���������m;��CQ�qdp��h����Qǈ�^����Y)��rj2ڶ�2�0ԹԪȟ�Eav���� ���Ζȃʓ�XGa��_�ڶR-�pI Ռ���i��(�΄r��R�!�tfz��[�����y0�����}8��\nT�7�*�a7�34|��3�>�Z�N�� �0 �1Ռ�C�c��G1*��] ��׳��ll���B��h�|�N��k��_pz|����� ��x'V�
k�,��j�ě%q���ӂ��¿����loa�D=Jw$Xy�hr)��,-���wŶ�݁s��H�D�����f���x�1�U �So���mSnƷ�����OGK|ݪ��ܡYi��� �-% �z��T�Lb���G	A��V���AP�z3P	d��&*���ı����0���W��5��EB�H��ψ�
��0��l`w��vxܳ+���c��kn�{{&�0�~z�XάɌѠ�����Fh|3�2$P�L�Z	ѡ@i�)�x����R5l߄���E�Ʋ�^?�E���H�P�� �k(7�w�2�O��H�GY�Rt�t����o{�����.��u��2����H"�$�w�m��H���ڔ�����쑶܎���q��o�B^K�{���z���'�Xk��*#�)CZB��C�^~��'�$�|4%�l��Y��3I�y���&���4�._fM�e`s�ܒ,3���)
C����n�o`a~|uu�f[�c�X�^@$ u��d�� N�ީ�ܲ����d�,Œ�V��Q�UX�|�\�,ho`gbnF_a*.����eƞ�a�JqUtpxj}ݱU�ՐSZ�lJS���,�RK�Ԝ�Ue^[��p�nx}p?��\b��f�-���L�5�c�Y�ADO;\�����۵���X�6���8��5-�"O�h<���Q��`nqczz��Ͽ��k�5�%��&v���ާ_.-nvt�~Px�?���pB3� �o�����`�N圆~^MA!T���U튆|UE.�t���Bm�I�5����
����߽�_ow�� �{;����j�U�-��U�֔0�jh �K��+�|<��a-��Յ�����6YCگ.�G�3��OJ��K!�) h~u�L�01�f. ��F�*@j, UgF��p40����&�6U�,��mx�m���������������=SS}�+.�g;������	�^�Χ���NBѡ(i|�	�_I��ݨ�!�u����ގW`ջg��}��ja�D h�1t4U/�j�������JC~5+��]�C�B!]˥X�0͏�)R͋�>��og �Q�IS�	�s���-�x��,9��bhݾ�G���_�o��tt���u?9�'۶G���ZQ\m�r������\�́����Rw^_��P��|"�};��z
��d�+	����WrhD��e��*|�@Rܰ`d�-�8��� C�#J�k�{X(	�㥋���`����F<GыK����� ?�wz=s�KEUf�,�l�_Xu{];�����;G�w�HA��=- i� �a��(?�@P@��@T�1#4�f˄Ӿ�EQ�@���q����Eh)�������@û�#��Q�k�<NF.U����Y��4|��i��tA}Uh��L:��T�[�iE�;�[�7��ʪ�5Җ:Iu�,M�V��-	>�J|=���Ʋ�of��h��%I��t���2QÊ�^��{Lt����s�Oe�?�E|=�|Y-bUf+��{��2��1z�@c�-����,���7
z�D�L+-P7WTt�NN,��<o�4|0M���efkE۬��Gf��L\�Y�hQ�ts�5��0rb���؛_]���Z^��xp/
 �k������4K�Ԍ�q8&�,�ˋW�A����wpe)�BK�J���p-;RǏ6cR�6Q^�\[��9���;���P�$L'������$�4�c�o~c��g�d����~��0=�KT�M��g���oy:;ǆ������������R ��|�˙�U��F� ��Z*�� @���Z���٠J/.��oWi-Y�y�Ez��� �w��w���9�#JEE�Q_17��k @gT3��1GH��U���`������h�J��>5�Zy�&�t���t��Y\�D)Oפ�JEL��H;̈&�F��x�w4*J���dubB����S>�W��i�O+Ѫ����e:nn
/7�~x�% ��.|�~�Ͻ��Y�)l0�U(n�`FE�b�b�s���M�H`B�d�,�����\�6=�%�jyO5� �Y��f�4�eJ�'[��*�.Jc@�|ޑ��Tk
S�a��&Q�A��\

`� ����ӵ(R���7���J�(Oɭ/�96|;��]�,kv��Tyi�H�ew����'����l��`��jw�����Cǣ���FO�TGNwSrUc���w5��Q2��t曩�S	�w夈|IV�^�e[�*�p�Dl5���hDq���G)�`�(Ӣ6���l 4�טR"Gc�?q@G�Z-6����4bcO������m:m�u�<�H��hV�T����=�\�l���H*Tz�b�A��$���RYa(_�c�
^�	�a�Did橞9�� ���:�E��=zf0C�96Kx�v�-�b-,�*���.�f� ��)����ɉ��.E��f��t*��t�{����R�)��BPVŭ�dʸr-�2��d�;Y��+��W��e���Ͼ����-�fA��OH�<��Lf�3�q/d�^O']*�SKӓ�
;T�21KK��$M<]Ga<�k`p�t��
�f�\=O`������$~qzz����gh/��r��7ܾ����b�N$2��z*��	&e�hۆ���;Dr{l�{�����v����W�|���/�ӄ�"�|�$Ҳ܁Uw��	(����JM��𺡡^��nj�@������fl�o,.]-f_Q3�9AZZ��#�$�Z���++�-��������o��	H������gw�~��7��ɥ����{��\Qh)�L�f��\�kٔ�j�M�����\ �uT�EG�B�`��T*���RZWj���[�l�}��7�{ǿ���C�O����te�5-k+�G��c��Y�@_����F
�7@/.Lϭ���*�a� �q%�R��Dr�*�H@����eB~	�e��-l�W�Lǻ�qwlq@c
�g��qE"�JN,����T����8�U�J�U����ہϻ�~?����zMOSz����S�B�	��茸�-Ёś0<���~��fnv��]����-cm��nD}fAbS,�5Eb�k�������"ďZ��~��v�-t)-2�Y@��H���ˬ�c�އI��w#�:��C6Ӱ�I�}�{�Xy�Ă����M��C@�8ló#���Ҽ����|�W����;���K@����F���%�~��j�#��.��5�q�R�I����$��~
�t� ���۶:�-�WW��:��T��k����^+ʣ��쓣�X9$,���`�pƜ('���l���NP�.#%Z{c�b�`ςof� 蕭�kS�%i�4��^,3�7��w� ��{�����	|DjU4}����;9������a F��sT�I�&U͏Ϲ�0�p��
��@S���ZԀ9X�<3�1cǦ���D=7Nˀ�>J�1P�V{�jy�t��6j����umoL��w�W����s/�2��Y�<vNuJQ����j(g�pt��t��$�����o�q^ɢ��K2%�Qٍ��מ�]~Dp�Q��gR�_�&��Ky)��f:�Z��Y��P��ߞ/��F2]O @�uT�Q��Pd�)-lT%Z��t���"5�x6�V W�@��I���N��m���XG����̲|F>��aRU$����T���ŭm?|F� �m��U Ó��~TrNl0�3��n[EoG�'jhqZZ�����M�=�3�N/(h ��s��[S��^@�TD>�O�X@�Q�"*�Fz&l�i�0��X~=�{.�z&�r��|� �f��%���ZZ2RsT�F��R^���W?}��׿��_o_|~﫯�Y��zz&z���v���LnX>�YxJ�z���f>��A\"����z�e=�7}MG�sH&QQ�5��Xg���շ4w��ޟ���~��;��v������~�i|b�j�.�V��n�NL� ��j8 h��(�Z^)�T�ű�8��9ѷ�%iL��U^�R�v��\��Tz�D^�D.KV&����#4V�_�4�!�ţ߰�8>��CU/X����s�F̉X:�Ԙ�1?��C�ty�v�'�IFY������@�!�� �`BQn��@	�2Y���\3�p�X�:���@k��<��G5�X�Ĝ��~�����c1����Z��b�A��v��;�mS�2��eB�4S�-�[��7�׿�Yϩ�a��&���9�����me��*������. ���t�͎��x4)���x���>��ｽ:t��{0Ӿ3^�*�Z��@��ĒR��2����n��kH�\N������ξg�`�`Ͻ�Xp���4t��oD͡�f%�] �^Ή7��FK�Ho��K��2 �����������(EPO@���<; h�׹d�ϱfHz
YϤjDI%�y��{�SgP�c��bv��-*���_�ǪV��U�өe�D��h!^WŅ�����ZU͎�S� 薉^���悡�~�f�/"�H�n),�4tn�M��wNֲb5�h%�먠��ڄ��>P� /�-��jH_W�Q�K�4��Z����m%��F� �"%��W\��Tp��ʚ�ʊ�֜�R�!�\��ޛ��)��F�1%�d�� ���JK�T&��|��4����W��R���Q'�	�&2CK���I<��n�uҵ4�Z��/t��H��+��Ӓ�J�| �����������\�䚂��M�p��\�����*�U~�i��3��$��i��ّ5�ۅ��!C��v�,��kw���e��H �p;|>������Џ�A(�?�G�����j��6m�:S��̈́��!o�¯g��۫�7זܞe�wrk�|��J&�E���7_R�zVp�5����BY1��`g���t�G�}��w���_o �o����oJ���+�qg����)�E��ޫ���i�q�����
 �9�xIGF_72����uL 4�(-�ʳ�AAWW�NbŦ<�����񯴣��/>�����O-f�iU*�ƺ��801Ӭ-a�6p	5"��4 �[��"���mf�ޗИY�x�*�\��t��R�GV�Y�$�\I.Q
+����G3�jE�����`A�W�e�J�Fsp�Nxt` /@п7@-<B�G�Z2I��D��#�K�L���뎭����F=S+#���Fa&��~.�g4VN��¢�B�>9��rl˾�8�w�}��F�L/�D�<�ȵ�q��y��ߴ�.��/��9�ؒ�߽p�9*z�2���U&W��z�7}�9�rZe茹@x�OʰrXV��*O�Tw.ͯno;v��\�x:���9�s��Py\�%��N=�_�6R�5^g�^*���Ot���3�j�kd�2A�E`n�o�j�kj�XŹm++�{�������' Z={�E�tnM&S�z6�:wY����a��� �CR���1��hP�Fh0��t�������z���A���7�q���J�Ө:�X�3�u��;+�դ�T�caZ���0K�3[�RC����ꞣ{���UR?Y'6J �D9ZK��2)��g�f](���y�������H��eV���L�V�6۾�~�w�7��3�9�mJy
C�&j� ��F> �z�w��Gt�=���55���N6���k�������=߬s��d�-Mͫ��
�MC˾��΂��c_F��:��2��S#I�Ǥ��ңM�~2��r6�T&�R>�]�t���ҫ$R3�k���c�b#�)�m�I���m��۷�[���T|.�m����ן�_{�u	�)���WN�c+�z ��Q,�:���A�z�ޣ��¼�"��[���r�k��4�ww�@�����\�ٚ���p�8��}�����ۆ�"04Њ�Y6���(��g��_ᇲK�A�`aڻ()1����H{;!�uE��rJAO�m���׿�r���Gj�_�G=-}Z���Ӣ�JÂ��W��fVZz��L]d��;���{����v��O������}e2U�Z+v��l!���}��V�|������,)�^T�(��:
����y����
'у4t�Q��-��UUV6���̬a�����?��}�J���o��`˵���-,4�o����Z�tb��J��j�)hl��!���W�7�7��Q5IWkq@\&��Yx�*E�.K�֧
�E�R.��z�H���YY���� ����F�0�-n��I& Y3�g��p߷��auk�{z0Q�I+Q"�Y h�i2R�X0_�������F�2�; �jNIo�s:7��]Л;��������RM��f�w��_����]f�L�ur]a�E�ii�XX�F�� v����Z�H]�!�j��f��wz�}3�ń�D��A�c�Pk�Q�Y��Ze�򢖹�E�/�}8��Φ�ar���?�"'��N/6��W�4�74�U�g�T%iJ�E�2����T��D�%JM]a�xK�hO����Ξ�����;'wn����p� ��w����LB�h=�N`�Fe�0"A,#:�%A���	�Cߴ��qopGR��ǂ�t�-�dd�D��:���w�����#=	![ˠk�L�0ќ����w�v}��e�Zq�.^��p�i����i��^���;{�c�F`�c��s�-�<��&ƫa��,���%��)�r`w4�u3��8j�3-�5�q�i��:8�mc���t��w\�����*�䩡th��|�k��u�w`���qvNȊ�r*��7��P�=ώo�6��+�+��+����v|�'�a,�O�j9��{=��Dz�Y�e�>��xV�S�����SY��*1�6?�._׭M)�L�1�������̌��@*�����P_]4Z��o�n����?�ޕǽ)�z]�?�#Q<�(cܾ���pE�Y��m��Gz���(���Y11���#��o�t^u�&���V��W��ևV7{V�������W�7mn/��u���KY��^TD�&#�K�(�&�~t� ����I�Ģ��ƽ����7V�<~�3\#pz���f�uio��_J'<��bZ�I1�&�]��\�E�7������\�4�����o��[����������ݱX���uM֪�fu�1.�Y�|O�{U�y��}V#
�*�TL;Ӏ�׍l���M=#XC���-������GU������ry�>
>|0���S`*/o���n�M4�KY�Uh,Q�F�8�ZƩ�x��p�7�'�[��)U
T&	����AA_,S�U'�J\d#ل�g࣑�5��#:PL�ᚇ9�uXn4�`7�.դXs��Ww�>�Ώ�@8ݎ��Aa���R�|�8��0rPR
� CI�zT�9��«&��xS�ED�%d�W�9���=��'�����=�c'����l�T�4��j)E#��蚔�ƪ�ŕ)���98�����Ό��\��C
��Ll�+J��x��_��aXF�J8,�DQ��XZ�����g�[e#=Y�si����I#�e���y� 8H,	��^�_��u�4�"1;^f䤘��VN�U�Q����6���`������������=`�so�m������d�u-��/���=!�nFK��x�1(�>G��AD��q2�d1*��g�AA/�v��GG'�w���F�{���3K�SM]�Þ�*��u.�s��x����s[F�a�y�p�����������Ã;G�'��C�}"�2�^�"�-c=Sv��Ǉ���^ 4(h�N@ֲh:aZCq��4�ұ��@�&@eoo�a���$ɽ���g��QE�r��F^6ֹ����^w;Z�z8�	�u�s^���������{�ؠ�(��������{;X�ԓͽ@���,����r�Og���"���\�S���hod2��e�����"u�&�J.�9�h�.&�8�rv�[�g�橑i����/*�h_�� � 9,��* ����U��%������Y��Z�����L����l�;�{h�t1h�ə��r�V�1�%���r��(�0/�(?2'����z��l0A����_�8s�>I��J&��H.NoYY^to�8?�M0<~�э��Kv��g	�B���ql��rx̣�r��2�d�_� ��餗S�e1BҘ)���^}Aa��ʶ�B����D�_c��~�շ?��K_�A_�.жU����"Y͹aU���\�z��s� �,K2	��/jiH>c��|UK�������:P����-L�l5�������/?�]����FƖ�Zk�Za�} ���*i����U�#j�ܚ����.�m�6ӹ�,�M
-��.|R&:��.��0���_��l-b�&��&�2�l��8���W��1X�	*.j�q�Yu��K@'JT�����WK���!I��qcڙm�D`�4�?�N�������x�"��һi[��9��RD�޽}����#���m.�����:� D�m� ^+!k�2j���~x���m "L3�{ �@>�9l����d�X�Cw���fZd��֞��Y��Ȋ�3����\s3Sr.K�a&��T�)Y��°7!on�+�u�{�����7E����"�l���h��%�V��O�����G��D���}�=���X*�ճ�4��
�#�N0w30�2
��Ƈi�"�0 4<���k	�i$����h,���4����BP�K~�����J �����X��mloyv��2��{fm�)�R���䵗���s�^��x�Ä+C�sp��m�k�h��b���m|ss�����Aٶj�Xj]����9�@-��E�ߗ�ιͭ�ۼ;��nx���ͮ��!�AD� @���/��x9�5��q�/��P54�� �'{��0��y��MƔ	|�5�q�����C���ݶ:��x#��L6�i�Έљ��3���/�9u�I����E�������д�1EWs�^�_yNp�=g�{��XF�w  ���9�[�l�o-��qֳ��w�x�	H���c�H���[[Yu�e��X�ܢ����qD��._`��*���*����Ix	X����xg��r��qTz����I�E�W@�d�F�LK�Gɴw�觓xE�=c[���)�h������#��߶���=<r�@y��>��v�ۄU%聆_�f���|!��2`���7�H!�Hm~i��d�����1��M}�x�믾�������۲yu��κ�ɩ!B2���F髅�W
���C̊��� ��������4� TZ�M��J��;���}��S��w�r����_c���M���m�7�ܾ{���8��x-�� ��z����5���JGjsvx��b� 
���'��4�,�P��V*9V�Ġ�vF#Wp���|�&�0[�k:�ř�$}JQO����.t"z}+����A�!�����QJ7<9���X�	3�Ñ��u�(��6�Հ0I����D,kv����# �\�x(���Φs���V�S2u"�A@2	�"��&>� %��������C�.Jk���þ�tO��4OI-Ydz	�z�mfG���[*�1-������M 4��H��0E�}9K�q���L��3��&��R�Rľ��;!�Me�	��'ƽ��Vb�)I��,�(%)�Ԇ��e�˅EG��ܝ=��}P������v=K��º���!����V�b�ԭ�H��Ń^"�?���i<�#J�%cEDQ0������D��#�=t����N��;9��d���o���;m[յZ�Yb����jf��::��F\@��cz�6�f_��1����;�v�}dy ٘�.J�w7Nll��<��5�snc�����˭iK���6���鵍���Ҿ.}[SYO���n�F���m?�oR��)>M�,�Xp;@b�7<i�B�ki[���щ��\W��Jd
��5]��p�'K6���Wgo�������П͡ ���"��A9WȧUd*r��e��tf��Ԉ�o(�>)��$�	1Ƣ�ZX�� ��x~e����;w�Ɲ��G��o�?��܅��p���d�ކ�ehiI�)�HE�J�E���[{�0��AD�g_]��F%ÓEi��daP� ,4]t#�s#��"�NKH-��;�0�=�88^�*&²�W3�R�q�9U����~)�v�{��~n8HxGg`wk{��9�w��4��]/H{#��R�<�K9��rY �3��������խ5��ͺB]cu���1�����/��/�/>���w�ݿ���/lh�jkV���hJ�c�YQe��4ܗ�i���.$�%����[F�y5*	}VCB1v
���Z�-���t��l����;CCS��]�3�ˮ_�����w��k��9���?���/���������kdh��~�퉩]	3��W]-@�U+ ЃKXOB �s�c�YQ�Q���q���R) ��U~�T_*�V&��� �	z�Qwh`wȡ�c��Q n�Slda�cBa�SA�������>��A;/�V[ƺ�,�b!Q�B��Ψ�iBt�-�Ć�y�H��a*�$47��QҹY��&֕5.,͸|�I �)���v�eM%2���0�B�ED1	@��<�AD�*9�����5߁'�"�~�e^[T՗���H*q��R�0��(l�)���9��\p�ڒ���ڎ������,1���!8��=��>��=���0��n:��tƩ4�k��Sʸ7%᡹�6A�l��X���BQS�K?0������`����[ێ�ա$������ȡh�Q��q@#�l "�Q�?�� b+�X�I��4�I��a74>�tgw��G���GV�ˇ�iR���N�[�X��� ���FmOgv�1����`�怩1|x���1�6�WR�+H���Oo�`��,v��7��z���Ҍ�⁕�ew ��hE���G�ͦ��)�
Va���a���8�(-hα��25R�&�|� ��Bl�}��K�������F�g���$&��$-j�Nlm���;�0�_�x �A��H��2^.�v~1��j��JD��We��Jx<=��	g��5�sC@;?ƿ��,�qyԳr�)�j5Z'g6./�O`�OA,�98As#�2���m���n���W]������ֲ����ʡ���m�ȍ�����33Y��Q1�V6�V2�bi67��4Ԩ�3ԛ�U����e����Qf�;;�K�E]u��}tN����:;?k��y���G���]�rt^�nolu�nX��V�I��Ө�f�^�a���}9�Ӌ�2(/e�?�gG��섁�~m���X96<�ӏU������}z����˃�weekW�@eIE�`+�K�$\2� �����e)��LzU�b
��7@��@D���#t,���uw��ls�3���^�L��?��G*�~w��v���gwn��Ï�aH���{�-m�m{^�ޗ�u���l�Z��'!RСUf�����1�4S/�M�J�\�<W���R.��":m��%Pʕ��^����8��A�-��g���[�õ3�P�1	&M���n��!K|� �Q?��)15B��<K�͹Qf��@�K�3'�Ȋ-�Z8(��@�`�����,s#/Z'�R)�e����Y7J�C�:,�$�ͳY�aI4*$(�C�5��� ��"}ZA�N�-���׷ms��VkF��b�Fk����.��WFz�D�����)�nzlr����kn��+��.�$�6]R�D�f�J�EjAYq�*)N��N�V�p�X
�~#��f*�d��jf�e`y~ËJ⁮�d�=~�v ac�.�o}.�߻�����t���s��h����ԓa�H������Q45�I&*܉Ǣ�b�$����l�3	�����>�@=�幢:�ؐ_��)�G�)�Զ�����0ϯ�sbPZ����|�P��>;/Ģ��v�kv}^[e�f�u/��7��q����;=#�lEF�vpy�1�>����jn��U$�j�0!������Ms�.����U,gj�AA/{]
w����%rR���o9G0�n�=m=0cxB����2e���hv0Z�z[����4�3D�/f�Oeѯ�强"e}AnK~B�H`$�q\jNx#?�5٥?��="���"���ا�����W%��i��]-��vϒgj���:wP�=�}�V>������ځM}�~`MS=��=ss?L��M{��DeoK�X{�hs�Xc�8������ɖ��֙����Ҿ�������ŕ�-'�l��,�(ioZ-�j
�J�Zf����p�0����I�-�nߐ�n�ׄ��N��_�d=�I{6��\��,�s��g1 ��<��Qd
WUi����h��U��n�'̾���{��p���W�����@g����u���Xf�*..NӦF�S�̊w�9/�_ɧ]�K�+�8��Q���Ӫ�s*�e��:�U=��U��q�X��o>���m�3�����R!~�������y�wrt���A������dauwq�wr��ן��ݣ��Vm)3��F��\��ܬ�ި��U�05�������呚�jA]Jxuҥ��UJ�3�菬b,Q%�Z�(���YF:���RT�O9.�`;��02�1�b�~����1��:Vv�M����#Pgn�o��]�H0�04<j��0�9Z���Q]i����+ӣ�zjM���:T�M�F��?������*�ױ�uX1�\��G{���ɍ�ᵡ���ʡ����������)��Ǝ׵���J날[�o�/����d��JgNg����n�Ӎ��z����\`n��^��S˫�����8������4C'�u����JV��*N��/�(��~7�}6C��Q7�v��A�˻� �m��M���9�0����y��;~�H����V\�͓Mb=������mc%�P�*$�����'��
wF"�D�1��n@Q� huGӂ7�Zl��m�(8}k�_�j�����ˏ/bG�ѯ��R������=._`չU�U���34l���-N��^q��^�| �����K��8js d�S�odw{&��T�������:�@�n��Z���t/��0�eCAH���ݶ��n�&��J*E�� E��;�? ���Էu��Ћ���*\�8j���J��/ԋm�sN'|^�%�r�㮜��.x=��B�7�7
Q�*��@ݭI��$�!�k���"��^��\p����ǒ"M�z"%��D
��$���E��ױ�:ms�k݃l��^v�p�nn�ll������ ��J%�T����"��L2%g�Wtw����/v����dZ��-Y�֔tkjZIr�5QiNH�$&�)愌����체̲����dcvQ��il^۳0�85�j�RX�R��ڮ��������R0�nljhusf�=�pÌp���r��o�'�	F�{)��YO�џ�b>�M{&��L6�t���4��x���Z�4FX�<:�W��dg��%�;�с��X��ۧ��@��G����ݥ�-�ͽ��Բ���$j�A����Z��\ʛ̰�TRE�>뺆\��|^M�����a��+�-DE��E����h���ͽ���ŝ���Ͼ��!��?|��������>������u����{'��,oMn�-�m��;G���=B
�����\��
�����s#��e�Z[ޚiYl�U)C*.U'��V|��~b_*I+O$�*��
a	5�51���
�`�-(��h�ʍ�j��h=��F˃@^�\^m�������`m��^��沾��R(ل��"!�������gb������c�{��C0s�~��oę�qz)E���DSK���E���;G��Q����6V{z����ý�'(�d� ���Vm��5Z�Q�	���^o4-��\�a�Y��Ҽ���E�-���S��캲�4I�*CZk-�j2v����O6N�4M�͎6N���e5X@M_����;�)�V�v�\k��@
8�M�kas�{|<�����6����=0Qu8f�������u�ۗ��*X6IC"1�\̈�X�Ư�pl$��d0@3�3�h0����X�z�=�U�-�{n}�mt���1��(1��
�3Z��"Q���Aѧ��c.c,WbٱZ�ns��P/Ph�z�&`�:�ǖ앝������0 =���lҗ�� V��6�{��^K�$ʌ��)4H,������ۭ�����Zf��U�Բ0b�a~������Y_ef����O�v��T&�|��wh~4�"?� ��Em��0r����t؋�>N弖N{)�r*�vE#aW禶�
��*�Ij!L�4}TPn�k�3��G�G#I�:?��DB�3��gH�H/�io'p?Q��z��w�svnpqq`a�gn�}r�y|�}�� 䳪�Rc
[�g��\�k����m����\]K������,�'��"��#��d&���F�1������2#[�g)M\��+7qeF�� O��f��-�e�QI׋Xf��2K�[S7?R1:�]S�[]�ii�n��m�Y���1�67F���K���~.��t&�L:سy���頣AD���|�@p*��z6��Y�ȢaNjnaQrRFyImG�����_ Y�͌�s��헟=���/�������UU�U�5�$g&e��y1Z�y���"��W觵���nSQ\e�E5���rVC�	A>�2rn`�e��1�٫����?=�o�/�Ì��������v����8�������N8�_���+��N��;G�̮���mM�W�@"��w������VI���]�^�]�W�)}󣰇�u�Vs��º�Ъ���3ҏJE�HN[e��	aeJJY��:IT��pP�Q�bA+Vz�� �\�#��"�	f>���O.���;1?&Ȩ%�Juo�@%�I+��!��C<�������̀\Ϙ���c�}��]@��&�$� �n��C���UGs���ݽ��К��.����탓��'w��o���,���m�cz4�Z�T+�z ���	F#5����:&�u�s����@�D�oq���e�r���5��S}�`����t�&�ms���-Ӄ�㝙M��<م,��LeQ���`k��8/�|a&��$V固ڇV6�^�Js�mNHl�x�غ�1�6�\�NTQ�L��d3�d�"hP� �x��|pǀa�LCI+h9�IՉK{f]�5sͶ�1�'*H�Hy��f���EtƋc�$1�PV��<aw R�x��[S㪚�T�"�"�m�s���b�H�0�:)%�v/(hx0��̓O=��&(�O��Z������Z��R��dW���W�:�l�+M���2s!W�V�w��o�@��;��(/'������D|�0��p�,k�T��n���Q�;+.O���B�A��t��9LD��<D��r��B��	Bs]Z�����K� ��y�#J��1�%�>��@?�$ ����S�^S��S�o�H؅9�u�5�\�f)Ps���:�]$g�dL����Rut���0���F�:J�a�B�����^�R��**[G�?	����A�hl#�g���`$����H��|�o�puB�V�PK@y����;�"$������f�u��8�X�^�Z���DE�U&�8�����*�(��F:��T�s��'�)HAg �b>��\��Y�7�9�d��^M���A���|����n�J�,���򖞞	���� L#z����{��|���_����>���g������P�Rs��˃�����JK�j����))׈�I��z�;Ŝ׋Qz�;���,zM�.���Q�8���c� @����7t�fz(f��J[[s�-9W���˻CS��9�и���+8Z|D��n������Ï?|�=؏�~���_=����?�g�??<l�u?����>������zGm�#�s�{��w��8�S�(QU��U ��:�4A��0;��>�:�<W/�UFT).THN��>)��.S���/[��)��B��ͷpXj|���C.i#�#Q�
�4�r�"��$C��B3�e��=���|��m`nP��14\�茀���X
5���:F_�`�H�1> ��Q�h�^ˡ�y����3L|��KXk�ubb��r|�ouk�枵���e�ww}`����-�ޥ-���z�ԐؐI,�k�HQ�<��Q��I�r�L|�Q��h��/���a�b��j�X�Y�sN[yqoEfC�� f�E4z����)�-����zUc��ڛY��̊�ř��MLc��֭��̼�:���9�a����.��3k��kv���=���9����)M��)�D�HQjb����p�r���\:�)J�����Gh�õ��jB������5�M�v8���Uss9-�]@�R�C�I�EĠ��[jB�$�f1%$�ϳu,,��P��j�c_��6��-��(9�kd��r.�qs2�:Ӡ͵��#��	���77�������IG`�0�_�\�=�s׵p�w<�,~FD�k|uM�R�+��J'�u����x��=��β˥���*+�ă �F�P����w��}�d5̱�G�ڴ�{����Ng��� :T�-����J��D�X�S,Yv+7�uم���W�At4?�Dx4!�qE�㲘'qO)�^H �J�\J�r�Y���vcAm��$ ��סw(��IT3�iq*J���&tD�.��#Qtd���6�9z:��ep�,�����z*�@��)D-��YK��	tm<[O��,-��#Qaj�%S��x%^ME�դP)��
7�t�P� RˋQ�i*&��&, �����Dq�V@	ˣ^+���}=��Z6����2�/�q^�a�W �P(	էi���>�ᾕ�~'��~6�b�0f�iI	�iֲ���щ������_�i?&.q��D������?��`e����[Y����93����BO�G�^$}���F�ۅ��:OҪ"�&^ӲΨ�g���z�e-��� �oa� �u�H������}��ɥ�����h|)�3�$��_��u/������g8�_�����6��-n��Ͽ�?������Onv��wtO���=��>�-N�h+� ��Z��J��iP}Bh��Y�>�1�FQ��#S���$ ��*ٹr��
T����% M)MV*V��̂���D�8L��7P����jt����g#�j�1�i�c�x�3���]�\46yZՀ�[���89���������]?��3���n1�Tb�"�T���XLɜY�ŌR�J*V1sI%���3�[�[۳���n��w�9};2*"2���w�=�@9�tT��3�C	EC)F}��y�"�� _`1�'�d�����rww��y �&_S���,���V�:�+?�����e��P��h��H����ى�U���ެ��,���L6��jKE����a@�P�E�w�O �
�/c{3]C�+���fi�kb,��/��u���:+ƅ6�LXh\+�Q� �҈�,J!`:��^^�������̉�֖�X{�٫������U��E1��]ͯ�Ǘ7'����L�5775�[��̏,��)�+�}s�����䫒���Q�a�Ǘ$�D��H#���\QE^VF\QD\���]UF^WF��K��򈋲�긛��p-���{x�����,��U=Q�]�k*���#�Iá=���<	S>�(I|��z^��_{����	����6���.��c���fq������W��p0pycs�n66G�ns���w�kƦ@�4��I?̳�1ԧ�bu�'W�:'�p�Y7�)�xq�zY����[�x/1��Q���h��5V����Х�̇+�����Dl�����j��՚s������4��&}���Ţ+��A�z���L���_�h��s�^]�W��� ڽ�T��oD�{e��d�G�)�28o�!X��pV�~(q���I	��[��[���d�`�D�.�_?�&�!��-��#�/��+y�@	�eQ���TO�p�E4�M���������۲�����{�Ȼ��[ʈ���G�����/)]�E��Iy�`�U�(���BBb!�a�K�����a���\/S� 3-�d3�Q�f�h������W̒(�N�Y�i342�
"L�y�k°,vX�a�����g�ź��guu{g����������{���!��o�a����׭���%%�6����elj�h* ��l�S��J>�\���{��y���l�:��ٖ�<�QC�Ý�H'�JQ�Z����]8�i6VV������΁��}o6:_�5uOV7��i��{��>�70=:������������
������������?}�����[����������O�����O�������V��TW�xk�`YekmcwqySK[������
�������{)�X� �H�+��U��*%te���xK~��� 
��B��!+%��LI��VDk�J��5��Q$����ba�fxHG��V��B��f���A@�J�]Acpp}}�����ݻ�����7x�'�¢A@��~�3rq`���R�l��b��W�nt�ڊ�{j^L����76��*_�Ͼ]Z��1��4�5�6Ѩ	�Yn1�-�{�t���4<YBw&�ad���2Gы�ڡ���}�=������e ��V�-�{P�SxvP�`x?����@g0�x�s�����홵�ީ���2��@Vd��Xn!�J�R���[�.�~p*,�r�)5�Fɧ�ML�GY�^����z����/Z6�6����GTe�p�0�I�,���{~ �fy�r��Uv7Utu�vv��9��3���捦���w��ƃ/��b?��~��ۿ���5�ޗ�G�a��5�������;��ƽ����!l|�z�%��nJ����Z���B�������Ƚ��{��_p��u�(�+a�~Q�o��?#$d��v̯#�1*��T]�F��1G9�5 ���Ԥ��(�>o+�i�}�D�_X��_�5�����,���:=?���<ًl�P4��6\m`a������{�{R�zG#����F�����o߬,�w5Z�<�@���������

�[߂k��Pp$�jZu���k+������B�0�oh���ԥb��t�y�(��'y�g��=دMاOݧ���T�|�H>���W���Ҿ'��I�N*�e�x�y��Bk�5'�:+�4���uRS�qwԱ���'���ro���;G��K�_�n�"�
�_Q����G�w��� ��>��=�ۇ���P*�������`/��_���g?8�zp��p/���>:�{t@�O�W�O�x�������r���H=�F�+H"���xA���gn|u����I��it�9vb����*|d�^�^���$%�,��l]Gy��jWsng�V�iV�._�C~��#�`ъM�2������͵��]�oެ���~�����_��������������w��g@���dO�Hii��]�w���+,P�4)VM�Mq��f�.dC{�$`טe�m��\��q��Z��GR��i��**N�9�J��]t2Ҝ]ua��VQ���=��|��u���Ui��Қ�����Ί��͝���}S/^���oj�ol�������lmy���W^^W_�����E�p{W�/PSV���UUT�������j:�5�=�&�w6w��/��kE
��N���W�"��'Ai\�����&	��f_w̴ʪqeJ ��R�k ��DY�J(VS�� hi_�gs��	hF�U�n����b.Vtf�����wya�#Z��vwwa�
���)ᠹAe���h8볯��+$BUy)gy5u���љ����������}�v����>����7�~���|��q{f�M��R~@A��(1�'�y���撂1\
�]E7kx�L�� d��d����K�s�E�	 �(�ُҀ ��N��а�-����Ck�; ���J������PX�+�*6���~F�������_�����?����l���F����@�ð�x>]��
c��jˤ:l�����Q��n~�㮊u]C�� \3���~���ƝWf.�T���nn-�tw>WW��%�$�C�����R��&��%��+N�'OگH>(G�n�(�+a,������I�_����xZH��xѳ��������녅�ޮ��IE�AY�e�v�
tb�>i\��`)����-.��Y��b��6�*A�eucjielz������9��j�Up����P=�j`zlbbhh��EgkU�`K�'메.�f��u�/��nͭ�`/ 5��qL����_�~���/�)�d��
�)+���ousfsw~kgz}��u���-(�.�ؕ�{��595���" 8h�+��n<��-hix������YU�zkz���Ŭ-��"�X�4�-�i~�)ɽ������}�O�R���� �+y��įdI{)��i$ɧ���|!�(�Y�rg��^��K�	\o&�T<=��>�vX���wX�|H�v>/޳��g�s??~�0a� ��0��)ᜆr����^�����S�IR���#��N����G@��S�)��(���SO�ǌ�C�����}�����c�����Vj��cN![R%.�]��8��?=��?;�����v��r�7Q�&3,�D3'�(�V��b��MV �^(�vi�5�?[U�t�5�����G&��|��\nX�J�N�dR�Wz<����Ҳ���ښ�V$�;��[{_�������YS����Uy<��yfI���ī������»3��a���9�|!�E@�,��ڌ~V�1�%������i�l��v��(%�Ayb�<uP��P��D3���T���ʚV_q��_��-i�y�����[Y`+6;+J*�+*� ��6g��Uc���*��2?��v�����]%GiQ������	z�5y^�����X<NgQmCgM}��������=��C#ͶR����Z)zD":�BT�����%�,ϿY�m��������K5���~9 �Q���AA��(��ve�Ą3�E�Z:�>{y�TA ���{����O�}���~���_�agwmp�C�BSա�'�h��s ��K�in�&A��d�XT����Vg��l|���ӧO��wX���}���>}�VX��zys}bi��e5�)C���D����R0'	��.>*���|r�SDr
�����Ԥ�xD?����np>�bN�G��[&_��N���@ {5=��9	��?�_l ��{8"c�W��_~�_~������?��?������_��Ej�4"���Jҕ�V^��A�gLs��s��u�:��tf��yW+w�� (@׿-"������츥Ʀti2K+^��>oV��ϴ�[R����|BI:�Bv\M;����Q5鐜xR�8�����J"�	�Q��� %��$��wRHe��kgV��7W[�L�+������tA-j��	p���e�a%�b�ଊk�W��M��,��_\\^\ZX}=��3=�|h�����ұ�W��j�H���z[~gE�@c�ps�`�g�ڲ�|�/���~"���٭-M��=k��CK�Ë�k/g����d75��Ή��E>�b%Y�ǧ�桟�Ω�
�R��J��fբή���읃{�[AK�`��>�����.�k>-T(k���N���X$�˝B�'��<;�x��y����/Չ_��~�L�B��G�рi 4���T��\�7]WY���fW�e��M@+��B��#��c���R�Q	ᘔx\F>�����
�1)鸌tBI9� �T�����=;$H�ǉ��WP��Hg5t��|JI=�$���������Z�i=�\&�|.�d&���|"�v.�~1�z5n�D��i6���NSD�i����޾?���On|��+_���ޟ�鍘3��\�e� �:ڡ��#�T 9����E��$�dD���;���A�f>.�|7L���{Y�'�|�3]�+�ux����2��_��6TW5UV6VT4�V48��eu 5��U�ilow��f��o!����5��Κ�m�kv�=�(����t�nqm~�[���xh%ݳ��[�ld��ȇ���TU9�I���i+�]֌lSv�ݐiQhr��
Ch�4�x*
CBgJ��,���0ߕ�ki����Ȱ��E��n�-PP ��6�/�P����
E�^_ g3,:c~FF��_ZZQW��180�T�VV\���{|h�o��\�VW�Ҫ� hPБAY\��S��c�����P�d��ƈt�*<�F?(Q?(V�I�Zz�ZT��x!@ӽL�)͏eJFcI9N 1ڍT0ťȨ+����.��[ 4؇O۽�M�T�	�2>fBfn�ħ��5�n���*�IX��%;e�:w��̛���e�	]��w�����MT@o{je��̨��KsH�m�P���H��?�Q=Dq n������	�mAK�=�&-�d���QdT[ۧ_OlmL��[�^Z*�y�OW�-���G*�rme҈�S?����������G?��?��O�g��?�ӿ;}P�P��
�S@r���9Dw�U-����q��g�l��E��q��xlrx��N.�ΌYk�
�\�R���V�j,~�@*P?P1o�WՌK*�E=LM��c�kj�W��*�%���j�+)���yNA>+'�ór�91LA5�Vg7�����VW?U����KJ\;�g]P�@ĝU�/h(���j�55�F����/����|�_݋����R^�c˫)-\��j*x�ITG�{t诮����I���ܑ���`�du��sO_o��P�T�y����n{KGQ�����/-�%���b�U���rn	^��zY���*+��_z��eV�KF��v|�%%�L�̤ޔ1�E����@��X��8lh�k"�TW��|���[A�Y]"���B/�3Ζ���&b��ᗊ'_��P%�F	�N�J��2	�+iB��|X���':�:35[��*��)�"?	ہÙq7dQ	�A�U���g��09���}Yɸ(�]V1�븗U��
z���}v��칤d��igŤ�"�i!ᜄ|NB	�Q�,0�M�jط�y7��kFΝ��tV��y1�s�@|>�w2�y:���V!�~!��	V2�ǶT�n$��o7�������~r��~r�?9�����g����]���F��6A�[}�$>�'<��<��8��zh�G�xϬ|Z@�h��7e�1��̲���Ez�"�g��d=��s�Z�#[o�ɶ[�&S��g,0�j��(�d�s���b������ȭ�Z�E6��kR�+��sΘP��Y몉��*�T�I�V��ю�J�E9� �f�!@G9h�>N��
:�A�sR�Mp2N��� �c����2*)��ȋw܊��p�α�kg��M �����1�ix:KaH*�<��+Ud�,m:O�k�B�Li̔��'8�����	DC ��eB�&�b-����k����8��m-���
����P))h t|� �9���-�OM�5��J��I���e�G@�R%ZOX${������*PВb�0�f�Y/3V���@KW���8@KNm�p��ۯw>|��")��o�����>nl;lm쩫 ��R�U�2��3���xW�������7K�继;�j2���J�`ǫ�������;��~���=�9��?, ��{��/jyN5�d k(n6P4�0!�2���8�k���X�T�6ŉx�����EYv�p����»w�og�7a����a�����XT_:�%U���A����/��o�����������?�����_���%�f����8ѭ�.�N�g@e��Ǎ�S��axN����:
ؘYY���Xe��#�y��芾�`_�ܕ�b%gIRr%IY�Rri9J\�:-O�.L˕'���X��������1��İ�)1:�3� ^-&�k�V��ae大jEI预-��Nɑ<�>M��e��yO��F�t�"U+#�ܜL�QG7h��<G����wyv��/��k_\��'�O��?�����sG�<�x�)W:_��X�>S�1�S��Y�,P��V���	ZI���T�4�(-C��.��F��#��H79[.�f�����|��цO�$=3%?�ÝQ��Ā�<�`_7�"�ӣ
2�g�n�7��<���t�m*�	yN2�M��1H��'�I������"z�6i�>u�.���~q��y�~%������(�%����TJ����s@;�
Ӯ�#2��gG���TQO)i�ed`�#=�)��E����tq�Q�����jn�������F�x�c���0Z���a�B�8.K�+�!z�%��DYCo97�D����3Y��Y��6q���D�T咢��3�����o�(��N<�	�� ��O���ON���^��؈su� ��">��:�ד�dP��1:v�3?�!�f�GZ�^��U����H��S}�*�Y(��ϻ�ɼ�N���M�hY�|q�Mp(�vn~Ũ�e�eϒ�4��7'ѡ��#��ǻQ��i_��ì�Kf��B��\Xk��(��,���|�/��@ӃҝB�}񑝂|�.�#�N��cl�;!�IJ�SRLye��̦�$�9Q�6���J���,e�Z�+�$��)2��0#����Pfl�t�8?=��'6�5Rv�J�6�y������Y@Q
���D)UB�jp�3>�	�`ص�B��0�Ȭ��Ҡ�U-���|�U��*El��U��2��XZ��}��Q��#�ʇe�{�J��%�W����*� ���$:S} �C�Cd,������r����M�|���)���Ç]�����o������~z�����7o��~�������������?�����?}�a��R�t+`��P*j<�c����^Ol��x�!�]�Z�������r�����6��V>��Fk�@)�.F�}��C�sXZ���f%���X��φ��CS�6��cz��*s����.J�q~}kryup~��u?˜Sʾ�Ę�����Zw��ڭ����_��W��ى�'�9q�������_��௵]VE��LE�R]��ԳZ�)=�}:�w*�s"�u\�<����0��FG7P�������o�Ob��<��/�)2J�k��&�k�;���[��m+@Y�_5�V�n��z�j�=��5��u�Wue�[ˇ��8�����USi_[�uWɫβ~�`Gy_Kis�`K�p;���d���uk�`K��&[|(\�����ESEwc�����`�ʩ��ݮ�RUF��{�����=�ž�����}����/bF\��+�3e������������U=u=�`p͊W-���iG��u+<�o���S��+�ktv��;�s�
%~1�A�:H>���07��*z�(r�"ሁ|T�8�aQ0��@if	�M
i���WY,��.Β�wZ�K��_�"~�K<�K=�A>�A
�M�&앧���*� ��e��jK~�IU*������i+�<
M�q���N��G⢖� SDtf��]-���Z{g���2��4�������Q��Pln�(l.���4�������/k]=u�
[G���o.�m,��ܦ��������̦���E�d>�]�d�B
�q�H�k��� h�W�le�#w~��O��Q���F��s���R��Q��t��m�Ue�ol��#�W8��؟o�B>�K�؆�؞99	vïw����v%A[���Ԫ�o���R  	|!��ù�žbd�2pf�f�������B]b��Y��q��n�Z�b6�\�|�&�j^,�^3	�D)��ŗ���������Z���'�~�B�g&��F? Lۈ6����̆���@J��Ab�g�%*�M��,&WW N0I����DЂ�����	9�4�<�P��+��#������,��nR�85O��/N�$�pr�)�|�W�3Kb��	&1=�����s��v�TN�Q�O����GU��J��J%�:��L(Y����T_�d��Rth��v��n@^��/V�%r 4��B��|,�g��p�e�L@3э���7�jE��mna|��:޷��(�
����-�]��\}�vmť�2�(�"JC�rk~By�_����*�SLt�8��#W��m����PΠ������[;s˳%~I���"G�W��2b�i�Lя&�H>��?�Os�u1�vFU�B*��7�㕫��ڧ_O��Y����h�������ٺ�>�5����Ӌj��Q�Y
�8�>��F���Wg�gG~�����iW�����/~b�ߝٗS��Q���l��f傁~BK?��}.�w��>�f��)�=���,�o̬.��֊
�|'[��H|U�<�,���꯫j�nmik�hmoj�}�V7��8��<�m�H{�Hk�@]�@C�j8���&�S[�]�0�U7�U?��v��n�y�hg-py��z���uK\p�ڊ��ʑ�򡖚�Ά����uc�UC��6��wLt���i1����~t0�4X��j]'��'�~u�؝�����׾��K���8t����u���˕��J�pS��벑���і�7]/'�^L<o��/a��z��q��f��r��j���u#l׍���K�j��~���
فO���%�>�+�گJګ�������c�q풑tV�ڳm���"��C�y�G
Ζ�B��ג@�_k�gf��dQ �����{)�igT��l�$�\�dU�Ʌ^��Kf�	L!ٜvQ��uT<��SQO*(���Fۓ�S��uע����~Z�C���u+|
�=u�#�['zZ�_B����e�>����B��`����u`b|ppb���ɗ͓�e��������s錓��F�|�c�4� �Z��]����qG�����+{�s��?�;�߮����{l��
��Bc�5����3���y< n�[��Ήp0�\�'Nn�S�l��|�&{w]vK)+�m�=4�@G_3���y����a9��,6�:̈
%_�`�iә��Y�3�g3h���&�E�Et�$�g���
KV{	t ��*M���U�y�dF9h�l�GV�+��F�"4G:�Q��h�s���QV���Yc�1]�a}�#�H&�D	�d�L.�|�l.�L�|�\�B.�R�J�z�Z>�|�\.�e.�/�Q.���R��h׭��6�5+ڛ�5'뺋}�͹�b�r�`�m/�~�q��q��|?(yX-�����j П���_�����5�����{er�&!
��(R���b%(h���f��t/J��F1@�Pa���2��$�RXl���nO�aE�67W6B�b�B)��VVGG�����f�7�6��6W���ߢ��[K]]���`yA��A�st/�-�{��Ei�Q�5�卥�#������=�"8��!�P���'�V*��~�D��V-��-p�7�#b������k~��q������[T�
�,����B}_��^x]@A�@휆qYG��Ou*M��%�9Jc��;������{��ԡ������~s��#�SS�MZ���U����ʽ�I=���1�ΦsO�Y��:�I- }E)�hi�z�b�� z~c��WB��ff�\��+��>�Ư04�]F��̢����L�W��G��>�ѫ��벋�]z@�Q�3�������Zr�L�ĥ�y���t0�_�.2��ڒU� �� dN�ң���*�J_d�{�-����b��H,մ�k����5����_f�#þ�J��G��4�������q{�_����a���_?wmէ�W�z���*u}��2�YV��fY�2r��ņ��t]@��kT��J�R�Qh��j�Z��l��t���)6|T^�IY�~�W��}Z�Wj�a��tHG>n���Q�M�;��im����|wۓJp$G$ �)�t�mܯ�I�3IG�h`���į4i_�R�I@�s*Bx��M�WZڝ�z�3�CNv�%�R����q��A~j�a���ex�6W{����+�T��R�V]��+�2�dfW�K��K�r+�+

*�9���*<��������'��8#+��d��dW�V��+r+�uO���|'����K�mf=u��2�-�%M��̔=���x�o�a�b^�[R�Ϟ���$K�-���@�C��.y���HB���^+�?v�Р[�<�('��y���ۄ�&w`�50ؒ��T��X�&ܢ�g�����"L_��^)@�;��"_�°��W��e���IiS��҅������ն�*e�	�i���I`-��\&?������x�r���$�[Ws�Oe$LOڟ��W@�[H�g!�P�Z�G���V�Q3츃r�F>f!�q�N��睬�vl�q1O:�lԓv�鬓~�E;�f��2���>�/㜟�g�� ;�g�0�TpoV
��r���oV�nEw�$��e�j�ѵ���&��B���7Co^VW}t��n�3彀,�H�T��䲠F�硯����3i�L���F�o�B�OL�ʨn����jd���l������`���^�οx��e�����P^��Y����yk���k||diuly������M�
�.>h^�WDu+�^s���VT����2Ӻ������3듵=��Y��]\�����YŢ��^ :T��DRX�p��2<b�[!��{:*�֧g߭̽]����Zٚ\ߚX]{�0�4ԧ+6�U�dh�팚c��J�%-�M�l�V���0Q�=w�ȑk�O�:q���{���������� ��[��Z�i=���}��:�c�3Nh�t�K*Izkk�����2tls���f�y�t"�N縘/G���<�O����~���Wz�
�@��*}��/�r��9
�gps5>��H���`�m�W��r�l���r��n6���y�P��	<l���q�y.�˅�!l�\��	{�J?�P��.⚊�RAeP�Q��5,�e��玞BvԵ�N�����B:�S��_P��峣u���4Zտ�+�m�]h4�*ڪ�5U��2���g.��5�~�U���z"7JU�w2P�f�����0����sS�ʟ���S$��� ����&_ֳ�*U�-���h��drM���2�F�ƞT>�����)��N�+C�W��Y�C��鴃�=�LC<�&<3I�^��"��j�`T3ŕFt�ƚ�/HE��%'j�0�4�pVB���|��
���g(O�yt��FFw3�1�t�y>�>���/�q��m6|^.��Cy�=�$�]�9|4�I|�d^��2C̉���`K���ɦ����7QS\��.[y�=�^��>�w�t�S��'�O�zr8�y����^��٘�/�]�'�S'�$�1���w��'i���d�� nh���X�@Zov4X_T�{�]=u�Mq��6>�(�d@�{ ��Y����"�k=���Xe�n��@���婢Ky�����
y�9�%���?��q�í������F~�>���<40�r���"G��W�Ҏg&���'2�Z�!;jc�2�h���V�2���u�� CD>��]��ι��|��^��z�g<@a�� �B���	��_��R"�R�+f�](a_,�^4%w���ޮ�ݮ�ܭ�>��F�(м���i������_�1�%�_�D�.Q�/�G�
Z�����(`y�L4������ac%QP�$9ɦ�y�Yե�boF�/��,�,�SY�]Y����yJ�UK�j-�PMʓS�"[��y���A_jeX�d �F97@D���3o�vP������١陉%�m�㧏�~�\�Vެ����V�x�{`̫(R�<|���R]\�[@�i^�+ax�`,���U���zky}��������(-���zsOwAyi���˹��7c��Mgê��5�2��d��0b=�g�R���S<Zw������ �̡I��:I�/(�/��ӕ�.Ze���ڙI.��t�E%1LO?���M� Fa�ǿ�.��SZ�{��}�c�|�5~LD&�ha�l�����EbC@��	t^��'����c@��Ð{��!u���>d�S�F�^��e+.@�e���fb��]��כ�d��,���s107��F�^��lY�(c	���c+f�����bc����G||�F��/R���q�x�ͻ󫴳{��~tz����ޢw��M�T���� 7P�����K�� M�I4����Q�}���6���r��~�`�	�M��K;-��/z���8���hOf0/�/�ر&��ږWgw��3�*��)�V��l����gՑ{e����LO��'��?�r �3pZ��z�q-霖� ��/�Ҕ����r%�����݄Xsj�,�W�_���Hq'�k:֓��8�49���`:�ˣ�)>ՅKs�I>эN�;S�n�Gd���"'@gzIt7��]���P�+�=�3*�K�{�/2��?[i�LU��`�\�f��f�̤O'��_Ά�?�[�����_X
�\�2:N�����t	�-�ͅ�v��>���y"#y�6y��/�v8�~1���.}�FXQ��'.&V3�R:��
����@i������e���fgo���5%���J�y2�]�h�<�,�0I�%�����Nb KPmQ7zL�U�W���&o_������&��-(�H��0:ӱ8�c�i�����)�75�NL���T7%�E����6&��J=P ��v�B?dc�1ۙ���6��h;�|ʁ��Y@���#��B{��;�ႝ��Yg�h7�Hp���,������^.�T�+�\*��1F�V�`��*���Z��Et�*�V
�3�W�f'�_�5����Q��^��N��N��N@��H�T���(�eJi� 
��E�1�B˻Ch���465' �$D��`�LB�ID2��˭E�V1�)	E"��"0졄b��_�x��Or"�1�^<�Ȕ�R\���7[[�;۳+�%u�������������ݏ��|��w�|����oޮ�Zy�6�vnx�7�4��,��2�K�q�E>Un���֖_mu�wU=���YY�zw盏;ߠ�vK�[S����]rW6S���3�j��yᗥ\�*R��yZC?*������YE���9T[1\�iq�-���ՙUS(HnA����f'zX	6ţ`���;zڕ��,��L����|IX��N���շ�9��VU̮����d�.��Nr"�kR�,�]���Z�9�ꂒfGMWQ�����������6��(\L��L�bJ��s�9��NuP�:�A!9h��`2\��"�X_���9�=����5���z��/��YB;�e#�m$����	N2�A�K�]T���C�p�E��2IWP;�T��`��;K�����N���ú���A�ݣ)��Ğ��I�2���CU�]��ּ�]SPTV�s��l��)�PA��T��Hq��.2�F�g$�(d'�l���,��N1�q&rD.�.�,���p@C<�� :k(G��F�謩qZZ��6gF�R�K|T�O��F�%�i��+��P��1�|eLݓ�H�k L'�?�'N�5R�(g��G9~i^F����N�Ҋ�̐��o�]�G~żt�+�;$J	lDf�E�<}EaA�]W��/�w4���w��=i0M���T�� q�G���4gl �1jCK!�H/�������"�ۈţ����L�1#�&�2�N9��TTeW��6V�<�Tu�+ڬ�vGe�������H�X������ҧ�� �M�2���r��'N> �s��	�N�#�����M���6n�_ɪ�ѵ����c���&[W��WͰa�*h��m.�i.�k-�<�����wG_T�</����^զ��im��o�'8YqN�3�����;��ȀрllY
)���]t�P�]7-�F�^�?���X>~��r�t�� RCh>��C{��>�d�p��N�9�\lh��g< ��ʰ�s��:�e"s���y������yaż�%����`a傋]��_
oV�nW���TI~tqpks{簄��K�C3}�� �c��˥wJķKŷ�ķ���~Yl�<f'��8h�2��^6��ż�P�$ј�F�F�]7�b�\�@%"�I(A� =b��B;� ��+�9=���BK�m�$+#ՅV����QL�ODq�E~���������D��@`5�܅������7�[�o�w?����������ań���w�6F�_�>/��[F닞�����wK��./�__�������oQ]�w���A��'W�_/Nz;*9v5�&�;�T�ݿWH��%:e�)����e]4rO(I��ie	g�����gv9�$#��a�t巘U�n��&{��>~����a$;T�$��U�UL��d�.��.f.d���f]V�s^���n�n�d� ��S#�|�e)��0�;����W���y�2��5�����~��כ�Qr��ͷ�#�i��#{�H}[uGyS�������K�;��P�I�UY����8^]d�zU�|�{b}ffsazlnrurbedx��}���dٹ������(k�*�"�����ۢ��	�H�(J$O��$�+򖻃�����+�gѸ��)W�0nݠ޼�tI.��n���޴}�)[��Lv8{��G�$M-y���+��&}xE��2�����$��"�*b��������|]ifB:�0���A��!u���W�?��_�s�
ԩ6��.�h)�5�fg�Z�@�fr�ļ���'���_���'�d��ݟIB�	3('2�Gd`�	���aE���bmsfV���-P2΂?/��z�'�8�0��&#?ɒ
�ӫl�����r�A�<D����R�iI�Th�ݩ8W*ޝ
��z��h����#�C؟�J�';��p.\��2R�D@9�G�zɢ"��*CY��hW^�d�Od��S���Q��-�������E�u��m��e���ue�H��; ��zb�_�!�$|�Mܗ��7d��p�@�t���(;�������j���i�m i�1.Q�WIU5v�Jo_C�HG�����PG��h+�:*G�jƻ�F��;K_��pv��<��<�[�`���9�.F��sDs���f�8i�vZ��n%G٨Qvr��m��9H����n�S+�p"+yofҞ�^e��v��<�`�v>�`u�O89�ܼ3^�IH}��	1�������{N�y?"�6q��>�g��1��8��g�8���J�J���J�ʹ�����KU�K��+A����Z��j) �A�4�VW������A���_��c���[%" ����Q@���j@AK|I�4�-W��e 萎&�Pd4 7d���� k2����="���w���\h�h��+pN�ՙMu��\Iv&Z�����lH�{��r������J�X��c��t�B��s�h��_�\�Bi�wv7�}�A�Z>��ߡ4�_oo�n�����������>}��_��;d�}���|�z���h�U�ܮ}|�r�S�ˠ;�d��h��	^!�'��D,�<��-*�{�c�0��k��d�eI�ı'5�wL�h;?�%HvR<�4�4�/M��}�� ��Ktӓ�T�����+ꫵuT�,��鬫F0�|:�Np]���~��^ۙ[ߙ���!櫮(hge���o��gi~jmei{c���ۏ�>|��'���v߽��y�9�:U�]%J���>.�>�yv����)�_P��c?�ˍ�Ϗ:�}z�O,�֍�-�l��n�̭��o��څMhW�6V�7��ڃ+#Y����'�1��)g�qǥ��$ѧEOn����V���ss�K�}o'z����?��|^a��$餱`�l���5=ճ/k'^�,���MN��YJ�"Y�9��q�<8�����K���������{x�yC��w׽��[��|3h먺����Ȋ=��}
J���\���2�/ZJz�W�z�9:00=<�4>8��������Uq'�O����Rd��P��0f��Ҁ�{8��H;�S/e��*����Z��ӭ�^6�K��p�)��ɗ�;�1�帓J�I	����P�R�������r1(n�9p���^2�GBhv���|��Z��%��pe�Mt���T0��Nr"KqR=�xj�i ����^�Kz��U��N����'���9�K?�Eڧ���$�>�F>>�LM��i~��L��ΒUeP�8���q)�pܘvP�z(� otQW�quj�*چ �fE��F�����N���M=t0P�'�x�K���I>�4CV]�op洗�:v��Yz���5�%�z����Y��w˓��0��}f.3�٩ �c=�x �`�f<�����Ѭ`���"Ż)�nT��s��t3/��>fof�^~��t�og �:ه�#�q7ﰓ�>h������� k r�ˠ���Š�O:!��q'���y ������y�J�K�` ���e�� �
XX��R��w�Zt�J��:YМ�ܞyLA���@׏�H�1����2�bɭ��a�*�XW��#��H E�f2=L��7�N�u�<v?�A�b9P�QJ����ܨ�7�'"�Ũ66�S��{�in&�ǧ���%���@�P>h��ć���0��4L���w��y61���2�MK)4���Ɔ;�G�fG'W��7��v�b��P-D����͏@h��~��E9���ztkX�!,��򋉡�b�Жζihpq� -uAQ(z���}MMAAW)ɮ��e\�QOi���dI_
��=���3����!���!d?��-�d+��{�;��2��Z1��쪠X��0g�8 ���=]�kkog7v�VWkF�ⳤ�4�s
f�)?02ѽ�*M ���������f��s+K�/�Ԭ�
�I5�0�X�$��8��$�"��1F  }�#�afztc�Yߙ�+��ʭ��XBj���Ř�YZ�T��>�S��n�O���a����^���������}�n����Λ�O�/�c{��w#��~�a��͡���4Ը�[7�ײ2=�����	�ͻ�ݭ��)S��I�rB�tD�|T��_�x@��O�pT�rEC��-/��gvv�`г��6=�������(�'����v�ȉ*Ԗ��o���l�2�?��i���v�߭���	6���g5��(�$3HE�3��F�>�I=�I;����+�s�������/�R/� ��4�H:�)��sA;G���VS.�WT�g�rE��li���T9Y��1�"���9��#͙:���N8���ehS��d΅�� ��%��x^��Dnᵼ(�<��_�e�ɦ1�T��ZyPu.#�F>����nb�[�L��9i'����ԉ�2�G3)����g�c�Ryf�WeC�gDg3�AP4ߵ��X�w��HJS@JG�XX4;�Ό�s����(�!�;e8�,�!K�K�x�$�-~��F;X� ����?u���@8��`L 4rt jS���㙝h�s�\��=X��|� ��!v�1�}v*����v�ņ }��=���C��n�	�O "����<'��Ny�C�r�8h���9�� ��g�x���E| ��2��
aX� \�X��Т� �r�j�w�Rp�t��Q�<�N�`�5�w�!@�LOL/�֏�
*4��з���wK���%*PД"9 Z^"T���� �L�PB��>��PLt(�t4&��AA<|�� \ƴ�g��8�`�W��Z؃։��l�n4�/@L �(����ө�X�@g�%�@��]B�SJ��y�L�Y�+�k��������޹�����卉��7k��Z>Ë+(��ƻ��w ��խ���ѥ�ޙ���^mQ!�*�9$4���Ǆ��B1yXo��yEl�*��n�(I���QO��Ǖi ���=☯�Q{��$�G�1�ձGeqgdiɎ���*��`vU����8B�@Y�ɯ����/��f�#}�(��W�ˇ�,m��n�ZX�P˽�g�iX��/��g{���17߾{�~��{T|�� ����73LH]V��hi����r�a�Ɓ|RE=�e��PϨ�,���fjj`m�����**o���zfeF�+�X��D퍭����ݷc�� �:�E#~���y4��cqf����VwQ�e�������o�n�[�ܙ�zf໙W?���#-K}-s����'��W�7�ַw�wvױ�(�[���t�MJ.q�@E���i-������{=����TPuq�m�򂮶覚����t̀Bof�DUEϗgwv7>~z���o?~���������	���͵�)}CI��~$��/�p(����kc�<0�P�d�j� ��.�ud���������{����=3�����e�?$�=*O9�"�VR����b�7GWe�txt�\?���Rd])���x{j�# �Nr�&ؓm�8r4#@����MHv�R�i�� HA�QۘG���$`4�KF�k?�姱}ly����(�Ňw���q����$Q�K��"�W��_J#+cNhbOj����G�R�+ٓ���� ���_�b�8�Ĳ,jUF�-Qy
��E@���#;宕x�B �e�ߵ�n[	wl�;V�{X���-=��|jg��8���+쩝�`?�;P��p;㱍��F�pҢ�'N*P��]��InV���b�9�O�X:�X*{��&;�q^�6�\z�W�g{
qH8;�j>��|>��us���!Q���q��8���=�dq��!l`tf�����= ��aE�g���h��.t1�t�}��{�\!��A>���+E�?(h �F��V��A��Q�2�A[��=��$\]�@׎V�t������X��R5 :����
5 ZV��|?�3����@g��@Y����C.i`4�R�XB8���҅ b�1�萎��f�|Nv�Sܬ��N�p�E�(W�竑�"��Gras�X�R�[��E%��d���T��:�E�w��<f��j��[�uA{CUf�7������>1�==��f�q���e����P�93h6)ɉ
qaA)������VCc)^$�E���2}�=\ϸ���S��ˑ�c�(n�����_�"�^��uA���޹8?�4�j�UY�O�+��W��kL�֊�zkGqj��A�f��^��X_4�.��-T�3<���%-�z���V�����.��Z�����E����n���(ۤ��f���h'��cJ�9J�vZE=�����]�Y�]�ZX11��?��f~damje ��\^���Ϭo/�[��\��7�i��Yq&C�̛���s��w�6ߢ<�;[��[����6�v��f����W��{�&�*G^��OM���,cI�W��-����Vvޭ�ߝ�^�u�E�W�Y��Yg3X0¸��ᬙUCS;;�\m����G�W]/[��t�S:|9��@��R׿������{�zm�-6`ښYۘ^�Y]o���V��;�A�R��KM����F�+m���t�t���S�ZY��nv;��9Uz��tf��d�iA�9y 5@ʿ���{��O��'��3r�M='Ѭ�m�ZW~�S[�?���E ��J�cl��h�x�H��"Fj:Ս�̀�47$3R��~l'.ٕ���':R`OHA�C��v�&i^:�'0Te;^�����N̓B��l֩�Aa�&�KU��
�)���8�W��=4���?�פ��Ni�t�+��Δ�l^�)�#��3�y9O<l�2b���<����m�f�M>d���HS; ���"��)�F��@Xh�h�|�B��3�P�`��r�hq���@D���i!>����$'�c��Q��r}��x�?7���~��F� � 8F;�t����3lr��>C����F���3 ��17 ���30����>S�9[�;[�E��R޹2��r>hѥ*��j��*��J> Eq�+�Ѡ�������W��&���*�u��G�X��z%����N(V�J��r�,I`	�,�������0Y>�t4���2���<�0jCt�s�0��^`��`O��Y��.fС=�4���D4�Ӂ�hj=<
 ���M�xڌs�H^	�-���Xd���1m2�C�vʨf�P@2�)f���@Uf�s�f5�$%�P<	�Eq�Ρ�<���|x]~�y�:@�1�2u���>��:���tQ�;�$W�;�*�wP�|�$>*#]7��C�/W��llL�/O�O��n,,5|"�Ob,�Z����-�4�<"[p+[|3S�䴪[���M�"�m� d�U#璑�b\U�(D��OK���奭������Bt��݅G˛�fFy�*�9-�qJ�LS����3J������sa�z(c\��h^Y���0=��9��ʬ��F�_M��ͮ ʧ7w@GOﬕ�Eerf��_���1��;���[�斚ǧ��߬opW7w6��g�޼�k/i���U�;�ތ�^\ZYZ[��h�9���,K[o�vޮ�?��"
�7�@��1�i��
O����������ج(��y�fc=8���_�2P�FZ+(���Z��WWޡ��(�4�ye}baux~�o~�uv��������.�C� �+C2l�1�Nf1Υ3"MRI�5��i��v�Lg��$=�K<#}���h�(f�4� aZ�M-;Ū��Y��ܦV��&��R�d�3����)IN�9ց���>�&�c���v\���AV���`�H����Ӊ��4/	N���$�q�A�Q�~t}�������g7�������m�����Nf������䃺T��ԉ{5��;�A����Z�^6/ţ�T��m�`V�9B�u��A�F�H��V�����x�L�n�]+L�j�]��[	!F?pP� b�����=�SXP�W��&�����B�Y�ܬX4 ���9�O��H>Қ��FHt�C����rR����lt���f�� (��@S��`!@vҎ�X �c�������揦�p�0Y�<�e��fhO`�u��}��V.� }�Jt�R#�\)�V%�
�Fz�N~�V^�@3�s>�8Vg�G�DuƄ*�
�=��_v# @?.R�hY�@�c�}L���2|,��M������43�Bn��iN�7�]LN���g:�Pu��[#D�PUo���	U����v�c7z.:��[��U2��	��-Bq#������Ŕ�d�\��OpH�6	�
bYNr�nTH%����y�ٍ��A/'�AKtP�)(��d�����j`t����[��eE�w���(��"��uh� uOH�a
����kik|�H�ŭ��͹�������]F@�Yl��؃��m%$��Q��^��FtO'����V�o�׵ �����Z�C5'V+U�u��A�.l�b�ѻ�?T�o���_N�Q� ��*�)%���~Z�:�D�G��g�,���<3?��t~�f������׵�ͯ!w��[�s머������r�󞒮^����������櫥)�U��(���l�_�]��]Zk��6�����%����[� �76��V{z���:#�l3��[Z\�<�o�PzҶ���ɹ��U$��v��}Xx��n����wIK;�e&X2A��l���_���x�~�Gy7S?1��<�728O�rQ�=�&P����::�[�K��3�/F'�z�흲`YD�s8��mʯ0��k}ҞLJ:��zjW	���:��Õ^���9|�㥒��8���Aq�AE�!E
����t7�K�������6��&���\(Zi^Wj�y6 ���i��j�hk�[`��=%��j�_1���mI�b)���8�8��X�;��"��7	�"=T��@#{�t7h,Iz]!0��2�.ʎ1K��	��z�H?�#�ᏧS��IGu�:��L֕,��\^x��ME�gH���2'�!��1Pd����3��N����( ��	Ì�증td��td2��gF��� ����8��}3p9T�����@ce�X1NZ���4��m�G�p(��')�� 5�N�p�/�����#N�1� Z41��k����a'㘇y��F� �F��Ԙ�>�f ��� ��.�I��4�����8�g���s.�	.V :���7��H�ї�$��U�kU�U⻵�{5��5��Z5�6�w!��f'�K�u ��*՝2��R�"�m��Q@_��+E�2��+���>6Z΀�!Ă��(��ǌ �T'�W��uq ����{\LdN�&,�i b��*(S��E���]L��a�,��D�Z1���$�b,2�&�@�Nx�p��N�����R��<เũnA�����y�(4Jn��'����H5{i:��Æ�^�n���?�' `Ž��9����ᎂ�bJ�"FϊHg�Og��Ӯh(W�T�U���xl�g�-�jq{�����vi|q��UmQ��Qar�8k��}]54�6![��-{bEj�O�H7JωO��T�RG���Q�Ǳ��0`_�\�y�vkg{����66��.����VSN*�����tTI>,#�V1�(��==�kۣ�;���ս���<���rzqz����{������*����grR���Z��g��v&7��7W��z����9��rj�lb��R�$[y� |h�ttn�]��vs{kve���'��4Վ.̡| X���9s}��$+*-Y�\�~���������y�-���rM�Q�V��-�^ݚ\ۙ��n�@�$;�����S�iY��Z��|���PWeϮ��>o�X]]�D.��fQ�jsy)^��Ԉ��9@��>=no�׺����F��l�)�q��4�vFt�6H��l	�S�zN�_~H�xL�?�"�W�"���CUnI�utx�5�� )nr_�v� ��l����h{Z�5%ҚmML�ci ����n���$GrX�_���g��9�Dt]3ю� ������Z�?6P�37���*����2]���4<�>����a�� ).�ײ� ��ټ�<a�YN��<ƶ���I/�ǹy��l��L��,E���X�|�-�&�´+�4Dgᶕp�J�g#��FQ6j����������vϔ���@��O�c!��` }�>rq ͱy����Ċ���=����p#�W=�7ng\( 5Q@2����y�\�#����6:2,r)h'�hsC��],��pҁ��4�# �݀f�I=�@t>�r� Р���`�(��R��r��N��RP�9� ;�!�D��E7k�w@D���1@3��^�a�8֖���J�8U��
�à"��B]�H,S3JT�RP�B���$����Ɗ�� ;�p*Й�S�X����t�4���1z�\��;�A��1�hl���ј�:$l],������b;�En0�^��BI{_�%7'�������}�/iy�G:�vNqӒ��h
l'9AA�>&����%)%z�4�����6xP���VWw�2h�{�ife�Y�lR�(h���b���td�����&*�
�X��X�^��]]ݞ�X�z�����2�]����rvV��P���2SKyѫ����׫3�����������]���+o�קVQ5`pH����fe�r��3-���zVM=� �T���I`��Ϗ�ұ���S�����tQ����滅��k[c�k}��냋�k�����67��;pY��/����no�/O��O2Tx�SX�W��ڳnf��e��fJ����!���r���dP4�z������- ��Ԕ����Z�Ѩ�U�K�K;�P·���ƪ{j��E^����Ŏٕ��f��Wց�kX�����W�|svJ�\D���]�bT����
���-ll�-.v��dV��2dw��KF�	#���-�  �e����ϥ3 U�j���njs��� O�g��J?���ԋ�'DQ��)t�kz�]�������ܶ�b]U.��N���\�x��3'i^	%�q��8p�N\�59�đeKyjO~jO{�֤8[
��8k<X�-���lJxbI��v��NB�������NEj���@R�$ܔPw��/,�嶺��5����M~e��Y��lSA���@oRЋ�uN]�����j��u�(�M����
�>��#��(0��(���tߌCx��A�>r�n �M�[f�mB3��v" G�+��=$�A;�7�޷��E �w
q��xl����{l'Dّ���� J9�I> �A8���D 5 �����wQ�]t ��|�B�~+�((h��v�+Z=;�C���J�6z�B��1�����t�A	-/D栜rPO;���.l��0���@��<�3� �+�"`��R��P��|�-�D��yD��i��U����cavji��[�
�b�(̮r�X���Q�2�D
ZZ�V�ID�P���к�6P9/�ޏ�,��M܅p�P�@�
y@�E~;�AdĎ�x>	x��t`1���1����`?�ЕAk�D.�lȑ��h�=���('z8`�ȟņ� y�@F���.O�蠂at���} 0z	�%�s�ZyE����x��j�y͛������ڱ���vcБ�!�JpV����e~chu�8�i]\_]�����v��ۍw;Kۀ��������Տ�k߁��������;�|���w;?��7��� ~�&��ǧ�AP� y K����*)�WՌ�Z�)鼖~^�3po�%d��}i}��'�������"�nn����푥���1Ks����ir������v���ek|�F���ϯO�_�ٙ�^�~�$Cp;�{'[z�@y-[t=Ot#O�0GF��;痖�z�+[[#K�Y�%����������?������Ņ���8R�0������~�|�a�Çŭ��W/#4Z�#��K����y�������3��������v|u��¯��j�9���b�Ɨ�8��*����&t](���G�ow^̎*��=�d:�p:�`:�(ZnG9g���x�KA�CU��y�L��"����&�����#���$��By�7��,����\�e|m6�{ť:���h%�X�Bz9ʖ��Iք,҆�vRJ����O�)HGے���xGB�Ζ�$��%�%.��Z/�`��[ь"�9�Ea�pʘ���sBKIu�Am�/��l�LQ���(nN��olQ3�׭Η�(����P��U����3����v:hX�)�A�I�v��`>�;�9T0p(|��M�Y�v�Dw��1��T6 >�J����� ��(��gJ�S�r�0��	���h�ᶴ+�3��Ζ�.�4�ڨ�K@�C t����W
/9�E}l���#5���p]��t��5G��\>�b��1G(h��;�!@#��SPF$;휃	v�ż��\�q/{�aN�y���y�Ͻ\̿V&���.q�:�!._��A{1��BW�/�H��HC��n1�4��������7�t�Ks��_��fW�1�
eJ�S���<*V'��Yey9Z�"��y>6;�f`Y8Bz+vE:�T���<�.:��0E|t��y?�!4%C^l�b$o]h?�@	J$-�s�!_�� a�94B�)e8�@��OB3�� ��C��{��t4�9�!@cQ;H��EB�����	'�up'p?�ٍ��=�%l�P��)��\�Ϩ.�Ϩ��ڊ�/��=u��My��<��0\��VԔ�L��_~���M��o"��}������ov?}����>/������� ���ݏH0n �����j{��K��Vgy׫��- \
4��)��0R�z�a��q��X��x���FQ�Q����Y�\�� k~}�Z���������ͭ�������>Řn(��~�9=�0:�����l��sam��7p�Ƈw#�3�1*��/~�'��/~�/z�-L4i���P�`��pc�g�Ȓ/sY{痖v�����xzk��eG�N���6�nn�D������MKW��y��b�Ǘ���D��|m�s�'��<�z���������٭/׈]"CY^�H������t��-&�CΓ�o�ޭ�{���zډډL&
��S�-ri�5�ޞ�b�U�nJ?�"��
�Ω��<=�J>�ğ��bM*mCI~{���:����S_<��z]���(�Ǜ��#��O)�G;H?�8ʎ��㡍t�[S ��!�F�y��4X��f`7·	���8/������G�U���B��&͜�$�� ~q$���S���u�&S���Y��*st�8�ʬ��z�����*R�x+����)v ����mi��N*��pK�cs��5��	T0R� \�P6�1�	g�wT-Ίq�|FuOP.:��hp��9(�c+.�4��@�;~�`qR��cn�1b�vC}�G���8/
�}��r��D!�N�	'礋{��9� 5��3 46IH=h� �C>@�)���}�˿������K$�eҘ�"�Z�T�L�Q�W�b*%�傈
�"��b�5?�R�s�T v�Lp�����8a�K�����+U���ظQ#@?��$�f&6��9��㘂^��(��Tkc��Aսr0��2����__�d�*�*y�@�er=L^��g��y�	N4�  �	^d��~L�b�Z��d�/����H8c�D�^6	H�	�$77��O!�
�n¹p$��%��<!&�ѕ�!b��x�;�\����ck���'����Y���?#��L�|4<)Hc�	�^���z��@�{E��Ft�J����B���(1�'�)8~�#���&��V2ؒ�X��)y���ш�
�M-�#S��}�C�cKS�hFnq�Fqf�* Th�Pl�������Y��]�	44���j���v�k{g�'7����94d���\�'G�ʔ�r��Eq�ě/v�|o[�������`��n�R8��~59it��n�t�3K���Rm�&u����ޥ����@��o��ڂ�|e�YYa����%�����oia������@�Ϭ��57��x���V>|�����b^���ym�,ͯ*��Lln�}�f��7��u��k�V�Ǣ-r�\[�0#���}|z�#� �����fO�?�� �E�:�Y��58?r�����<�7P�Xx'޽�\V=aj�	��M��X墠)��ans�*�</��&�<ȳ���<z�8
�|RK>�"%9ӵM�٭�ƆRi�]�QD	�FZ����M���;f�C#9��W�b�L���1��@fOmG�S#l� ���8�t�q��'���8'�SR�O��`��d�p���ɮ���-�ILv�eu4����8NNqQѐI"9y4'���7��������~}h"΁�P#Ǳ�D�A�B�P�����351:�^ ed���y6@���t"\΅�"�ҏL8$������-D0�8Ԍ�K��ȡaM�w&�E:��O)''�2��L�PR�d��LT��cD�i�
�'̌#�Oz���cv�	�th���9�X�3Z7x��:e�̽���KUIUzb��Z��W�i|r1�TL��0�elF�K���$�zEr��iP�H]"�Z¿TʿRοD��6��
�*
�\���ݪ���)�4jc����+	��f�z�cU?%F��o�%�E
V�BT+�� h�Ŗz�������8@c�^�d !|�O�,4�A�h݇�?��Q�N�'L�	��8�C������tt� �zRt�1Z�ׇ���#�CGb#��hFۡ+�6 H�Ļ�9���r� �9�14o���^���L�c���!�ϧ�xL����|Z`t�@����`R>6n���ղgy��&o�@pp�fx���ԫ��ᥥ��7++�+�Skk3�������듫� ���Z�{뺻�{^��j��koz��a�u�����b��t�`O�XO�P{�@K�`k�P;�ͣ]�-M��[G����ַ�?|��������껯W�?,�}�?9�5��:��:��26�2:�6:�>>�0��4�_���rva��{�����u#���&�W��u5����FiR> �N���5���k_uTtA��f~�����;���;>����~��������k ��뵍ΑᖱW���c�գϫG�P���a������w��6�F��A��H-�P�>�e����mS�=���K��_-,������:����&�׋�����b:�J��M.�6�,�v��D-� :���ZA3�:�+a�i�Q5ႁ�0��"q��[f�����g]�!_*�^0�/ZH����&�����X*���@/�C�gl#)ډö�#�)���� �]��]�ѡ�E��`���-)`Q��'��r���d7!�(Z�-lAKɁ��ɠ.�b�n���4���Ϙ��"����q�EF�'���)?qS�z�hۆ��F|�>s���D82
(l�ѐ�0pG|w g�	�G��	p�H���ۀ��f|����D�5񱅄ε?;��$x4h'��P�:��tAC�u?X(4�}���b]5�NZ�!@���w �F���T!���r؎��O�yg]�sv��A�4�JK��Q�*f�-�����%�oO�SdN�ą�x�|w�ObQ �� �T+K��=��-�(\+���`W+D7� ���U���>hzeF�D/���L�TOp��S����<�Tc"Zq�Tq�H��K4�2��֠.�H,���Ɩ��,z�KŸ�0��A��|F:q���2P�]��{��,[�A�B���^�+L��CX�ֆ��YX��5#y��G�%�9�'�<�7���87�,r���Bs�)�c:��C�
�9��x=3|(��P���	�L�/t�⡇�t�r�~��lhi~��czB�"��\�Wo蘒[u���Z�E碜w['���<��p��������5��5�/k^���Y���n+j���T{������5�m��k{��^���V����{Z*<�Ձ�z+�]�0�\?��4�Z����uK�`s�`SM=��֊�Y�H����`[{�����&��kk�ý�=M�Y�;�{^��4���y�9�_��Y���<<�\�;�@n�N����諯�*�@�6��blxbu������\Co�����H[�PW��ͥ��0b�c^�L�����i���|����wo�W�^�t5Uu�4��7�{X>�R>���E�x�S�[�-j.�(�+�,��$pvJrg��|����e67i���=M���[���-�������w7����ʪ��Vg�[_��Y,'��Iv����O����)i	g�H�NR_����vji^�O{%�c�3��fR��r�L�`�]���.�R/��2�b<��ȧaCP��H�x�S�3�(2�6Ltbӌ�H�	�ٙ
�:��N�w� �$�]���ƥz�j���C�4
� ��&�H�E3��!@F��3�]�$Љ����E�q#:�c=(]Qh�8�Ċ�w�� .- 5�Ay�dD�iQ���t���X�E�km$*g"��(�fr��JP�?���p�gh7%�D4�NHr�V�1��GG�/�䥣�~��^53@A��BhF�;��e�4�R��Y�l �'7�����V����2a�-�R� �&(��:Kb�59ǚbrl^��Ku�)6��K�$ɚ�IQ���̮���5��A��Jٍrѵ2��
`�FPx�B���UKP��y(YR(�~_��Sc�/JG��Z]| Z��Z
�q�"�T�,U�˕�">����*?Z�t� �j��:^0��H/cn������vFJ[�M��I������B���@��`8F���:6�に	�
"�_��C
W�p��\ϡ0;.��!:��LN��NG�p`4�_$9��u0@#a��p�a�pa$(*Q�47V���yx��	��;*���!��P���q��ЯJ�2�6ػ�	6�=#�Z:7��=�圕3.*���Lլ�یb{�̕��dI���(wN��8'=�e�")�E陨<�>��TJ�
)Z�F�6�<Z�A��:�_�Ub�{�/*���7`UT����"G��������Zs_O��U�{fq`~���԰'����
��]�@�O,/�,M7���.������o�Z�-8p��g�}z]Q�џc.u�}�zi�����뙙�mY�} SWd��uZ����o~yf}{vm(�|t(�ؖUR`,��*�5�YZ�\�x=7�l*<9r�ȧz�|���RH}z��hk(y573������ޣv�n�ȕƶ�p���ʤ��{zqd��NqYʿ�?2�5Uu-h��������D�\ZV���pw���Z��)��Q"$75΂SE��$�h����|z�KZ�g��s���k�����yi�rR�d%�-$����/Z�pa�T�˅��&|\1?�I
��A;?q!gt���@�.���
� ��7�XD�--֎���S`�-0��35$���h���=x`t����J�6.eG��16`=v$��������q�$'z���� Ghc�4���NR����%�)�d1���C9�4��D˲�̧v�!�w1⽬X�Kx��ډ`1V�3p���J|j%G���V* 娳���!����$��`g�_��5��C�Vл�=(G�CC����W
h'
��#V&�-����#VB��q��>ic���/:����j=�X�l!R�D���h-bU7j��(�}i����������a���j��T�@���Q�-gYK��%�b���((e0���z��*��2!H鐚:ߪ�T����ղ���ǵ��Yl���[�|��Ӄ3� МjmR��~T�/W�F��%*v�ZQ��P�QTQ3Dg/�4� [o�D4p�0&�w`!҅��H{��(F-���"l��C�5P�m�͠�Бn���� D4%���R�FNHl�xQe�#��ьe���Y�p1�v2�kL�ý����1c*$y����<i�!�љ^�xQfo�)\re@%��n>��c�٬ Rʴ �3��}?B-5�H�9�E��q�$<�2��Q:�\� [��9hq`:uVK;��]����s�N)�#{eҀL����G��K���+��%*�Zm�X�i��_���^�27S$Ux�rO��A+���r��\��<r�'�~x`hayby�wb �g2��Fzf���w������ף�o��QT���j�����D�Щ}��7c�����R��V�G%��e����jjlncsu�����Bsg�?[�K}b��'�����!�|v~ty(<����߭��+|�O�-�mx��0���=1�+.`ۥ��|7\\��IvR�N�.ί���N���XY��*m/1���$q�8b!��"�7�,墒|I˸�A�L�k�Wt�p����jxm�7����%�+O[V�_k�t���J?[⣉(x)�F9���'yz@�|PK8b��6���F�F-���3#�Ky�����Y)��_*b��F1$�L=]H5}�B�d#���CR����e>��>�$�c�d�1p��yh`@�g|(�#���)`�,��h����!�5���M�AE��(��(�	CgZ�;5͓��BKɑw}v���'����<"rX;��"�����A��(�pR����@�8+r���Щ�'���gv*�`�.�	�2��t�NtS��!L���D �#-D�3
� Y����%u���Я���n8�E!�i.�aG�7B�dd�0���87z�3V���# 2�Y��6%up�[p�%7�D�V�B�.�1���l;��Z?3������������ǿ��?~���|���b������������_?~��fr���9�_�R�4%Da�� ����)�(�_/も�|�0-@���UF�*ck�����q�ű�4;4;X>Vū��W��� ����*#J�e����EE^0��#� ��A��C�V�p�\�΀?h�`4����	Xum�O�� \@3X�!�ʊr�!��������|c.���@j����!����|v�`��C�����E�eh?�n{�W]�Q$x܀�a�w�������7s;�}�/�WZǛ�f{�5�2`-�8���G!.�@g��x�8~)߯1T�J���8��^�F�b',�yFG:&O<#��31�>���x"G���X[���<0��{�+7-�U�eJ}L���wӅ^6�����1y^׃R�c;9�L�	zߋ�޹y ���Dic�֞稩j�Y�XB��k;[`�۳��(�_N�El��}�����ѥeа��r�C�s����ơ��뫫owQ������B��Z�Ti<�������N���]?6�?����k��2�2 �b�\��h��_�]l���4'R�i�:����8��D��*�/�'Q8貎2�C�wP���e17T����8�.Օ�(��8Wa�^�S��X�4Rǋ�[K;�Vvvv�;���@�+/�QX� ]�0<�B�E�ST�E�r�@9j��Jg_�K
���D�>�&�cc���5$�J��O���S��??�g�a��>>�O9o"�3/���ׁI��洇z������@>G�A>�y�@� :c�
Ӓ\x0 5��8 �v\�E�a�
��1���`�E�L�h�Н��Aɦ�"��:�m��"b��Nt��<�t�-�B<\�'
kCH� ���7@A���Y�7?�7��A��!@�C+
�z�x
�B�d'6�@MG���6�wF���bR\4�X!����d�[L�1F#��	#����0S�n��<�븃rq�!5��LDj���y���}�Ή*����i���9�]*��|����~�������������_���VV�fgW'�,,.����_������_1^������w�/�;�|e,K	9��*�`��dɵ�GA��J!��_-���UIС�*�X���ї�zyn`���u9 :�Jt~P�|X���	Ъ�
 ZTI��X"�4rqx�`���È��)� |`qv�3o�D���G���N 2�F� �$P��<JB�������%�����@�к�Ͼ$�ᩑ?��n	������i�oа ����쀯퇙_�b�Є	�l79�1َ�'^>�%VT����w�o���o?}���������������~ijc��us��
O���B�p@>cC-�I��$�����}"�G�^]��m��Ho�W��0#㬞��b�q##3�|�>#X`,�K|��ưQ)&���9XT;�bc`td*ӉZ��Nr���vj�%XQ������Ҭ�2P�;�bQ*���s�c��#e�9΂�W�@����������5��nzyutn���[c3��[eɫ���������>�'�e��슢Κ�兕�w�X*Wl�����Tcw��Ɣ�S��,��N�
趬�W��f�A>��/��}^�����J�''� ��U=4�$��ND���0�6�b�)	�  �ꙙz��:��627U�Y�+��Qo(��%&z������ʑ��������S�i��¬������k�>,o���Xoh)����u� [��|$�U8���: �ܯJڧ�ГO��b�{2���d�6�.��j?�Of&U��_G~r��?9�?9��?9������=�G���, t��p�N�d�����"���v��A��v�S`�3sh�$bhlU7R����P3@4hm�(|���*HZ��t1�h8Z0���9։��@��k���=Б6����pq���86��K�H�Ё��i:�"|��<hg8���4EU�P�xV����QK� h������6J���ق�mC����(�~�v*��i%� 4��C+���zj������o����������3���Q�|��9����X��̴���'-�VNd�W.K5�X�qVJO��~��������o�����ϭtu��K,f��S�v���`���+o�����o�?���t���O��s�U
{5�����	%)uʈ*���}���W%P��ͮ�!���< �z��_�O�����_��*Ӡ�WE
I�B�#!�c��*nl��;T�	C`bH�"~��@1�X|"
�@�s..����g���sC�e7����2=b�[�r�@�2�l��(.=�z����W�r����H��J�.A�����8}x��� |�B� �4/������S�O�B0�|�in.�-a��5��S�������~������������~x��㻝��w�ۚy7�)Q�\H;�h+�=�0��+J�
�������EcU���:��(դ �����<g��TOIҢ������7mc�6�H���w�����<8˾{�sړ�[�Y�.	����?ͻw�u���	�m�>#xtV�ړ��'��
#Nr�憟cƑm9o�Prѵ����驕�������ŵ��uT�wumkae}fqetf���@iKe�p���ܛ$�_�LY[j�E������yO����n���ow߽��~�ӻ��WW��L�uy�9�[�r���%������Ϯ��m,���l/,�]Y�܀{ q]��e��uYs^��2����!�����Hp�����S(����Hճ/��N�c��H�3-��Ss�K����K�5>�U�^�~13���دQ��͝�7�e-~GMfzW�=8����*#���S%�#:���z���\���RǺ� ���	g�R�f��5��O�� ��N��>�?8�������z��!U������� h�30��)9� 鎍E�T,����	�,��2�H���he
rw �3�,2(@��<+�<��4�+�64�˸���0��A���|�Iu0$��@�)��u�y�l�'���8yd����Lʀ�I����
�sg�t���� u��e �S�0���I��XkR�g3��4'
�B���T�����H�D5�F���04;@�3��̀��~�Bh��?��~���ńW!	oG~��JsӸn��#�Ey��&�Y3����>a�(�6ѡݟO:XH9�O<c�?.R�*�	�)��dk@���������N�O�Դ����Kn�Y&V���)��i	)�"�RRZ�2Ka�f��fo{m������t����O��FW#����y���`  ��IDAT�Zգ
��JTK ��F�)h ��^꽸4;�0\;^+�3&UkW��cɒ�K����"�X�M
��WL�PŃ�Ɔ �Do�����.2���zN`4-�� 	��j
��C�7B>
�J�m��U���g+��rj��ʖ���&_�E���0�����n�%�z5���ã3�W�;g��m4H����?R}�X�#�V���!C*K��zQ��,�K(v���qb��懯?}���~�; ����v߿������=��5��6���X��p!��Z�5��uch�u ���:ZP��ZJ^7y^�
�!F_��^0r.�8��ⶹ��������K���]a�i�ӣ��#§���������<�,��EsnOw��j�������L���N���L�P��9!�,�"�@����lٖI��,�l'TUda޵�Qz��{߽�NO~�;y���o���k��=�)��+O��=�~RȞ�k�鯼w����Ӝ����?���(��+��~{�Gq������ -@ҿ���6�baf��X�| ��=^��B S9�p����vqijn=���67�k��X���??_��%�f�L�Mxw��}+��U0`4�ڷ�w-�f�}Kc�Ú3����Ǐ�@��A/��ٷ��__��$3nH�[#�Wsc��]�a��oiO����5'�^u�ʳR5������1��;��x{�?<?q��O�~\�[���c�#����gkca�?��^����u�������[o���.Q��H�6��兛��&�yYw����O$΍4\ ��� )��S��	�G�W�Vn�;�C���?���/^z�������{�������W��Ko�|�/g����8�}s�^*bOq��E!�MaG�c�P��<g�}�i I1��	`{�T� ��RX��1��1��)�1���`:�a�DG��" .����<�X�m!h�|�
����氎��Q}M�sq8�g����7̍��w��n����f7H<�@�o�9(�(�r�9�a䑴FmM��U=����7�i�_�p&vAK	MbU���zǦg�j2� L1y�x@�P|�^�{���L�΋�LCFs9h6�o�͂v��$�!���yu�T�=���L>ȗ�]� ��It~�(�Aa�˅�WEoK�8c�k��D�r�l�O����/~��/��?6���Ԅ䔘�l�!/5%/%�8-5נOөs��d�<:"27:�v���*y�����_�0�������/=�mf[�<�R�P�P݌�X{�V��$<\{�N��p�fڕ�$y]���^�����L_�@]\S&�(R���3�JY<�8*cQA+0Ǝ,�B�"D? (M�SBHP�/s!� h���/ M|�r�@oL��0�kY�ʪ,ӓ�[S�����5�gsٷ�^\�~��*	�e�K�C:+l�e�-��.�&���Z�����nY��R �p-��d��	�����Q�M������uFG8PD���E�>��b���Y����z��mmo�%��{bv�~����G�#-#�ѶUi4�e�i4���4�*F�K��q&�+��M��<sҩ�l�Ǚڏ�c���j_p�8�k�i��j�+����J����*���J,|Wj��LѮޮ��WR�?J}��W�"���(��C��C~d�a"���A�n�&��f��Bע�d��� h�ʺ?�%�89X[_�|���#[K>�cYr��W��(>L��67= �zq�����{���9�R�g���������)�k��%͓�}.?) �˕a���o8����57��||<#�m�{��M�NB�?$\����?��v��7o�b�A��cv���v$I����Oq�ߋ~3�I7�N���+kp�+�OW���lm��;\�z���he*r��b2��@��y&އ����V�%��^N��QV29�#)��U�k�_���E|X�nQ��y�2C���?���_�����������~i�_�������ao�v�ߧy �w����>.��r��&�ӂ3}�
�rDF'	��`
�-�R@c05���H5.��98�.B��D}�1��i�+�U� �.
�F}�"�Żj�c��U��Z�,��Ϛwγ���\Y���,\�+�+<��|�i:P�\�)<b�h�2�E��$Vvހc]���)N\�&:cʳ�l:7��	-�mS�3������~ߠ��RD��XǢ���&��L�d`~�;}k�-��R�Ԡ��GG��P�#�ErVɶZ݃c����s��Ic��y�W
���_.�_)�V$y�(�o�^�4���_�U����ů����g����t:�J��[�lA���uGa^���0"���J�����׵�Ni��?�����\k�,�J_���a8[�?\��>T�}�! �l��IT�������T�t�ր���]�<�j9*��$�C��X��{$�߉+ d&��1�	$���򧃬��g�Oxq�,Qp�y'��?s|b]I��Ȑ�Jgm��֧����dg,�@����@o�2���no�no�rK]S���9j'K�'�0����	�Q�9o�h,�a�r�	��Z�RkJ�]���������?���o�]���K�c%*KJ�Bo/��7��B���<5p��N�a]�Ħ�٢U����Λ�w���Ig2�G34'��Ύ~�oqy���m��'L���*~'�`�ҥ�f�V�v�hW�pO�k�f)���x+Uz;M�f���T��Q���H忖�Ǭ�4ٞTՑ����w����pE�@I�ʊwy�X[Y�\�~��� :���Y�:��n�����7k��i?HSɎ7vt�N�z��ܔm��Ü=7.�� ܁�Ŷ�q�Ö��	��^O̼��<9�1�^
L���ն&ݸ�K��BM߀�Ĳ;^�F��eC����O��^"�{)<\�*Qz�8��I�ɥ;��U��B��MM�+�0�^Ӈ��G^H�[��v�OM,��\�%ϲ۷�uG��Y�OO=|r��2�ZW�d:��,Q|S侤���^����}?!�t��T���]�I_U��lRW��0
�#>4��]�ߛ/��S/���߾t������G���҇�������{���Q�)�������P|�q��5���'�(R�"�{���@�r�gP���H��	�͜��+.��v��ˌ�PȠ�9��o����*@)����UCmH�`,���P�� 0J	�\��`���ml�?�t��Ӆ��1��M�ʉ��@S�����'�������5#. �t�0d�]Y�;9[����:�-F�^�7�%������7P�J�p�FbI�l�9�["+;o�/�����ZS���o�;h��^`�i�k�z�=�.��G��[Sâ��=��$�_]$y�X�Qq�,�
�K��I�6�. ���ׇ�&
r�Ó�w�S��-�eK��H��G�.m���}�[�J���?}�|��)��]�jcBN���F��=Vw�6�l]蝂��3��]چ��$� }���VNV$\-7H+�b*��ʎ�S.�(��3���*�XU&n`,�x�i;��K����U�
`:�q�X��T�����5�r��m}�����Սg���͕���e�6��J���j�x�X}R���5�HjV�ll�R��.�?�e�#i���Icl+8=��q�&�!�p�)�S!4ǠNb8�[��AG,�jk��ŕ�յ�oks}scmscee���sGOdf���噵�hgh.h�Ο@[����;!jKJq�1Z
:�Z[\�u��~#����,���������M�ʺ{myhi"њw:E~8Su0Mu8K{0CM��C�՟d(>N�HW�O��KS|��8��;��9��۟.�8�tهi�)3���}��ڃ���R5֒����9��h^0`4�iಟ�R�y��흝-|?,/�D��XN��Ԙs�����ep�����ѩ'����:�&�'g�z�f;'����[[�t��T��t�����i	���{[�G�O�L/���wO�>�d[n��N$�xB�~�xw���������R��'��H�� �P��t�%��y�}�A�z����7B�&��O�j��,U̝;�=��u����N̎O��u�m���*��N�W(�J�)�(9%8�t����;���k?H�|5	�+:���2&�Q��-�Y|G��b���C*r/�����'����K��oN|�ߞ��=�����K��Ϳ;�73�_�@�6��g
G:���~���~S�Q�(�"�� ��h`(�3�H�0H��4�I��7�peވ[�*�w2��h4�<�͝�'��Y������,��h9NR@�G����Ȝ\�qw��v�nV�����\��m�$lL�=x(Alr�*$�l@��1%��C��58dym۷�9������2���-Vo�޳0#�O?����?�x�ti}����OǆX�a�FfI�3ر� ����g��[s����eBVZ(�O�B�f)ʪJ��|29���������Z�7����z�@
\F] y���lq�Jb/dG_����������T7�h�������sr�y�_�a����������,��WD%G�嚘�51��O��_ ��$7I8?�?�U�]��K� ��KB@�'b��ʔ��t]I�Ҧ[���%�s:�5:1�Ӡ.KQ8$�y/G�]uզ$tV]X�աmV�@7�e� G��,�&5��y057�l���ono���&��;���`��#���������k�П��WW�����^�Ĩ�>u1�%��v;�#M�"��חD�� �9�0��44�+�1��h6:ʔ�840@��|g�?t@�v�?[rϡ4+E���µl r��eh�\o��	�h��Ձ�9��::����1��4�Y������Ż��9��W'\��{�-7��@�d��t�5L�d�VbN�9�K
��l���d�)-�:rel�ܒ���*m9�/e҅����BxELg�,�ն�h{��*ʭ���;�3�]�/yg���&�e0xql���j��d5��pB�9Ce+L*����d��W�Pu��U��%μҒ��j�����d���q:�mf�)CX�iJ	-H��r�"���9��l�Mk������\�=2C��{9[{1K}1K{)Ww.[}*[u0]�7��n/y7Q�n���[��,x+��~BxH�<˖|����U��Q9s��2�U3��lO�Ymj��~P��RWS�p�J���Fp�p�U����.|76��������d@g]���fܤ�+Ry���Ez���Q<G��)�|?O��Q��3/����̏^:�/���Ao\�����t~��9����w���Wx����V2��S��<ֺ�Z(�iLF�#��&IҠ�M�����!H�k6�;�	�LG�3��e: }�"�j�bQ_��EA�[�s�D����@�$¢�2�{���� �Æ����wM�-9/�(9@�C������QD�ѹ�V��Ѐ�3���������R:1�-���9C�����������k[�������=9��Sj�3�cfػ�����ٳgϟ?_�9�ͭ�ue�aJux���B�>IV�V]�7?9�U�VV�z����u{sU���6�^+���/������	#�Ү�ܤ~�O?��'���N[y}e��d�SW��_���i���o~�˭��Rk�"�Zd�W��Ŝ�џ���q���p�>EU��`���8
�v���ZñjL#<T�p�*�terPE��<)�2 �+��9t"G����JMi1�=v��ʍ�UE�Eݕ���{E��T�Cw�U\�*�X�W��94!v�7�~�zF:=�D�Z���МV�?8�][�����m?]���S��ql�����ߪ���\k����e����KO�z��I+ 4�@"#1������4��,{�Ȣ1�(FƷHx69���+&��@XPR6�ax`��ǵYWq�`5t��eך�v�ƨ��1�;�k�D���L�î���� htw`qm�3�a��Pz�m��1�����ݡa����2���l�{dj.i�W��F]OkC߽��u�w+;0���~u�mد�i�ᯰ��W7p���m���4�o��8����-��w�O5}w�{5�wU?yR���:8�>9�7778�0��A0�vz��;&�owwU޿[���8�~�a�����5����<l��l��k��h�yR�� ��qc���������0��n�A�P[�p[i��������Xܪ�|\��Y���Im�ê�ʞ֪��5#�F��ݷ���݁���fֽ�0&y�K]��N��''$v�{��KY�����G��w�h��Pu�X�n��sdO��VfU&���=��ުV�SaPƵ7�Κ?Ї���{-I�A���95��Mk��:@;�`�bF��y ���L��T��&��|��Bɏ.��x�_
?�{��73B��
�U�v�|�x@gP�@�݅W�]�g@ł���<H`&b�IBAc"1����_�
��X*�h����\���ae2Pk���d4���/3�����F�����h�)/r� ��F�Qoy251����������@��P�3� ����څ�$� -4Ŗ<l��y�׷`蹼�ǎ�ضZ)k @K-�)��!׬}}m�,E������1�#5�цR����q���S�����wc���5�$C�h`(�#c݋�]�Jb��ib�f �.����j�˕}�Ƈ9��
�o(^Α�V ��1�.5\N�[ �~���7_ݹݖ�cL�M��;�����/�wtvky�_"���>:SU�BWFe�
7�/��� �Ӎ ���emn�4�A�gz*z��u�A��'뒏U�T%|R�<�TE�ղ$IErLU�ʩ�
mii���JS��p{�e*�t��t��Yd�K�Ƕ��j�/��K�e�:���f+'����gAP�dkR�qn�DXc"L��;��|��J�5�YW��n�lz'3����ƪ�7�\�[�O�	,/x�#������"u�	�}�N�EL��)�9�U���>+�AX�4�4��
�
�&�]���i�e�8;����s�v Z�dV�uN��K�e��lX��\��9�R�Lg�#(���Irh�@g��3Hj�`�������@G�?ڮV�1<�2��fU�����Ź ���v�t6wa٣����w�z[��G`7�ښ�<����F��[��[a��^i��4 ;w�?q��h.{��4��4��������^3{��|���Y�ܪe[�,7kMM���
ssYI[#t5�w �@���{����@�����܅�p;U��ͷ+�������t������H۞ە}wk۪��ۛ;nw�(�e���h������Ip���ʾ���[�+4�>rv���9�J�I��J��Δ��M�Hf8S��V:�s�Y�������y��;1�'����������T���1��NG;��bO�RY{񕄈�ǅ��(؝,=_�]M�[��u�0|� �~�
��	���?�"?b0��M���D��sx��_�}+/�B�;E����5��P>�g
�]|�+�4�±Ƚ9���8��$����3f�$����mD��W��d� p1^؊��X#����i@����&�y���\��+6<��E�	� եm���u#lj�Ư��������Ͽ
Jŵ �ֳ���b��X!�p�R0I-#��? d�oeu�蝛Ȫ�%l��-�ƥ��}0]Y[Y[!2��ݝ�X �C�h�3���{yyǻ������O���̷
6��D��3�D-���������Ԃ��)��%O����s��)R���/L�S ?a�_5i"A��տ��/�\�ɚ�\�ZG�:�j���n㝡��_��׿��o��ų�ћ�
YA�0���Z]����S�fw�.!�)S�X�9��.�Pa�w���T.��@e 4 4 ZS�r�h+R�[��{ViY��b�Y��I}�֞ft�i�	���Q}�X}�Hy�Z�x�s��s� ��6�5��x�w,�U�#�h�6�M�Z�*�����@�	�V`��&��)��҆߻���篬��^��"F�j�I��@�MEb-:��4 �s��f�Uçc�*r�Lw��-.���g{�]�7
DeGؔ�%�9����I�=��i�����7��827;8=52���F]#��b1�ُ8�lۙ`��*h,X�����Tr�0�<�o�#r(�6�̩�;�v�ΞM��螝�l�x��Ks�OZ��yie�i���9׫�2+��2��K��T�$�^Opf&�e�;2�˳Ӫ�%�	��/�=I�����58Ӓ�2�K3����YIepl*>�$;֙gό�����x'�[�#�P�o���9�bl)1�4�hG��,�c�J�'���?J�௱%��δ���Xg�ΑS������)�G�6ڙ�/�I�-�n��7P)�I�y)5FCyQlIN��ڞ)��*,)
k������o0����*N�j�I�|ە*��!�U74��=���������'{��[��������n��7�b�*�\ՉS�qC�q���q)g�xSw�����_1D�I��)H�T�R�٢�%�u9bV��-	��'L���!�ذ�tć4�C��+���~H��w	ѭQ�I�{�{La��@C�-��?B�1��Чi��3L�ya���lّ��,�*r�� [.���}���u�.�	8�5�������&nk`�y6�,���1��*D_��'��1���`N
Ǿ�N��ה�OOM��$��t��;Zk���(�BhS��jh��!����6���5?���X�đ�����6�mO�Z����a�>� �WW�|ޮ�i��6¤�٢�Ae�Iw�{0��X__F��~��3��J���C!�F7��0X�R6&����G��Ӛk�OW��S��'}=G�f�|O��rI��,�.K�����_}�tT_�wi������B�_c����7�}��_���_}���g��uzs�4�A'l�?_w�� ��ܜќ����$q�f7�_�[	�r�o��B��ݡ�xTЕ)���+��N}ler�]s���k�y��,hV�� �OY�9;F)OP�c&�Q���Y~Φ�`��`Q���fW_�(�!�i���k���q��8������o� �Q��y�|l���泧OI�z�����f�Ô�"^����X�7��ICG�(g�ԑd�,�3�7���nnx��f�K}Kc��B]i �Q>p�-U$��\zor�o�;0��9>^r�)��Zr�a������M��D��8:��!��F^��3�+���C*.Qq!�b�R��(�z�#��������4%ڒ�%��R��S��+K��F��˭�2�N�ôb2[�ܮ[R�v�v�ҡV95�ʷ�8S:� �q��ۃ7�c�T������pk4t�p8l�6-��V�V8��v|��@W!��d��=�b�VlU�>�7���c6ߢ#��b�A�M˷Ëy��Ϩx��h� ��"�Q�ҊPF	������D�\e��4��:�1��$E��"{��?��+(Ilc�[�S����;����o����{��ׯ���qlo7eXn�Y�K�KxR�Wǟޯ>�f\�z�+	�7�'���z��՞T�� \Q�Up�;i
:N�0}l����"�o�H?����(��o���3�8��^b �?4�P|m���a*�v��8�D���O2l�s��tԮEp�*"51H�ǎq��\�yKU�\��Ͷ��1 �`C�X>�	YO48�Mޏ��������~h����0�LGa��U�g�LF]O����Ǐ���z|��;�%��r�V��+Sb6�[�������E��\�b���Ȓ���M�����2K��J
�{]� �ǖ抛ʄƄPJ�`FE�9�7M�]�Ix�����ٳ��-׺��`��n�����YEv�¦�m����q=�@`>��xv6����L�۹�r%od���T�v���;�鯾�|iɝ�[Tcs<x������z�z���{�������~��/���ig*T�juS����	g�С����ܮi�1::���Q7$_�I>U��#�J⎗&\.O������-�qM�Wi�YZq�Q�fէ��f�	��8�=e�@�d5`��a��Iz����h�ZT,�KV�U�
 ��V�-�fQ��Om���?ܪ���UV��g�o������������ڄѐ����qWgL��Cu�sd@Acxqhp�aV1qV��"kB�M�����4�9o`ܵ�p��z�YHcT.`�<-`U
�1r6���tkx��`��N��(YT��c�[��]�㎖������4h���r�.�� �h��L%(Qcz:)���	�v�"	���\"���� �T듖��I��)�����8k�ʦ��r�J�Tk�ce�G��_H�=��d��D�	�N�L��K$B�l�U��E�����In�:��
-b���$)Y���.����m"�S��I��+:v���m�6�G���`R/鴰����Y ��R�5�*���
�"�Xg�#��B��㒠"�MS��.I=�!ٝ,|+I�V�`WB��Ԩ����֢��u	����������]�o��ۗ��͟�����_�}�{�3뷌�ƌ��Į���<ޡث{���H࿮��ٲ���[�)�Ы�� ��x%`�s�Ѣ�
�~b�ǉh*���M���|� �E�.o�#&�@�>2G�}l��8h�U��q:�3�:�t�0���7���#�C@#�Hj��]�Fo�5
��ia�� �Q���@j2	_�9
�䃚�\��Q_��(�8\ ���:UXڲP����J�k*259��]����jC�S�]���FC#���:6��j�[�G].�
k�S<�tLOfTb�����������i��
 ڳ�2�4���0��P	��Dk��¬�R���U��[��ۛ�9��.���C
O+6?�Zn�@�O�w�Нs���7�į_�w�J������>hp�����ŝ�{Y�Y7�˷\�;�py�f����������w?��s���Z�[��7h�j�N�&��џ���OU��wϏ ���'G��kU�I��NV'p���T��=^�x�"CX�[��ڜoh�Ī�1�Ӭ��:N��P�Cf�aJuȬ>BkO�1��`�SV�J�>l��ϳ��%�h0�a5Wm���r���7RmI��ҒkK�O���g���]�	�8���(�1r����O�fI��<� �",D5��v�N����BX!�Ū�M#=c���
���'��x�g�ʟ�P0	����E� L�2����̻a�f�g�۵ΜHc,���Q�sVI��Gs�lsy����<��Ł��$�D�cLHY��g��1�q� �AM��ѩ@È��� +�{��K�U�j�JZ��N�WBd�$�� �X|�hs���,�'���H�*�MP��F�E�,�����Xx�L`�E`�qD���[�K�����/�&�\�����:����%x-R��U 4�FI=I���	�ޔ̠��E8�sŨ),�cb�3.8�	z0���C�V�M}3��~��G�!�}#o�N��{TA�������]��?�y�O�O�~�?������~s�6�ܔ;]��Րbd���!�&F�m�z=��7QB%�4]o��85"�lָ �jE���0��3�>�"8/�>���C�F�+�Ѩȏh�>:r?��G�Tt��Q��r�*:��>j
9i9C }ъe�A���j���$c��	X���{c�&'0��2̓��%�6oF"S�zƀ<B^x3.P����5<�a���|�`�',#�b͆0��g��2iU��f�f�>޳<�����Ӥ��i�j�#V���S^/NqV��.WC�#�9I� ıp���l�@���A>�L�g6���:�?m8�dbcج��	��߿|~�v��0���v�X�%��0����i	���~O`yqe�{a1�������7�Kv�)�ug-��rĒ����_}e�7'�$��?x�a���tc�����~��O��_���?~�=W^�n�Q��+#�����/4&��MnH�5;fH�ѩ鱱����*Mc����c���U�b�ǥ���OU�Ue�*����s���3&�I���D�e�
ş�������(�;:F�NZ�OZ��Y�QZ"�y�R�a����1����e�p|�E4s��
	��a�-.ܒ(�d��ޙ�\� �9ͅ��o�Мk��~���w(���f]�q:�M�f�Lt@3����Α��Pڵ0;��͹p�ֱ���Q��:%�$��<V��H�*��(��p&�d
���z��A�Z�(=FnNɻ[�hn�T�5�5���U�)��|A���s��!	����!�d'��W�/�&@K,Iŭu=s3����;�0iiq�ht/��c� h 1�eV�&�� �8�
[n�H�_C,W��Ş�"n��4V�E��z%+��dM�H�F����DL���W��V\K	^��\�\��
wZ�6��;h6)<�$��1��;G�`���V�}��,v��e����fB�\�]}ĵ$�����>kc��>��+���}�//��������w����������#o�+��囅�ui�kE��h���q�7�v�'�.�ia���Jp� �8�� ���m��B�G��}���пLp�����
�3�� �f��cj�}E����Χ��W�( 4'��2X��� ��f &a4���/�>W�g-@g,�ƅB���:K,:Jz\��<�f�p�*3K�S���is8��T�9į�
�!|��Z����2%�F)x�8��j[tͻq�|iey�3�|X���c%X`�U%��cmi���>ts��3{g��Bs:�,0�R)l�Tga�� �wye·�^o�d�a4�)�"�������a�j��|��k��Y��������UOm�M�=�<�����@��O�z|����ڷ��l��(]�V�D40zO��-�jjT�9����=�|���������l��7����⼻�ֽ���/>������_�ܸCӕ��Z��F�Zù���) huS���g�QA��*�/Wc���őp�*-��zTE��>O]�~�V����݃F����=IW_��~���}Mr�}C�ǹ��P���1F��6+�:��3ʣ���8kQ]�j.ٴ�c�hFem�^`TAV�5���Ul��&
,�S�������?��~��쨱����<�:����W-r074��Eɳj$V}z��}ql��^X,������|��(O���Vm8CmȑNX��[t-TEGc��ZCe��Ra���C��:����ca���z��gl�S�]�1c9���5c���O�X���'�k�P%�k$�����Z�&d7;��f�� ` ilf�V��XɊ�D��%��b��y�g�P"�av�F� �@�J���}0 h����T07g {��>��a�G�o�x,Sdǋœ�h�<�:83�9��X1���.�"�u a��\�Ԯ��5�#83 ��8� �U.�,Ѐ��H	�6tN5�X'���N�hO��C� 8)��){�f�W=��	W���?��Gߍ��;����?�gw���׾����~�'e���9OR�)�'�oņ�J�g�/���ij�:��_��<�� lA~r뽞�Ï��?1�}d
Fh� �|���7��7#��7�៌!���@�C�!`��'���`'(\�s�8-p��iLξ�˩��g�3t@�+z��΂F��
&8� ��WG�I�~8�e.��4	��N�Q�
4hU��~Π��W@_�ė�⫌<����*:,̃nX��3���΅��&3�sX�����6����G�V�	���p�ʒ�c465&��J�E�`�홟���9@�)��1�f�Ѳ0Z�eR �K+�1������?9���@�=۞^Y4�r���a h�%6���3;���}���Ə2Իr�o�*ߺ./��K���*��Ϸ{ڻ3s�me_l>]x=s����������'=C��[����g?�쳍���L�"�V�h�<W�
��ؔz�!]�X�>=���kkU��WjGk�q��:�`&���L�V�.�H��dF�ş�d�����>J�n���_��������������o��?_}�����Es�Q�� �O����'i�9���G�/Yq��K,�>.�hW8:ۣ����ƄXa����s�9��� :��<�k�+֋�|�B�"#�^FF\_��Cx��j�ld��6���{8���ӓ�7�uEIJ�^i�S����L|\�F�R>�21�Ɩ����%r�:��c�<R��K����Y+*���X�wN?L`�"\�KU���=N3B�n�Y�I[�"�,�E.ca��[~^��b�g�,���̈{ѵ�2dpn4��@�h�X��XΔxu9�C_���t���HGV:��
s�E1kr,�*��Hc`(�ef��£!WYX�ʚxo ��sA�r��+T�hn���p �8j�&�8G*:7	pa���o֚#��A �!d��Q���K�3�W�cX��R��[��*��p��x�{ɒ�S�{�#/"�곧[
9P�m�".������+��^	�p_���_?�η�ʳ����6�5_�]����+?�v\��d��)��5׊c�j�dV�:�-YA�����V1+ի��Y�M��M!������h�'��#3��6G|`y��
����`@3Hf��'in�>1��_�W�%0��&�F_����= R/�b8�:���������m�D�u�N����E��ˤ�)'��t4"_>lCrBg!*hF
zG�Ƅ������I��a��49�Qk�h1�A�<�>�� �]���ha���!�r��8�R7ޞ�5;��� �[J"L� Zy��^�%�&E�5�oiҵ�Zz��2-LL^U[>:7�[Y]�~��|�oi,�<W�j�{�[�r�)h,,�gѝ�Ҽ�z���w������S;�.Ņ��t<��7�o�dޮm��O���ٱ���}�t���g�+[�s���ӟ=�^��a�PeT��M)gj@D'�/צ(�w�%-��&\�C�����5�#��Õ�@烕IG�S�U�\+O�,K�T��ԧ��c&ɑb���.��?�[/��?~�/������/��z�������d���J}�� �q�Pu���/�:�Ӓӌ�<� @_uh/ZU��J��^F_����/^b����p&Ia5ݙ���>Pumm�M/Mѵ�X���RPd��R.���,�"Fx�X�-��fY�kƳ������瘰����_r�7������eU䤔���cر�ɬ�E'3��8�-GaUQ��PE��fT<sJ�h74���������w0ݞ fp��H�d�QK٘{|��`p�$8���U%�J����~ 4K�
�M8P�r�%&Β^�~{iu�$�����h�7���� ��`�X ��-�	:c
Au��A� ._�Z���T0�Ii /�)�'�H�`N�qG���s��3tpE2Ɯ�:L���B�@sX�T6��7�\n���D8
=���� ��6�%���U�V��� ���0�`��W8��4��p(E�~�dO�doB���klIr�mӳ���Qu�;'Ͼz����O�v���$�o�o?}�\�]�Ә�P��ͥw��M����PF��Ԥ@���+�;���B���@���6�|���-A�й0Ќʺ���EW]>\|�8ƭ�
��-|(4V��ha���t�
�@�'3��a��J���94�q��ΙB���T8�d�i3�RN1��N�1*��)��4;��:o���7\3Y0JD|�^$t��ȯY�!��0FWY�prsM=~`4����1�t���JLk�j-�SX-� z��m��H-7	L�%�-RP�zKV��(4�u�޴E�4�(,�y�U��5)�C.�H��=�5_טS���ǃ��@`umcmkӵ�i鿟�LS��jZ�_O��p�^�_^�\�d�h�(]�+G�v���lŞ<�Uk�X^ݽ��ϞV�Ueu�=��m�,���,��o?�����d{���� ��ӭ��V�R�Y#�jL:�|>_�t�6YQ���&�k	 =�V�.���փ|��"~_y����ӕ�W* �IQ@ ��Yr�Hx�:�;'_{�o��K�g����ٞ��7��������?^9P������r��ôt�Y��8�)�-9kQ\�k � ���h�H�<K+�.XPe�\�Eu��D0��������2N��������6uf5hR���� }Ů"I��`�6�#�$��GImɍ�Ϟ=���O?}�����6���tݷ��MN&&����í�w,�邦��Ҵ�FcyGm���֑���C�u�����Q	h��҈Mi�3#��)s	�`hh~c}~u�T�+���]�Ȫ��Wߛy������F`���j�5��q�����8G\�5.�<%�,9ޑ`�Q��|0�ĵ�|�ts{~㱅ќ�,9�?A������(~i\�Z�������B�,V���@�؅���MRv����A�	�;� 3@̿ye��7������=��`��ۇ+����_��i��Ĉ�C:��;G�s�(��b#�q �%@g�Mzނro�>���]��!K�KU������(E�'Q�� �XsU�Ȼs�����T����O5�e���.��O�7��*25v��7�m���w�S�-ڣ�#{uA��]���KqQl��� #����> |-d 	r*�GQ�>f
F0��+
��(H��4���>d4����1�>�rM�}�6�Y`4���'�U-\�8�#�ӥ0j��)y�Fc'�ERS;E� ���� ��Î#��A�� а=l�ۆ�9��dd g����"c�E��->OI ���*����3z��\Sn���� �I�S���UT\�������n���RS_�����4Γ��cٴ'S��� ����i�#M�`F]�%JjTe��ƽ���u�+'�T��5�鄪���.�2�_X�\�̛j�x&9�J��([�%�&+����yWJC���UodJwe��Q�+	���[�n7�7�e��>���?@/M����� �?��'O�?@�,o|��O�m��a���5��F�������Р�w ����{�����Z���`U���������/�'��"��/Y')�q���Qz&-�o>��K�����������}�/���K�|�o.ڗ��Ĥ9ʪ��
��G�A�x�I��H �>�H��T��:��@a���C��<���+�T��6���Y3̷��=>��:t��f�(�*���{I�NHI�(�5V��61�5,�h�ښ}n��&���O��� ͛�X��������l<ǥR֟m.?[�n��g�sknϦ߻X~���շ��N�O<i�j(jȋ��2�ͣˮi�LiMi��$ z60�41iŢ�b̓Ʊ5�����뛟mn}�t����6|K�S]=��c������1���g��O��2\n����Ϟ����؟��7�6�͊(FN*+%	.q �7��3����J!��.�4gHX��
�c9��b� %�+ɒ��YRS8 �E����A4��"jAӘ��(pNΩ�����B�΄,8�L��@P���a��������,#>A�x�M� ��	E6��,VW�q9K�/Y�^�xwB�ޘ�Ê��w���[?�~�kw�\]OGo1��[o�o�?�h���o}�x��"���WrjOL�;	�w��ʫ��*g��, �|tp=�0b�e�d�g�FS�L�@M��4�?��"N0��?yK�l����1��Yx�	���paV����I,b~��U�α{ $ ��|SkU0��`�%�r�á�1s��Ac8�ہ���x��9��i���F-��	v$�s��,#9O�XlA6EZ��{-�&g�����E׸k��T_nea�%)�,�sb�3���}�_��{�A`��`�dZ�L���(Z�6%r��-�oL�s-&�5
g���*:��p�7�X�n�>�ј�`H
o�i��z��3���<�o�l~�<8=�[Y��nx���W��-��V����_K��%~=St�{1QPv���Yr���cO{�[8n���3���/>'��lxhܽ����b��=�t�
 Y�p�)�	k/�$�jsvVTYZ����R֧\�3��=X���
,�@��d� R��+�I��'X�yZy13�o�}륿���w���������؏��O~�Ү�~'��c�!F���E}��B!�?1���g���6�E���Q,��YZv��6q�U��[F�p��׳���W�c��6��lE��N�)5	�(`�
��FGk��,�L�m�7�7�d~�f������VV7�}��o�nn�h�A���6Vq[��\Ս͵-,沼����ͬL��߿4���6�Y70�8��:��.ψ2�x�&����kv~cce���3��@'�[��g�7�>��|�����^��(���>���po�1hz�s��t�KLJ����R$ς�^ y��p��-��'L���,ʾ��a� J�������©�O��BV� 4��E��Θ�F��8$Gè t�C���豅�'NT���;����� dQ�(F���	8=7o��Y1�7 �)3�$����b��\@� �7Tf�JrO�)>2H���-;wJu�-�~t׹8pg{��Og;~6���D���MwG�L{e{���<16;�#ቷ�߉ �?��Sņ��<�3:Ҋ.�y��p|���Ci9�Q
�0�,��]�D�q�&�� �# QI�:�c�B$���a(��N�U�k�Y0�Λ�Y��"�@>8��r�F_<I��o�������a�M��sv����?a
@*D;X��0dq���E��0 7)�zP�'Mh�<��O��'<���K�2Kd�Uݝmc�]�3cK��\��3������h�\��]Y_�zg=��%�ѡ�҂pSt�
�Ðׯ
e%J��Ӻ��|k\����+��a��j�_4K�ZattZi��w�;��z��(h1-d4Rc<(���	��/������������?�����Uee��̒��)z�dw��X��R��\g���.�8����:� �����@���_����s!��6����W����5������g�������zЋ�c��5�K���k� �� Ї*NU%@�CJbN�R`�qV}��5�t���ÿ�����Ͼ�g�v��7���+�f߫{��&�!F}�Q�|>nUe��Z�>`�IN��3+?򁒢�����fa<�N�ˬ��&:����Kk@g�x~?�I��?�ֳ�E�d����lP����
���W�Ԛ`6!������D`ӵ��M�����FR���WW|~�[�`Խ��_��`��x�n���r��Y�ѻ<��x�n���;�����9���Vs����7�k��MR��l�jwyg��<�k��5�`����W1(c?X=e0�Z���	`�b�2�Ƣ.i��n0E���:�Om#j�2���F�	��p�`)Lʽ�p��9J`�.Ò: c9/$hۋfDvD)0	��Ψa�;w!�2M̿D���AV� :�;0���b�!�a�76��5ܬc;j/vW�W�:�4����������}Gd��-:��2�DZ
���Sx��o�i�����{·�A{��j.�d���C5KC���w#�|C��MCJ��(r�%��΢c��v��v�	?4�#��Jk�Ζ�u�(�ip��.��K0��Ϩb�IE���'5e��mm%	���f1|.P�G(�q*
���9VtF3�Y2J��
�"V�-M����p���/Y$8A��ч����������@��5_qHៗl�4E!�ё��#�Y�'L�ǊC�5�&���9�c�(GMXH�&�UC�_/�s�����u�u�,�g���H�B�	�
SNS5s��v�r`cÿ��]�6V@�@��������v�W̨��c1����y��9�����hn�]�Rn��/�ҋ�,Ĭ�^e�]^\�Z[y�5�_�(3J-�HZ%0ieEz뭺��9xl�����O?}���}��� t@c�;����gj���Ѳ�����rU�L���H��i�C�#����>��e���H�/�m��_�0__������@%�m�Z��5��z�5L�N<Ә"�R]��6��hznvb�5��.��'_�M ���gj�ϕ��ae1Ѕg���iZ%,��9��}�/������+���o����eЁ��F�Atn�A>�(�R 4(h`4����@���8n�oɪ�l�L�0֐q��˽����Y�`!:=^�~��}`(�����ӵ��Ş��hVç$ m.c��Eb�WW��u,,M�` �(� Ñ����3��4<����4��8��48?�7338;�16������;}}O&&����ffM����z�}rzhq�Y_�=5?����h��3.��S�nON,�'�^h�s`n7���vM��&�ǖf��&�:&F<~<1�;=�?;�3=10?w�33yo���S-4��(E0W�xj 4� �1<����?����"�W�2��o2 �;���<`�AM���%�dr����K\��hrf��'D�!P����P�R�9�)0��oQ�fk/������ݮ���P�#2�DX��`a@�G��J�+c�ؕ�9�;�������zSK�� �P���x��Q{tA{D�DWg�-�뛩�VG۽���n߶�T\ϥcI�{��?�^���7^z�z��n�Yrs��4|�����+��B�L0?,�r�ͬ/x�z�۞���nW��:����$-;͊1X�A����W�:���a��P�{s�A�o��bg��0
�X�~����M§"���2tn�׋'� ����h#:p�,��A�����L �O��� e�3�gҝ3C�u�*���4��}��w�]��4�'"��3�˔&��SRJپ�9�*E��3�6�4H�i����db	f��>{�e�j�aP��������n�y��k��2-�C�b%���Mb�6V*��PX�,Z��2��ɵ��F�����a[[O�n�don/��u/���*>LW��#{;W��u�٢Ej���陱��n��u���_��g?�pø�_���~��_�䧟}����k�F�˫sΆ��j��A{�*�Xm±���u���ɲ��G��X���8)�T�lH�T��B�����'�>Z�p�L\Y{�E��	Vu��]��𝆏d��s���v��z���ta�_��?T�9X�9JiOZ��l��V�1�A}���� �@瓔���iF�9�/��+v,�b�S9�Z&���������7237<�8�"%�Ȃ�k�0��_�����,���\��T�,� VBŪ���wn��M,�A��\�=����λ���7�;��+yt���������}��[���j�=_X�ϋ�%E[2�K�7�'�S2:Sa��:�ą�M-M�3��%����Q���I��X!���F@�dߪ��;6�dr�������C�7�;�W�ߵ�֧W�t�T�)���d%�v��V�\�6f[jJ���k,�X�#���f��H������5����cW���Nny|��(r�OD�_���ܔE� b�rrNa0ˁj����:LK!Ap�9ԁ3����e+�.����U�>��0�L�E|݊Nj���!Tt����U��v`{m20g�e	3J����?�UB0����F���6���R6��[��h��綸�L����t(E�n���[�ӻ"��U���1�y��$�i���G��μ���7^�^�a��DZ��i��f����(�5Z`S�r e�]dQ�����c+K�	�Ӎ姛0�[\��M>�Y���sTt';�I8��bN;�0_nK�9�xlyq~�3曽9zO�ƀ��� ��� h�t!v�U��
��y~.3߂�'� �\sU�@����.�\D�9�9��O���`�G�(�44Ftpw��'� |�ASQg(hx��Zg	�aZ�E����jzhiѷ����u���m �;�
������0:�_�cnGO�آ����v ��>��ʮ��khm,BaV�� �7q�9��FK��%Ql���!��5�r��}b�L�b���M�4���K˫=�K)��e`�Ʈ<��ʷr%{�`�m�h��<i(���V4T4��W�F�����/����Ͽ���������y���B�����[X�5V��b��u�������'�uI��'\4烮�@_�K<T�?\�x�!�`m�@���E���]̨O��Kl4ߡ��'ޟ�Gy�u�յ��\�
ڪ9eӂ�@������Gh1�Q
����u� �sV����� �Y�Ȫ�}2��7�� �A��Ͷvvִ=윞���@{�א�뛁u_�����!�~t�
��*��G%��S�K-��=s$rF^��ܮ����w4���~A�����"#���#�t<�6�VG��#�z�11�d3Ƅ����at"ߔ�s����@����;8������0Z���
�d�k7��HtPq�u]Z�(+L���bE�X	�&��El,�-0�yEq`��z~Q|.\Lcj"��h�"��k8��E�L�h[b6	�p���l""~�;Lf��A��<\nU3!;Jit@Ù�Y>�\R�b����I(� GX<���w|�z�)�Y*�� E�HCͱM�������y_`xi�x�aƔ68|
n
�� bq�E�$0��X�;�U�s�\�W�u��э�zgTn��d��x	��mMЫ�ӯ�����!����G>�4�V\�(>��D��Ɋ���):	��T�&���c˒D.��T`Z���u���=7���f�ۥ�5������َ����&1��F�!�\���AX�E��@=��-z�6�+��9?l(�~�=��T%Q"DfrEKp������;����,�#�9RsNR�c�)�	�sǻm����@/�Q83��C@�#OS`1��y�)���Q��A\�M\`�M�8��Ճqm︔���gkN�b}���&���!�77ml��6�� и�4.�!�t���Rk�����qql���jM ��� ���)�����p�OkM������]����K/�;'��|^��0��ŕe trC�Y��s�@�]������ʓ�ؠ�hs���f�6Z�lOן�����n}S��_c?�ɏ��_����@O�M����V���Ξ���xm}��j���Cu�C5q�k�9@�� �v͍.VT���4&oH:R�t��p��p�"�du��J :�	߬�<�U"��E{�V�2��1�Ӭ��<ƨ����,Y��
Jj 4�h���Cf�aJt��r�>K�p�B����`\\]�����C^�kmÿ��w��^�4ؕ���˞<�Y���2�a���z��<���L�ȣX�|�Ͱ�e�Q�>�lP����]_�ι�sK��s�-�h�01�L4��-��h����#W?K�Ѫ`
���Y�U�
�I7=��hz�Xfo�\v�� �����F�0�Q���.Ҥᛵ�ZHi.� �;>����0���b� �ii8��dEZ7��?1�>��*ſFc� ���w�.@�SМ��;|$�`�M��W"�^!���.� �f�, ���ux�(H,3w8 �N���A�0G�1wVt���^����&��Ԇ�g3G3O��*�+#K����kf�Qz��=���.R ��q8�ޙ��������f��2�M�����`��5t��7����2b%H��
vkBw���!=����.�w��jC��E�K�}��ܗ ?�����PΤUZ2�hS�#�>WlU�w64~4���l签��Q�wx�;�sƗ�����?��f���F�ZJ���-x�,W���ЪK�*�Zqo�,o���ku�oq:��	7)�������wu�W���R���_#E[%��mF����@!�%ҢS�(�-�~�8�1��9���f���dG�#�-r�g8��`'i 4��`��@�֚f��"����?x0��}29�ȍdb��h\)ԡ	�+�4�� �qtz�� �[_����5��Ӳ+�~�(Ktv�i.������^��Hw�5Wrj�8�E�g�2�`�[;47�����tXS	�. �T_��u����b�[��{
T�uaL�,#���˔S��ѽ��(���/�n�����>����կ~��~������<(h�g��9;�:ZX��|�Rt>Z�?Yw�.Y]��:܎�^X�w�TɛR/�'�AA�I @(��0\�H�,���}���D����$�ׂ7@,C_�����	����똢r�Qed@�O�@g	�g`4 �3�s ��s��i%�է5�v�VpY`�8"�����z{tq�ڔ���?z�5�8��zZ��W�Vqe,Ϡ�1[�` �;��E�Y5��X���ė�l�����K�ӳ��]ݩ��S/aU|�����%�`D���Q��h.�}<���MfN,��8�����WV&��7z��\0�x��2��ʸ�K�ȾY�{'c�+�F�p���%��u�%H�
P�\�&���A�bf
�PG�
��:�x�v��M�:��Ѩ�9�ΌL�
��b�}(�m�KV�dCM
s�|av���	��pcpf8?���r:_$�n8�%*��Ǝ58.�(�5*G���ɽ��{���Qa4tH�zt��b�(��w~��I[ �F'x�W&�I��	����[]����շ�ͨ��]7�M֜0�Ɖ?���@q@/>l�I�O�MT�W�N�ɘ��j��f����񠶠���%(�HF�H�����LjIGk�����~ۍ憞�澾֡�ǓSC��I�f��>�gK�� ?�����<E�"��'���nb�4r�����yFu0���J�UF��9-dհ�*�
@.��*���(������%��� ;#�����L|�AC���5��."�^~D<֕�n3S�Rr����IZ3Fj�ֆ-v���M�=�cz�D 4p����VVp�h��k�},���h�S?>5�)~5kt�9�sj�����s+��*�(�좥 ��F�����^]o�P��6�b�X�oQøDͦ�?�7�v7�6���s������>Ή�U�{3_�f�rO�D�&!4]]q����./9��^���Y��|k�53�����۳͍_������~�����~63�07�����x\�O�qI5��j��Jݑj\��hM, �Rm��&���$t-��.��6$��7�7�5 �?�����L�P����W �+��3f�q��EuƮF���iA)��[�'l��V�i{4�>_w����D�(	��g�����v윣%W0C'��x�{<��ZY�.Y��'�fn=�c�⵴F�j�lB�����cp�5��T%έ�Y[�oM�~�F^�@u�W�-�g���qZ#�Fͭщ�Y7H!2�Onv�[�4��` +��?��X�t�Ǖ�r
=Ԣ	���m��X1k��^��[,2Z�ge�`;�᜞%�N(�uǐd��`�I���"�9"����E�983I��H;��f� 2z��̭\��J�!�)�����8��7_ �ڄ�Eݺ3���_� ��=���\H��d����Ŝ��d&Q}X���;��h&�	̲jAD�M)��ì)�KL*���
��B���G�`$a�D�9�Z9��1!����,f}�ܦ/n��?i������֞��ݏw�3J=[�6f�M�E�)�	��eq��Εf�m���JsK����~���_�%�*�-�����rZ(%}����ݞ�I����Q��(-N��W19ɥ����{nyy&�T���oVC��vy�vu�E-f������%���	�b1 �%۽�H��|\M m>�¢���n�K�c-���̴��5V�j��_f�X)�b�T�!���(al����r	L ��A5�mI\9�G8��yzg
4��+ ��iCx�)�ׂ��O��:
t⽑�9���#[Y��s�a]� |������g��9����b�}q��D�-&і�;7�'Ѐk�ˮ▒p#*��tT-���K��-����1j�h�/5�`W���p ߕ�����y���٩%?�h�l#��.,�t.��k��ž��z#W�F���\,��V�x�2�/�K���)�,(Υ�v|��_}�;�� �?��Zx��������W?�����V���～e ��شkia�5Qv�άIP�E�.W��U������k��;������s�UH�gk��%pq����>��;Y�x	tY��D�DG�1�O�a��U�9:R+�YǭhΎ�XS�l���'&�g�G(9 �-9�J ����A�iF~��_��|&1�ve�kq~y�X�x�n�ovq�k���q=�V%��6i�E�gs*���1c⺐� �w�7��js(PXp~<С(�l�p�&̪�9b���jgm�@׼{qc{���ʧ��Ց��L�f?9���c� e�<��p�#k�cu&�yrh��p��gn>�2q�C P�Յ��p;F���cZA��&%�7_���� n.~�2��#5G7xg���`:�OHC��J�S �h�`
a+�o��8���F��y�%.Z�Zh;�wWm��z9PzSa�YL�4;�#�͑��S�od���pÁ��P����x���!�^���<:&���pj`�3�2�j(M�d䠈#�aIl����ݒ'%�-&�%6�,��؝ww�������'�qN�����b�7S���� ��K+�ѹ�{�7�o���y��I͓�lK��fӝ��G�#O&�:V?�S���Z[��̶�eTgW[GM,O��o�t%ZU�j�S5���n�=��1I|�.ܬ�R��t�< @�^[��.I	�&��w�5�X�Ub[|z=չ06��bx;��\_�/--R����h 4g0P���Ċ��G��L���,�=�j���F��˪͗0Z�
�-�ќ+�	\:�Q�˗�Q�l ������bD���#09����Qz[P�C8GcaR��&h9Bx�q�~��Pn�!Z��8�)�$�v�M��8��,�~�?0��<���np��p���{��': �2 4�h�{mO��gV�l[�ȚaS_�Dp	 4�\g�.���c���:��������9-E�^�FnN��;�Z� ���-�2X~��hh�����y��r� ��s�{rħ�1�y1�tC\\|��b]��A�/�;�����/��)�W�K�����?�����oA���_?}�9 ���dhtn~�Q_svE��.>�Fw�\}�.�H]��Z=�V5� ���\���Tڐp�x���Tǁ�>X
�be��B/���lW}u�9��|�Q��8#?aU���NX��-
 �!V�Fa����9
�����S,�l�%�DΨ�1���Q�y-5f�ǽ,��	 ����&�ʛ��6êH��3�t�4éMf����^�p�f=�%/�}5垹?|?�'bv����׍�5Vp1\:VL�#��2&����߻
��g`i(�4�O�t�@��9��~�mG;�fA���A�D�y���Ş�I��:�,��зC�"�)�I�
�?�E<-���
���RvX�����X?��k��\����b"�,��	 V���t�e�lr�,�̭D;`p8:L��� ��y�ŷ�7���و�Ny�
��'�"8�} �G�n�s�B�2�0ϩ�ɹ2���t�u��p�hN���p�aպҼ{����+@���Bi[%@D+hC�%�a�����ly�;�374�<�˟��}���������ޖ��YqL|4�T��2���mmo<������%��}�������O�׷?����688��-��L�gg���u޶�U��F;qq�ڞ�3+���ہ�ˏ&;�}��=t$����O���S�s�&E�s"Ɛ����a��__���߶E�AF_�@f1�g�%���m�����a@m��럟+h,��t���������1߿���m�{77��k��e�_~���
���k�ն�PF	��8�1k��]vŪ�2�߽@qE���1�}܌)?�Y0�Ø�B"��8�A�2�;���6ΘCO��O�aX4�"���ň`#�$�o7��?d��%�'�\�Pe�b*%�����u<X��ƖO<#��ft͎���\�t*�>��c��胆oC@i2�M�%��ⲯ}jDgN�x�x,<>�?�'%�UEQ�������E(<�H`�h���V�콮y#W�z��\�[��7�e��ʕ�7j.ӆ�I�0�0&�`ʷ���z�'~��F��7���g_~���t}e���D�1�g-�����_����-��_���LMΏOܿ����{p���*9�*:�>�X�z_�����qjb���3\�O�0;.�p~f�o���W&k4���8tM,��C�	G�.T��Y%��p�oi
�����Y�=��NZ �2������b6�� ��F����Yx����X��Y���|F��(��FG'4������E�Ԓgv�=;�0:5���)��)�)m"c��*�JŅq�#:ϑ���A����[Zz0֝U�+f����o�=6Y�Ƙ;kBC��#��Q	2��vh���T�Pw}����1� %���%�7��_�gxpN�U��x�ur�o~�q�ZZ-f�,��q��Dq���4��V�Wޞԥ������YxgA/C�@&�1	7C�)�3� Y* h"W�Pؒ\x�8"���W 19C�^��^��h����6a�]l�ou=	��z����Lb"�k83�4k�T �$>W	�*/��Qm�/Pumk��;}Tl�ũQ��p{�oqusu{{ek÷����u#WV=k+[[[�n/o��|c�m�]=�i�&�ܞ��58�ȞnϺ�w�;[�߾�����3������k��a�h�'���q�H`�n�7T?��nnm=�|���Q�Try6߬���)��5���g@��u��%ʤ��!�hbn��^��.^^ߘ��mU"Jl_�`$
cdBF��D?��=�¶��8C�9��v��d���* hh��%$���ί�����&�~���)�������m<ߚ^���-�c���_��0�sP`����1'����E'�|��fp���ĊC�ðw7�^2��7���� ИJn��>nFF�%夡A�ѡRh�Ǖ�蝟[t�38���53��׮s�k�2�y1Y�ԕ�B�E�P��hv|�����=�!����5���� 諔(�֤��] �'��ۣ]Rc<��mA�$Ο&N81*	��|xk`ffr�=��vy�܍c��R�l��E�7��I�-`zO��(L%\�Fȥ*uLa>[Uqs�w�'����G�;�ҿ�闟=}�������tm�k?��/���~�����W_�����~�ydx�n���-��o6��[��Uq�Z��*��U�*�T�>����&�`]����s��⺜�dMB��L�TgY��)�bc� �	 �&}�J�B�+�9ո��zK�?��"N��O��02�,<��
�(�9��'�H�#f�a��;AK�r�Et>er>�KV�eV�$�ߩ�l���q�-M��������,vUY���T\Q&����TI��D�9�3�2+o7?�^�Y왞�;�[t�"1�y,(h�G�N=�%�K�EFD+CL1"KZR=����+�ee8IEc� g�4)LD�X��l��$��[Y�vs�;�9ٗbI��D;��O\���Q�;��QA%�\`��PFn��h�o�*���Jd�Ur�
I�&��GР�ÉC�$*�d�����*yDq�x�J�j������Lr��b�}47M�."���$J@���> g���N�7Bތ����3�mxl9��;���D�6wϮ��7��k���G#�Z�^dQ�(�ܒ�dv�K"�4���51�15�5�8����}kk��X<��n�t�MUw>2�j`Z�:''�WW7��>X[^�̭f��zk~e��I�?���b�����@s�=c�;�6���i�9�&A�n?}}Ƅo���C?�]�\�x����<��� ��������������X}W��8:�"�[�cmi�Fۻ�f�f:'f��gG����i��sf*��	7k@C�7�D�v��y�+���ޙ������N�F�����|��k��ȓH*�<%�x;Vruއ~',8���@/3���9�f��2�p\a&l!�p�Y�K��N�bX��4G�SP���8��8�Q���	�f���7�nUv?aܖ[�������d�	}gp�N�b�@��Y�=Z�ǞLζO͵MN��>��)�l�^�p�����������ߵT;�Dh���U ��	IG�������H�hmz��e��{j�wj�w&�?<m�|;[�J���)��y�W����,��S,�����Bc�Y5����PǤ$fW:k;������QJL�����~���~��/[�~���p\����?�ɗw`p`��w�������ag���(�R/�ӟ���P�W����au�>ѵ��u��)���@/-�Lw;�JЗ�S�7%�7��>����?^�p�*!�4F\�@�? 9{�v�ȃ���c$�M���}��MXYv��RbP٧-rLD���ex_ªЪ+�:���U��n��?n��h����V��92*��+5w��eһe�U�{�����2iu��j�)�f2�κ���O�;:4����@p	��0V	����=��kfU�Isͨ��ǖ^��$�5�H<)�[0`k�(/�e��.���hapry�������{S�Y��op�.؁FǢv&�' Ќ�Rϓ��x�я���{�;aq���8�$�ҡ&� Q4(\`"��hU�2��mB0���O����N����s1s8���{,q�`JBA�� ��h��KFrh�0�=0���U+<x���s�?�t��CfAI��-�$ݟ�[��o��a*�d���&4+EtL�=�iν���h>_˓'	E�̪������Y@�N���}tC��052?>2'��X;�ɚuk[�����ZZ�$��������ͧ�����K�9�&)iS��Պ����G<�����2)�F�Lgջ6Vpy��-��--q1ic�\��z0;������,�xo>�ł���EltzCQc��A�\��̽���w���'��3n����wv&��BmU^aeBGR�Hwoa�}z�~�E��,1&+
��Я�o��� �[��#L� ��&�;K�9}���pL� ��&+��᷀�����D�x!�8W��4
���S&tXs��v�"4�$��ƣ!�&�Y�����y!9q!���E�K&�Zr�,:O��=-4��uQxQ��"�h�%]c�38�̚��r6��iI�h�^0�;��Lʘ҂���MC}]jLpH8�kS���W��Y!N&����,�Z��A����*-�gǼS�}�@�z��M���"��ˬ�cV�[��S ;f�	1���)��Q҂좆��ۏ{�}�/�����!�����Dh�p��z:33791�z�������[o4��*j�/�D\�~�\��R�~��Z��u������M8
�!��Y4vnv�o���U"nH�ܔ�>\� ���BE<�4FV#u�AA���X ��9 ta�I#H�H`�#�ü���_=P�GM��f���8%>n���ѧII賴�k�^dd8E�"Lx�ttZ�=�-�ȚD[c��bZ���5���#�1���#���ѵ��Z+�u*�S�oѥ�	�LJ��a�D4F���e,�eY�ш�P�#F9Lܦ��
����2$�9ȡQ�4�i:TМ��26�������ʳ��������G1��(�t�2Y;U�#�	����aq+rηK�����	����eR2o���9:s����*��]�QpQ����癈Kt8��@��*�{ A"��C���CK�\y�?4�K�3sG��qd�s���{��
j1��b�;d4'����8�a(Q0�YR�f�9@��aY���ጊl,�MJ�oL/��O����s��"O�+Є����1�l�膿N{2ʋ�E��b�T�dw�\k�+��@��\F�	�7'3�w<ޅn󯮌̏'� ���řd�V`�on@g����@�jÍj8��Z��:ZO���5s�"-V��ġ&��N,�I��g��95`p\��0<7�洎vL�У����o�+�L4���sN[`���la��gT1h�<�>��������Ir%+6'�:!�2'����.���~�Um��AJ�)�[���1���4��$/}�&�9��~)��a@��"-|�-*�g� �)�^�&�5'���)�R �8��i\�R�W��W�
īI\�v�"�
*X�3��XiI�Yb��)C�՗��%gM"��)	P�J�`�iN)V��!4V�Ŏ��Sx�0.�<~�ϣe"J+7ǫ��)�H�vw�|w����W�T *@տ?ʗ�\ R�Q�@�eT�1k�1�v+������4�P�X�T_O̬wTߪn�U���gjrqm���}���~��/�կ`�۟��_|��>�b}m{~�5=5?48v����"cJrBY-k��H�����>[��W�~�R�N�bw�|O�jo�voM�5��z�Y�h�����\���)iL�ܐr�!�Pm< z_U��ʘ�U����ȲX�Sǹ8pN�р��q��?m�8C	��J@����cF�)Z|��d�'h	0���	Jv�Q ���1X	�)oc:���\�k�D'Y��:�DWS�m�PuViz��>��A��%[t'W�mՏW��b���j*��Ry�U�d�F��E!��Zԑx��Ǣs
�P�*����/2R�r4�'Œ��t�3�!2`J&	ɱ�`Ji��W�u���<d<�o�;�6�0���4�@��w����$��D�e	�hd����9��><*��g.���Ԁ��h�,1=ď��$sw e�x0Z�r���� Ќ��<!��������'Ƽ�\��(�c�7�Ox>f$� Y:]+���&�O֙��#&�LI�h%�2����.o��^_�orxn,�֨(�M�0v�&�����
�u色(.�(�R,�V���u΍{H����t��2����*�8�a�c6������Tbh�6��.+6��--�zV��G���ULk&��sc�\z�s�OTjTE��ԽjP� ���u/��H�  ��N�1�;O*Á�����:����J3�NtCO�!yϳ����)Tv~�?=IJhm��6g}ު�7F���A#�ZH�(-�r&#�8.�t�J�����I�"h���&t3�ƺE��%?Er�NPQ��H�RXR
ϳ4����S�3ꐂ쀖��6X�<6�,��l����.D)�b2"���S�y��GL��a�c���;Ж�=`g�4�:-%�:v@��Z;��pZx�.�x��b\6�/��MQ�Ѕ`V���ҋf�%��Qq�(�� h�� ])�N&�apՌ�N�azDh����d�� ]�V���|�k��׍�W��oӺ׋���(���F��~���2+�)�R��b�ˌ'�"��Bqz���Zfg�e����?��������^ .��Lvw�>|��ƍ���x�V�Zh�^��\/�R�,W}P�|�B��R�v�bW� �n� �Q}ܾ:=��s)���vnM������!kL�ڐ|3	��>���B@�/����Ju2�\LVE�X0��*t��>���؇��)h�.������q�>m!QVD3��D��cd�\n�G[��N��LY]�n�������K�yǮ}�����u��(.lʏ�H��K���_��-�ӥ�,�i��U$��Z�l+�0��~���+V������R ���J�F?<�¡cAbV?nn����VW�����30;F�r�M�cx6�C�����[��LB2@,�i,���v�7�B>C;C]C2�[���o:8�Q�`
�'����s&� ���T>"s�ϙC��(jg�9$��բ�㲁���|W9�Zh��W(�jx2��炠��pE�x�S��H4^����>��$�ī0�7�o ��P��	�'�lrinv�c��r�se`�]O��`<�
b���U"*�{a҇�ZY�P��#�*�AC5��ϻY>�q�k�@��^�H{�$�B��u2�z�p���
��	�t�=��-d1�(�����@��'�� a�-�[� ��ުk�mi�KL*���%���l*���q�\�.�/�%Z5�����V7��X^�r//w��M�a�ͭ��g`Ж�'�4�z.G�y1�RJ#��j*&�$��V}��m��S���~F}K�rk�%Jy�,9Na*�9�*�����mƖ ��$���G��Q��5Bf�)��j+_e��Xy+_c��[�d61`�`
�)4H8�m�/���,�@���� ��;��F��%RЃ�c����&:�w�7�f�ݒ��7
n[,R^pք�>m��g�$ |_1cN��p�F�0�<5����&�:���J`�\�5{�G����\	��M��GER�J^+�s�~�X
��ҼM)w��-�P�8C�/��Nj".E��W/^��G�ԙI��������h����s���qWgGoWgߍ[7s��k|�9]vd�M�����)��-��P�!�~�Z��J�n5*h�uq�^ ��!�(��~G�SZg��`8ِȹ8>���_{�Z�J/������,�ڐ�$`�nf����B�KI��s�9c*�U}�U���X������p����D>����5�T6YR�"�\�VݪQ�6�NV�К�{��o����O������������w�\�3Y�>ה2Ш�W�sV�
K�I6q�S��K�`N�N��������*�����`Hgn���@Z���;	#�p:�����yטu֏uGg������G�dE�dZ�70l��$|��5�И��A��I�v��&�0.� G�����L�Q�;2��^i��'��KvB�v�s`�����H`)��Wp��t:0�7tM�0�����9 ʜ
�C@�S������܌">u�~~.�0�Η�a/ ��͗_c�zM�=s+[��c��j������V����������*#@˭iC��b�����p� ªyT��NX�u��ouߋ,A$��%�*4/������2 z�3�U�Ik�lXI �
��gk@O�)}p�xj=����Ҫ��Z�0kH���o�N./���� �]��������uc�{ve��MUq����Ӎ��6�=媾����g��)��Z*4�"i�Q�,�1%�������}ޱ��B�������h,�ײ�57*��^2��PX��+�dWp��=K�9�zt� D��3<�[xJ�8<�M�E�hIV^�=2�!�u�t��&[��Td8��
g��4d4)j
��N�Koa���D�+�v:s��)J�B㠈ۄ��PXF�r�웱k�6��j� �wf2#�ΤR9� �8��\.�f���DQ61��V�9����k9Q��^+V�R����Ѐi`�&囔�u��b�[f�[F�.��m�bO���Q}��+П��]
�>~l���'�^��E
c�ⳮ�X���Һ�,sΩ�S��`%U�����N��rՇ*���e�w`�R��F�^�������?��n0�n@��)R�nzf|p����L\w�>�h}�١:�*��ċ5���xyY�̩�p�i��@L���`n�EO)� �u���(ʳ�H����*\�zx���pu2��6Y�S�┛*Q>?����]�2�Q��|�Ͼ�W��?��w�����{��O������Gu���ڂ���Ѧ��u�u�js��z�<�&RXDp6�{а�V�v'֍�xG�q�� %�a$<�22�3	:�^�[�t�7j�'g;�C���Ew������6F����t8��N�M�	�6�1�	��l�M
�ĭ��$$���&�r3���
)8�	�"�&°�@�8�C悗�� M��\�>�$$�:<f�����s>|lh|�C����U��6q\�pq��K�y�=!���wr􆑏�= چ>��=+�� u�z_ �#0ɯ3�������*z0�WW �@�4gn�	6k�*�'雸����ǧHV�Eͣu2�п0����>��v[U0F�(�W���	���E�BAEQ�Ss�,�`ZY�8��4���8:�HdT�li��y7��k��S*3j�U$���3�( 4'�A��닥q֫mnrfy�
��g����m����Nc�ob=�ͭ�U�h�ʜ �bbK�zn�-������'W���3�GK��W�tNN�y��u�>�ެ+�>oV��@_�b�7�%� �l`|C�������g���L8H�Gd�#"��W�/(�,pD�`��d:�	��8+_g�@�R��B�ߡ�D1il`���95�M�,�<.#X9O+��"*� �#z�Q�x����8CcC'	8�M��NS�x�0�D���iF9DQv��&�d�)���#���� �׌R���^5�^�T���: z7�~�E)��e��oT6i/��"G���P&��������d�s!�F^�褊8y\N�4C�)�.6Ԯ�R�9��:%@��*Ԁ�*�oW*8��A}��1{k����.�����	g��M���DA��M��:{J$u������G��mH>\c @_�F@�$�M�y�N)��nYL -�+h�_�,A�XsުCFӈ��6\l�������#Y�b�\�Pė�2K�l���6��6a�4�]� y�o^������e��?yo�������]o|��+��DO�q�)��.��Vk���*�P��Tb�E9���M�A���=s���% �4Ι ���<���D�Ő�#R�X7`w��r�ܩ�m�1�[���ޞ#hTR,����
}�V����[�����a��R��48�̭�t��7����0�wV�Fb��
�v���
H��;L-�)Jx��Ap-8?�%���z"�)|$�(VpɊ6�@�!h�kq��0�;��u1��މ�a-��'�m���|���<������7�zgWp�?�~2֓hO�cbl�w&Gf��D*��ݩ��pJu��L��8@/��M���IZJ��X ZcK�-�_W6�Gܓ*6>���42�_�ygi}yusÿ櫸S)��#,��D�L��z�T�Ί��!��03hvY�1������o����Ji҉��Ո���:f·�Xq�W&�K�}$�)J:�v�k���f<��\�i�X�cF�=�--�|B� �I΂h&�i����kuZ�����U�U:�Yy~V�{Sn�gee��bn���8`(�34N$ Qp�X͎�$@c����%dx26Bg��t{D~	�)�;��rQy��ጴ8#鲨���t� ��*�"!:v� #��	�#�OA��Ih? VhH�T��ĉ�:�Ѩ�_<qX' ����$�4�	 �����( �/�a0��D��	�����n��!��(H��[��ʗ��B���������^$@�(_���˅�X,{�R�\,{դx�X�	0-�Q��E+�aT�1�)�A��bM�YR"�	�b�Ξ-ʋ�w�İiZ&I��#hu�M}ޡ8h��J޶Iv�*��)S�*'V��U�@�ֽW�#�߯��4%p��4��'k����=��� �`����'����(ѩJTR�Dd� ��i�cŸ�5  �����rSX�̅�]�i�γĭ�M]$x޶)ì*�]eWKm*m�:�D�_m��5��u�%��g�٣�^�/���?~�����H�A��)2e��}���蝲t���s�VnOc⭺Xg�:�L�T���2�Ll�Da��/<����C�+Xc����!��HM:s0�9|@"~�Â@���4H-�R&]�fF�"M�Pp	.#�L��A���c�%�i���(C;epEeZiU,�r��38@C	`�� �	��8i��`�7�y�:AhB�FK�A��V��!q �ݣ���0M�w����v�d��X��v�D�����L�BS�?�Lb-$4Q�������U��E2F���Xѓ�C
Fi���@�q���E��fG��8ZL�Ƹ�Z��������M���f&C��iM �}07�8��b"()VPb �щUES+���- ��w&ښ��_�ՑTREO�kc���ͱ��Ԓ��j1˴�ͯ��@�n�=���QA��W�ҰbM񍪩�e������lQ��4V%��R�M��{އA�F�ӫ)�sbR��i��mr����㉹�cSSs�^��V��z=^?����m�z�w6�����s��ѥ�
JTd�����8)����,�yWW�|�Zk$s��٭�R�.�e\�{�Q 4K���T��1NQ���^*(,�b��%��JaK��N��n��n���BX_&����+E�2a�S�R"�٣�V��* ��>�P<,u�c/���}���\�%Ni���	ΐGR���屝`K�Ξ�kb��	��	���q8	�nt�Q�X��L�Ѽ0�7 ��;�3Pܜ!�C<�P`E�,�GIl" �EF�a.��\�$x�H�z٬�a��GF�+f�+f��&9��e�����7)�f��0��U�ef�������o�0kS�Ô���%�g`�z����k��Kw9�o�(v�*�,��Y� ��~�.�UZ�wAA���kL�_�!�Xc҅�4Yc���'G�,�%���Ƥ��G1�:�I�Xei�ҩ@�&@�,���{�P�u	t���R&�uF+�^jL�&�v���
ڮ	��`�˳�Ev�̮�:T ��rmIm|sM|g]�\����t�;���o]�x��懷��A'�|��ޏ��䣷kr��{��[y�7�o7$8*4��j t�M����z�(R(�-z�I��c;&�� �B�&p���4���!:]��c#�H�^0;
�%&���4����ʢp~@Wv����r("lr�3����T²�oaG�΀NͰ�}�.Q�� pN[���L�z��% 9C�ƸfR��YH$	�����\u�����$d1�:sZQ�U5"�Y��4&���X����&�lx�����;�����sr���P�򜊺F�x��[cC���<O�?�^b�
�N����m�}��UO ��:��,�aFY-�nRW�=p�����v��ʊ�a&q0=��o�O���W���������Bjenh���I|�R�̉����0�ٳg+��#w��%�R�;��m��A>��4�)2j���kz92������啥���� �3��<A�vc3c7�36��s���S"��,]�J����"�� �%4B�֚
 	� Hh���D@��̒]���U��� ��o�nogh��O�?����Ϸ�u7k���&5���������j(<��|�Ƃ2�͹�S��6_n��\��s[��{�.,�nn��(e�/����G��,%u��c�ؓ'�(����ܨ�2Wlҥ[T0��R��tak�,��O3e���L����{XrTM�;e&��t���S��绅W=i�AM���Av�^:�L�R�5#��f�H���Vr�^�� �6�j�5�{i]�2G��! �h�+����,��qe�i�;4��0�4�hN�����nl�D	�e��,��|n,��'�(~k>Ic-}*���(h+Ep�J�� ��Ì�8��?( �oV24WJ�0�޲hH/[� 4���Q��I�Q��I�y�
�|ˢ`�V�oW�ޱ+����0�&�*��m�s�q��]�����A���To���mT��@��V�-����4�Ւ�6�[�?���iW�']�v_Wv}�+�s[ӎa��=�|W �Q'l���Q�Ic��T�eij5r�L�b.���c��$0uI�`hh�!�k'�����^��E���r��R��uO^LA��j�2�F[\��j��j/��m��=�=�ǒ#?z|���w_�������G�{��;��o϶X�w=���C�E�-��Mi-:�#W�d�`hR���,����4-\)Y�5FC�5�cM���F��NSN�h|�����X��Kt��0,M��`(����vHSxz<��A�'F3o8iOhnLM�O��bԘ�����������,���Ӫqd1��:p�E=��Q�AgT3N���ig:8�������9�q.f��><^�H1�)�P�GL��W���N1�W:�E� ���C)p��\�]Q�{(����쮑��B�^�<����Ѳ��@��#�1B��M�`Qi\���}=<�X^�K2�@��#ՖU�j]��ٸ�bx���$�$;m�6ɒLٶ��k�`����Ov;M7�꫼=uKA�3��rh�Ѿ������Lr����a�B8�mV�k7{�͆b���[��q3���?�T�N�v(l�T�6��g-Y"�^lɖ�
��-�f�[k�00��>\Z���T^��߿�F���	AS1�[�h+ԙ�J�Je�f���z�{��'O��;���-�xH"�2	t>�Ź�.lKZ�M���%*�S��Lu��FyO��A�v�E?^�����d�s�k
�j�f���k���e]�R0�R'�^-�s����'�i̐r��͢���kV�(n�y9hV1��C�i��z{L|`/����
>Y�����l�ASyf"%*�E��S��%�[���ؠ� ���:Eb'S>�/�O�R�o�oU�5 4D��V��UP� 5�g���i�j�m#Ӱ����y����|�P�k'#|;���M��m��-���C��S��[
{�#��� F�(ޮQ�ר��mP��{��Z3�oѱO��2 ��t�}ԙ����?��]]#@��LB ��?c�O��?i�>ݘ#��CA+<��� e��B�p�O����K�h*+V�y� -ጦ$��f��P����NU�G@k���Z���,s}VS�Ň7*�C޿�lY�^�.�~��|��}����l���O����bu��p��=��͊��׻;
��Z :߫�W+�d#���N1 �N�����|:�l�0A.�Q�Ag
0p@ز� ��-��h�/��M���n%�h�@�C�c�T'���<�� ��6�F�"�2�]`\�2��_����[8tq�Ј^�qt�#��y�,��	l����"��z�zhL�$6s����Fa�3�2���m�_�%��9@���8)�3L�w��q#�N�)���F�����֜���6����Мo�}���N����r]��<��Y#u��6�'1d�[���֌��J(h0q3y�2�s�I<�IN����_l�̈́���=_tg&���t�(9eAD'3��m�� �����<��ף���Ɣos1^E����A�Q{�,9m�3K���ʑ�եp8t���l/��A�?���v@�K��Z�������~�:d)4�[�fS�Zt"S^��<��,���֑A��r�!���i"\�Ƃۻ�`�n�����;no�����9rs}7��W";���h����:��#�F��脮D@]�y$E5�:��V�� hҎ6e9u�*�%��i?}_���/��.��j2F�5��Z�lO��P-�����
g����Q����9��>�ZCM�Mx�D3Y`�m��)��B!t�&3y3�B� XB������>�W.g$�(Q)n�9:���v�:�)LuBAK���Ш�/ �f���J9��E��A�R��=����&9�FC;�^2�^���~Ìe0��wl*�
�!���w�j|⯯��o��)}�.~�!z�%���?�U}�N���;�J���zջڷ4o6��jR�ۤ��k�@P�	�՞����C��a>��Y߄c�Z�}�|��cݗ�ID7d}ܨ�V�h�%�G*���!�G4��o@1a��:�Y���!���h!4�|ک8K�)�2Ҙ�Ψ�ȫ˼T�aj̫o���kX��|��o&z��݊-e��]m�[漱��퇭OG��}��ە�o\kiͳ7�J�5����e.)�2:SO
�9�L53�<��Dw��h\<�d��@���.V|+Ag�&�(ZmYj����Y,3J���ca��d�3��݇�v�\�>#	�9��8!���m@s	���M �"��J�b�R�G|�:�_.8�N>ɐT9��EC������K}G��4-�\~�u�1'�[��gٱ������&⤦��
�"�-�-�ڨ��G:m��H�L�K����}�����opy���!��R���j�����̤/2�Y]��I�ҝ7I�[d�����ǳ��J(�
�ύH-���rp+R\Y�������B0roq2�Jw�H;'��8c����a��B`�����"Ҿ���V�m|80��9.B���8�O�h���bҗ�4�]^�����	���v7c�Ӿ����:sB��Q���$V���xúnT6��6I�]N�y֬LOō��G��V7�g箵T'Ve$u�5�ޅ����� n����O�����;��pd5L�����Kjg!��	��ꝋXa��4t�g������W˯T+�u��y?�ܐ�ث�,U��7�˿���O����'��_���W����Kǡ���Z��ze]��X-*��f�EJ��{9Ѝ�Id �,���$M��=f|f"��E4Hd�h0��n����L;^6P�N�(����XT���<��	wDfM��)��I��d0:�jX�1Q�]���Y�E����7K�_/��R&y�B
{	���e�-�8�D/ɹ���I�?_��ao:�`��f�k&	�p�L搿i��f��f�j�b����tK��H��*߯Q�!�[��I>�ݠz�^@���tt��&��[(�Yަ��3��v>������u�%�,:�^�YG�g]Eu�trq4�L��z��!S]�� Hh�[*���]4�>47$�w�@@���e�U�����V{wʩ9��P�$
���0 t�K%�֪��,���:��>��R��Q6���|���ۿ���{�f���{��h��t�|���]�~����ʛ=W������uj�G�vK!P.ѐp���H�$W=#�l�K��4Fd�ij��o`E����b$���|'�	��� �,09�E̅J�_ M=8���tl���0n*�,��5&�3wn௴��t���4�m'�|p�L�<mH@�	��T�:�	4��s��?aG�,�g�/ؘ�|Le��&c��As ������A��-�<�l����c:���.<F��'���Z~%ؘ�.�J�V7>tkq����^��q1�J+%;T"g^����յˋ-����E�f�y���E�l˫��?���h}��ʜ�VC��F���C���t��;w������:Η�O)���I�����tTݽ939��4��6��>��zoq:�^�^V �>�X]z���2v/٠:c���؝�X�:�<+�mh~�Y[y���py����lwErU���?�Y�B���X��g�g.24$I6��AK�ݘ�흛����U�]0*�L�z}��r��u��ov�����-ײ�L��wf&k��l~poheitu���[f��N�i��rR>hic��(��:�j�"ϫ(�Q����{u�1�v��K��{�o�/����o���o|�7��K�?����������r���x]�@���Ai��^���Q|�5ǤZ^,�u33��g,�S
��Ę���̒�9�;+@^�S,���E�f-:!-F�&"��|6%1��N�O�y��Y30-0*Sb�)9���hM��GZ�3m	�{�$~�re�W�D����Y.�_1��$y�"��7��4�^�H@�W̒�m�7�Jhdhj���ﻵ���&}�%�_��^q�_s�淽�����n�x�Z���|��1�~�^	4à�!��Ւ�A�
�mYّ@��3�x�E ���=���1�u�j�����?i���Ƭ��r��ٚz�ҫ�)e���	�\b ���?�u� 5���r@�6�q+�7 �#6	$<�`�vvZ�4�UG	�UB�F�R�=���:}U]nm�����G��������2����_,<��ʣϧ����|�j��'����T�v\�5d�Ԓ|ֹe$��2 W�a��(�@c��j��PA��e��1�sȁC�3 �E�C@3�M�e����`���,}1�/0l���H{���'iI�t�e��� �1���-Q�0��ϴ�N&{�x�)c<����)$=̩4��&�(���<���'⒙*i�3�-����Wl�F	@�y�*� ;��C?��}��1��f��<�T��:�qiOG���5�/42�5mu��q%�R�`R$X��G�hV�;���+o��ܔ팅�9�Zeqf����>x�v�7�[�f�H 4���⅞2J��A��DV}�x��)�E���9�.�]W� f8ˮ�8/7ً�<��2U�Q���EE^�n}��L��!�Ê��*�-4+�s�yw	Tp^�Q�.N��L Lҳfj��4xww�V�y{�K��4haS&�3uU�7�/w�	�q&:4	ެ8oP$���rە�{eOs��p��#����jbIFr��r����Vk�������-�ҝb��8�Q𠜄n�ܣ�U�P5�k��:ew�f�>s���:;�������7��k�o��������_�������?���od�~oԑ?Ә?ܘ�Ѩ��H�jd�n��N��4)hV�q.�8)c-�И����t�Ⱔ|hL<L��֥E;ǣ�y�9�4CB� φ)�3����D�M)Oi��bN�`N��Ӊ��d�s�:��':�EA��(�.��(��Z�[e�7�7��T�@�W�oT�_1ɿQ%�}� ���0MC��4K9�����h�3D�M�_ȹa��e���T@>C;�l Ͱ��rg����5�w�TL>g�]�~�)��&��F%��f���i-������w�LBigy�£C@Oo�ه\��ܳ��v~�Y�a{�O�rڜ�IKޙ�\Q}��6�Vx�zDg0���G�X]*�Z2�:C���dv�hh��'���v
� "�B�in5��ju^��ڬ�u9�Ƃ��k7zM�Ԯ��'��`7Ïz�C���j��9�M�7�M��j�Y^��-�8!���/V�c.9B3��� @Lf��#Q��Uw�Rp�!w\ �J��!2"�aNT�*�}#�i����!K�����3����q���F���{���wYI%ً-�/��{��W"�	$Fs@��TI�ێ�|gST���`ܹ���vτ�����bn����_Z���M�wFsk~w����Kž����9e�1��`b�YK~[3s��/���=ѐ�P�	��5�N���gl��E�Y�d̅�O��c�'���]x�,:i���R��T�3�|��VZ��Yr�(9c��7��+����J�gK�gʄ��s���5�O��N�i���OEG�i?-��Yy�1s���h Т�a	-du�Yy�$<k��p�]�g��h���E��R�zQvE�M�`�H�ʎ7���\��J�f�,A? ět�f}�!/�"/�,'�T�dʊ3i�mzګXW>Ц�)9[��!���.١��g
����^ua���N]נ�ݜ=ژ��^r9�G�����_�ÿ�Ɵ�?��O`���O���������'���lC�|��Ѧ�-��UE�*�#U8h�HrP�@è�@O�F* �0 �S4���Q�6�Y�i��EO=n��:>aD�aeؔ�I%����*/|\��1�����P̨�Z��6P;�)�I00"F����R��Y�(��
ޥ�)��+尗�%�TɿY%y�(�z�� m������fD~�$����߰J�u)�s� �- �U��ЭQ�y�V�v���:	�:�{��w��j��v{�;��wUo4���w[� 4��w[�~؞���/&��_f	�}�%rq���|Uo���΂�����%�Hk޹�<IC��^��V+]r�� M^]���uN�j�4VFӱ�����⌋����1�u�B��R�Z�V�Aw�-D��&G�[��h����Z}IC���rM{i[�����`�������ő���������޾>K����bE��R�V�Q)�RNg�[��L�$[�,0�s���97d�NmjM6��+�d�9pa�Qta&���-���5p��DO���a?b�1�+w�U8Z"Q�q��w憃q,�P��A�9%؉��e���#��)��͎%@�84atvT�Ɗ���i�aU�9.	�`�q��оL�pw���|�~��ex����<�w��`_��*���3���N��V14)x<��C���U�4`Ծ�LbHK�����(e��Ax�$BC�_�z�I|Z�|�(8fH?i�NT~?Tpf�IS�� �e&dl%C�A�-J@�Ӳ�Ϫ�!��@>��č����
�/.;Z�*�Ń�0��$Y�#1�=�N�h��`��7�2N�k(J�-�;�J��r�YhM)B�Es����x2�l*t&(��A�П3�ϙ�G�b�����q@�i�P�W!s*2<��^��V�Ш�Ӝ;�v9�k*���ٿ���?������������~��������?=���g���]������eժ�j��%�i��&�a���ޚ��1^�QK����OL	�?�J�ԔN�Z�y�st��1��6%�4ğ0&7$�,3$��5�.�QC }�L��S�����״��̀r�1����d;!�<�	��{łw�)��m��]K ��214��UB�7��0
_2��i�>_������0��\����7�
j��<��]�7�7��W�7<��\���S�~�Z�V��z�;���p�{�Y�D41��R Ƿ�2�ߞ@��#�H{���dp���G���#^QG��N4�U����#����Zr�4ꅵY���W@�vc#o 4[Al�h37SR'���8h�p�ig)$3
Mv��
��S�~Υ���v�
�ά�*�˻^_X�p��Z\�Uu��=8�02�<����@M_��떱�F���Rq]�Ś�l�F�Q1:KqUl�5EV���,�4˪@�4�1�.=cU${�$�q6��h�{�����$�C��L��h6�I�p��!����3ڀ����/��(�ģ��i(�D"va�h�h���	D���I�e�cG&4~�6���}�c�~�I:�:�l�	�}�r4�8�i�����qI�A�F���c=c��dp������D1�3�:8���y�`����wp.�|3�����p٧-Ԥ����T	��鼼�bJ��Q0@��������&�tP	�ߩ}�Q$8}a9F�#�����Mz�T�+�&��q@����#�L�ñ�,�\�$Q�bk��l�,�
��=������{�Ἤx�֠�?��p! ͵���'�\��흵RO�Rؤh?N��쪳6�1����Z�M
�a@+=�jMt�����n�����My�?����K����7~��k?�����k?|����:������Ϊ��k=-��e�G����2�� �4{Yv�s�0FS
��f�3ӡ�-�
�`;6]�F���'M�7f�E���X�4I(E'L���1���0Rf�y��`O��l 4qPN4�(k*�s��Y�/�4�(9fV~�j�[%�7*䯔�_-��^*}�4���	�V��5т�V��ua��@SL����i�C,��V��"w�M���O��U��U�t���U�^�*߬!F�00
��z%��Dggh����z ���Y\A���]���	����!�C���G����'l���m���O7dq@�}*���t��O�Ƌ8�.�`���u�]�i߀/�X(�)�K~x�);� C!��fۀ����A�V<�W�Q��W�}�.�����r��eh赴���{�����7���fй>��:C��hH}��/���7MId3SP�����Il<���(Q�i��)3��*��G,f��ŤCYmG1�󵠛�]2�,>J���$'���J%����X���3�Q���ƹ��!���0��ᅲ~�qlI��E_p⼀/�>2��P7��8"�K�%F��!vԜD>�G�r'�@PWHpG��F�4H4��0�10�HwA���_'~�z�.�(�5�9Sc�`ǇC�1��[#��D��p���$ۭ��
o��YGv� ;�ʏ{�^�{dYG`x�In����?�K$�C33�Zif&�G��4��a� �-��r�}�&l�lj	(���U2�=��y��#o.�<l�!$?1����a�0��ŏ(������[�0R��I:��c<�(�$B�c��ћ䀾\�36fշ��-[��mv[�G��ӿz��y�q�
.e��&������/�l����^�5�ݨ�l�w�k���,��H�
ݒdJqO�y1Cy����F�q�DQ�3t��p��\Xr%r�Q��{a5��;��Le��H2&1%���
6�C�]�$':R�Dk2�2y6l4�줄v�?��%I��#f�wJ�h�w���R�k�W���(M�zY�+O���T|~�R {�$!O�Y��U��M��
�l�w�j��m��&:���N��v	��N��t~ͣ 2@Ϳ �ߨU�U�~�N���Z��s@�(ͷ�3�ۑ��V�w!�[3�ݚ}��P�Vrk�!�A��G��[�ܢ��S]$�����ږ�f�GM٧�3%9��Y�:-'�z����g�{�WI�vN%-�ɢ}�Ӗzj�c��̼Ҥ�����v��Ort<��Kw��.%t��6�ί˽X���RI�������
c[������rYS�պ����:C�Rʜ*�S�f#�K�=H;�,��u����SPiM�6�����
��%�k@^qT'�4�KDIcDM��w�N$��Og#������`+����ύ���+JB9���F���L'�BOt�홺Lt�8�9�_�	
:�.��E���e|�ܤ]�t"��%
�zX����O'��Y���i��ꬅV����Y��Jb�����C�� ���"mE��r�<�/��8d5x��Hi�=H����`#j=L�>�q�n�&y�xxA8�Cw���U�`ǛD猔k-"���x�8 %��
���THT��N��]� ����t�ə\�S�
CCB�\0���63��5Wؘ�ǝ�OCQ�4��`���T�8�&J�
R-�)6A�]}g��dT�B��E��6�K2�[v��0e[D�����fq�[�
u�B�CJX�,�Y��_,���Z����.������6���D�=s�ϒ+;�	������Ͼ�W?����5�Svv�z�n�Fn:ۋl��k^e�[�t�T�S�
e�Ч�	/J�3+��a�2�RAg�I����@#w�DI�if ��B���R#j"������pn0��K�Z����:'�(�sME��Z�F�r��3�������(� Я�Q��W�`�7+�W��,���%�&��d�vB'd��� �!���&y�.z�!y�-�|~�Z��W��f��Z|Q�ݠ�_����o5Q�;LA��e �ޑ@��#�X{����p�p˿6���9�t������ "����[)����|I}��N�Q��x|���3�4���Ф6��
&;��\�t-��Pz�Y��q���O�z�P��iN9-u����:3ë/�/(��/�-�X��6�R}nQ]���lH��N�TDg�J�F�AوOy2u�H�n�E�̞1�z{�ANL�N��D9�j^��C�pLl�j�PN�vT�؜C`�Bʘg��1���;��l,���`�@f�;�!����Ŧ��s�A��1�2�a8`���Q���9"�A�P���%Ȳ�U�1P���jC��7�G�{����e�fn�	�N����O����8���3��x�� d�7�%�K��ޡ��J�Lb�[��x�xS %���m�9��aP�iN�Ɲ�_{�R��]o�&���+�*61v�ܥ�t���DVI���5��gO��
�8)1�B� j]XQLc0&���HW��f��_�'�"{~Shc�҈���\�Ne��2�M"��S�b�a�����JE�e�!S�4�!O�J�-�b%Z�$�ř���9�8ޮ@��8�çeaO����I�T@K��� ��)ϩ�\�˴6t�T��n��?���+���-֌�K��]N;R">~ה��x����kf��*�[
L�E^y�G*�R�&�K ��T�Y���Rě(��S3rp��^��rց.�7p�ؗ�_�q�ƤcF���Ч��o��YQAP�i�Jj�]�.[ӓ,h������_�GA�䊑��*�s-��ki��H^+��^)�+��R)�9ް(�4�_7+^1�	�U¯�4�a��M�w�7-��84��m�����~����wܪ������jͻu�w�4o�4B�;�*0�c���!��|B�g �;�?l��Ug. M�F� �oe|���]�g�
>aÃ�莂�� �s����l�Y}�&ӫ��yN������lH������=T9������V ͤ�)Ũ�g�?�3�&[��v�\1M�ꐥ���̣Sz3u����l���Y����f�D�с�P�����u�-���||00Fs�^8��"F�@�Ga�f!mC��w�ў�|�H��;���X-����)��M���&���<�;vv�?�E�y��l�
/���S�@c��q"|b/ڑ���f���P U�kUb(K��"���'G$Pˍ�=a�Lw��w�3 +�"�881�A��}�I8t���izˡ��|9��$������UcXo�?7<C���M1AM��ʬ�mx�p���w����Vv��=z �7��لr����0�ޥ�w)���fn�&'��-��"�*��z<V!Ji�M*�)�޼�G�7����]�ʢ�z��NN|SC�R�v�O�J�i,S ]-^J�خR�t�ݶ��W�J���s���v�[��$�*�C�rh�z�z��ݩ�wߚ�n��rf*�*�EY?^/�)pa4Ǆ�OZ-.^��*�(sxJ:J��L�U�b'���"��n'@CA�/���^oh�x��T��8amVYc������顶��_,���|���n=n��Xׯƺ�n��/ƻ#�VԎ�[;;�9sJk5�5*--�D�/l%2���7CABK	|Ę���/�B顁��}�a ��xVl �Am���d-(θL3)x��CD�P;P�li�"&���BDsM���2�h�2��A�5ɾs-��b�[�w�ڷMڷ����*����fP�j�}�B����oh��f�Z�Q:��B|�dB�{N%�-���-���+�:����x�ޭV}P�~�N�~����{����M�V����`��?h#��>��?�yQ�Fk��76W��G]�뤝E�;?�*$�ܞ�ag��ւs����윦 Z_�T��r�L�Izb�D�fUB��h� h:zD1�M����O�J���NE�[�c��yHg�Ұ 6 ���OR�R]�['uk�n�ңUyu���[���"�h8\�s��!y-�Y��]
�i
���8�@L*���Z�~OtOI%�!/b+a���1|cG�����ӤL!)����� Ll_��<g4�/v� 8�rB-�Nͤ����R-�W���+ d#C-m�M��%,�j�}h��q��Ri3rY��s	|�D3\p�PXG�6��������#��ς��)���.	{��*�/\�!�L��(EC�GKr˙�����^5�Э��ґ��g�i(��N식�X�it#�1㛼�ؗW���P�v���C�<�{��4��Z���on#�����/��&��lS_-�.�9tzg^�����^hm/��$�]��Y[^Svs�V�H��L��v�z4ϟ�$=LtP �D6e~��󡕍'����2�&���{��NS
�'�a�������`� y�y��"���7��?u��nлs�V��&7�񠠑���^k�ĝ��z��os&0�:ܪ�g�����ғV�I��MBDQJOr��ŋCQA�?�)���j�:�6�JCNUSamw�݁��G�ٻ;���.<x6{��L������^�P��`�㻎�ە5-������
}Y�&ک�G'��¨�bkC��п�����S��;H��V##IVBXrD&eа�3'�(��|CJ'�h(�(�T�X9���+H3�q��B �i.�h!��8�" ����K�oU�ު$:�^�|ߖ�F���f�����(r�4 :�ѯ�e,k�����XV�a���8԰o9U��(MһV��v��6���xT��*?� Ӳw��wk��*	�Ԫ����4(�mT�4I�f}�M���L�߀|���C��0zmcytm�=�(�*:�{�HO�g�E�f.�#-� ��!7�>K�Ugz���C�!��@�.�U�K>h��"Xd�4ZԊ;:@�S���4j9��cf�{��^�]X�SKr��i�a��� �b��,u�EE��pqX�?5YVq����ST����6���e�WTr*X@6�?@�>)�)�D��_��F�i�z2J�� .�ӁM���3T����D���Ϗ��3��z� :���p��w�o�N��s�P3�0�Y.6٘!���؅ә��"�P8���;i�E�824�.��.�џ�x(�9���0�Ot�OO�-<��ǽ`숫�&���-�Bdss;�����k�H`go����ӝ��zm_�¡�[��|�d�;W��.�oT�j��[��>_l���׫z�&u�U�dW*�Ym=��i�^�����..��6V������Ͽ�90_e��K((�(�
{�qЏ.�k:����������'ѧ�C�cj�>�r�� �d�K:����}Z�ȓ\�F4�ۍ���=��
�nMl��xӭJ�|싧�d�)��uU=�����n(��yr{����^���m�I�b���m�B���bNx�
uh�Q��<J��G��jr�6�[�j�K;{��[&n�������?h]{ܵ4�>5�0t��{�����ܘs�Z��U*Y +XϜ��=I+���-���RJ�5��i�����0@�XG�a��HK����Ɯt�H��u�i��=�5R��D���ô����M+����"Z`DvԤ�~���b�e�WJ�/�H`/��i�w���������4ۻRHAi/W	_3I_3H^3���L�w,,I�I�=��/��v������)��W���C��.�_:�?pJ��}�-��K�F�U�tt��:���j �&�͙0�n��ԙ��Nr2k/�ߙe>���(h˰�	;�?����O�X�]}6tVm&�s�W��P�8Z��EoK�$O4���"������gYՌ"΍���	"��5>��T6A�J���q��x1:J�&C�&/�ȣ��I$��r=S�Ree�����:����$�I�{Д��d,�p���OXK��=��/UxF^��v�|"k�J`��"��oT��f>��M�B)�1	Fl�ۿ�
�ĠF������ �������ƀv$.3ơnp�r���0br�l�����I߹O�qōO^%�y�P!�2�_�-a��VƉ8��	�_��gE��7f�A�9Ұ΅GA��o�ؑY�a����o�&��n�>l��9�h·�َ��w"g3�+�[���6��oz�����J�mz��Ή-P��.6=��DFm�E����\��O��ˁ����CIeWS���\8����ߞ^���$4J����v��g�H`(�Rg��n�J̷�ų/��{���Kn���|�^�B���]�ͅ��E��q����7�F��6���@tg�`���Jd�x�)����F�C"���5{o׎���~<�������o�v7b���
+-&p�L� �8�fa���7E�F�Iu��oX kF~m�պ���|g��Ʈʮ�;�\����rܻ��e��54v��j�*k��j2r�*��/�L�DR�4����u�$�/B��%k�h)5r��G�bc�]L�+6՛j��A�⹃�8K�t�H����+s�Rl�0�s@�P4ti�L�}�l�#�c�MvĬ��J���%�K�qU��k�/��`<����~�
b��%�ѐ�l�0��*!���A�A�m��/l��Y'��/4&��4g%�+��I�2|I�U�6e%4�N�i>���ȫ��W���w�4�m�}�Q��&���Q�~��'���m�|��_w���=�=ޖ'n�~�^�\]{lv
۲Ow��Ih���%�����\stv�^_-׹�*��)�J��wȠ�h��Qy.Xh��<c���v&�z:v��qΥ�Y���Ʒd�j����1�&9ɿ�⒃���v�I�;)�g�WG!��g��3�o2�.��f�x7���\�VCZrљ�&Ž��+)\�Y=�C��L?A��?Q�E�qbB`�Xrg
�aY��IGx.�Q|9�q1�&�j{�B*wl	t�;�#�<��%"3���\�p��7;�aܡg�m�D���q��|@}ғNy<��,Ez�]Z�@9�U3��i|=�G�6\9����0���w&��O�u�Y[�gk���4m�c�E���z8��߫(ɑ���˯uO��J`Ydgwik�}�)7˒-����E��^i�F՘�� %�jɼ��ZYZG}!t݃ie�آw?l�n�<ћ���ʒ��FR��^��sTޘ��|���nhru���U�#�hP9�q:�[�=�������ϟ}��;OvGW�����F`�6�̚e��n���q�����KҲ�e�����V��8�k%�h�Դ*�U�Q��0�2^�ڃ����T�6U�5�:Z�>ZXX	��{�����̙�R����Oڥ/��\��f%��j�jjh��R�/�ϭj�hk��n��m�^�^�m��m�bo*�j�/��)���<Z-�쐃�)���h��8>K���H��J�)3�w�,`���3Za�"Ag�Y(��9���jF�@��8aL�@c����
$9�P��xR(F �X��/�|})n4�4>O���^Y�]���HA�],z����bB�k2n|���*�&�+�+�����,K��[�Y%~�R���'Չ}RcnJm͚6�&UƧV�K�8+1��ϊM���5I�HK�Sj��M��M�6�~T���z���z5H��&�{*HiZ����њ:�����Nv\��Fq��/Nn�:{eyg;s?}i�"�����juY^E�S�s+�B3w5��xm�l�ԍd����D�FA��܉A����e ����\���E4�� 8 ����,Ω�	�,���Q"0�!�k�ǹԴ觃�r�n`A�8�M�������v�Ư�;�Ng�yJ*$��С��|6Hǧ{�K�'���X�B�Wc����Ca
�����`�^E�W�v{�f�ʱ%�)
";�eI�rT�$�#��G�#�<�}"5ss��N[)���'e���[�u�P|r\�1�^F};abuS80�OC|䰦�(�ءo���3r@cK���j�e�D=n��y�����^�t.B� :rmw[VvB���͐���Na�X�Uَ�]����2ps�?y��Z�����b*yNT�y0ymV�]�f֪��L��Gh���f�`��B/3t�=\ۉFw����u�&�9O`�$[�i�L��ꍉ��H<�g��u�F�Ys*���X ��خ-i�,D6���>����ޏ-��+[,i,�H�M.qf�=�[���";�E��%{��R#1gHٹ����UJ��-���#=cF�E���t�n:�؏E�v6"���~EU��*#�B+3z������Phdk9��xʨ<jÎ��l}Urqz(h����<g��R�j���,��6�j��zmvY].4ueC>Kks.Ug�y5Y.��)�9B��G�Nph �� z�^���P�(%�U̇�QApm�
��$��)��F���X�-�g�IЌ�;nJ8f9L��G���lH�6�b�ֽC�Jd=t� Gh���51J߿��N���b�+%�K���k���a2���R�Uү��d%)����U.��A��v��ڜ��������'%ǳ�OT�Tq�jՉ��bө��b۹K����s9���sJw��F i�ŵfܠ�P��N��;�����4��۬�>����6�_��|�U�i����4Hx���Ϗ��8y$m9g;�?�������n��YK���|YCvF�Vϲ�gx�
�L┓sé�v/ :C>��|N"�y9��B�Q��}�� ��C��5�r<�3�/���u��b��R�ơx�%�@̲.� ,����<?�4�-�CJa�$�]8/w��~I���`2��g���c�$�)~ğP�C��\��[ß����@o�A��ɇ�����R�§�Y�3M�H;.�a����`A�M���p��86C��� ��xJ�|����>�f��}O�(n����64G��t�6��8(�TH�&b_B33�d��8 4>qk�n4���`�\�Gx����ūS^�$�Jl��v��û�[�@���I.��RM������Zd;����݈n��kZ�2x�x�xA���= �fW�X��;ܹ��w@�堯i�GZ���\��2��C�F#K���2�Q�b��d�"ݔQ�^;@��\�����;if%�
���ЮV;��-<ơB;��>w���࣍I�#'�$�`���>X���ف`mG�˅�"�EU.�fdX/���R�SZ�p�i�Ȭ�ѺT��^�D����Z(�t�[n�XT�f� �VE��v����k�7��Zl'��|I�#�8�J�D;%W %���zY�K��R�
�K�Q���h�<꼚�|�.ߣ�/�G���dP���.ËH⭔�鴙�gqL��^:sK��oW\�ͨᤨ&����L
�j3��-7+ꇆN�!�@&5'|f��7�SycE����Pƨc�r:�b�
�n+���we��� ����7��CA�t]Ȉ,&]&�T�߮$þY��R����WJ�_/�S"��Av�6/���At��iᕓ��g.W�lO���5�VO�@�Ƞa�^i��K��955r�7��I*w�]w��2�S�rqWNʍ���+X+�n��{���h�hZ1�U��m�?n���=���B Z�Z|�+荍���1�SԞs���Ӯ�O�Y G[�ǭyG��$uY��-��Eє��v��;��~
M�,?1|dh�7
c.���`e)�]�7DQ����^�TC/>����d8�O����F@�d|�etp*�l�,�:}q�,a��x�#��b���YL��ǀ5���F�|���}X��{ю4���Ѹ6;�j�;����h��G@��,�%%'S�2vR���,�O�G�����aq.֜0?���wf4G	f�$�1N�"���)+&&�������,�p#	?�ԯ4QT?~�J����{����0��Q��"�a�w���>�v">���_��勐&ڔRga���nJ�n��&5(ҭR���n�&Tm��1_x�g�تC�Ó�s �Ӽ*QMF�M�d�Z�Rk����k�0v!}��ߒ��fX��6bQ�R�jh��� 3*�-b�g�� �o�L��m�#��uw_S��|�x栳�V+rh��Eu:���@he+��#�Q��xt�7�]s-������u��.,i��@$�٬��T�5
�Re��:.Mo��10z޿^7�-4e�Z5BKV�ݎ�H(����]���5
�NdU�,J�I�n�i�ׯw�V�w��iMw^>j�fa˳�+y�D����_��l�45�Nڶd�"�A#�P��j�V��V뼔	G�T��:,�"h���|��t��n�Q��E{p�)�/�I3�)��E�z���(jL�̜vĘJU�ך�pLRE�x���
BS��iP	4��@��ό	��F���ȱG1�֦�PQ�n,�/�`I�lX�+��^M{�D��u�7���YLn�]M��u��/���S_-�^.y�\�=���Vͅ�´j��˧�.;z�ʐ��tq~�}?:�߄��_���������W_���?|�����峕����x�F��:�̛XT���K�vf���?�W��F����4��w���m�?n��Ik��y�u�����0�nkket��MО�	h���Q�I[�ɶ��M��z}f�N��Т�r@S4�x@g(h�o��q�s������.S��h6bp����e3�T|AyB�:A	�$<�]
��F~�ęM���G�t�i��S�fqQ<����‾�T<��@�B`�N=k�	\Y�u�A-�<e~	��M���<�g�����(L���ٙ��v�0�K��~;�]�/�iu8(���& ���m�AP�H5�Yf��%Hc���e^��w���/��/����D^l��D���,b؅� �1�4����p^ Ά���Nr�c{��折ÚS����(����#Ͽ��︼�x\�Nz8�楣?ahʽ�48�����n7*��t�hH7��ڗ�Q(��6-N�?5(�d&X)&����Lܬ�C!L���Ϋ�ksk�h0�}�����*�ך��-M�oGp�ES��]6�I�f�&�ۄB����|>�.ފ����,	�l���9=�*�9�Z�.�綶n�4޼9����C��f02���]So��Ω֜�G#�_`%���1�kh��vd�9
;Gz�����4��抡��N1k��;��6��ORU�Ig�*��X=�u�;�/�2K3�\Ӝ*ў�R�s�@g0u�,F��s�@j��
Ս���$�<�I��rWL�.2wc�^��(�b�)��h�� ͟�
S.�&�V��\��s��Y4q�,�O�EǍ�h�����j
�?�,� T�Y7���8��3dM�6�8!��QJ���SQ��Չ�B�,�)��z�:����rF�;dG���-�Q,���K�@�ׯ�~�z>��_-�UIt�n��#{FBmZٳy��ϖ�7�������������7_��������~���_<������������W��W��W����W4�j,5���)y5��fUJG槍�jP��A��z��4�oT�eK%� @�|Җs�%_�Z�?���G*� ��\>SB����Zr�� ��Ɯ�Z��-W:�

���X�YO���w�J�n����<wS���s��0���'H�(�?�P�l���� �(O�;��e���#�	��@-4�����d��[��4�?<):�`�S�B���l cN�~S��g�1�F$�.9j>'5/L��a��/��A8�5�e�8�4'c?�d���sJxX�o��q	�����:��M���r|'沱5HcP�&�;g4w�c����'�?�)�>E@��A�k&)m$t��ԯdi�h*�z�Ρ[�z��lG֜�����°1'@���n��b�_hhmz>t��Bh�{�=���߁�n�kV�5���r�5�z�e1eKF!W�&%F]�CAA{.`��OM�I��r��ҍ���P��ވ�g�5��
å����pz�7�����&!�,�JF���n���B���҄֘�lV�K�|\b�U}��bq����x}��f�_/�z4��1c�[������8��Y~֨Rx���o���ZZ�܎�b+ᕇ�/<�w��Fw	У+��m�I���6�<�W��vc���Cގ�G+�O°��J��&I�.�Lz��R���)>3�?5	>�h=Y�KN$ďR)w>�)* ��h�l��2}e���VsXC2Cx%�h�,���)�z�`�Y�N-�&�(�p #�}�F�u�=* Zܐ+�ˎ�)��&j���ޗr��X���������&%R�єD3���}8;�
�)�Fg��8�J�Q��qǟ��y���M���W�_-�J�7�	ު��\, ��QJ��~�z������%;2��
����#�����
�[�_����[��?�}��?TW��tT[-��������q���٩ş?��W������(k��Pp��粫NZY�VԘ�۩td|ڤ��F���y��G��?n!��=���my�����x�~����]�C��#�$�!̥��ܟ��|؜}�5?�9WՔ�o��z�j�T��[�c��F�	�]��W��C��h��f��	ű1�J��e3�R2���i�'H�����v)��/8f��'�2��jA9.c4)S���-�P(7���M�"H���	�$�:ޥ�.�0i�A���Z���q��'��@��>#�-Kd����X�v��f�&�μ4��M� ��ˡ�sq=����
���(,Hc�����Z���4�M8����8!3B�1qmDU;hc7K\9���M�f�e�Sf��
4s�Ӿ�]�aq ��99��r�!��v1����,����3�;�8ʹ���I���B�Bd�,r@�u7�3�9"��H3k-7��#/ }k�> ���J�4v��$�K����)��f0
@�����K���@�\0����hx'�\�潬�(��Ҭ��W/�V���<}݋�.������r�N)*Þ�1ٷ�]��ݑ��K����䑠m��ǕւD���J�g+�iU��K�w6�����ؓ��g�{O��bluZ����3z�%�Y�b��ח�. �;�����`tto{k'�ۉ@V�wb�������^��Ί$��I|�
1?4���2ymB� ~��2���$`�3#�%8��d�L�3Cl���T��慹(up2�R ���l�bha�GDg�gt�p,OpkN�R��3"~�U���&[x\)e�I��USS ����,�3SlU�,*�]�t�%���JB��J҄�
��y�(�
lQ����,��BsO-4�	Mx�I�f��D�<�"�7	Ιip���,��=fU}�j��Wh���ŢWJį�y-�kW� 藮_�Jٔ~f�&�䟼���{��J~���&�D�?�򗿞�v�jK�U�]���ӤR�<=I��S��˽ZXb.�5y[�'��o���M�����񨧺IYU�~�^�m��tf}ܤ�+h�&�_5�~Ԝ��6��mٟu�m�=ٞ/k+~>�{svp���Mڕ�=�μ��
~֑�� :�Hs.4��F���ۥ��ڥd:�4O�Oav.	�D�
�㄀��p�7W�x��k�<X߇�����2�3�Xr�X6�;bl��K���D(y)ebb�E�Ʊ��9���>|�\�a��P�		��q���3EFw��(F�ϥ1�C�uaC���h�8M C��w�/KS�Iͤ%��Cn�z`ܗ�'�����5 �l�:Et��eCj�P������:�\�����f\�r�r�Ø���`�\5ٙĦ��L�s���=�fm ��9��#i��8:�0
YAA�K��F��2�cD�Frw��o�K���5̝�X ����JJ$t��Mj��֥h$��"a_0pk�ȜA��h���|<��6 �H�-Z���wlx-����B[#�ӹ�����V���e�!���;~窧0Ǭ�j�\��l?�~����� z|}*ӒǦ��[3ͦ*n��F7�+�5��^fʯ�߹�ۛ���¤�Q ��	E�`S
-YE�ʑ�Y(��Pde+��l��}�(�<����BQ])n

��۱��.d4�`6.,��L�������?2]�x��ZJeG�V�)3R66�AS�Q��33��F^c��YU�i�h�=s���@�HGQ�50:�!Ob+	P���x*1��:�6)ͅ��N�%�M�D�Lj�]l+�;3ҭ�$�ѪH�����|�Y���r��k�ݷ��G��L�.�M�ݙ�sw�~�P���kY��M�j�Y'4c(���܅M��,I�)�ޜ�B�]'���v-pnQ��F�ά��-4v�*{Z��B0i$��	@ǻTP�߹��v��٫�2
�(�RB!w߸�R�|%���¿�R��'.%$�^K�����?�ꏿ����~f|�e�6U�f{�k���3��B�411C,�Q(.9�LL���]�[�,6uն�ͬ�����+������'��5-��F���TM�2�=�F�_7�`��'m9G:�0@�j�(�(���ҍnl���1�坅 4��u����	���r,��Vx���R�&sSHMɗ�r�qB6Tx	G�p�ҨK��&����8(�?K;�]����.9�����v0��a@�s��h���v�,6`%�5�8���A$���@��;���Kv(@�E�V����:
skR�<�ԃ�6�f�s�l0�@L;�4 `1����GFRB0] �-�S�'A7�RԃtxT��8;���s�`����}ؒ��_p=��\�%��@�s��)s��l��ah���|��|�!���ԒN��(����Lwj3�_6(Jo��C���w2�f�<�9��@D[�絩�& ��E�jz��&��N�Т��j[�O���f`��q�Ф�`屒$�a�6��:"���1�}�4��+��lGqj�.ͤ��w�_^���\
ͭ�����݉۾]�bwoo'�]��Y�H��ĩ��Spw��j�(\\S%����:�9�e���^$�����o-��$fu��]�Z�J[v�x���6����z��{]���VV�[����p�5�-Y��L]u񃕹�H������V�㑪�z��Re������F������v+zg��z�1|��l�"Z�ʆc�Jt�* ����-�����mM:�����3yKb�&�d(�G���� ��i"�	��Y���T=�rs�o*2{{��a����Tb�R[�:��t��ޜ�u{�΄|!8�G~�Dv��b�x�h��+�]m#m%�%�V!L�4��| 4���*ԣ=gC�T�w��\蝺������1����q[�pc���͉���\dE��<y����ɏ�^*�v���2��r��%d/_�r]�z����B���'?� ?�y<�J��D�W��˯�������)�V�\��\[o)/��M�떒��֪�M5�{ښ�VOU������*��5mFm���V;ro�׿�ۯ����W|���oh�47	/5�U���5e��)�-Y�f�̇k�;�Q$o/Xb
zuuzjc�>�u_<�E�8>�.��&L��o+�k�S6�e�g��i�+�o����J�\�Q�=
��C`g����qw9�r��[p�/.
� 61�*5w��R��d�T,�f �<�l��������:����?�W�.ٲl�~�~���-1��w�X8`�]!u��6�ҡ�ũv���#�98����؝J�P�
n3	�i9Drt��Y���H���Gl���]E\0Z,���)Ҏ��EƈFqČ�sN��)e8c�A�����'��f���crd��f�#IZ_�����N�q����8N�^h��&Q��+���@��#.o�_9�7]��/06�'��r"G.�?
֐0�m?�K�f��qy*��G�>�j��
#�FJw(ŖL���a�h�X�@�w��Д�`�֝>OM��*<��d���^�r$
�-��fi-E)Fe�E�n�-h�ov�NO���8���"O�";�0���E�@���!
"Q�ȹ�<z��V���:�2#äͰ讠iY��}�����>	톆�
�B�J`Qjmz����Vpo>h���,T�/�++Zkz/n!�}�����Hdի\W�-N�G�Cۻ[����b��$�V$0f
�z�1;�m`sp"��أ���N{���^�P��+���zrY��^&�Gf �g�T��ޙP t���� |��?5�s�ɡA=Kt@��ʻ�T��i�<ͮ��[���_�Ǿ<<�Y>����خ{n6��|����n0�,������O�x���/�|�9ΓgO�};����Ah|u�s�Y��T�,��vIj�
���*�r�EWy�;�_��К�Q��<cyZ�#����w����������hq�u۝��K�4;�e;fV��X��J��e�7J$/]|�j*	�k·�d�+�+�|l�'��Oꎨ��F���;pY=�
���1��d--���v7�vw�wmj��F�[�� =w�j��Zf�3������]�-:S���U��-8ْF���n���-�Xk���K�����	�����ʐq�*�,8�Up����n����M�����Z=pLDv�4�9��W��r�3�nm�G�tȤ6��!��l�>m��V  ��IDAT��ײ��e��+�{��^�TIh~6�7�B۠���M1z���~<j����cĹU\�$�:�C��;TQR����:��ZکJ���32��n
Vdq:0���*ɮ����u�&:n�tߘ��&��8}�1i^��l�])�i2�9�7+���M�6��H6:h5~�l�-uS��\9F� �8;�Tl��<ٮ�zs��,�K'�ˡ8�y���1��صC7��E�va6q�E�b���j�'C���/��g	Nݴ���A�l����Ϛ9���ؒ���	O�X,��I�c��<dc��p�Y~iN%Z�t�T`��h�r��ޯ]F�X�c��3>�%0cÉ��[�Ot`���㑵�^d��n�ݤ�g�lJ�K������# �?^�mv=�O7h �!��"��5���O�"�E�0H�y�Ȝo��A�ؘ�`��h-���������A��������͍����-�?�N�F����w��bQ$��ƛ5�Ὗ��˃��G7\�沖��������S���_|������m��]���bK�����o��ݝ��ImU.Ch���r��ku���5\�o;:X��n�[s5�+�g�V�LEw�����\��ؤ�e���l��[��vb�����&�I+�,'픓c�y�H Y�|�l(��f�qt;Lګ�#kh ��;����{���u�^0T7T:�5񴙖��7OW#O  @߿��>�>8؈Ʀ����S�������ԣ�<��c;{�1�'	S��f �V6���=�}r��lǿ�1�>��w(E�D���iipT��m���;���ޓg����Oh�`����r����O�<y���'� �͝;����2�K�fS�4���X��b�;%�w+�P�/]O��~�D�v���b�_T���&��{{m��/���vw�Z�nk�m��@qA����q_�� ���M߾�����	��ecC3��qF��?�?x��6��9����#-Y?k%4 �Ik��s�E ���
�6�%݅��x�݇y�t]����	������l�G�t�U������ͱ)�d�Xw�XG�x[�]��Z��.@����.U2 �T$;�bg�g�w:��]�3��;�\3`V;d�6)�5���j��g���Ɏ�a�ΥM���Y�f�����|8�M�N84�qvY�<��S,����M%���k'�S�}���D6@�S��R$;5{��1�j5�4y<��|PX�#��aqL�x$��"����T�jD�m}wqx�p�F��Zt �ٴl��8�BQ��}�P�^v��J����&J2��Zc���سp������;5��x)l�[����]@F���@�o�IV��"�Y��ͥ�����{n�.�d��Ls���S�a;��.���%-������ !q��DCA�9,��s��@X�r�ig�9�&���TX]x�����[}�]��1�^w�m��X��K�hZw���1��7NǞy9� �
�����j`w;� �m����\�M}��\�(lzx�^�׷B�뫞��4�&աZUr�:ӕ���H�Y�-�.��]����h{/L渋E�l �9(���bQ���"�^c���.���(t�ou��|�T|d#�k�Ve$[�i֌�G�6vcO��	O?��y�s�D!ܠ�={����it�k���T���C��e�X��A�Ҙ-�e����Vd��Z�ܜY	�6#۫�`�܈�Q$�v�><T�����\. m����e�Vl�-�5L�ֱ�Z4�=~/ŜA^+˗�2rĹ�{�R���ѐܱ��w�[��Θ4"����@���c+���v�x�=�҇���K��[d��̪^��Np������V4:��=��\]�V7��\
D�ǆB�� њ�CQ��� ^\x��[ߚY��n��"[�Xl�]식I�TEK�ʡ�T��|`u7m
�9���]
m �`?��n�;�p�a�P$���G�cp���rd�v�p�o���k�w/�*��� 4��b���7K��)�8r�ړ��ʌY��"����ٓ/ݎ��Rc{Mӥ�̮Zǝ��N���v��%�̅ԳI�b����o���ѿ�U���Uk��j�<�;�\����,��-�O��':��/*�K��41�1l���
Nu�S�����?n�=ޒ�>����u5:�7;���{��r,��w�$�w���-�f:��z�X撉��t�.ͭMq������a���{(��O��O׆��J�Uʒ�%��;�c[�oǾ�Ŧ�[/C���i!����hW]j�%u+�Y�l�f^$��5�}J�aW��2*﵎��CO#[{k5�,ja7]��2�v�ou:p���/��_�?���_�-D�m��)В�"i�E�7Ɩw�#Oß�-xhg}t��ޭN�YL�hK,:�p�C�x����{��*�Y��+m鸼x�Z�|s��b��wק�C�X�M�BYx�k�'(F𲧓��5��rh�R�*�3����s�g�7x�>�=]Y�Y���X�� �SFsyh�0��"��D4O
�A|��`g�?�g
��,��٩�92��vV�B��[�A�'�ؓ�����ӭ��չ�hY{�]T36I�'���������:��Y�C�ݕi�.�Wڱ�~�ʜ!�k��.i�� �| ��o��L>ʰ\��۵�������Ѻ�^�M�3E�	�[m�X�Ŷ�B���wE�W��N��~4�y"��6�U-1:aU��2G]QxwrL�WB���w��8�,ŚY��q{���c����3�݃T��ۅ�Z�vPV��6���h��o��n��6��V}�Ҙ�V'�)�@Z�JC��f�*@���"�S�5�bs~�[ӛ>�n3�\�ͳ_�ش7��&pi%��<o9�J8X{�+٤;c! ��	;\�ր�	n�Y���X:�d�3�@r*n4Ml���~�zmðښ�j�*@c_J���'6�#Owgez��]|<؉��������l��BXQ 1\v߽5�0?����(��[_������4��pov��ဥ������gru]<LH����ѵ�K�W�ܢtq@S�@cSJMY�w[W�>z����6�3k�ӫ+3�p"|N-/ͭm�B��{�O�X��Ćק3�*>,����b�k�����o��R�-<�A\���1��?�����ۺ�����&��ʵ���[-����VGۅ�'��ª�������=������Px��Eol�_lS���菴� П�do�9�Z o-\?Tг[�U���3]?��iW�G�9��~ښw���BC��V����x5�ŝ����ʔ���?��>��/bO7ζ]t*��z4�s��>E����wbϾ���g_������ʽG�ȪHs��s�Q��;x��^�7]Y�mt��d�M�k�!7��#�3}�'`�J���g����{n���Llwkw}{��Wc�i5h�m��Z���q`3|������ቕ��)�2٥L���;2+��g"[x�h�����q���\)��N���SWk�m�<�_]�_�5uS�Ԥ�D�g�$]�l�8��J�gĿ���l��Yߤ��$�*�(�L
3yK*�c��/󓐢gy�r�ݜ{���=	�F+�X�EC{���Kn�����f��ď\�3�5�45�E1��ہkg悤�J��ִ����Q�&2�H�.��6�.��������wП���}�<�̇�,�v�}6間�����ivZ4�z�qe�)�}zh#F#�c׽�I+�*Qc�֜��A(�E`ty�s�]T�-��T��g�<	6��(Ϯ�ڥ*�D�Phm��u;A��n����4�B�$vEQC�L:�2íZ�
W�ܪ՘r;ﬅI�O�V�w��+�����:7֧}��� 7���5��#B�4#���V��kz�Z�Wb(�}������Mw��&-ZZ��Ŧ�w^�36@��pl9�3;��.0�^m�@��v"4��p�S��gH\�[%q�4μ+uUs���hd)���kM0jN[��C'���Aup�W�S�;iQ^��$�K��'���0y���g/zK�6�������q?�PͲ�E��ڇ7Wc�탽��=4Q�A����"ݜ�fʔZ�������5p+LM˽�ǚ�˸��u�ګQ�R+�ҫ���*�=������Q��=����Ǘx<�a<�y�0Ţ��\�=~#ݼ�������/�s��ꌭ�����s{mUs��V����ٍ-z)�(.2�d-���n*��b�U)!@�U&{�\�V���r�G6}�U>�tMK����_��#�J��_�.l�TO>|�/��܆��n������EUN_�@���p��������sy�2K[Ԛ���9'�r>m�m���6�I��ݟgQ���C��E|�7 �qG�'����o+8۠��뵵Y �ڕW��1���yr����嗟�ų�'�ō�%�Yj;�a)�ݥ:u4�v~vs��ݧ�Ob{����y��M=���R��//N@���y5Eŷr9�OzO��ܳ����,ښ��D
�s*��	M�-����Lxos{g5�Vwǥ�P>����2�۪bې?����Fb����B{*������u)��^�R4�.�gO��v�ę͉���Va�S�hW��/w.L-oGW��͐�������n�$�)<So{�3����>o���g���Cu@�	؞� l�oô MQ�C�Q{�����v`wg)�9�� u60� R���у͙��=*�$�L~��4�x(��C��S$KR�c?pF~����M�����A�Wt�5�.��ڕrk��ő�X8����&j���� ��,B�[�W�/7��Yd؋��١��h:;; ;&)h��`U╹�n-F��8oE]w���L�VoϺR}u|m~%{F�������w���N4v����g������eE�m�L]�5w�"�����n6�@%�S ���w�a22>u�2�94j�ReSf:��+�6��#���͛�j��D��Yv������=�۽��VC[������q��cܸ/������F.z*GE�97�*���u&����gmy�Ra�k��Bo�����1jE�C��ͭơ�Bsv��V��$q��Q���e��8�*�Vm�(t_�����z$]��3kO�i��@�S�ɓ�����(%��H�;���w����vd=����Saς��w��8t(���Y�N����=6�g]��`9�_/ms�V钭�T���Z�t>�]ڎ��7'�K�J���2�*��Wi���4N�f�)����[##K���H,���ߞ����%�Q����*N3�����+!r�E���Ω�,�T�+�����̴���Ҭ��l���^����4��۝�5��5~����R	�Ί�˔o�˿U.?��;S,��&����?�v'v�ysT��7o��L����k�3c��Jo��Y�|�7�{��������[��֮�-�9��)-��MY��di�s-k�~g�M�^Y�_{X1`u��������μ;r~�F"�Xk. -��Px�J�V�,���;����?}����� �Ih���\��u(�ڀ�b�^i+z����b��3lFt���go�Z5)�R����5C��7ެK5i��4��$��䀶I�,�s�S����M�������,��v���s��3��)��ע��;H��F�8�r�kew�6��خ���ĥWZe� S�A�'��'F�b�@���1H�p`z}�Zz٢$Z� ���<����~�z�?�6}��:4Z�%�O|:o�Be׌>��|l�16_��R[�b��t&F�A��S<� ��͠	�)���`�b,��F�X��jtKJr2���S[�|r��/6]�|)�$����'-),И�z3F�qp���,K2��5;����sa�'�+�қ`KOv�h^�C�_S�ؿ�����ohn�e�~�����>nz4X�S#2�i�V;������8�4B ��VY�E_����\
o��7k7�n�N�-�Q{WCa��&Or�6ђ�f.j���ӈ��޳��a��Z`#�d+�l��Y����+@3�9�0Šm����,���w��X�����p��a�Jt5�������2��+T�d�Qx�$:o�_0��*TI���
(М�*��"������Z&t�'W�,�S�3/T*ϙ�qF��r�ethnk�hh788~�����p��X�pv���lv�н���zG�A�`�|)�]��=���涿w���a����y8� ��W��[s����m����at屡�B��<f�Y��!�#EC5
�L�����&��6��}vXk�EG-Ω�Ɂd�w���i%��K��mr�����R^uE�)#ɦI��ӬYE�t;ШDvbہ�Ӄ h\���Y}ڤ8c��1�1	.X��V����������GV�\Cdog9�+��H�g�ە���U�̞Q��IC�;�Pm���F�И��������8�*��o�%��S�ru��ۣ#�� �h8��߉MF���n����K寗J_/��V"{�B�F�y��xn|���W_n��7����Wy���U����/h��fG�?�hr�u�u̎��ͯ��������n�ms���W;����3�4�9'���;����^[�]yhrI{��v�D�L�C+RG���\IC ��� h��[��} ݜ����nlo��[�=�ޮP8e"�}%�-�z�{o� � B[�Nh��4z��m�"s���@R�+(�&P�ȭF��J/Xe)6e�C)r�`�F��J�:�S#sR2�	aq#��P���߮�9
��^��P�6«5����y�:�5�m����3 W���F}��l]������H9
R��X���'7c�P������6:�����+u�Fe�Do�V2��X�n���m��G�M2�6
�VZKe�.����Cې�k[�3���T��"�ҁ�=eH:i8�u�AҞ2	�"K~��og����Zw�EV�!��	y:�����zd;���n�yܦ�HX�0�w.>�\Na�k:��)VZ�4�&J�8tژ �&v�Ɩ440�A���f�EGH왦�Ʃ��Q ^���Θ=��z����k�)��I%Y)��T[F����r�Ǥւ�I�����.ΪI���z�6|+�������/�Ͼ�=�b0���{&��W�T`_�1�t�ƈc>�����&M�CI{���ڢ��裊�:��b"��[�[;k���m�!��{�}��b�"��퉍��FGJ��\ա�å�@�1���8�,����CS��V�;=5�����V���$���4��gQ\0dʬWoL����Ҹ�R���w6��Dq_4<���;�o���@f�ۊ<��V'66��a��Aؿ��]���=ۍ��� ��ŭ���3V-ye��B��2�R�cf���檤������z6ْ�׶��G}u�-R{f�C{�A"��˥y� �Мsnb#L3k�� d,��V�Ow�y���=�j�e>�NyNvb��Ѝ����F�I�FqYf�͌�"����ކ���k�[���4�6�-G�(w��#��ަ�q.5R�j<�ᴙf���Ȏ���̲�&ՙ*Mre��� "�Q���M\���Rś��%߼"|�D�����B�`����Ϸ�{M�m�J��Ñ���@��i�|�3�*�`�CP����������������ܮ��&���\���m�P���T�����˃UCNq7�-��ӎlR��'�/��r���[�rT�t�w�v�q֝Xtw-J�m{sr��%O��"�$hE��cC�;(LO�R�v�;;� �����"K���+R�*�%�����򥚋2��8gb),J�[�������j}�M���*��l�4?ll�uި�R����dY�9���m�$k֥���&.�
Jt�V�)���m�%����r�)�4���ݎ�B��3ݡ����@>��urk���խ�'�h;�_4��3kӗ�B�0�&#dh��`hc{'	o�����&5�G��lrJZ#��ƩG��w��T��,Դ�օ0J�y����)hp��Q��h��lw�q���<+a�<դH�d�MW:��E��wv�S�Z�*ѐ|�L>��y�g6����sۋ/���x�/5�MMf+b��Z-��P�E^zA��Cw��rF}6��d�Zd��^�DQ��o�?��~aevF�JU)U���$�ݠ8Za��>3���e��Vr���L�C��~��E�Y�zu������|p�iH*�?��M�أ�����r\ |�LEMi��`�������Z`f3�n�&�hl�*��)��zb��Q��~mM���В�gdu�f�ĶûQD�R 4��kzx7�LW	S����)TF�W��y���,�5c_�ݥu4��3�w�y��7<4�(���ey�S�LG��>؅N� �`t�������3�qw�m�&��q�R��|������f���vw�n������?toaVn���NZ�@3���VT�P�F��M��̔�QU�GU)��>2���R�n��m� ��\���۞�ϗ��!`��g��|��G(־�Q�ȃ�__+iq'V���x;>u��K���"�I���۳Cª,4rxb'L�;	�W���2v�"M�($���5�9� ��ٌ��uB���,7ʵ΋f����r�ʌ-��8ф�t3	Oؤ�,���I~̨8^%��̸\gG� J�<���ۡޅ�3�߹.�B�j��kE)o�>4kΗ��S������o��Z���=����������	�G��ã t�����܎-����W.��hn�n��m΃�o˓�^�55H��ؘ[*`��\��u��)���f�m���5YJo�ʑ_��5�ۀZۆ����H$
����-�הf��*��rT��;ˋh�h��(��FݙY,�g Аc�L˪��j	Mφ��ǋ[�D�3�iV��q����������퉎�s�k�������[[�K�[CuwL�N��&M�HRl�4k�����`0�s�>��(���y�J��t�ga� ۋ�Tl�q��	����Y&�ȪH%?IvVu�Tpkk��F��fq� znc����H!��VMf�}8th_`�s�Ue��J�e�K�R\���
'G�a������\[V��M+gSi�'�\�,<��
4���`ή�Ӽ�tn�hdnc;�M"��_�?��]�xP.��y�L�=#՘�=?�i���'nóUU�o�矘N��Ư4榛�ΚRPy(��L0����F���}����������Ck���'���p4Bs�C#��o��v�֣"���,i��1�:w�������%��AY�)y�5��������+��nK�����*�<��=^Y���'�(��О7�(\�ɢ<c@;��R~1��u��S���7;=����G��[�t��)�gM2 ⼝V����I|�J�R�[�Z?��4����<������Eyq��Ui'D:��B(?a��ͤ�dA_D~��Q�TX��t<�[v�-��(s�J��M�3FibU��Z�;56��1���lm������g�;FG��sj�q���&�+ė�U��I�yk����ofv�X��}[����+K��ͷ��2Θ�l�+���^4����-��H�>q1hS�ϪR?6�NV)sk�������UN���.�Y��;kS�Y�"S���ɵ`d#��1�HX��`T�ε+ ����[��!?*���N�nDTI��hf
ZR�oAc�V)z�KV~u �� ���H��-�%;� ;o�$��9�돗�ojB����/g�� �(08E�2�O�z�gɑ*	��Z:4�� �y��o'2�[S�Z~X�$@S:������%�|c��/v��o~w����vcv� �?а�{�a�N�����_��W�_<}�����zd��ܴ��C{R����BE����������a�K�s�|oё�fG�v��P�G�sO7d	j� ���:��big�#_t5��v	���6At"6[�s�[f�[-�*����<��@�A`toN�>��Ћ�r�W�dW
�Y���+�ؗ{[�[���nSmY�����?����_>y���γ�o/�
���(�A���9^����`�hS�G'���MΑ�3��V�����7n5�-�+�)��%�RS�t��`hf(l3�9��0Ϛ��֧��{��N�l8Q��_(�
��V���VY�4�צ�:+��6)a1�@��qf�V���9�0d$�Ƈ�����&�B�7�1U�\�f"@�\�X%l��M��<:��L=��[��!�DhH�����-GC��^��滳�M�s&�I'm"����.�*�e֛��;�σ�7��8#%���聢�>q��4�<�9�!3��5�bW��}u|k=��^��,=�\���H�Ip)6��7J,��4��O4?��y�r#��#O:a&@��yI'�?��X����*��<�����p����V%�e$4P���0����,R�oV��m��JN�A�*/�3�s�X�:k�2Q[tD ҁO@�dT�Ve^jv�ovZov�nwԚRK�.\��)��� \<��<�-98�	hAa�� �ا�3��e�s��r%�a�;Έ1ٔ�Uk��m������k4�����d&W�.�+��rP�f��X֋sU�D�6�J�u���{k���*m��pV���ҭ�g�X�B�vy��K�'�����R>5&}f&4�U2KN�i����3>�/!����2�9��P�d������� ��s�]�����tٔ珢>�j����]�����{�{��U��&9d8�G#e_Xte�� �-�����E ���Z$���C�;?٬J1���i(h!�������y)���l�i�->b"�� <j�5��#�{pgη�������2���U�;e�7K�o��/wd�.�35��0���o�����'��j��d�{�ٓ����#ccã{������_<߸�tի��K$m9���Ϸ^T?��z�4���βt�~�⣥�좮�s=c�a-\H֖{�%�L�^T����Tz�xjW[׃K�Ⱥky}mvyqbyuvckqskzm�{êw�%v�ԙ��i,]E@p 	� L�n ��ll��T��,���1\?�<r�4��o�Ә䠃���������Γ�)��
N�,w>���~����0���do� ��n|��Xȵb�3�ڌ��@�?0ٝcR���a�].�������p��o��Xܘ�/���tj���ּ��z�м����c˹�eZ��H������;槗��E�����krZޟB����dS�g���߿Φ�B���[�=�H�(���b�7�4�M�sVe�)�x�w.���O��to�C��Q��ܚ[��݈�Y�2��5���T��7U��I=On���8�n,-.G�"����
�b���L~4��Y}e~�~r���#7�ӭJ�=���j.�R��f-^�
���h��}`zx���3��'�%�N�!G���|���$a|}B�B�%*����%����Ҍ�>k�ZM�U��IZJZK�ăbd'��Q�P�K��.�D����6Ǎ���ɨ�"8kNG�'�,��+��J����I���*�9d�6���a��V�3���G�{���{iN����'��C��,Ɩ��L�����dU$�I��R=�{jyΘP��W�x���e��c�8Z !�V�L1gb���lXbyօ2��
�!��aK��Y�0u���\*����,A�qj�ԉ��������V(��Y���}uB[&9�ҳ�������xeq%�G7V.�X���jÀ�DK��V�Jx��� �X���Đ�3A>���2R#D^�ҧe|͹}cQw����̇���x�i��L�u�Pф@
�:'}K:WQ�U�Vx�@��*9j��������&U�Q��}lm��������V���d�W*�R�V��U��N������ރ/�#�X�������g?ߍF^���={�y`c���H���~����Ñfw���E*��9�L�>�T�����T�`����|#��A���J��t�8hY�֜�my�r��Y��j�Z�Ƚ�Pso�7�XX[���p4��6�L.��&���nX�lJ9�;��M�����Չ%��fh�Z�ZEw8Ϯ��Mqj�\�[��Օ��/"�����x�άY�s�,��������"���ꜳͣ,��别.e9]7�VB�T�bPګw'������jW����bh�e+�]����m�t�g��/l�<�
�C��[3+�S�h`ֶ|���r�M-��2W��]	�W�B3�>���֚/��L��{o�*̺d����~bx���C��Jp�u˪�PR�$6-
�5�*�<pkܿ��Ԁ�bu���"��"
E���Ln�̍����F��ю��Rhr>nm/wT�Y�V�ƔS�3��ɵ��k�媖�2�0�D>_TQ.�8�X)}R�]�`�+�i�
6�C+����������T3�y�y5�b+z��n���h�жUު���7"�hi�扵ͻ���fW���utJb���Z�`�}#� �A9C��Kz����na�{����]@3Y��`t�Y�X!�P��d��[dl,HȢh�%��	S�q����y��f	ZdIV�:
�6 U��ҽR@�)�s��D)6e�YA��(9o��q�L�'M���Kf�QJb��..�� �ϒ��,��@cpĔH9�-�D�Be�H(�NG����r�"�\��b��㆛B�H��0h2����H�* �ϚĸZ�ȣ��t%�hx�$�س'p�]'����aV�)��l�Fj�|srl���(Av0��6?�A�N�r<s��x���v�����@�zhu���|������ɣ	��2ܨ�.��.�����f%uzX猿��gbKK�D6�ƒ{gl ҘS,�[�l֌�&WRx������ ������)�r^}I�]��P�㙣U���YFl!��0J��:�����욟�/h��V�~�J�F��2�O�y��9�����w��ln�UΖ��_�������h�?��`��ģ�Յ ������nO���U&���� �[�w�E=��ɇ���X2<pH��Nw�3@g��3�<��#�Gq��:�[�s��׺�� ���Ց��K�b���x�΃ō������*�U�q�\���
�.�;�˪,�/�B�+����,�]+p鄮l��ҽ������}_d�g�Eg�H�9�������~`g��
8>�Y�W�2E��4K��Tb�;�̍Ф[����E�l�9Wn�f��7��O�}-0mov�"Jۤ�:(j��������\�����х����j`��;�:����'�|K����f˝��[}ӫ����������*5()ϙU�b��|ط��i�(,Vl=& Z���l��9W���//��AQ�[��Sʊ�T�<�*J��R��"�����"Y%";�(�,�.�!�zx�/���F�+�^�����X\\S6\�>��w�b���~��$L&=N*11E���`]�M�`�g�F�K��Rp��eWX��I�E!��K;��ŵhx5@w���$1��'(��[��}�Ӿ����ݙ	KW���$�j�9�0��_�6�����Z��V*�g�x�(��0�[k���Alqh\!	mk*[eF@+��ғ�B�Xq.1�u��f�s�/K��)�T����P�JH���E��
2h'xO�gy
i�	���4%�0&ѧ����B���FhfY��L2Nj\�*�$.���8)>�__F�n�"@�@�z�Q�4��x���`�|$�����DkZ��r.Ƒ��AhE�ur�[i���n!=�D?�=�(�o�=v<^<@R�v�apl5+�����=c�l^�rg���:G��l�琣�@��>�E�^P���/xkzT�x� ����m2ڱ�n�/R��=������X���k�����+�E�B�M���������mE�����ڔ*=��+�@39���_[Lv6�݉��B�f|bLg��by�r]��^F�F6���~������߯T�cP�V*x�L
@���ܮ�l/.�����޿��o�(�����_BD�����/����m'fn����-2Q{�q�|�-_�Q\6�po��IH	���3��
Nw�~ڝ�I7��;��m�皡��55��j�֓w��{wi�zyx���e���Y��xb�:0�3ؐm��.�_����n<�����*�ǧ�,��{��y�l�C't�2�����ӭHl#��v�NkP�,Z�9�����F`=B�Ǜ����w�lYb��m�-+�r�}��_	��������U5�T�)Gc�x����m����6�ܪ�F?=��	y>���̎��:wg淢�H`fe��SP`ˣ!x�_^.�T\�X�W�V)�opju��iRe�i�M�n�h�]ӌ2 z~s���Lf���)'�d�P4��R���9H�@hѿ�=ҭ���n�nWK�:�=����q���^R}�dl�Z�\���B�&�kY�ȣ������h�Ax%��X�QZ���ؠh�G\��;��x;��Q���0(.)�Fu�[A�ÁQ_`η1�<��*�[:Sf�p����b8�kvs���#�1יfW�Z5J���ݖ��%m�*S��2[dʓڮ^n�u��ߜ����W"�ɭ��5�hc�����3��j�� /�X6����dB��`�d�0	"˚v�L�M��F:q�6���&�=&���5�c��\0ZhƎ-�x�(:/x���!/��� ùh�/���(a� /��B��ғ��y%�� ��V���I�[c�v�7��D�ڒX�A��JD��m4Y�|\����@8�/E�X(D���;)�bpg��I�p΋O�D����c���|��F��,�s&�,�V�����oq-��1z-Y�F�X�)vy*e;��7�hvs��F�����tc&���4��2g9�"����8�[��D�����	�)|5�Ζ��#�ӣ�R�M��gCAs@�c����ݹq��0Ւ�j�i\�Ό��m�)�W8�[.�-F�%���N�����I�ڔ����&��ok�rp���u��yi�[�7�$��	ޭ��pd'^�ߨ��F�ל��ζ� ��O������Ͽ�ů���������/����݉�;�F��6���b쎷��I��+���T�@`��0I���v��)<r��'�w~ܑ���|K. ���k�(��z�����ō��{E�\�5Sn)r�ߟ��^o<��w�Ut�]<��<�_k��1�(׫Nmn����N����R�Z���ن�#C����ptuk���KcT�z���{v~%^�ژ_��lWZU<H9�A	���k�K�[��u�L��֪�Y��ֲ3���ږojm�z�U�M@�hM�̂F��Ƽ���@�� �v����\ ���>M,x;��wn��8��>87�g+�j���m��i�܂o��~}��2�����} 4�t�f6�TQ�
%������~:��J��8 ��=�:�F�خ�d~���G��������gk�O�b���O�Vc�}�r�,ͬL�ʒ;ˍ7��̑V��
-�BK�-|���l�lG��5}��i �ꕓLc�5PK�biCf�K�dW�Z�T��y
cX�����F�o>�1X^�����������F��J%�)RXb�;7͘/�\N��Z�i6m��fB�r�K/]����6!��|���%2�"�)�Pb|I'L��b�\�2Ӫ���yD=��>�ʱ~o��N��+3�u>�J����x{2v���h^��bh>4��^
��o��㝔���lJ�E3F�4��d���xs��p%Lbzչ��;ⓘβ�P:'���`I��i`�5����E��d
���
0���g����;k9jY��$���-4�8�)7��9eH��3��,�?c��M߳hSMއ�#++sk� �8��T�dRشl�q���G+3�>�xy�x�9٤���,
9��Įϯ.��X�L	GhEG��H0Qv��f*��<O<1<v4�N)��#gha�9*�˼
��u��)u�E����^&7E���8��� M!�>@�C���1c�$�?��[W>0?��jrwmE�2~�T�f��J�+�i���92��{]۱����Z��z㷿��/�����~���_/�,�/�}��������^G��j�,�]�|�5�TGAbە�>ϣ�9���Z�dIm�݅Go^���蓞��֎ �\u�*�.�Z���/j�~��_�W�+ó}��,�Y�:�ݝ���i����݉��`,�j?8{���X��i�?���δ_�_yf��-�s���Vl�,愜�9gd�P�9�9�(Q�(&1g*K�m��x�c��ﵫ(��9k��}��r>���^�v�]����`�v^�~��<�<?0z��.X�vl�5廯���?'�\���M\])�k�k��.<l��Vj+���R�_N�����:O?"��/{qe�g�CN)D�Jf��%UX���U�e<� t�9E|�2ߩ���Z]�ꅍQ�T�H��ʓ��?��_��x��b��.k�s}|��������YZ�L�0̯�ߟ���f�y�����6�x}��ӕ�e؃R{!��e�n���\���.�f �ӫ�ɛ���c��(F��,����T��~��<R�7/������j�<ǔ�n"�1x-������SS�w��==���ȃoV��'�%��<�)�K���\�v�����lJ�k,������um������c�z�1₼16fJ�s�����@�_�f&�� wo)r_���?�(�5�4w��X�2��(���N��\���JϱO�#3��~�<����.3/�B K��Zr��A��=K��]��]4_�`J��m1L'|g=b�[EY4�����qW)@3��G���Q�U
��#D'�\�����b�ؠ9�k��ͩg)buX��e+�bs�	A��Bh���_kbh�6�{�a�$Fg��(�\ls�{��� %@ڿ�!��#gJ��R��ig)�9}�9l8L�3* �Er_[��h�oޙ�%\_�^�v�J��
�]ǝ���>�/.ߛ��)�.�E�^>�_3�����bO��	,��GO��W�JM��e�_b�Έ�Ly^��ϷIUt���} ��>��dLz��R����m���&�/,��/<zroi�,��f+�r��Գ�oF���GZ�'��"/p�ޚ�Y\YX!��j�?o��X#۪ �[5y�5y���4_l���y0��Z����_���'O��@���~���o>;=S�W/�?Y��D�qqJX~,Vx"A~��r�Lk�e�$\X���p�~�-l+;�^~���3 }���p��d��|P��Q��2�[��5�C����<��N�UYUb�PH:�@�x�ӯ^���ϡg/�-��ӷtAC���v�<�vfu��x�E!4r�G-[Ԏ��է�+�&��z�Yĥey�B)��:;5�h�6y����*ʳqɃ�ɣ�kŵ���'��u ���ܵ��Jk�Вo숌<Z[z�lau�m �6HD��Xb�M]`��Y�[|�>�>��(4� z�ūW?�@��������zud��W��1���
�E��ű�ak��3�sͲ�=�<�L��N>ŁC�6���ɱ�;'�Ǳ�e�ꞇ���'g�\�V�:�$�z��?�*������G� <~������O��/_~h��᪓�@�w����l*R8�� ����P*��į]_\�YZ�+vsL�t*���\�ė4g2�y��U�0�UQ���30N�^=�U��GϞ�[��v�Ge��#|g��l��[r�,9��L3�K4���D�n�G��I���2���"��|�8�&�z�,L�1||�s��c�W���d�f�M�d�M2�_ȃ�%�4��X�%�c ̈́�LqR'j@�˦�TKz��8� ���T������eC)T�
�TN ��v!?�ndFp�4[�C��u��D#��)�A70�sFrk�X�kJ�\A��n>�y�f"$��2&n2xw�H��E%l0.F�d�M����`hȏ< %��J.���(��)���~���'s�f���M��@�wzuf��L����k����\c	�b� �B���/��{jnόШd�����{JSi�Y̼g˹d&�?��O�k��,/s�<�_y��|����C�'�(I3q3,|�I�_X�a<���]�.�65 M~G�&b�����A���kQՇ���A��֣��Ǵ�j��u�M ���U���QpI�-0��gG����]����������a�o�W?�4�����O�{~j���'?�z��2m�k��E͊KQձ��HD~"�)Q"N4��1�$�_�={�r��o���Qq���H{�ᶒ�-Ň�E�8�>��|�4�Vd�j���l�ɳ�GK��&9̬�*r_�2��ǵ?��ӏ?����K��
@����Ku޻;��x�ً�����;�P��ƾVW£
\}�kO��O/Oґ�E ��H�R{�d���'˷��l�z%%�Qy����*t����.?%�^y�>�4w}��Z���bwnL>y@�=^��VCI��*XeE����ޅgOV�>]|��w���XL�&�W��<{���K��̬�/�L޽75bM����Վ�u�"����1o�Gh�b��=z���%�hO�>^^��u�+���yyخZyJ�I��.�ά����/�t�3$%_3���蟙��p���������������ڽ����V�I@gS�\K^�)��6����\��c
urK<0��<�0��M�I�!?��a}rI���3��J~v�(U8�'�G��w�֟�/��!7j�&��[`�#2�P*Ôk��KJ��[�Yf@'W ����`m	F������v�]b�0��EYC,2R�����P� {t.�]T���"���)lfd`�	��`B&*�p�����#D4�I~�k�-t ��	���p�	���o<폘�Fs)��h"5ͺ�(tɘv�)h�9�i4G��2�=��Ac�2�)֜?�aE�3FR	Rp]��cf,8kD���QƖ�R��'����:��4��@���u�p��dn�_b~���6�ŦbkKp|����?b�?[�]�\{���y���ڝ�����!� Oöɒ�BX YX�f1���� 4*Yy�hx�A��NHə_� o��M�C�bk�m4�)[�~�������\]Ԗc��aY�|�*|��4<h�q��&+B�<�2���|��Pi�]�NFÉ>C~4~��&���i!����=Zs�8�P�V�h6�n��|��#��o���=�7������?��Ͽ�ݿ?~��?P�GO�w���^��GO�F����z��0;�VUE�%I�ٰ�h\}$�<S���5��@���X9�;+�u��(�����&��>Rq=2 Z��K�W{�=����hyy�As����ɩb﵁��?��ǒ��=Y�Y�K�wk}�[ӳ̍`}eam����RO�a�M.�w���>e����Nc�FB)
�}Ǧ�����X=���-s�ɇ�%ke��-�ct���������k�oP�j{u�����WpE�P��^�FY)[R��z����|�cqm����r��1俳����9�οz��WϞ�|tfԞ�����c��w#x%���EF)߬ܺ�`�9 G ����W�=��p�UV��*/�K:�o�=y�F��1y����ݙ�����M�2*����1�jP�u.������Q�M��k��q���H�P��+*�j�9�o�ɰu�ůw?\]��s&=<�(��%�`�B��y�J,@I8ũ�*	�ZX#_>b�ށ���?7F�;x~����i�*׌Ю��._�h��6�-\�T�E�~w`��S���as+K����iy�%����:��i�+$�u���ǚ@� f1nfV���"�s������a	��'�F�4�2��Ȱ��J4I��0<"�e~��ܦ`����2�d ��%c
ʒ�bnI� k�Af��.�.A����择�� ��/R���
1̆ e��ʡt:�M��^6^B[LArO\Fd�,^1�a&����1F���O�4�M&5�/��M�04��@6��Chy�ycv3X'�Ϩr�DƗ�[|O��`T��_�B��W�R&���M4�|Y:y-M�pX�MhK��bAZe���[��D��������7���<� ��[�2��38V���^��.����ң8��/�q��{r����,3�oRF�uN,.�wN �;�e�&�o�P�U���boA��|�,�n���`[�Vg��v��W����4��͛��w���h�wj�N�׉[�u<��tP�x������'��^�$�(lK�;п��-���?��e�����X�%TR�(�I柌������'�h~��{�&��܃���@_�(;�Y@b�hh�����S�\�|���V���O�=^]\y�3�,��
Kq���A?}	�1"j��r$��H�������%����;��5�*�EƷ6���ש������t~m<~-,��D��ff���0��K#�w����Ƿ��m�-cÓpt�_G^Z[��s���R�o��_'&�|s�p�)\	V�x�Wfj�>cM�.�\��澩�u�K�O�=�ߓ'�V'�ֻ�%6s�������啵����Io�t�I��l���hz��b G~u��Ǐ��޸��o5��W���>ZZ!?D���-̴��U��YF��t3֢0�(�5Ist����G��IBUs��ZA�IZҴO�}<���ؕ{͞6�9RoK��M�N��5����g��q�Q�es�my�yϗ�ً*�#\��i��L��<�{�BF��N��sK��Õ��Y�Kq�my���+7�B~npqb���ҋ���{�vC�3��^D%���3��|N�����+b�?������ ��]���~f;8� �#&S�8���W�%;�!�N�A94�D�F��7"6���!I�`I
	.�z�pNY�1bzEx�&c���"D6_N�\��^��F��[���ZD ��W	pd�4/F�Ɣ�Ƌ��ě�����Eef[��-��T*	-陦T$���	v�n��0�7��iɀ�0!N&�8�)0	�vγ�L�c�[]�s0��2���/!�1X�c����$�J��T��#��%;��U��[JR���]}�!���S����/>]��(��-�%+גť���\-�r)��jO�>�2���	V����������B���i�(5�����%�G)���M��k�f)�b��i�o@��\`��]i���ʽ����ֱ���Wo.�V���j>0�7������wu�۵9_y��*G���d��a�޽=�׿ �?��Oz������#��w��?��������y kmm��
���ٰ�H����}��t����g�I83?zc�ᶋ�Q@�^������E#j Z��tYt����3�k�k�s�3=�;���rsQ���a�G�=~L��M�6zm�X������s�S����!X/�UbkEp�l}��x%��Y�Y�j��"5W��+�ǖ�ͭ��F�--=��W�e�<>� �#Cc�!�71�0қT�
Te��+�1�䍅��{�6�fy��xez�!�v06�Ӌ��C=�T�ܤiypbu��T�������]��:C�ϋ�:3��4<=f��yf�¡���[\�^%���j�+��%�Lc���|����cҘFo���ŭy:q6y~HN�57���k�Q�L�(]+!�c��LM{����J������������gӏ^��?'&jv�|@��b�&F�t�E�i�E���qqi��b3(4�&��?X\�L��/�L,̷��\/��ˡs��9N�Y�hZ\�%������>�\[�;�k���EǵG�#s3��0_��5.�9t6�e#�Fg_��4h#K�#|��1,\�P�"|XP�b���p��Y!W�-ӄ����~��m_ә��@H�lIG�l�!�b$,c(FZ��5C�9ˆ̗�)B[(�t�h��
��6�w�@[��H�0���R�LK�V�k����l=)�T��2�e�S�̩\k�\*-Ϛ�D��ܻ`��A������PY9TF�USF�	�3 �$J]6�0�;1QdmXsr(�Т�����N-���7�#y�.�W@ơ����'Wt�랍Ń%w8������)���`��?�7��������5��|Z��I����XM�����������駯��E`}fe}hv������ hx�B����U�NO���<XxX㩗�eJ �	D4�c�͵�f���L�QPl/츓\~���0��hti�{fB���D#ۡl1��hӹ�5Y��NY�9u��]�@�Po���x�ǿ����������p�O:����w���������3�K�ӳ��he�_�U���U��U��j��x��-���с�ǹ��^~���XG){��`� ��dYJ���*R�]������]z>�B~\yr~2�SS*�Y�mn�^["?JcM��t�(��Ul=�S��O-�O.,�ݮ��H��"�*2|���:(22����'%�B�������Ⓡ+Of�V��_/����m!-[��C7��VP-2�zw>�Dlb�Jd)�߼yg��8�L�xs�V��DF)6M|xx������*|��[���2	�+]C��7&X
/����#&����fh�_�XX}��2:;30:T�i�/׉9�⊰39�����å�,�0	��<^���3��Eƒ�cZܧ��㘴<�0�ʃ�eѹ�`.�a0��0a�Ƀk'7͜@��I��<��\�w�=~��>0�ѹَ�WT�b�Q\6�xȻs@3�H���k��9P/���5ӽ�3�D�Kk8A�Gu+W'ȣ�r��yt���66ה�����[��.�E��ǧ�w����b�&��W8�$���XsP�h�K ͼ)�n5؄�|�V�pa�E6��y���aɠ���Z3�:nf�5a�� �2�`��I� U�Q"��Qk�:jC�YB�?"��$+��5��dިu�@g�T��LZDY�e����Ǟ�A��_ &���I���Y��ek:ߖ�����4H@gp(B��l ��N��L)i��@y:�J�SY:�G���2���n�KJmK$�<�UQ�"�ٛ^^[�\��e��.��#����(�L�@�����,*;גãxR������b=h��ŋ�~|��W/V��<��c���������Of������/~z�#3���.B׃�bw}�Q���e��6�e���{7 hp����Ew3]N)�)~1�˷���r��%�V���wږ���CZ�T�XZ���^?N��lo��7���5r7��6鲷�s���9E����)/�������?�����������G������ۃpg��>��sm�����T׵�.V���/D������>��?�P��s�u4�d��Y�Y�Dgٱ�r�� ���ñ���| Z�9e��b����������"�akܪ�� >�Uk�rmbzdayrie|a���;�%5�lu���������s�w���7�մZB)��*��^�ף�� #Jݞz`o��K1����pahn���½金k�p�h�](���T���m`jzx~et~qxf�ox��Q#���fuc2�=>uwv	e��N�v�[�r�Rd�з��'&qhxz��������.��p{v���%iq^d��Pn�Ϸ78�v_���3�04=wcb��vo���O�9��c�s�"�~�����*H7��hf���&������Z�]SKy&1y�&b �ϳs���x��. ��V	�R�u}p~ek�)�\MX�'�6���L߽�u>�@/�Z�9�k��\��F��x�5#�5��ޖ�u�#p�0����ĭn���g����h��X�8#��jɣ�fW'�Ϯ<!�@'o-'#��=1�8�p,p%)7��h�Ȗ+@�4��1��X��tf����$��g̀��]$�;���,^�)He�~�-E�3�J�5_F�� xJ���s��l�l�\��{�RT⤟�U�Jçfpɲ;Ϟ��y�,�!�̢{�%�gR�$q�Y��N7a.�s
��gI^��LW3�J��P����%u�YӐ�G�A{�ؖ.��H�T!Hm� �7�3FB2kj�=#�F�Ad�5Sj�[3d�lHL[2jg�`4c�Ⱦ�c��l�*C˭����F���5���ݝ^]�6q_e+�12��Ne2K�YT�L.�+��� ��ŵ&��7���W/����?�x��l+_�w���
�=���K���+�#��KdRqL�LcV�9;�B �w���2y� M~/����}C��U{���^��{-�~��mw�o,=�~�j��+�	9�I������`���a�t��Og#��]#�Cλ�����O�����ZV������DϓG?��ȍ0�O��?b��O��w����w��������]�v����%?6y���V6s�cQ�w���	����>�,8�,�%�7 =�0re�M���(�Ov������`[Ɂ��ñ��A%�#S:DEI����C����M�����K��U�ZN*-������ѫ�S}�J�Zj�K,�R��w}���D��D�����UN)��DD�+����;��s�&��F�ⷮ���EV����wW���w��%�U{5R�Dj��B�M,�ե>}h�f��d�����~S���i�Ъ G����{]��ۆnjÔ�"�٤p�Uv8���C�[����E�2�P��
�L���F'��=HܼZ��*�J�U"��x�������ح[�k=u�Ȭ�SB.��[���oʗ�*Mm��{0����{3+f��k�������[���LM� �K�o��ly|:�g�A(���\{�f^c��	�5ϔ_q��NέÞ�/�;?>���oNL�^���&ٛjy6.
�Tȳ�pmٸ����t&+�-S`��PIKGs��hσ��+���^�|`&eQJ@s�6�L��u_˽ћ�K�����
�3�V'������$�ْXp��g��p��ڲQ!ǖƁ&�A���d�7�=�q���td�[I�X�N����p`_��E$�����i����Q��� :�	��t:
�3`k tp�G��9�K�S���8�YA3E���0ot�;��4��r���@�#��YV�NC�؊� J�aQ�L�s�Z9���-�gHmRk�ґ��g!��2�YrG�Ė�gFͳ��
1KH��Ȝ���Q\���wd��7E�����5$�s$4Gf�)Mrm��>>������T6yK|����J���
k�2g"˒�([6֏؞'��*Jem�ܝ��!'z�y�%�
�G~�.-���"�+�S�#����+�C�Ki.��&$����Xr�V!���3���
����g/מ��<y����/�ן���g/6n�L,�����l���J>y�(�3�mc�;���f�f3a�Vc�Gf޷f�e��ߤ��tM��a7'�����_A�����������o��?��(������W?�N/޺������3>q/�in���gc��o�o��Z��g���x}������7�{��͜�R �Tw�D3��[7�	)r��[Z�TŶ�*�ɘ��^����*���|�Li-ȧ�|Nsk�>d�\+�J����R�rj��ڐ+���
�Ln�HlJ1U\�4T=�@]ح�kaB����f��@f���QJM�)�B�]�p� �Cڂ�EN2T�̅�:	�	}��.�:��XNU�y-�>k��An)��R�d��-J����a*�id&r�Cb�bk��\���\t��������XJn��QHj� ��f|U�$�G·��oR
�ej��)�\�K�l�3�94�q�N����+Tk����Չ�P@��(�f�5Oh��A�ʱ1��ɽ����<�XH�hZ"abB�@^{0�3<�~���[*E%��R���E�� >��hH��.�[A2G!�#[d�)	��2��p
F�:�{�L�A�Aȉ�c�Q�9�;��޻6>90�a��H�ƀ%V[�Z���%�lYls��z�	\N��r�P�/!���Ȗ�J�%���,����6D	4�u�J'�9�H?�Ȗ��:��3�8Ka��V`	�݃Y� Mb	X�R�AF�s9��-�0�qN	gQ��΄s*�Ӆ��bk�%��`=q�l:\f�	���ı�Q0�W:�c�i��,�Af����*&,p��'G��S:r��\1������!L^�t.v��y���GV�-SmG"i�!�#gDb#�(w�hN�]YL�z�n?|82K6���pamln�����3
��]��r"dG��l�DN�Ec�p��h���k���ρ�̮�JB��V�>�n�~��c�7����*�;�"~ג'1��W���]\}�����Gę&>2q�ɝ���^�z���L�9�����V]���@�tgm�6=��]s�+���b�o��J�l3qާ�`�a�,�,�h�E��j�����97���b�����׿�#��[�kO��Wɯ���~������?����W/~���{0����[����H�2,MM�*�;�P~�`�����ls�(��;�܃���={�a���Q~���ܕ��]��:��r�ǂ�Kv��),pKK݊g~!�V�����*SY�J�Hn*�"�\�JF僆b���*�1Z`����'�HE���D6�ȦPJU	-��J�6!�p�Bwp� %�3[!��<1��?Z%�T�I�&G�(ȷ�V��V*�r+\c����Hb�m"��Z@������H␡'�$j#w��r��R��H���g��6��`_LzB��s�C�!-Yd&r�DAU��Z5]��jd�
�������pD(���<x�X�b+���OT�c����r�N�͵���\�Zl�.��axj��"�Vb(�I��N��9`4.$�d'4�Z 	�$.Q)��(�a��Qb`�R�Q��5�qm��2�Z<1%!��X\��T�i��J��Rj(��{��MB-�5�ýB[��炏�$�-\F�1*Ӹ�Ÿ��Y p1��!8��|jP�.!`�����Y2��L)�� �%�s��
�Ee|I��%`B�#3<}��Y��Ig3��Clzn�&���`������	'7��ו�سl�y;��������������B���N���";���鳍�̷�l9j[.P[@� TY�ն<����!289�..��B[;��%����`7���F�O����� E��4�@��J ��Q�z���ԍ����O,v��{;��Xc��5�e����B�z�$7��/�奎�������;�K�>��.C�WA#3�ó��f����ޙZ�59�{,��Ya�Q���X\f�AXB؂k"ξ�Ql@a*&�ɛ@�K�����!��ٷ|���ɏ��ͭM-��h#>�^}N'�F��^����}��Cq���61��m�p��m7�}d�;n����YE������r�3��;8ro��~�������?��_���?���o���|�������ӏ�����O��_�h����?�e}qyj���͡ޞ�.������c��0Y�W��$
�&U��7I��f�f��ͅ�Z������g���;Y@_�<�]y���Xgё���m�Z��G��ӆ����T]j�!=E���I��MExI���K�lH�ؔzA�rA�v�)�.�|S�9M�9�����D�KM�٦�SM�h/��\F�iM�)M�)M�im�Ym�Y}6�'��t�t��5�P�L#�˧�6�R��ϝl�p�k�N7��h@z����7\���]@�$֓��4��D��S�O7\:�x�t�E��&�dS�ɦ��M�g�Q��R����v�������ԓ�h�"���x��c��H[�)guh�&����j�;S�=Y�w��s��s��w�6�D}:j���ܱ�'�.!D�cu����������^������KG���={�����Ǜ0�'ӎ5d��;^�?V%�NVs/h�g2��I�ed;��|J�a�Ok/��^<�A[�7��0�紗�j.�n����g�-�OC��>�6��4a�Dg1v(B�K���9��k������������o�k��0]fj�Dε�2ʲ/��0Q)gt�Njϝ�\8��t���i��ȅS�p���`�k.]֥\h�xAGD>,�U��t���/���0t�����ϟ��4��"J19/�S����X'h��!����I�E�� ��]D+��P�'d�]&�71`6.�ѧ��_�����Q���e:v�������K��r���e>
MBs
t�p��2�O�SҌ��73�)馴�ן�#��`n�#���pԐJ>�aL�6e�(C��iHCb�1�4ef����-�Ae�ӳL�٦�,c�%�k��քg�y}뙼J"�G;r-Y�0۔�k����B5T'c��NcOOC{[�Ǟ�+I�JR��[���3-�Q8�Vx �Kn���m�	馺�$�w�=p�w�(p���M���ޛ7��oدX��[z�L�]����їp���ǡx���S��(����k.kl��o^O޽�12��`�o����č�ӃgnO�ߞ��3=wsjf��d�����mKw��a�Ԩ:��}���P��E�����Lߵr���l"h+-�f�o�xH��9�Ss�i�<S+KU�pD�BuIk��������������kLC�����/��?����!\f�A����{���ѻ#���z����:��Յ�Kc���1�! �Y�tޛT���UG�g�K͍]�̏Ƃ������.wV��8�Yr�����b0�P��@B�ϗ�ϑ�5u���k�����П�J��t	�F	�/��О�Bs�s��_�#���9�9���§�s{4��B�h.|������C����Ou�?�\�>l<�_�Æ35������>j:��� l8�A���OPw���3֟���"���ܮ��;jO�9���̮�S8�Q�YԳ���Κ��TXs�ê3T�~�
����s��Q����N�8���$�<����ӻkN#��������ʾ�v������U��$�������*P��eg�+=�����c$,:���m*:���ȖD��Sp�m�G��%Ǒ�n�w�m*:�n������R�����.<�K�wo�ZrrK�w�o.dB��]�g7�ڶ��RrS��l)9��������z��Ц�#�������T��I��n.=BRJ�l);J�D�g����1�y��;T�<(��n*<��l->��������H��)8�N����E��>���*�}@��[���@�,:�"z�d�G-:���л�����R@�����G6�0�����B��/�yK����͘Ƃ��
�#�.���Խ���ʽ�[���R���KվU|��r�[��!�7o+���އJ�W�^Ԍ~"�V�E��_�{Q
�Ami"�[�o�.����_C��E#�Q��vɁ����U��/�����D��e�as!��B6s��5Nr"����{�Gv��Zx �^xp����{Ň�ؒ�{�w[Q6��wU{7����o/>���n�� J���}�!�j�{%�sx[�ARJ��*�Qth���Yx�=�ɝ��g~V���8�����)��OnS�Vx�`k�!t٦gth[��m�c���>*���Z��Z��Fq�>�ro�l_���
ɗ��=�OK������֮�3�
��it`G��%�o/d�b4whg����~Q�}�X�a��}VI�Q������{ ��+�k���+M=1�k��!�れ��3��N�]r��ꓛ���6��m�y��{���dnsHXXo���4��Nq�3��1s��9f�\T�Pe�mAW������ʭ�����|��?��g��!������������󗷮^�o��5892z������1�L�e�pafD�}Xv N������-�p��A�n.�%����6 �?ޡ�a�w��t���(;�Uv������#�:
���	��Q.#�޸���1��0�@X����y{���}��=9����sI���
����/|y_�9G��W�������ĕ��Sw�'�'�cgR�����"�;�lD>rd@gd�����ؑ������b���J�MeB�r>��~d�A�}k��֜������ٟX���ns߷dC����3�7��6��o�����K����e��iD��M��C��gHG�]�����O��S��S��M��Esa��"��dơ�m�)�/oiJ���py�6�M�67^��pz���;�gޮ=�V͹��ο]����Ȍ�65]�K���t	UmoJ%ŵ�[5�	$B�i[u)�j.n�]ޢKۤI�2�Kķ�ӑy3�B��S�R�y��2����!ͥMM75����՜ߢ'���)��ݐ�U����xB��5�i8˾|���b��I{ᝦs�4��w�.�����ۍg�j8���H/b6ם�T{ns�Y��M�V��wQ��[u�Y{ꭆSoןy��<�	ɤa�P�/k����4�/U'�����V��Eՙ_T��e�iT���"�����DA���Qw�������=�/ugP}���CN��g�[s�Yw� �	ѧ��=����[�s�@�l"�0^vB�h��"^�T�	G����YC=8�;��~�7]�oi.n�]ڡ��U{q�����B�6�G�{�˘��)��l�Y��7��Twfk��-u�1�H�b�HG�-�0j��ty[#YKd95��h��ѐ��>�������qtk#9E4�Qj@��
�8Y����ԝM9�4�mu�;js�Ve!�^��^M��l$��Z���:usmʖڋ�i����0/�4��v5�쨽��:��J·�O�ğUK��U�kT�X�����:վz՞jѧ���5�?ȿ֟��������[F�9�:�m+�]o��0�w(�-V�v�x�K����j���~n�s�rM��Zy��1��S]Y�s�����������L�/>y�ÿ����߿G�.?��u��@W��+�w�ݺ��o�T��M��K�V��)��ɿM�����Ƞ�I����`R}�����k��_#���sc��t��vV��|裝��;���1�n��o��kV�oQ��$���'��U���}1��7a�o#�o�x)����{��o�"�*�K%U�!_�_�D_���}2!)l���3�!I���ȿ
*���g^�g���O\���\y�9�'n>�C{<�O�b�>v
>�}h�~��C��~d��:x$�.��.��!�>u�>q!$~`�O�ߧ8����ּ��D>�r��A|�}K�ns�n*w�9w�%o�9�=S�C֛���vs��3�3fC8����Q����n�����ɾLel�gm�g lĶs��w�`�rv�r?�Q/�3Ym5eA�д5o��:��n!)�lܝ4)졍����G����-��m�,�Gd�)s�%ځ�t�:�"�9�Q�m�r���3 Aq6D%L�
U��Ȗ�V�ْ��6em2�o6�m1b�i��R�!ѥo3d"�9a{�J�5����i���i�� '�p�v���Ie-l�[0i��]��w��wH���-��͆�����/u)��S��^���2�o�SI���M�,t�Ȝ����T�6�����%�m�fn�2޵�obCK:�L*���h�N���I��%f�0���<L2�bO";LY;�]XQ9wXu�Q��t���ȹ��a��Ԡo�%�0&�!�
�����i�l7�3e�ġ]�,! ��LK.#�C�{F�Nw�)�=c.Y�X��v����CΦ)�t�̬
�#���m�&,K,�<L/Ħ �j́�L����*��3����١a�hzf���Ӑ��E�����Y�[ρ��(��$������i��h�0�t���%h~�"t~��Bo#�s�h z����)B���l��[i�{4���;HI3�e|sQ�W/+��y�겪�����To���FC-wn߇�oݾu���`owߵޫW��z�����5��UYE��V��O��b
py_�������&@Q��֢m��#̯zOL]���P®���ꋽ5g��OuF��.����h���h8���t@��B�̿K*�c ��r_|C��P�)���!p=�&.��
I��Ⱦ�I�/#�**�""�3�",�>J��>o�˰�p��h��$��ʙP��O�G��W�O���}����~�>��1�Чn��x��	y?s�"��fY��}�R�q�?sI?uK~�hB`4�n;������}d��|h�#}��pc��p]�v[9 �V�.3�L�;�m�q�Y�F ��/Y�(�Y�D\Ed����Eߣ��CXx0!ȶ��*�Y P#o�KM��N���X4�v�w��D/"�.!Ƃ�	@�g��
^ �R�vg����C����a�nŵdC:m!��l"!5
�!�8(���4R��D�$�t5o��8 )\� 1�l��
4�j�Јpm�(ǥ����b�0E�R0��5a7C�w�D�Y��9�����2�KA3�v�1o�	��j�}ǘ�!;�w��o��6e@�3�5���8��1RbT�a�`�abB`�r����9�l9�X����\�ǤA����"8k���v�1������x �" 53��.�ef&!��p�v`����c��;�� 3@K��8���q
P�}��ƴ����+A�XK�h>��O Yc��V���Ėӹ����N$�(L>�6�ųq��;!�Xt�([�n7&&�o�%�sِL�������92$��4F6��޾��ֈ�3ie1	�|L5*DC[�-N�Vo�[���#t�s��m�t޻h��C�����:��ۅ;�;�������V�9��c+UZ*ˌ5G��x|!/--��4�75�5�f��F�ZZ=�F�D9,������o�d� 7 :}��+�	�����%o���w�Sm��+��ڍ�AO���wВ���ޚ=�,���]䋅��m/8����p��0�M@�w[���vK����pK�D>`Mx��a!]�W��7&cR�k��uL�����!D�̤|M$EF�$OH�MX�uH�eP
}���/�<(g(�!��)�|1���}�#�Z�:��>r�@������=n��8��#�ң��-G
�	��" �S'�j�Y�8f�փ������0�'.	��!-@6�׌�t��M��q�ߧx�7�eL9$Bv[0�&��� �2X��R�?�	a$p�Ẃ�S��D"W8cK�K����#��=Ħ �nP�Y�v暧�_L �BX�r2@'xE6`���\���K�1m� �R�]v�^d`M���"���`
�4��׳  Gaޘ�
;(B7Ӧ\�}���)�fm���B:"�2 �bi�Y�)���t��|f+��ћ��-��:���Z&��$(3�$�p�	h�<�lwp@j��Q�e(��|�.�� ���v
w�Ż\`���)e�
9aSI���`���d>��E6`G�B��g�M0t~�zX�{@$�����h���Ȧz��b�Q��� �9$άD�Q�aͮ�p��������9^��c�M�� �y��X��N6���a�;&�,?&$����qw8��ݼ���Ͷ<"�dBj���r�u��i'h�����d��[ 2�3м�%�`��\��p�~f��D���R�QmLP��2i�؉����O��>3+��8��@QP(SK2���Ҽ2w��_�f�g���������~� �U{[��ZU�$e{[@�֢�-%����:kem��{�3s��]���������`4t���>�SFnw�iSC�j�'h� o!���"mj.8ܜlV�n5p�B�%5B��p��YW�ѬX4C�e�H?K�b�� �2Z�M��|�������e@FL6�z�,�Ag0������4q��A3���7�s�,�« �?�H��*��/}J̀�p����!��uY�X���%p��4!5X��������!Ņ>��(��k���e4��dw��r6����C�Z��Bq\���3�1f)b2����5�:{�9.l���0�N1�B$��8Ũ�`�������$B\<�Hm0��p\�@	c �;mB��e�Q	�]p�
0��l�,p�p�0[2��2�5���!bL�>f��\L�	¹����5����Ǯ_��;A3ĺ�7s��1-��v��[t�	%�&6�
��,�	����\ /؁��#�Q�`�c���!�q�
n��I�bИLb�1�Ĉb�1{Ĉ�a�P���N�%��Cd��]#�L2�@GY���0,
�|Q���Bn��F]��9)W�a.��.!�b�����9A��������ô����	I��n�!0��,��Ve�w���G.j@�P��L���Z)�*2x;�| z���������#�Ѐ5M`|��[�|py�S@#.�l�o��b�>3{D8�8��>v�{h�^Jp���=%"�@��K����F�Uȉ\KĮ7KT�b�Y!r�yթ~�I��HH�7,�6�BYA��T�oQ�Z��-��fL3w���u���L���{'��$|8=40���u�ft���>�Uv���DW!t�Cm���'��i�<�í�6�]p��t>Ң��o.<o�9�PRE�5'����� �ftL@�* �	������@���7����*$a������8��boD�m5��oBJ��������� �E,���s��8��F�0������� ���쁯O��Ag��/�R�3����?��� \F
�N�h;����'.9\i���hr�oܳ��k�}:[�{l�O��Ol"���
#a`m&�5�,�Y�!���S�����؀��wc�3�4�DY�^-�i�+�I$E���V�%"�#�;���f��5�!\T�Zb�\]X�,�o�;AjF)r�3�9�m�����L�����;f����L[2�À�4�����6� ��q?�Ep���F�	Xc��8׀2s�~;�h�����ё�u���m5��1�˼�J����َ��cB�'�z@M|Xb�<"��Y&W8�P��A$���$C�;�Zq��8��sȉ��2� ����2�A���<�
�"w��ۉ�2��0]l�=F�Tΰ�w���o�n�N:�=k6�z�ʑ��I��>�	����c�ɎJ�{���%�v��K��'[���u��(����L���E��	���4��
BdD$��Q���{^�n�����
��Bp���mN�y��%p�%ـ{�����a*`�>�y�[9�Zy�-�C��8->n�x�����9��t�Y���Wy�-��$����L�X4�k�'jU��ۋ���5n.(z�u�t��4 }g��2h�vUeuV^ꩼ�]q���lW���S� ��xg ��������Eħ�(�Y:��6\����X��XR�ȡ���+@��s\��VG7�ޞ&���1p�ˠ!tP��&$�:(c:�ѯ-�* �� ����Y��@����� ���Kne��E�\f��s׆�,#X�?Bƕ0qrW����z��&n�DX"�P�X�q�c~n�|�Q���B�P۸Ȁ�o��/�"wBH��t���M�%k�"�=D"��8ַ�{�v>,h\���,����X���|�	
LU�3z�D�cC\B��kd��41lY�6��q��Ȗtᥲ�#� �Aěc.W�dD�1p@��zM��ּ��X�Iد�Jf"�txӠ-+�#��M\�a o��`�G}c3X���(�t	�۸3�^m�hf��c�HB�s�#� L��a���&�c�F]<�"q����M �,�رcqv��}�,E�(f��3�s����UF��n�bf�D�<Pa߇.އL/&3�5���&�ٳ�3��(���͠BF�;�B����$07U0R����Ж)&�5B���Ʉ��,��q�Ba�ˮ��ܤ���$~�)ej6�E3:I�%��v1�3��vy�Dn1���W#os�7D&f�A�i�Y@�f�5���i�#'�c�\�v�'v�4�3+�����I�t�>w��x� ϗ~	\I�+F�0_d?���8�:��k'��/���Z��&_{�w箚��ݕ9]����J�w��,:�Qx�� "~t{��m���$�MD4o%���$y���s�C�]B@L���7&�7�&����}1�o#�}�ڄ�dG!�+�GT{C
hH�]X���L0V"ϗ~̈��3�����s��숓��?�J��H�8���n"8�_zd,��/#d}�}��/?s
A^q� R�)�7�A�
P��!�B���3��	�PP�� ʠ0�i>��qTN�����1�k�{��0!j �7��\���rR-�u�4�g��!�������8��M"�Z�%�8�=�"���&@fr���'�)�9�d ��e�^ެ�̶���G(3$��?d& �n:�qE6�t�q���f����Ll ,�K���,�� |1���z+)�L��!���bb�H��6+�0,�썎����G5��#=��M8�A`|`���q���!A3s�����D��؈�!2(�8�� ��^B1�p�r0� [����!~e�?���!����R�6�ǀ����s��ˢa�h��n:!3���c� �}d�
^�K�!��ܸ�E=�i��!�,4��{��O�a��}������W���,��N��.f�XË�	Aq���4$�"e݌�����<Ԁ�<��v2v�I^b*0�!X�q@(c�^~��	*�=(7���8ΈǙ�'B��� ��5$�{�<V�Y ���cߵ�?u���}d�n^�-�y�������֟(N �~]p�S�-
�V�f���V5p
�B�ڊ/��IZzƙ��-��,ݠoY���������Ҕ����:��w�m/<�Vp�U}�M�:�^ v��(>�Vx�5�x��d��ds�����	�c��'���	�ф�HB�}��p\y$�@��x���C�'�Ĕ��
�`Xv("�.�Py8,#����B�C���䩩�������@Xu0� �@~h�_�7 ������{}R�ٗ���'���J����qK�o]�+�����'�z�%�o ����I�v�vї���>�	��l|p��	�F:R��O)�'`.l,�\+�+^r��|�姀2��l����<�*����?6s>�p?�j#�V�8�0�L���l�lBT��Ds?%���X����ﱣ,16��î�b?h����kt�f�	!���|s��O%{����2`
'��L�s��C��k%$�>��*�"6��D�3 g�\���Ղ��(N��즲wS��,Ć�H(�Ә��%�#ٚ�o&��6�g�D�n�Ƈ��m�)z�D>��{����;ͨ�d#�rv�1g��dA9�7�A"�L�|h�Õ��0���ޅ!�?�l8�cg1� G���_N,�Ƽ��5������7�#B:3��L3��Fr2�3�j�''f�S��b��M�q�>d����Iǘ��L���pZ�`�`ULc�L%(N���Ń��W�iA�>v�N2�Bl�����EB�B��!���>�G@zȌ���FN�KL�Q?�V�~�����2<n�֑�� 4sS{�'`nX���ęq��)������{`k�=®�6���F�L��/�R8Οy���0���6J��~� yf����EhQ�[���E�ζ���I[z�o�����f�n*멖�ԉ���U��2NgEV[ifgx��^t���R��bK��f"x��Q��U��^v���\2�bk����3���j�'㊳	��X����(Yp&��y�%�/4��O_l.>�(��SQՉ��TXq<$?T~�0$;��(��#�����x	ʞ���E
�GO �a��_�}@z,(;旟��Oq�';������DA�!��_uУ8��HNxd�|��n��x�S��%���G�<�r����#^�~�l�K��!�oC]��N)��C�u��i*��!9����E�I�8e߹���%��D�Fd~E�7�o�"�~eB_Z�_P�/h>9D�P�k��K+�+
)�&��!��}�|�c DqF������/�h.�{�"F$��-"N�^�愱7"����CNT���������t/���G��SȘ1���ƅ>�v���>u�d��։MLv!؋����K�lMlB�$1N�^y{�0?��:��=� �A����҆i���@�I�Y�u���󾴐�G�0l{���-9�� b��y�Y8{`,qS.��NF0�|�o�E�
~d�AO���60�c���j�'6a��"�`�F�C0���b��Ϝ�=.&��gg�#���\�?wr1�ƈl��>!<D��K@����Mk}���[�\�/�I(�q�l���p�b�**$M�q��h!�(Hֆ>9HG
f�9#$ұ$Ȅ8$����
���z����_�I�?w��7�_�e�=!'Y!Xl��d��'NKy��ݧ��o<bd�G�%�
*AN���O���A��1�[��3�;٠����.
�O��6(X�bo�3;�7!X��An[��;�8Ā�5��7�)��ܰ@0��/|B�s� "�x��W1D���큽Q���컄���@��`��`��P���n/:�V��L[��̶֒*u����0����+�[����ƫ�=�}�o���6��k
���U��2H�V*n+A��`_��+dmU��ZA�X�,�'Jxͥ�D17Y�I��˅���^���F�Z��8�`���J�\#��T�:j��Rqk���Z�\�)V�i��5�DYn�4+V����$+3BEy�
AKMn�<3R�ĜDif�0'VƉWd�K�
Ik]^����'�D]n�,=Pe�J�ɚ�pYv�"#\��/�ƫ�m�ʶu�F���V^p*S���^U�/ER�ّʬp/ِ*O�^p�P0#X���%jR%Y�JQ{#r^��!DP0�_��V�8UY��T_1�4_i��첧ʋW���.�)��Kq����IO;�g����|�M~�)'�2��s�/8�/�ԗ����y�
�To�Ew!t�W����3v�9��Gu��>�Q�v�N8�'�ҴHiz��8�xV���[yʮ8�-8�P�q�q+���7yr╨^���/�p*k�-���g�K/��y���P��ӭD�>�q��Sr��CG��chڭ8�QB'=��}'ݪc)�;���6�yO��S~�!;a��I�Т�풣6�	���S�2�r�O���Q��{;ə+G�42H�3q�9�h1�_�фyCc�B��B�Et�.Gx�FC26ŕl�#����B�:$�;��m��v1t�!9�s���#v�1��Cvԣ<�VvI��I&:�|g�p�,[j��%#������ ��)/�I�G���߻%g��^�q7�	��O}ܯ>�Q@߻G�rD���Z�A�H�O;�K�i�I���O�߭8��GU(�"�!�8(�;�xI����!���ahc9H���d�p�Nx�"Le��K�jB'���>�1�)������J�|p���=�C�Gq�_pE��$��!@x�A�w�!����sZj����2��
��~��^T�ԧb�v� V
�܎�ܒCn�A�q8�gx$N֞qa���``�x�q�u�`P�~�d�G��%��������y��A�����q$	H���5YE'#�3q婘�dTt,">����&%gr����Z�.��������崖���]��O���s����D�mO���J�;�vO���o��tTo���	�����]Gu�[���k����X���������Z:5��F���`j��w�v�����X:u�n���r�X�]K���a��)K���U�k�j�5���v��U[�l�kn�I��&�%!M���E_���57�$j��6�����fcS�l�����Ioh�5$Mmf���T�l�M��K����ֶPMqmC��*TW�+T��H�-�UU�u�.GEL[�+�4��+#������T��k���`}q���VE�kb�����PmU��KÍ������(P!���\�ԡ�|_��S�v�*ExY�E=����L�(T�Jd�B����[�J��z��Y^��������&Ԇ�T�5���bF��$�XmPyK���]Zݢ�L6��ehJ"���:��@�,���+�%2g��xSE\��u�j�1H�	�i6"��j0��u��҈�,�Qy+P�ڏY�Զ��a��X�.�ە2O��_&��j������B體�J�"��`��Y��U׶Z�:l���H�FKõ�� PM2{JT���hc~�N�)ի�ը'?X���k����W�ȑ������Gq\�
��tRl�r_Uq�Q�)�
��u�P�./
֫}5���P-�Wr_��_��C�Kܥo�}���2�Q�Q�+�
��h��[
)cu�@��W.TB<W�,T!��%%�:tC�y�Q��[YkRE됹�����Tah�:T����݅�@ʖ47*����k��-e�A����
4]ܢU�*���S$W���@`Wc���Be�
)5�F��J��O4)��\W��_���}e�dcmUҬ)hn��I�=Ehqy�N��*��Yv%�]�n���!�&ˢ$�E�M��\wǥ��J�\�Z�l�����J��L�����r�9nU�W-��,����,�"�.Cz�+?˝��+�!����P��j��"����/D)��/��
���0�-I�0vE�^�l����Us�(R%�V˛PO~�V�������2��K�Z�(Hs*�������%f��/ڤ��4���]t�#I�)�;���4��C|��8e�.y�K��Qfxi.Y�K��pC꼀*ǧ@��Key^B���
���bN0?7�̋*�q5'"ϋ��1�0!�EE9a./.6����J�ȗ$�ĉB����%�*�@���ɉ�۷c7o��\�W��+��K�u{�UkK?�ճJ^5'���^]�G�������^}�K�5F{L�NC��Ż�����Nks����m���P�1�f�u���rڨP�
�[#]�`'겆��V����k7;[�=��؛u�k���r;��.G�ۉ��:��vy��P�#�n��:B�`������o+�p��iw��ӎ�ksx[���L���3X�t��k	�:f:n4E���ҙ�z*���H�')������57��H����0yZ�hΙ4zZ-�
E���l��fG����\-sX��5�Z���֢rKLoKR�����*�s�YQ�=A��6��b���5�/�y���@��Ь�6��hk6"FK�lk6�%����V�1�#�lF:�4�[L�V���bMڛ��$m�ZܭN:��e3m�QT���Vw����<g���ewvڐqg�j��BsB�9:i2ŌƄ��b57[-Dk��$�3Z�G�i�R��َY"CN��1�%j���Zs�l��Z��)��G�ڰ�E=f}@��oԆ��	�K�6���ͺ�A5"�&�1D�ڠ�g��q:La�>l�,A�("z�W�9nBh�!�34S�<�`JR���1�m6��ͺ��=�k6�G4!C���q]C�Q�օ꛰x0��.��j��ИԦEI�1AYZlt�yt	�&��&t�VJ5���a܈��c&mܬ��"�f"c���Q�6�1&���P�������N�&��EMz�R���5 rBua��@c���)���D�D�}u�}}DW��Ŵ���QC]��>Z_���W�+���Ց��pmu��:�XW��ܘ4�u���jc����.��J4U&��c�p ����T�S7K�n�τl�V3Zi�i TU�!�/d��V�$'L����ï��F4T�WÁ�j����PME��:��I4UD�T�F�J�U�Z8su	MC���ë�7V�+�u屚�xUq�\,V��å���p[!�C��TW�+�c��C�����p9���������PaU��2\R����ַT7��C�-��m�u�e�����Ś�����ڎ���T�[��R��o0^i���j�j���^c�H��0s��P��`���G߀������Bs�Uc�=��m��1!l�2�t電����Pw�Hgc�K��mn�0���[ډZ;,-�Ts��'�P�ٜh��[�h3k�$;h�H�BRZ��DZ��V*�B��:o����G�]�&_B�EJ���=	S���$�D�a0i	�h�1yC(5�&����6{cf_�HZ!D"��@�NX�1�/�'aP�6�|u����o��(��WO��wG5�`�3���7zCZ���rTl�fw�3ث�����쪳z)O�s�<�?�uk)w�o�}M���2��&�_���=���u����������{"F_���	ʟ��	{ �F큈��0�@���i_����(�X�1+����-oZDm��1���H�(��ŭ���j�a��W���g�苢B��7�c6D�����=d�M����%0:�g�B��&#��իqG0@�-d�[�b����Ӥ�i��%h��� �h�}�O�S� �	Y14o����\>=��hm^��Cb����W-NΈ�.��eT��o0{��Oo�h�|��]M���HY{ �6���D1v�;B!�3��;l�z0v3���D���tP�s���j~����0��!�ů��>���1d	���&�X�C���Y��5�k�d�<Z��Sa�Xla�٧G�0�����m��ְ���Z\�6���i�PT�٢�֠�C�tƬ��~J�¡W����<{��
[p����c���������bG��0:��̛'�5�u�:�Ӈqi<��β[q�U]M���:O�%�Cd�y5�lj}����YQ뫪�V�y�ዠ���
�ᣠfXJs�C�8j��8�џ�����0(:F!�Q{Ԋ9q%�R���"f�C@��3�	6hC��`��Wo
5���@���Ó�D�~�NS�3aІ�F���p�>�do�og�`�k��&*�`�jm�#�d7�#��X�+��׹c��Hu ��5���e�H�7YG���77Z��V�����V�m���W�;�]]e��r����]���Sf�p�����=u��Zw]��6�є���e�4?sk|�sb�kr�kl���D�ݱĝ������p�����;�[7�ׯn^ݸ�y3|톿���o��w��3���������vC==�.O{������Fw�9�Z�-��6G3"펎.7�d��F[۝m��D3�l��j�tw��@p xG�'��m�p�m�%Z-͎֤#�cq:��'-IW{���7������6'��-��CFP;1G��hh!��Z]�[s�F=ш%53q�ߧqy}a�
��'W�E��C���W"}���6':L��N���n[�������F����tv�Z:l�.To����=�-��w-�IO�+z��P"�D�����
Ƣ�ǫu�VC(b��\����Pk������ho!=����[� T���~`:���/ZĴ�ɉ:�1Z$)I7i7Fc0�4�X��M�"1ut��:H+I��(�Rh��B�٢qg8� L�a�.{�`�����íqz��ݍt�+h�<M�=k$ �@F���C1;*���-q$㮖�'�7EB�����qŒ�P5�1.�13G�d�vW�=��p�Eb�h����-'��#���4az[Z}m�X���@��:ۣaks��ނ���-��X��k0ۛh���1;�&���v1�p`h��3`�=:X�p3L��5�*� c��E ����kFm0��OO��Z2�0�>�'L��7@{�V�y6�.w�~d@=�l؂�1�Ȋs��~r��#��x��	��*��h.d��L������D��-�<>��m`�{�l�ӭ�,�9��;���悱$�ݭ��tv���ˢ����58�vO#1�.-eo�:�P��P
v��iԹj��Z�I�?\\���`=2`�(��rj1^O���CV���x�f���0z�&\>8
>��o@�'����	h�>�.�~�&roR������[��Y��Vh�r����QC�)w��Sk�����5o�5��
��z�����pA:�����y|����1��BM_m�[�C��`y,T��KF�["��`]2�5�Zb��X]<^m���U���e���PwU��*�U�mj��&���tm�ڶ.]{����~��U����կ��7�y�ZO~���?�j��_?B�׿~L��:��_=B���^�Zz�|���Ϧ�<�~�j�����/�x2���̓��G���+cO��f�L�\���59v������٩s�7a�gn�M���]�Y���D��M@K����p����������!D�W'�=�}�h�ţ����� )�4��<��ח'P�������3o.�-/?y4�R���={�������DO��=�����O?���r����2�����|B2/���c��/�-�"Z|�t�@+���g��NM�� �ߘ�>�ppa�����������^<[x�xvyq���������}6\]c�ޙ��=�p}~�h{�|�7?=�.�ޝ�����pmerq����������������]�7�sg�)�mqvdi���4?�8?��D"�	*���9>�?z�bt���Mtr|t`��������Gk��������'k�kK�Z�;�so�o����`��;}#�W�\81M�./���ML�������Ź{s�w&�o����[c�=���:1v����C��fi��L�ă����kKח'W�0���{���q��R�ۨm�&&!�5;u{c�'� ������SwgO�ݹ}����7ov��}��\A����G����!�ћ(��D-�,��̍ q�v��;(�ݼ�~c���^�����ё�R��۝w��o�l�z-~m �2�e�7�7:60|���;�C�{��d��A�[7��7D �J�5x��3؍̃7�{��}=��pGg������Nd&5��9�2x��;�ۯ�F��'�G���޺�}c�}��K�v��z�z��}]с+̓�; d )=�l�������u�;�|�=�a��{}è�VZ�u��Dx�B�o#�I�#���!��d~nt\�ww�{���W�Wc7n%o�l�>��v5�ȭ�ͬ#u�/|�/��]�M�vF���\i��i���tEz�B(���=�r�n���mw���kn}p�X_�{` t����@���7p5�Ǩ������~%t�j��`������B=].��͆<vx�}��+}�+W]���[{����~劯�����l��cn;CW;÷�b7{�^�VW`�/2����l���w:mכMw���α��hop�/:����������y�u���u����{�����Z��p\��
ݍ�I'��[��u���'���?����Ͽ��������?����Ͽ�������?���2PP�    IEND�B`�PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   �IgU�lp��       jsons/user_defined.json�_k�0ſ��sll�����F`	�Y�2°l���'�+!��Y����f�}�t��]�9���*�B�W�{�jmT��r^[I��)��^�R�V�N�îx�[m6�;�)�N�[w�t���a�t`u�k)U$)/"J8��8b�J�	���k�s�z�+_:�vm/�>�r">n�=������N����mSol�C<�M����[��h�	Βಋ��=0�j�9t
��A�V7���8c,��/�D��)X��6�T��k����mz:BO��u������ ���D��ݰ~2�'��|=ȧ#|:��i����/g�g�N���d�/�>jv?Õ��r�~�ZHNi�L�2z�UO�(RV��(M�,�JV�	��3)d%����)�	Ma�ӷ3J8�|~Fa0Ki�!D1�$�����g2B���|oL��7޽1���7PK
   �IgU����  �                  cirkitFile.jsonPK
   tFgU!�+�� �� /             J  images/0fc7fbbe-b47a-4373-9472-5e3944978531.pngPK
   1�_U���R�$  �/  /             �� images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   �IgU�lp��                 �� jsons/user_defined.jsonPK      <  ��   