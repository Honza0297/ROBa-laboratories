PK   �h_U�׶|�  ��     cirkitFile.jsonŝ[o��ǿ�����R�܇zK�5��F]���r���r���RC߽sȵDi�5�s��,������3r�/I�>��lڰ��}�l�+�Vɭk�G7>���]�]w�����n��/p�v�w!-��]��n-Ea\�*���S��,-x���*c�/-[g����Ջ�'�8���e�O�Km�SJ�:H�yk���օ4Z	��p����Sp�)�����9V,�H�w��I��-�H=�>�ď!��H�86�"��H�8�?��#��H�8�?��O �H�v�G�'P>ǌ�Ba�f����$�I�@R/��K$�I���r�QW"��D�'��I$ɟB��)$
ɟB��)$
ɟB��i$ɟF��i$�XG��i$ɟA�g��$ɟA�g��$ɟA�g��Y$ɟE�g��Y$v�����+��[���&�bCd�QY�j-0Y������B�l�ys!�K�%�{^8�A�E���BzQ$e�$^�K�%���^z���_&i���hf43�Ŝ�bN�i(�4s�9Ŝ�bNC1����P,h(4����H1U�q3P,aV�qCC���X�P,h(�4K�%ŒhFL�%M,�4K�%Œ�bEC���X�P�h(V4+�Ŋ�bEC���X�P�i(�4k�5Śh��bMC���X�Plh(64�ņ�bCC�!�f����Plh(�4[�-Ŗ�bKC��&�Ko�߷^z[��Js����ޥ7K����Ǿs]���؆C׺���'�"H�H/�ċ&�bH�X/9uD����h�e4�2���aF�0����P�i(�D1��bNC1����P�i(�4s�9ł�bAC� �J�P,h(4�ł�bAC���X�P,i(�D3b�%Œ�bIC���X�P�h(V4+�ŊhaGC���X�P�h(V4k�5Ś�bMC���X�O�P�i(�4k�ņ�bCC�����Plh(6D�l4�Ŗ�bKC�����Pli(�ߤx���o���x/�^�_�_?u��=ֵ��\��c݆�z�qe��z�nZ�����KT�IS�<��>��/S'T�z�E��qya�ț�7��g�p��L��ȪԬH�Ȫ�u�Qx�����溴����Q�
3Y�h�i�s�J��4�\Hy��W�*�`s�����L{/�y��^�-%L�����a�F��)���w���k�i�]�!F��SA�},�yn wT	��l	��8t�D8� ����f"�¦�̑���¦;_����E	���E	fzaay(�܅����`�J|	�C&� ؑ�N��C�}xb����T<�t�=�a�5�1&��#����h��s�(dq�iq0$dq,R�c�B��aeXB�ǒP�P��"�`9dX�D�%��#%�D�%�cI�X9�D�%�cI�X�D�%Q�m,�bb�F}X��CMb��
,�˩�r*��J,�˩D�.�Sb#�Ē(�$J,�K���$*,�
K���$*,�
K���$j,�K�ƒ��$j,���ƒ��$j,�K���h�$,�K���h�$,�K���h�$Z,�K�Œh�$Z,�����Y���i�e�ŏ�,[�-~>�d��~�<��=�G�{�\_��bV(TZ�me�V��m�wi����ARi$f��Ar�(8(x��/(((��u��($($($($($(((((T_iP(P(P(P(PhPhPhPhPhP辝@�A�A�Aa@a@a@a@a@a@a����E��gAaAaAa���.!�3�͹���m� �����,Q��x��5���4�'^N
�O���9��Qfuw�۸"l �S��_BwU?����NM�h�&q4���m6���k�y��Yo�}���Uy��*SY�.-*m�*W��Wk��w{�s~���_3����M�:艙\oFx�w׹x�K�m��B�ա��w�-�m���z�[�����1XW��9���P�>��u�$���o��o�����r�}��}h��u�	����C��\u�������P��;��=W�q�QI���%�WY4����Z��Trv�ՊIs��tvlO(��Kr�WZp��D�+�Ҳr.-�g,��,����]��Y4ꭒ��c���8�aO�u[n±ߧJĢ�x�ݬ�AD�� Yd>�H3��E�-bl�F�	3���E�-|la#�G��j�l\S>�)ה�k��5e�������>��6�y��W�y��W�yU>��y�$g�6m2�*;�p�6�y��W)=k2l�dgU�*�5�y��W�y��W�yU>�b�u��с|�R�l"���3�l^�켎�3:uF'�������2;���*5��r��d������t��l�=<ئ{�����`����6�Ãm���t���m�=ܛ�{�7M����U�=|l�y�'=���<�]� �������u?ϹN�����+o���uR����B�A���q�(s�Rk�N+�W+������n��	�?����A�����eZ1��X��4��̴�^�J�Z���C�d��� Ӕ��܃r�U)��6��{����8Np���4�.��e�SǜM+��7&E�
�_o���ϱM����k����quXQaD��R�Bl
�f�,+Ep��)^��m�7��y�ν�2U!�D\��`�L�t��*U	�Mxy�i�a\�JUŁ<ͭ�㤋�eE�bS�q6W��������m} L7��s�?�������c�zl��+c�ۦ������v�b+�媪7a���(UY�BVe)gE��ǅYQ��U�4�eF))�rE\��"
RG�r;7.�b�-� ʊO�m�<��.6zY�4�^���i��j�(_�e\#�e!s>�4��,��N�9/�U8OT9^'��_�Cw���o_����}w������r�/nCV]s��M��_������_�h�4�~�\��pӆ]p]��cgC�߅M(�F�W�*��?a-��ty��OV�q�xӯ~��w���ͯ��Kv�.�}ص߻Ic��w����߻�k�鰥_��@u�[-�V|�
�6fBi5^2'���Yre�Lj��iɍ31<���%ࢽ�%K�~>_�*�F�3&��Yf��'d�	��%;:V��1��Lw1�������	�ͷx�����=�]�,�Պpg�5�w7�9�uhN��O���'�ײ�s����R�\?�?=W~~�6�]y�{'o��u������g�`�����q|f��.m�����^��8�ڭ?�k�^g�uߑ�-:���x���vo]w�����:�ͪ7�[0���=��z?����9�WS�Rƾ��|y�ǋ@����q7B����-��|(:>5���2>���>�&Jٓ��I�c�\�����N�1������A=����y>v<ϧ��Y2����'K��Rff��Ϣ��tKi;�	i�t�	b�4)m�e��e�=M&N�sHf��$K�L�O�l��=�랎}0y�7�7��qI��qb�W�}P�/�����m~h�^w���o���PK
   �h_U�׶|�  ��                   cirkitFile.jsonPK      =   %    