PK   JvqU%V�  �Q    cirkitFile.json�]o�X����Bsk��qH�ng?���40�ً$ hK��XYY�to����H��f����f�ӑx^?*�J|�s�|Z�������������ե4�w�q�qx�h�X}����C��q��nu�I�]�~��-���asuHc��*��f]��*�x-Ew]IQVq;t]h��u���|���+�Y!�bf�*��43XB_��
���V��7f�B裙�����`U}gf�*�~mf�*�e/�f�D�J{�{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K$
{�4K�s+-|_��?n���~]n��	ۢ�t����*��ͺ�-���m��qe<1����^w��8I����^w���^w����dvU[3�^�K{�6K$
{�6K$
{�6K$
{�6K$/j?�5K$
{�5K$
{�5K$
���V��k�H��]�D���N�D���N�D���N�D���N�D�k{�4K$
{�4K$
{�4K$
{�4K$
�⪽v���i������Y�k�Y"Q�k�Y"Q�k�Y"�v�%��v�%��v�%��v�%��v�%pk�^;{�4K$
{�4K$
{�4K$
{�4K�>�k�Y"Q�k�Y"Q�k�L�����X��͋gW�7�q�%�#�n�?儥�.$A4v����.�%���J',]�+6v;�NX��!���l�P:a��9���J',]��gc�ءt�҅�ecײ�C鄥}�Ʈcc��	K�5�5;�NX:����΂��O�Q���m/`!���a�|���U8~��`���Y�p�`���	̧����n���Og:���'0��ц���O`>�]�v,��|:/��>X>��tF?|��,��|�� ��?X>��t%?�}��%�?J��|���8~��`���u3p�`���	̧�v�������O�����'0�������O`>]���,��|�:����O`>]W��,��|�"��?X>��t-#?z�=�
��?*��|���Q8~��`��ӕ�p�`���	̧kv�������OW����'0�������O`>]��Ư���'0��M����O`>]U��,��|� ��?X>����?z����5�?j��|�i�8~��`��Ӿp�`���	̧;�������O{�����'0�vIa�������O������'0�v�����O`>���,��|���?X>����?z�9����?��|�i�(8~��`��ӮWp�`���	̧���������O;����`���ip�`���	̧����������en;q��/s�yo����M�r�̰?o�9��wg��󦛙�ϻef?os�9��?en�X�Θw��r�3o��W�xc��v��o̾�nV���7�*w����o�gR�xc����o̿��>���7�S'��˘�}lr�[�x��7���e�o�k����;ۨ%w�1}g���7��lC������m�;�z�h,��-3�wA4~|���3��"w�1}g;K䞸�w��C�xc��vP�o5>����7�;ޘ�����7뫟;ޘ�^��������ۘјјј�1�Zc����k����5�_k��c̿֘�1�:c�u������3�_���j�&W�uh�Z�P���(�밾��&6�o\�}������J��:�z]Ǣ���7�:ic��o����q|:�ׇ��qu��r6��V���oJ(�d� ��W�"H(���
z?�!���ޢ`� ��w="H(��
zo�!�����a� �0�A�J$W�����m�
7�ƻgV�+ޔR��ALX���SJa�	1a5\�"N)��)Ą����R��BL��7w�����R�lCLX/���LX/�:N)��>Ą����Rg@LX��:N)�q�Ą��
��Rgs@LX��:N)�q�Ą��
��R��@LX��:N)�qĄ����R�ALX��:N)�qZ��]�.�cu���8��)]V�k��SJa�;1au���8��9nЭ��7X���8b��x��qJ)�s!&��&w{��V�)�0Η���:�`u�R
�N�	����R�BLX�X_R�_H|��WW����*.��?_����q�`�П�S�U��z��k���g�`\=XŅ5�.���w�b"��*.��<�%��]��x��k:Gq��y7.&������\�*WVqa�y�.\����������
�ՃU\XuN��1�q\.��C�s�}b�亜l����%>�˅V|hu��Ol}ܗ����y���80Z�չ�>��qa.��C�k|b���\hŇV�b���Ǎ�Њ��)񉭏#s�Z]�[W�B+>�����Ƃ�/s�Z]��[_�B+>����'�NwĜn�����Ǘ�>�̅V|hu�Ol}|�����Z>����2Z��5�>���e.��C�k+}b���\hŇV׈���Ǘ�Њ��u����/s�Z]��31�Ǘ�Њ��=����/s�Z]C�[_�B+>���'�N���+����ǗU>�̅V|hum�Ol}|����j�����2Z��^	>���e.��C�=|b���\hŇV{W���Ǘ�Њ���p�m���\hŇV{����Ǘ�Њ��D񉭏/s�Z���[_�B+>�ڣ�'�N+ɜ������Ǘ�>�̅V|h�g�Ol}|����j�#����2Z��N>���e.��C���|b���\hŇV{j�Ķ��e.��C���|b���\hŇV{����Ǘ�Њ��j󉭏/s�Z�9�[_�B+>��;�'�N]>��|����Ǘ5>�̅V|h���Ol}|����jOF����2Z��ޒ>���e.��C�=2]b}|����j�O����2Z�՞�>���e.��2���:�f�,���TY�&�����;Se��v��B��L���ֹ[�#*�3Uz>�f��L�.m��+����֪�2L/m`�+����6��2L/mƙ+�`&��v�̕a�xi/�\&��v\̕a�xi_��o]&��v̕�N%�,��՛oj�+�d���u�2L/m�+�d��Fl�2L/mw�+�3�xi�\&��v�ʕa�xiO�\��d���Q�2L/�ϔ+;&��6.ʕa�xi{�\&��6�ɕa�xi��\&�#���>�dqd�82Y�,n�,n�,n�,n�,n�,n�,n��lL�L�LwLwLwLwLwLw���X5m�/�:4E-q(��z]��uX_me�����H��SX�ˡ�]��㮨�u,��J�z롓6Ƹ�>ˋT��|e�ӡ�;����������v{:7O��������Z"H(��d"H(��w"H(���"H(���"H(���"H(���"H(���"H(���"H(L����Um�lcu[��M)���&Ä�n��7����V�+��R�n3LX��SJa�Q�0au���8��[�w�͝�cu���8���V�K��SJa���0au���8���V�K��SJa����q��WX���4#�a⮤p�R�:^au�R
���	��V�)�0M	b��:^au�R
�d%�	��5V�)�0M�b��:^cu�R
�/���&�]��x��qJ)L��&���X���4Îa��x��qJ)Ls��[?Xo�:N)�iV"Ä����R��K2L��M��&V���SJa��0au���8��	�V�#V�)�0M�e��:�:�����|ֵ�V����*.���u,�U��z��k�g�
hU0�����Y9Z�����&���Y�8$��΃\�:k�D��U\X�9�K\gM�x��k�g�hU0�����Y�8Z������~�)�V���*.�:'���8.Z�չ�>�ur]N���w�����B+>�:��'�>�˅V|huμOl}����������0Z��5>��qb.��C�k1|b���\hŇVה���Ǒ�Њ���񉭏+s�Z]��sc�Ǘ�Њ��U򉭏/s�Z]s�[�;bN��||Y���J_�B+>���'�>�̅V|hu-�Ol}|�����D����2Z�յ�>���e.��C�kD}b���\hŇV׺���Ǘ�Њ���������\hŇV����Ǘ�Њ�������/s�Z]�[�يN�}|Y���*_�B+>��6�'�>�̅V|h�ǀOl}|����j�����2Z�՞>���e.��C��+|b���\hŇV{p�Ķ��e.��C��D|b���\hŇV{����Ǘ�Њ��v񉭏/s�Z�Q�[��dNK�||Y���j_�B+>��3�'�>�̅V|h���Ol}|����j'����2Z��^T>���e.��C�=�\b���2Z���`>���e.��C�=�|b���\hŇV{����Ǘ�Њ���󉭏/s�Z��[�.Nm>||Y���_�B+>����'�>�̅V|h�'�Ol}|����joI����2Z���.��>�̅V|h�קOl}|����j�R����2Zym���n3Uz�f�,t��TY�㝩��y;Se�Wv��Bw��}���ҙ*=�s�J^&{�6}͕a�wik�\&��60͕arxi��\&��6�̕�j0��K�T��0Y��d���K;.��0Y���a�.��K���@�L/m��+�d���u�2L/m�+�d��Fl�2L/mw�+�3Y��X���K�m��0Y���U��`�xi�\&���gʕ����K��0Y��=P���K����0Y���M��ő��]�`�82Y�,�L�L�L�L�L�L�L��e6&�[&�[&�;&�;&�;&�;&�;&���fq���I�e���8C{�.��:����������_����)���Pʮ��qW��:�p%E����Ic�}��E*OY>_�����_n�~��yuY^�>�ۻ���p������p�l���ׯ-��	p�{e�z{�ڤl����Ǹ��?�����b�:������?�����}?�������'>�����;�m����>�v�|:������V{o	��%���`�0K�񦵑�,ƛ�F
�Do�)�a��n�0K�񦽑�,ƛ�F
�D')�a�t`�0K�i҂�lՓ(�@����5�4����P��]#L3?�@���5�4����R��]#L�_�@=�τ����|(�%P^�a��c� �k	�W�F�fY9��:NI:K�`��m	T[�F��HY9�j[�֮�YZV��V�٫]#L�Ĭ@y���j��L5+P^+���5�4W����
��v�0�ֳr ���]#L��@=��zj�ӌE+POk���5�4g��A\Q%.����]#L�>�@=��zj���S+POk���5�4��z���PO�a�|k� �i�S�F���Z9�{T�M*��6@=�k�i����PO�a�Cm� �i�]#L���@=�@=�k�7.�5�����&=��������ď��/���?�O`��ϚrzH�X>���߀�7�h|�,��|���߬;����|�� 8~������	��Y�?N��'0_�g�8=$~,��|��5������|��,F��v 0�Є:��!�BpB�����N&�Pg��1��L(4��ڥcH;�PhB�qLǐv%0�Є:[��!�L`B�	u�7Cڝ��B�,u:��C�	�&��ti�
M���մO�	�&ԥti�
M��0��wL�[&�O)i�R�>&�P���1�}
L(4�.ݡcH��PhB]gDǐ�)0�Є�F��!�S`B�	u}Cڧ��B��4:��O�	�&�uu�ڧ��B�@:��O�	�&���ti�
M�k1�⳻��]�O�h�R�>&�P���1�}
L(4��ߥcH��PhB]{Lǐ�)0�Є�n��!�S`B�	u�7Cڧ��B�zu8�5�S`B�	u�=Cڧ��Bj� :��O�	�&�ti�
M����+Q�(�O�i�R�>&�P�b�1�}
L(4����cH��PhB�GBǐ�)0�Є�K��!�S`B�	�Æ�)0�Є�Æ�!�S`B�	��Cڧ��Bj� :��O�	�&ԾGti�
M�=�����e�Oih���>&�P{e�1�}
L(4����cH��PhB�QFǐ�)0�Є�_�a�}
L(4����cH��PhB�kGǐ�)0�|�0s�Y����ބ��g=s7�4���D�?�e��]�q��wh�����^���cN@k�7a����|۳\k�7����|k�\k&�w��0�Bk&�7���f�|/�\k&�wO��f�|����4k&�w�0-[3q�L�[����Ys��M��51����
Xs�cK��51�{��
�O�%r��H�����92WϚ��8r��9��"W�����&r��9��!W����r��8�� W����Mr��8oӟ+`��h��hv��L��L��L��Ll���Z3��fbk��֚��5[�k&��Ll���Y3��fbg��Κ��5�odb���Ie���8C{�.��:�������[Wz_4��AX�ˡ�]��㮨�u,��J�z롓6Ƹ��������X}����C��V��V/	����Jm��/��J?u�i�OL?m����Z��#E=V�`ѣE=^t��RG����(uD�#JQ�RG�:�����tD5��JGT:�����tD�#jQ�ZG��+����uD�#jQ�FG4:����h��#��FG4:"ꈨ#���:"�8�IGDuD���huD�#Z��VG�chuD�#Z��NGt:����H��V��S�˛��$��Hyt?������ӧ'U���Cb���$��^�s"���7�Z����z����S3\mo4��ȭ�k{�'�u�0>%�inn�'�b�;�7�������X�e����6�U�7��i�l��v1^Qʔ>�mSt�,��롭��2��Z��>��m��	��B�����������#4��'5��_�Ӑ�>��p<|�O��X���տ�K�;��?��z;�������{��?+��!���'�U���w�����������NO�m����n��>v������ݬ.O	3�E�����N����[ O{Br���o IB�p�۟���ׅ�����_��]վjR8��Oi�j]�w�*cQn�U�nJ)�wÐ�`#������'}�����1/��X���~�*eFz�����;��(��Us���ۋ�оz
�~|B����҈�4�^Q-�����Lw�D��D[.<�,���F�K#�|D��L
��Od��O����3������|��v�����q��.<Q.���F��'��G|C)������vz|�������oz�Z8~�&L�?�~><3O��'�I���<���'���T~�
KC��\<>S��G��&.<�.��F�aaD)K#��u<K��'����o��/���؞'���f��QU��i��I�ux��v���p|�p|�p�,�?��?�m�o���/���xg�Y�y��;;?�wv~Tx��᝝?�.�����������?����ۅ㛅���˅������};���������f���x7���+y���4�?���?U;����D��ðI/�?�L���%_�5ۋZ�W�ly����+7m%�t��6�b+�\�.Y�]�v����xm᫳�ޗ�u6�����j�UA���i�{����Y��w�:�,���/��
��6�����iĒ]���u���7]Qo�6��:TŶ��*��u�U�<b/r��{�����)��x"��S�������f�D�)�VU�P,��1.W�]|y��~sz�����ػ���wzd�¯�|>����p�n���>����t�������NY~�f�ӛ���oV�oVH����Y]�I���x�a��������(���<#�}-e�:��]�����H�����G�a?����ӻQ�ӛ7oVz��/�􉿎U�N�|���O�On��O�[���g�JU�쨷�߬>����~x~�����}@����7X�2H}ó�pY=}����3��0yI�h�����e���=���b**)�����o��s��n�xx����������W��PK   1�_U���R�$  �/  /   images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.png�xwT�[�/�E��@�HUHh�����KhbBK�EDDJT���T�f�Hiҥ�4�ҥ#��y�������u׺k�?γ����3�7{f�={�0�S��t�			������NBB:y��H���J?��̛��r@#9=|ݐ�H	����D'OU��S,�2[��s?Bë�	Or��z�����Q:� �5���O�?)�Ŀ��L�9E��yζjF(�u/l}]�]n��y����a��<MU��a��L�8�o�~r �?qN��,���L\y���['��w~�4Xm��6>�q|lμO}BX{���V	��~�����'��`p$&vL��EK��e��$Гm�J֒��:������j�s��@sV�G6f��o>:�/8��g�l����ڳg[ܷ:�J,�[ڝ�o1K��K�?��d��1�˂��wjq�Y�	٧q��Y/�^��>�u�C��-dZ}6�v�}gm�&[�b�!��_�ZӜ4��cS�����Nz:�kLA4A��[nkm�ܭ��ٽ[L՝�ae�ܥy'Gz��{���!�(�3��e�������~�0���'Sj�m�T"�l)c��8[�S��%P>�%�������f���m{��^�1�u|~���Y(c���#��J���jf�V���x������z ːHI�U��n�S�ć�	�4�(2��{����V0?X�V��on�	u^\rʫ�.���p�����'�w�b?�ܛo�R�w��}ՠ�>�%\��0o?�[���;�tZL)=�ks���}w ����u�P���+H%#I��'�X�wa��<��)�,�!;�@��iS0#�������S���9k��{؉��3{�U����Űi��ka
6�
Q��$��DSFkț>%�N�Gǲz:��)'uU�q����+0��7s9�v��kx��\�Av͠��
��[W�:��c��;��2�}�ž3S.��.�F���B*�'��v�*C�x�t�	����.��Nɑ�G*C����o'�[���w��\֐���ܳ>���XU��xf̙}��R:Cg�?ޮ�����#��m�1���`������79˼#�?��E�,e��`�$�"�}�ӑO�d��_w4�l>	���n?0u����=e���'e�r�;��eUV�Q�f��s�ndtÉt��h¹�ՑK�E�
n6硆 \��^�-=�ї��}���v�şV�ɴ�W��,n�Qfi%$�m�ݺw�ZR��@��.��8�bu�]Q3qI/\c�+[٫����hz'/���"�ތ5�B˜��O�7Wt��yP�G_{1�kR�$nB��y�)iV+�q\`G[�8�\Y,5�z���=���cg�wU�Kmù��g��ۼ�b>c1}��=���;��ObW}�`/ɛn�ԗ>�0{=�?������o���"��8N8�H-},&�}��ڧ��ע����P���>�����*�)�(��{�Z!��J�B=Ź��T/,m��Ge�K�M� r�*_F}���ñ�1uӘ˧�E�|�����0�3/MO�v��W�]��/V�tK52$;jq��OFZmjD�����#r�[< �%Ϧ�)C=�%YU��JlZ��T�gMS-��mR�,IȄ)�f_�&�f���8j?:�|<R�nx o>��rpК;�NJ�>4j��sI��}W3�[իb5�m�ޓ̆4p�����#�U{���`r�7B���Td93�_h�[N�`2R�ly�<9��ᔭ�����x��'���;����׸1/���:�s[�Tꚕ0j�P_I�B�K����T�շU-d>�1!�d�������`���a5�	��%-��Cxd�:Zw���eV`Q�aM�)��w�qC�A�M�3��樷�z�n��*�ƾ�I%���`��k���
��A�}ٮ6߱1]=7����G��7��L�����&#�uƓ]~��Hu���×��DV��G����"� ��+�ކ���_�M�(��pΣ{L-v$z���I�Z�ԏt�Z[pʏ�������&�����xJ�N�}��9�`r4���Aw �B��*�a�������])(�%��Mޖ������>y4���#tor�{6��s��רܲ�;EQ���F� c����OyuW�Q�>g�	��������K҇��"?����\|�rwѽ>�W�h�E�ɹA�]=5"��j���nL#]�Io�k��EdK��x�a��O~�.eg.01�0�u�6l ��������H5�/�+R�W�,Xŗ� ^����vV�����U�Y�'���׎���2������o�f0F�����@$GoK{P����F2�C]���>��3Ԕ3ߑ*j�˷l�%���A%̠� ���z|Jƺ}㶦�\E�ݖR�]�/�&�J���v~���'6�kn�r~wj|��>}�t��G:�%`�vG}��x����VoE�A/)���	���ŘJ�2�#��oH�_yQ�����]�)��8�S����(r��ȼ��C�7��;�gߨ�b.%��A��k)P�X���jJ�\F1L���w]�f�����ݵ�֮�K�־ǲ�Π��R)e��p�����S��F���g5�9���0d��>�ɞR��p�H�JUW�K~�{�R�~<�\H��͐b��9�������o���a9U�����WFk^7�R�H>�>���rwj7���nz�G��"1�𒅓���G�5/ɠ9�����AV]�߉0u��:��]�J��0o��7e���F���v��BO��d�?d���z]��yX��W(EW�"q��������g���'W�D�S4/_�Y}6Y6'�d�gu9���ΔhI
�or��t�qu�.�/�IY��kL��<�����+?�X����q$��(�P=�!q?GhH<�V��v�Qò�X�S���\6wGR��F��4�v�1�����|v�$z��Pee����~7����@QtN_0���z���B�xcaԔ��]A�GA�Y_�����u��������?�hb�-��p�Z��q����
'W�k�-�{� �^�A�d�.f�I�A����oCC8p���mج���\cO�f��֑��=��zwŉq���s��^�E�刏~�ڤ�e�]�)��|�~�?��������
��R��u������L�d�6�7:����4��Lڴ+Q�����i�܅�-���Ν��OC����&2R�����{su��%���*y _��j���A�fA�55*�pnR:�w7^SQ�YJ��8(.Ms8\��i5%�n!0�.q�-�G�XQb���[{8�'d�6��W��.�$�ߴ�=���n[ZQr��;������q�Fd?S�q\�xh ��b�kٹ�A����Q}8um@�$�>B���l&��FF��-��I�_aR����/bU�Ձ \��`v�p������#���C8!=8�H{y���:.N;y.s	]]7e�=?��O��焐��RT�$�!8#=`�>�h,�G��.�H�usq��p���p*�b���B�B" U/1.�K�r;�HE�bK�랇�DX���[�,䊱���%@X_���}�;�
��8�y8��p��apWOy.."���sv���'��/�!�svv��������5!��FH��'�T�B�xp�����n��/s��H4ҙ(�%b��E�����_\`����kq���p@�����8�&�_��ϖ���#��+��lz�*�\g�!v�;�/���AH��dP	��
�FI�A`I��BI �"��t�z�\�3(b��GZ!F�I�``;0H\R��J���0iQ1)1��� �1�]	C�yVgPvD(�$J
CJ�$$$DA�(II.#	B�a2`$�,.��e����b�a��tp��#��\�1��m�)�%&$�4�E@<.v����L����3�JJJ��E�R�"Ғ`i�	�!1X�^<C���-̙9D#`�������A�<\1&��hy�3γ��d�����@AE�� �"����D\���I�����?I�N��ݬ�%�������2F������v�����X@`��M�¼�v\a!��\���!��~��$$�E$đ 0�N���(���
$)e'!*�D"�ܿ�`]Q�0�=яD_w�/_q��c�n�U����w'�DE@r���
��Z9�����)ĜE.�?B1
�3������J�V򷒿����o%+��JɥSHb�M,�f�͘�e9\[]�W�E�S�*���pӰ����4��I[\��;/xh�^���qY��N%GB�H��r�������k�P�Ǎ�ٷ���x�6$�4��,Δ��TN]�5d��Cs���5���O��&�L���3�sO��S/�z��&)[�*�;P�h�s�'��f�������<l��"�l�޹Y]zE@7�Vn�zS���\�_�*���d*�U*p?M�+Z�����Ene mt.��)�RLJʻ�tbbB13�ٌM���U�	����k�{y2��K#��r���:!qn�>�t�'`4h�8��ɘ�h�4��A��P&A�责}�J1�,fUxτpw�i1,if��		��l���*4�iu���B�۞0��f��5'ǥK紀��мQ��������nyc~~���=�O�2?����H�h)oI��<���Iψt�{.����~y������
P;�����ֺ��\|��8�ł����-5�Ŀ}�۴i�n�tZv�`3���Z�Vin �ǝT�;���צ�H���lۏ�3�\�h�r���s`��ٴ4sʁ���Ecn�x�?��ǥ>�|�A]���S����v���|ٲ>�ǋQ	�s�l 9�o�n�@�=��ج���k紁���G�%�d�%�#"4>+{���ޣ��ʷ��n��%O�nj�P�ސ7}joiL�Ο�=�����<.�.���Y5=mv�7)�J�آ'�s�ٜ�S5A��S�uд�ɒKI��?53�\�>�Yn�<��I�L7��Re���S?���r`����{\9@9�_]]��(�5v���{����p�hS��Ʊ=��[��cE�:����Bc�#���Ȳ�FVE�}BF���5����ٗoV�7����<ud@1'�ǝv ��
�D��`W��&�F�<r�C���٪cen;�{�uo;��ʎF�	�#��^\h��R&�7�gV�ֻk��8���E8³N��m͗���1�����?��H��ٔ���i�[��_��8Ɖ-������\�d������!���Cd+Z�z��Џ:�~�8��,B�+켺��ɮ>�\����2�������b�Z��!�
ۡ��k�{t�
�KG��kޝ�
��b�sh����?F���]s��Oy��.��}���F��Mrx�w<�S"�+Z=uf���JzFo=�4��j�خx��E����jRlS����O�	�����f��Sq�ml�߿٨ur�������)uJ�޶+>����R�&�gVw�B+���gq�ŉv��F�6G��u�=.�vWo�EU7�l6�Um��ѕ�ӂpU,���8߈��:^�D��m� ����<�FO����l~´1}�u������W��1�q�~�X״�T�ï|*|1BSy�	M��4�e-eɍ�9�`QJ&ܱ���
���߭�o~-�׶i7=5���ݟK�'`�����f;�	� ι�n{�+���E��Q[#o|�Y#\9)�r�c�Ř����<���F��R͇٘F��.��&����R��n� eNx��2��Y�m/��u�N}	��3���h��H�Kn��3;������v=ab?��mhǇU���R�>i/�v !k�=��斋��aA-Z�[K�Z����MgO�b��a6_�_�n����1otnx�'�^*|Tڿ��q�0�h����bt�^����N�ڱ�iW�q8�Q%���k��ې���O��[á�4R�2S��̎o���ۦ��ծJV7D�t�A�KS`��騣�@��)��X�#.��e�ǃ�VS�t��J�(�H�(���ٵ��_u����(١L�:6��Kl��B`���0h)GE�o�C�KD��<WVy ��~_1?�����⍓ki	�hA��>���Hu��D߈|U\uYF�Jk�ӵv&0��Te$���,3�j|W�����5\�&*��R8g���(���rIV�������� LS��2�1 G�u����b�x��o�F��2��^��xt /��ɰU����ݣ���Nⴋ��y�:��]�I��7�)֐�RG_Ex��އ7�WOw̓c�oj�	�w �}/��oo߀���K�{��z�A�G"�����=�St8h��,'>v�[B�j�Ι#)��*�
��J�Ժ������8{.BW
�v%�3wf�R����:�z�� �Px�>�1w��\]_�ݘ~3h�@k��Z�˼��,�J��p:�EY�Pl���kq� ����K9ױˆ��־Q�G�IV�2w{Y���)��Ө&&��H~+�bk�?�[��6�2p�;i�6GQxS����{��ŷ]�ĔU2��m��iG'Bd2>6 �j9���8��˾t�.'���V>gF`ތԳA��5n^��\X����87툣�E|�o�����B�\힋J��3��K6�h#|���k�kP��6�0�	�%��$J�83�I��9�ɳ&�i��ӳ�����y���
1�"�$�l"O+Jn�h�cM�14���~1-TAv�>k6��6�[ZJ��cf�oy@N�s�ڃ
>5��{����M��Xe|����FU����k**���qOǦ�Ve�kF>IR����@��pW�Eo��ճ[�^`���זk|�]~�S�@l3�枇x�K����5���3���p?�����4�\�C>��a��v/+�ɵ��Eɰ��x����pfF�b��L�	2���_҈x$���`p�[@t��c:��� *�xgf«lw#�2Xv���,�&����O�}FhK�pQ�Z(���}i�&0�}���1�ݙ��Q��8�W�s��e6�/v�tj�(6�������P�H߈�o!���s� C�AF����d�q�t�Cu�"�95ܧ&g�u��5ߎ����QK1�䣇c��	�Ў��[�~+�>4��y{8ۈO�'�i����^��E��^0��5���tUgh�~�?��|�nQ�D�Z#i]���fLBD��_{����w�5M�����@bֱ��ղV�A�!U��o�-��Q��*�R�[O΢k���$�或������tGG��Wh�IR֘Xq���I^��x�lu�;q��ʹ_�PssQ|u�Jx|�PL?PIa��Zγ���[,�����Ws`RGl\_�	����{�;�~�?Z�m]��r�XR	���Y+��F�ιO��=��?ֵ��O�c6�TY�TdF��Qޛ˗��J6i�#�:bL���0�ey�{��d��K�im��a�y?//��4���b�'>���Լ��}�)T~o�%+�#��Ot�����Q�$�#Q֨�Z���g��1��Y@S����:뼛(�A��4��ؿ��-+%���A(���5 �	S$�i�Ѷ	���Ly�+.>�b��5��x��	�E��ј`(���j����>-.�m�X
**��ȶ�������O�do�U~t��z��2���Wx�ֱ '�eܥ ��v� 5�$D��|}G�|��Ec�[rˌd
[(�����e�I@���X�0 s�kD�$��}s�s��.@�=�a����%�d;ތ \��� S�;��G��R�=#ޤ��+����g�PXȋ�HG�UR�1�A����N��ϛ���t�!I<�x�D��e�1�-ª�ౖ�}⥨\��YO(y�h^ѭ�zM�ޚ�ˎ�g�%��8�+������_���+��c�������kHد�����Mz����3z\��AKޭ��{-z-:'T��������X�� ��S�����
��g�Y�at8>H{���ep�����o�-%�j�������}��	�1��^�/\����I{_e���bn�Q%����!iL9�/j�V���6�Oܯ�iW��T�����/rs���e�ݔ�͓ٷ��X*qjՀ�09��ӂ�r2yoQ�����	�����$�Fb"6c[�cH�������ik��Ҹ�'�!���9�u{N	����N��u�ǎ&ZtuN��M�)$�˧E���=��Lk��[**�G��ς+`���M	��g�2�Ï���"+eX£�(4VR��f�������m�
2È���eB�~�M�Q�O�qeV�Ӏ���oV��v\���	�l b��;��k��
��\֜��SG�e����ڎ���)���2�~{�X�x�~����9�C��4'��#��c�uKv"M.����~���������d��4}S0V�.\�F����A�8�˻�5�.'�F7��;ت#:�ɭ�� �r�����[U��� E�я�E�3�Ap����rS������xŴ����)�^��.y�h��hܻmⰮY�?��M	�y7�d~���C��Ïɮ𑚳p���o��'[s�"*А��a
"�{VĐ��5!�����n�O���X�˽����W\�3���m�u���՚GJ�]�����i�u+�X~��1FR+�.�<>��ܗ�D`~�7������iܵ��"T/�(?�2s�m��4�_v�S����Y�x@�x*�{Hc���t^�X�=�P���G��w'���5�E�O/�9;��6�A�-��(�JYf(�j6��9m�U�����[��R���w䆗����6�vA�Aݬ 8\U�'�]�|c�G¢�g�3���u�t ����pP3��?:�6" �c��j�̽�g~	���D��#��;n��~�?�m���o5�%��`]d�� (�4��|.dzHOɐUUs�%���k�/�움f���� ��F\�2Q<Xvw����*��mm�Y��zWu�O��	3+�)m�����3���3S����wM��½�̗v|�/�qgh-�֗G	K>@�����q|�Bn;���3�W��"�Qk�̯4�+N+������6�E�g ���4P��mO�#T\��6?�}���պ"���p�+�=�� H�=*Yz��5Y�8��u��T���z0i#T�$*�}AaϢ��1f���"T�[�|��
u*�t,3ɤ��W�/C�d�M8�ļW8kk��(�}�� PK   JvqU!T��-  R     jsons/user_defined.json��AO�0��
ʹ��6eko�]vBNhBM�K]R������qVƄ�Ip��ޗg����V�ށ}SP���	֡�Ԉ�8�Tq��RǊ����P�w5��%������a/�Y|7CE�$�R	��<V�P�T���4!e��\���8>��Zt�����*�m7e;�z�����[򵨗�6�80���ڦ�MC�1�3�R�[k��-��,�M�i�Ə��z�,���ơϹ*�q��|�,�D�=ݝ�ލ%�i̦���l.��u�������bo�����ҚG*Yӂ��xc����u܌_PK
   JvqU%V�  �Q                  cirkitFile.jsonPK
   1�_U���R�$  �/  /             �  images/29bbd443-10d8-4ebd-b903-e4bb25b9bd96.pngPK
   JvqU!T��-  R               �D  jsons/user_defined.jsonPK      �   SF    